magic
tech gf180mcuD
magscale 1 10
timestamp 1702247546
<< metal1 >>
rect 13458 57038 13470 57090
rect 13522 57087 13534 57090
rect 14578 57087 14590 57090
rect 13522 57041 14590 57087
rect 13522 57038 13534 57041
rect 14578 57038 14590 57041
rect 14642 57038 14654 57090
rect 27122 57038 27134 57090
rect 27186 57087 27198 57090
rect 28354 57087 28366 57090
rect 27186 57041 28366 57087
rect 27186 57038 27198 57041
rect 28354 57038 28366 57041
rect 28418 57038 28430 57090
rect 1344 56474 48608 56508
rect 1344 56422 19838 56474
rect 19890 56422 19942 56474
rect 19994 56422 20046 56474
rect 20098 56422 48608 56474
rect 1344 56388 48608 56422
rect 3838 56306 3890 56318
rect 3838 56242 3890 56254
rect 5518 56306 5570 56318
rect 5518 56242 5570 56254
rect 6974 56306 7026 56318
rect 6974 56242 7026 56254
rect 8542 56306 8594 56318
rect 8542 56242 8594 56254
rect 10110 56306 10162 56318
rect 10110 56242 10162 56254
rect 11678 56306 11730 56318
rect 11678 56242 11730 56254
rect 12574 56306 12626 56318
rect 12574 56242 12626 56254
rect 13470 56306 13522 56318
rect 13470 56242 13522 56254
rect 15374 56306 15426 56318
rect 15374 56242 15426 56254
rect 22094 56306 22146 56318
rect 22094 56242 22146 56254
rect 27470 56306 27522 56318
rect 27470 56242 27522 56254
rect 28366 56306 28418 56318
rect 28366 56242 28418 56254
rect 40798 56306 40850 56318
rect 40798 56242 40850 56254
rect 44606 56306 44658 56318
rect 44606 56242 44658 56254
rect 47406 56306 47458 56318
rect 47406 56242 47458 56254
rect 42814 56194 42866 56206
rect 25330 56142 25342 56194
rect 25394 56142 25406 56194
rect 42814 56130 42866 56142
rect 47854 56082 47906 56094
rect 16034 56030 16046 56082
rect 16098 56030 16110 56082
rect 16930 56030 16942 56082
rect 16994 56030 17006 56082
rect 21074 56030 21086 56082
rect 21138 56030 21150 56082
rect 27122 56030 27134 56082
rect 27186 56030 27198 56082
rect 31602 56030 31614 56082
rect 31666 56030 31678 56082
rect 35074 56030 35086 56082
rect 35138 56030 35150 56082
rect 38770 56030 38782 56082
rect 38834 56030 38846 56082
rect 39778 56030 39790 56082
rect 39842 56030 39854 56082
rect 43810 56030 43822 56082
rect 43874 56030 43886 56082
rect 46834 56030 46846 56082
rect 46898 56030 46910 56082
rect 47618 56030 47630 56082
rect 47682 56030 47694 56082
rect 47854 56018 47906 56030
rect 48190 56082 48242 56094
rect 48190 56018 48242 56030
rect 42926 55970 42978 55982
rect 17714 55918 17726 55970
rect 17778 55918 17790 55970
rect 19842 55918 19854 55970
rect 19906 55918 19918 55970
rect 30146 55918 30158 55970
rect 30210 55918 30222 55970
rect 32162 55918 32174 55970
rect 32226 55918 32238 55970
rect 34290 55918 34302 55970
rect 34354 55918 34366 55970
rect 35970 55918 35982 55970
rect 36034 55918 36046 55970
rect 38098 55918 38110 55970
rect 38162 55918 38174 55970
rect 42926 55906 42978 55918
rect 43038 55858 43090 55870
rect 43038 55794 43090 55806
rect 46510 55858 46562 55870
rect 46510 55794 46562 55806
rect 46846 55858 46898 55870
rect 47618 55806 47630 55858
rect 47682 55806 47694 55858
rect 46846 55794 46898 55806
rect 1344 55690 48608 55724
rect 1344 55638 4478 55690
rect 4530 55638 4582 55690
rect 4634 55638 4686 55690
rect 4738 55638 35198 55690
rect 35250 55638 35302 55690
rect 35354 55638 35406 55690
rect 35458 55638 48608 55690
rect 1344 55604 48608 55638
rect 22206 55522 22258 55534
rect 22206 55458 22258 55470
rect 34190 55410 34242 55422
rect 43598 55410 43650 55422
rect 17490 55358 17502 55410
rect 17554 55358 17566 55410
rect 20738 55358 20750 55410
rect 20802 55358 20814 55410
rect 27010 55358 27022 55410
rect 27074 55358 27086 55410
rect 32834 55358 32846 55410
rect 32898 55358 32910 55410
rect 42018 55358 42030 55410
rect 42082 55358 42094 55410
rect 45266 55358 45278 55410
rect 45330 55358 45342 55410
rect 47394 55358 47406 55410
rect 47458 55358 47470 55410
rect 34190 55346 34242 55358
rect 43598 55346 43650 55358
rect 9662 55298 9714 55310
rect 13806 55298 13858 55310
rect 23438 55298 23490 55310
rect 36878 55298 36930 55310
rect 9874 55246 9886 55298
rect 9938 55246 9950 55298
rect 10770 55246 10782 55298
rect 10834 55246 10846 55298
rect 14578 55246 14590 55298
rect 14642 55246 14654 55298
rect 17938 55246 17950 55298
rect 18002 55246 18014 55298
rect 22866 55246 22878 55298
rect 22930 55246 22942 55298
rect 24098 55246 24110 55298
rect 24162 55246 24174 55298
rect 30034 55246 30046 55298
rect 30098 55246 30110 55298
rect 33170 55246 33182 55298
rect 33234 55246 33246 55298
rect 9662 55234 9714 55246
rect 13806 55234 13858 55246
rect 23438 55234 23490 55246
rect 36878 55234 36930 55246
rect 37214 55298 37266 55310
rect 38446 55298 38498 55310
rect 42702 55298 42754 55310
rect 37986 55246 37998 55298
rect 38050 55246 38062 55298
rect 39106 55246 39118 55298
rect 39170 55246 39182 55298
rect 37214 55234 37266 55246
rect 38446 55234 38498 55246
rect 42702 55234 42754 55246
rect 43374 55298 43426 55310
rect 44034 55246 44046 55298
rect 44098 55246 44110 55298
rect 48066 55246 48078 55298
rect 48130 55246 48142 55298
rect 43374 55234 43426 55246
rect 9326 55186 9378 55198
rect 11678 55186 11730 55198
rect 10098 55134 10110 55186
rect 10162 55134 10174 55186
rect 9326 55122 9378 55134
rect 11678 55122 11730 55134
rect 13470 55186 13522 55198
rect 13470 55122 13522 55134
rect 14030 55186 14082 55198
rect 21870 55186 21922 55198
rect 15362 55134 15374 55186
rect 15426 55134 15438 55186
rect 18610 55134 18622 55186
rect 18674 55134 18686 55186
rect 14030 55122 14082 55134
rect 21870 55122 21922 55134
rect 22318 55186 22370 55198
rect 22318 55122 22370 55134
rect 23102 55186 23154 55198
rect 23102 55122 23154 55134
rect 23774 55186 23826 55198
rect 27582 55186 27634 55198
rect 24882 55134 24894 55186
rect 24946 55134 24958 55186
rect 23774 55122 23826 55134
rect 27582 55122 27634 55134
rect 28030 55186 28082 55198
rect 28030 55122 28082 55134
rect 28366 55186 28418 55198
rect 28366 55122 28418 55134
rect 28590 55186 28642 55198
rect 28590 55122 28642 55134
rect 29150 55186 29202 55198
rect 36206 55186 36258 55198
rect 30706 55134 30718 55186
rect 30770 55134 30782 55186
rect 29150 55122 29202 55134
rect 36206 55122 36258 55134
rect 36318 55186 36370 55198
rect 36318 55122 36370 55134
rect 37550 55186 37602 55198
rect 43038 55186 43090 55198
rect 39890 55134 39902 55186
rect 39954 55134 39966 55186
rect 37550 55122 37602 55134
rect 43038 55122 43090 55134
rect 44942 55186 44994 55198
rect 44942 55122 44994 55134
rect 9438 55074 9490 55086
rect 11454 55074 11506 55086
rect 10882 55022 10894 55074
rect 10946 55022 10958 55074
rect 9438 55010 9490 55022
rect 11454 55010 11506 55022
rect 11566 55074 11618 55086
rect 11566 55010 11618 55022
rect 12238 55074 12290 55086
rect 12238 55010 12290 55022
rect 13694 55074 13746 55086
rect 13694 55010 13746 55022
rect 22206 55074 22258 55086
rect 22206 55010 22258 55022
rect 22542 55074 22594 55086
rect 22542 55010 22594 55022
rect 22654 55074 22706 55086
rect 22654 55010 22706 55022
rect 23662 55074 23714 55086
rect 23662 55010 23714 55022
rect 27246 55074 27298 55086
rect 27246 55010 27298 55022
rect 27470 55074 27522 55086
rect 27470 55010 27522 55022
rect 28254 55074 28306 55086
rect 28254 55010 28306 55022
rect 36542 55074 36594 55086
rect 36542 55010 36594 55022
rect 37102 55074 37154 55086
rect 37102 55010 37154 55022
rect 42478 55074 42530 55086
rect 42478 55010 42530 55022
rect 42590 55074 42642 55086
rect 42590 55010 42642 55022
rect 43710 55074 43762 55086
rect 43710 55010 43762 55022
rect 44270 55074 44322 55086
rect 44270 55010 44322 55022
rect 44830 55074 44882 55086
rect 44830 55010 44882 55022
rect 1344 54906 48608 54940
rect 1344 54854 19838 54906
rect 19890 54854 19942 54906
rect 19994 54854 20046 54906
rect 20098 54854 48608 54906
rect 1344 54820 48608 54854
rect 18622 54738 18674 54750
rect 11666 54686 11678 54738
rect 11730 54686 11742 54738
rect 18622 54674 18674 54686
rect 39342 54738 39394 54750
rect 39342 54674 39394 54686
rect 40238 54738 40290 54750
rect 40238 54674 40290 54686
rect 41246 54738 41298 54750
rect 41246 54674 41298 54686
rect 45726 54738 45778 54750
rect 45726 54674 45778 54686
rect 48190 54738 48242 54750
rect 48190 54674 48242 54686
rect 41022 54626 41074 54638
rect 6850 54574 6862 54626
rect 6914 54574 6926 54626
rect 9874 54574 9886 54626
rect 9938 54574 9950 54626
rect 13906 54574 13918 54626
rect 13970 54574 13982 54626
rect 30146 54574 30158 54626
rect 30210 54574 30222 54626
rect 37090 54574 37102 54626
rect 37154 54574 37166 54626
rect 43586 54574 43598 54626
rect 43650 54574 43662 54626
rect 41022 54562 41074 54574
rect 39230 54514 39282 54526
rect 6178 54462 6190 54514
rect 6242 54462 6254 54514
rect 10322 54462 10334 54514
rect 10386 54462 10398 54514
rect 11106 54462 11118 54514
rect 11170 54462 11182 54514
rect 12786 54462 12798 54514
rect 12850 54462 12862 54514
rect 13122 54462 13134 54514
rect 13186 54462 13198 54514
rect 19058 54462 19070 54514
rect 19122 54462 19134 54514
rect 22530 54462 22542 54514
rect 22594 54462 22606 54514
rect 23874 54462 23886 54514
rect 23938 54462 23950 54514
rect 25778 54462 25790 54514
rect 25842 54462 25854 54514
rect 27122 54462 27134 54514
rect 27186 54462 27198 54514
rect 30930 54462 30942 54514
rect 30994 54462 31006 54514
rect 35858 54462 35870 54514
rect 35922 54462 35934 54514
rect 38658 54462 38670 54514
rect 38722 54462 38734 54514
rect 39230 54450 39282 54462
rect 39454 54514 39506 54526
rect 39454 54450 39506 54462
rect 39678 54514 39730 54526
rect 39678 54450 39730 54462
rect 40910 54514 40962 54526
rect 47854 54514 47906 54526
rect 44258 54462 44270 54514
rect 44322 54462 44334 54514
rect 44706 54462 44718 54514
rect 44770 54462 44782 54514
rect 40910 54450 40962 54462
rect 47854 54450 47906 54462
rect 12574 54402 12626 54414
rect 16494 54402 16546 54414
rect 8978 54350 8990 54402
rect 9042 54350 9054 54402
rect 16034 54350 16046 54402
rect 16098 54350 16110 54402
rect 12574 54338 12626 54350
rect 16494 54338 16546 54350
rect 17726 54402 17778 54414
rect 17726 54338 17778 54350
rect 18286 54402 18338 54414
rect 18286 54338 18338 54350
rect 18734 54402 18786 54414
rect 26238 54402 26290 54414
rect 27694 54402 27746 54414
rect 31390 54402 31442 54414
rect 19842 54350 19854 54402
rect 19906 54350 19918 54402
rect 21970 54350 21982 54402
rect 22034 54350 22046 54402
rect 22642 54350 22654 54402
rect 22706 54350 22718 54402
rect 25442 54350 25454 54402
rect 25506 54350 25518 54402
rect 26898 54350 26910 54402
rect 26962 54350 26974 54402
rect 28018 54350 28030 54402
rect 28082 54350 28094 54402
rect 18734 54338 18786 54350
rect 26238 54338 26290 54350
rect 27694 54338 27746 54350
rect 31390 54338 31442 54350
rect 31838 54402 31890 54414
rect 31838 54338 31890 54350
rect 32510 54402 32562 54414
rect 40350 54402 40402 54414
rect 33058 54350 33070 54402
rect 33122 54350 33134 54402
rect 35186 54350 35198 54402
rect 35250 54350 35262 54402
rect 41458 54350 41470 54402
rect 41522 54350 41534 54402
rect 32510 54338 32562 54350
rect 40350 54338 40402 54350
rect 12462 54290 12514 54302
rect 24098 54238 24110 54290
rect 24162 54238 24174 54290
rect 12462 54226 12514 54238
rect 1344 54122 48608 54156
rect 1344 54070 4478 54122
rect 4530 54070 4582 54122
rect 4634 54070 4686 54122
rect 4738 54070 35198 54122
rect 35250 54070 35302 54122
rect 35354 54070 35406 54122
rect 35458 54070 48608 54122
rect 1344 54036 48608 54070
rect 10334 53954 10386 53966
rect 10334 53890 10386 53902
rect 16046 53954 16098 53966
rect 16046 53890 16098 53902
rect 22990 53954 23042 53966
rect 22990 53890 23042 53902
rect 23326 53954 23378 53966
rect 23326 53890 23378 53902
rect 9662 53842 9714 53854
rect 9662 53778 9714 53790
rect 10222 53842 10274 53854
rect 10222 53778 10274 53790
rect 14030 53842 14082 53854
rect 24222 53842 24274 53854
rect 21858 53790 21870 53842
rect 21922 53790 21934 53842
rect 14030 53778 14082 53790
rect 24222 53778 24274 53790
rect 25118 53842 25170 53854
rect 25118 53778 25170 53790
rect 27694 53842 27746 53854
rect 27694 53778 27746 53790
rect 29262 53842 29314 53854
rect 41346 53790 41358 53842
rect 41410 53790 41422 53842
rect 45266 53790 45278 53842
rect 45330 53790 45342 53842
rect 29262 53778 29314 53790
rect 14702 53730 14754 53742
rect 24334 53730 24386 53742
rect 9986 53678 9998 53730
rect 10050 53678 10062 53730
rect 12226 53678 12238 53730
rect 12290 53678 12302 53730
rect 16034 53678 16046 53730
rect 16098 53678 16110 53730
rect 17938 53678 17950 53730
rect 18002 53678 18014 53730
rect 22194 53678 22206 53730
rect 22258 53678 22270 53730
rect 14702 53666 14754 53678
rect 24334 53666 24386 53678
rect 24782 53730 24834 53742
rect 24782 53666 24834 53678
rect 25342 53730 25394 53742
rect 25342 53666 25394 53678
rect 25566 53730 25618 53742
rect 25566 53666 25618 53678
rect 26014 53730 26066 53742
rect 26014 53666 26066 53678
rect 26126 53730 26178 53742
rect 28030 53730 28082 53742
rect 27234 53678 27246 53730
rect 27298 53678 27310 53730
rect 26126 53666 26178 53678
rect 28030 53666 28082 53678
rect 29150 53730 29202 53742
rect 29150 53666 29202 53678
rect 32958 53730 33010 53742
rect 37214 53730 37266 53742
rect 33618 53678 33630 53730
rect 33682 53678 33694 53730
rect 32958 53666 33010 53678
rect 37214 53666 37266 53678
rect 37326 53730 37378 53742
rect 44942 53730 44994 53742
rect 37650 53678 37662 53730
rect 37714 53678 37726 53730
rect 38434 53678 38446 53730
rect 38498 53678 38510 53730
rect 39218 53678 39230 53730
rect 39282 53678 39294 53730
rect 41682 53678 41694 53730
rect 41746 53678 41758 53730
rect 47394 53678 47406 53730
rect 47458 53678 47470 53730
rect 48066 53678 48078 53730
rect 48130 53678 48142 53730
rect 37326 53666 37378 53678
rect 44942 53666 44994 53678
rect 9550 53618 9602 53630
rect 14142 53618 14194 53630
rect 10882 53566 10894 53618
rect 10946 53566 10958 53618
rect 12450 53566 12462 53618
rect 12514 53566 12526 53618
rect 9550 53554 9602 53566
rect 14142 53554 14194 53566
rect 14926 53618 14978 53630
rect 14926 53554 14978 53566
rect 15038 53618 15090 53630
rect 15038 53554 15090 53566
rect 16382 53618 16434 53630
rect 22430 53618 22482 53630
rect 22082 53566 22094 53618
rect 22146 53566 22158 53618
rect 16382 53554 16434 53566
rect 22430 53554 22482 53566
rect 23774 53618 23826 53630
rect 23774 53554 23826 53566
rect 25006 53618 25058 53630
rect 25006 53554 25058 53566
rect 27582 53618 27634 53630
rect 27582 53554 27634 53566
rect 28254 53618 28306 53630
rect 28254 53554 28306 53566
rect 28366 53618 28418 53630
rect 28366 53554 28418 53566
rect 30830 53618 30882 53630
rect 30830 53554 30882 53566
rect 31054 53618 31106 53630
rect 31054 53554 31106 53566
rect 31390 53618 31442 53630
rect 31390 53554 31442 53566
rect 37438 53618 37490 53630
rect 37438 53554 37490 53566
rect 9214 53506 9266 53518
rect 13582 53506 13634 53518
rect 10994 53454 11006 53506
rect 11058 53454 11070 53506
rect 9214 53442 9266 53454
rect 13582 53442 13634 53454
rect 13918 53506 13970 53518
rect 13918 53442 13970 53454
rect 14366 53506 14418 53518
rect 14366 53442 14418 53454
rect 15598 53506 15650 53518
rect 15598 53442 15650 53454
rect 18958 53506 19010 53518
rect 18958 53442 19010 53454
rect 21646 53506 21698 53518
rect 21646 53442 21698 53454
rect 22654 53506 22706 53518
rect 22654 53442 22706 53454
rect 23102 53506 23154 53518
rect 23102 53442 23154 53454
rect 24110 53506 24162 53518
rect 24110 53442 24162 53454
rect 25902 53506 25954 53518
rect 25902 53442 25954 53454
rect 26350 53506 26402 53518
rect 26350 53442 26402 53454
rect 27022 53506 27074 53518
rect 27022 53442 27074 53454
rect 27806 53506 27858 53518
rect 27806 53442 27858 53454
rect 29374 53506 29426 53518
rect 29374 53442 29426 53454
rect 29598 53506 29650 53518
rect 29598 53442 29650 53454
rect 30270 53506 30322 53518
rect 30270 53442 30322 53454
rect 31278 53506 31330 53518
rect 31278 53442 31330 53454
rect 33294 53506 33346 53518
rect 33294 53442 33346 53454
rect 34638 53506 34690 53518
rect 34638 53442 34690 53454
rect 37102 53506 37154 53518
rect 37102 53442 37154 53454
rect 38110 53506 38162 53518
rect 38110 53442 38162 53454
rect 42702 53506 42754 53518
rect 42702 53442 42754 53454
rect 1344 53338 48608 53372
rect 1344 53286 19838 53338
rect 19890 53286 19942 53338
rect 19994 53286 20046 53338
rect 20098 53286 48608 53338
rect 1344 53252 48608 53286
rect 15822 53170 15874 53182
rect 15822 53106 15874 53118
rect 16382 53170 16434 53182
rect 16382 53106 16434 53118
rect 20526 53170 20578 53182
rect 20526 53106 20578 53118
rect 22542 53170 22594 53182
rect 22542 53106 22594 53118
rect 23214 53170 23266 53182
rect 23214 53106 23266 53118
rect 23438 53170 23490 53182
rect 23438 53106 23490 53118
rect 24222 53170 24274 53182
rect 24222 53106 24274 53118
rect 25790 53170 25842 53182
rect 25790 53106 25842 53118
rect 27470 53170 27522 53182
rect 27470 53106 27522 53118
rect 37438 53170 37490 53182
rect 39454 53170 39506 53182
rect 38994 53118 39006 53170
rect 39058 53118 39070 53170
rect 37438 53106 37490 53118
rect 39454 53106 39506 53118
rect 41918 53170 41970 53182
rect 41918 53106 41970 53118
rect 45614 53170 45666 53182
rect 45614 53106 45666 53118
rect 7422 53058 7474 53070
rect 23102 53058 23154 53070
rect 12002 53006 12014 53058
rect 12066 53006 12078 53058
rect 7422 52994 7474 53006
rect 23102 52994 23154 53006
rect 29374 53058 29426 53070
rect 29374 52994 29426 53006
rect 31726 53058 31778 53070
rect 34290 53006 34302 53058
rect 34354 53006 34366 53058
rect 38210 53006 38222 53058
rect 38274 53006 38286 53058
rect 31726 52994 31778 53006
rect 7198 52946 7250 52958
rect 4162 52894 4174 52946
rect 4226 52894 4238 52946
rect 7198 52882 7250 52894
rect 7534 52946 7586 52958
rect 7534 52882 7586 52894
rect 7982 52946 8034 52958
rect 15374 52946 15426 52958
rect 11218 52894 11230 52946
rect 11282 52894 11294 52946
rect 7982 52882 8034 52894
rect 15374 52882 15426 52894
rect 15710 52946 15762 52958
rect 15710 52882 15762 52894
rect 16046 52946 16098 52958
rect 16046 52882 16098 52894
rect 16270 52946 16322 52958
rect 16270 52882 16322 52894
rect 16494 52946 16546 52958
rect 22430 52946 22482 52958
rect 16818 52894 16830 52946
rect 16882 52894 16894 52946
rect 19618 52894 19630 52946
rect 19682 52894 19694 52946
rect 16494 52882 16546 52894
rect 22430 52882 22482 52894
rect 25342 52946 25394 52958
rect 25342 52882 25394 52894
rect 29262 52946 29314 52958
rect 29262 52882 29314 52894
rect 29598 52946 29650 52958
rect 36206 52946 36258 52958
rect 31042 52894 31054 52946
rect 31106 52894 31118 52946
rect 35186 52894 35198 52946
rect 35250 52894 35262 52946
rect 29598 52882 29650 52894
rect 36206 52882 36258 52894
rect 36766 52946 36818 52958
rect 36766 52882 36818 52894
rect 36990 52946 37042 52958
rect 36990 52882 37042 52894
rect 37662 52946 37714 52958
rect 40014 52946 40066 52958
rect 37986 52894 37998 52946
rect 38050 52894 38062 52946
rect 38882 52894 38894 52946
rect 38946 52894 38958 52946
rect 41346 52894 41358 52946
rect 41410 52894 41422 52946
rect 44594 52894 44606 52946
rect 44658 52894 44670 52946
rect 47954 52894 47966 52946
rect 48018 52894 48030 52946
rect 37662 52882 37714 52894
rect 40014 52882 40066 52894
rect 14590 52834 14642 52846
rect 4834 52782 4846 52834
rect 4898 52782 4910 52834
rect 6962 52782 6974 52834
rect 7026 52782 7038 52834
rect 14130 52782 14142 52834
rect 14194 52782 14206 52834
rect 14590 52770 14642 52782
rect 17502 52834 17554 52846
rect 17502 52770 17554 52782
rect 23774 52834 23826 52846
rect 33854 52834 33906 52846
rect 30818 52782 30830 52834
rect 30882 52782 30894 52834
rect 23774 52770 23826 52782
rect 33854 52770 33906 52782
rect 35870 52834 35922 52846
rect 35870 52770 35922 52782
rect 37550 52834 37602 52846
rect 37550 52770 37602 52782
rect 43822 52834 43874 52846
rect 47518 52834 47570 52846
rect 44146 52782 44158 52834
rect 44210 52782 44222 52834
rect 43822 52770 43874 52782
rect 47518 52770 47570 52782
rect 22542 52722 22594 52734
rect 23762 52670 23774 52722
rect 23826 52719 23838 52722
rect 24098 52719 24110 52722
rect 23826 52673 24110 52719
rect 23826 52670 23838 52673
rect 24098 52670 24110 52673
rect 24162 52670 24174 52722
rect 22542 52658 22594 52670
rect 1344 52554 48608 52588
rect 1344 52502 4478 52554
rect 4530 52502 4582 52554
rect 4634 52502 4686 52554
rect 4738 52502 35198 52554
rect 35250 52502 35302 52554
rect 35354 52502 35406 52554
rect 35458 52502 48608 52554
rect 1344 52468 48608 52502
rect 6750 52386 6802 52398
rect 6750 52322 6802 52334
rect 27358 52386 27410 52398
rect 27358 52322 27410 52334
rect 38670 52386 38722 52398
rect 38670 52322 38722 52334
rect 39678 52386 39730 52398
rect 39678 52322 39730 52334
rect 46622 52386 46674 52398
rect 46622 52322 46674 52334
rect 6078 52274 6130 52286
rect 6078 52210 6130 52222
rect 7646 52274 7698 52286
rect 7646 52210 7698 52222
rect 8206 52274 8258 52286
rect 8206 52210 8258 52222
rect 8990 52274 9042 52286
rect 11118 52274 11170 52286
rect 34750 52274 34802 52286
rect 10322 52222 10334 52274
rect 10386 52222 10398 52274
rect 15474 52222 15486 52274
rect 15538 52222 15550 52274
rect 25218 52222 25230 52274
rect 25282 52222 25294 52274
rect 26786 52222 26798 52274
rect 26850 52222 26862 52274
rect 31602 52222 31614 52274
rect 31666 52222 31678 52274
rect 8990 52210 9042 52222
rect 11118 52210 11170 52222
rect 34750 52210 34802 52222
rect 35534 52274 35586 52286
rect 35534 52210 35586 52222
rect 36430 52274 36482 52286
rect 36430 52210 36482 52222
rect 38558 52274 38610 52286
rect 38558 52210 38610 52222
rect 5966 52162 6018 52174
rect 5966 52098 6018 52110
rect 6862 52162 6914 52174
rect 14030 52162 14082 52174
rect 22654 52162 22706 52174
rect 7186 52110 7198 52162
rect 7250 52110 7262 52162
rect 9650 52110 9662 52162
rect 9714 52110 9726 52162
rect 17602 52110 17614 52162
rect 17666 52110 17678 52162
rect 18274 52110 18286 52162
rect 18338 52110 18350 52162
rect 20066 52110 20078 52162
rect 20130 52110 20142 52162
rect 22306 52110 22318 52162
rect 22370 52110 22382 52162
rect 6862 52098 6914 52110
rect 14030 52098 14082 52110
rect 22654 52098 22706 52110
rect 23326 52162 23378 52174
rect 24222 52162 24274 52174
rect 29262 52162 29314 52174
rect 30158 52162 30210 52174
rect 23538 52110 23550 52162
rect 23602 52110 23614 52162
rect 26450 52110 26462 52162
rect 26514 52110 26526 52162
rect 27234 52110 27246 52162
rect 27298 52110 27310 52162
rect 29474 52110 29486 52162
rect 29538 52110 29550 52162
rect 23326 52098 23378 52110
rect 24222 52098 24274 52110
rect 29262 52098 29314 52110
rect 30158 52098 30210 52110
rect 30830 52162 30882 52174
rect 32286 52162 32338 52174
rect 31378 52110 31390 52162
rect 31442 52110 31454 52162
rect 30830 52098 30882 52110
rect 32286 52098 32338 52110
rect 32734 52162 32786 52174
rect 35646 52162 35698 52174
rect 32946 52110 32958 52162
rect 33010 52110 33022 52162
rect 35074 52110 35086 52162
rect 35138 52110 35150 52162
rect 32734 52098 32786 52110
rect 35646 52098 35698 52110
rect 37102 52162 37154 52174
rect 39118 52162 39170 52174
rect 41694 52162 41746 52174
rect 37426 52110 37438 52162
rect 37490 52110 37502 52162
rect 38322 52110 38334 52162
rect 38386 52110 38398 52162
rect 40450 52110 40462 52162
rect 40514 52110 40526 52162
rect 41234 52110 41246 52162
rect 41298 52110 41310 52162
rect 37102 52098 37154 52110
rect 39118 52098 39170 52110
rect 41694 52098 41746 52110
rect 42478 52162 42530 52174
rect 44258 52110 44270 52162
rect 44322 52110 44334 52162
rect 45602 52110 45614 52162
rect 45666 52110 45678 52162
rect 42478 52098 42530 52110
rect 5630 52050 5682 52062
rect 5630 51986 5682 51998
rect 6190 52050 6242 52062
rect 6190 51986 6242 51998
rect 9326 52050 9378 52062
rect 9326 51986 9378 51998
rect 10446 52050 10498 52062
rect 10446 51986 10498 51998
rect 10670 52050 10722 52062
rect 10670 51986 10722 51998
rect 19630 52050 19682 52062
rect 19630 51986 19682 51998
rect 19742 52050 19794 52062
rect 19742 51986 19794 51998
rect 20414 52050 20466 52062
rect 20414 51986 20466 51998
rect 25342 52050 25394 52062
rect 25342 51986 25394 51998
rect 25566 52050 25618 52062
rect 25566 51986 25618 51998
rect 33630 52050 33682 52062
rect 33630 51986 33682 51998
rect 36990 52050 37042 52062
rect 36990 51986 37042 51998
rect 39790 52050 39842 52062
rect 43486 52050 43538 52062
rect 40226 51998 40238 52050
rect 40290 51998 40302 52050
rect 42130 51998 42142 52050
rect 42194 51998 42206 52050
rect 39790 51986 39842 51998
rect 43486 51986 43538 51998
rect 43934 52050 43986 52062
rect 44818 51998 44830 52050
rect 44882 51998 44894 52050
rect 43934 51986 43986 51998
rect 6750 51938 6802 51950
rect 6750 51874 6802 51886
rect 7534 51938 7586 51950
rect 7534 51874 7586 51886
rect 7758 51938 7810 51950
rect 7758 51874 7810 51886
rect 8094 51938 8146 51950
rect 8094 51874 8146 51886
rect 9438 51938 9490 51950
rect 9438 51874 9490 51886
rect 14142 51938 14194 51950
rect 14142 51874 14194 51886
rect 14366 51938 14418 51950
rect 14366 51874 14418 51886
rect 19406 51938 19458 51950
rect 19406 51874 19458 51886
rect 20302 51938 20354 51950
rect 21646 51938 21698 51950
rect 21298 51886 21310 51938
rect 21362 51886 21374 51938
rect 20302 51874 20354 51886
rect 21646 51874 21698 51886
rect 22766 51938 22818 51950
rect 22766 51874 22818 51886
rect 22878 51938 22930 51950
rect 22878 51874 22930 51886
rect 35422 51938 35474 51950
rect 42926 51938 42978 51950
rect 40338 51886 40350 51938
rect 40402 51886 40414 51938
rect 35422 51874 35474 51886
rect 42926 51874 42978 51886
rect 44046 51938 44098 51950
rect 44046 51874 44098 51886
rect 45166 51938 45218 51950
rect 45166 51874 45218 51886
rect 1344 51770 48608 51804
rect 1344 51718 19838 51770
rect 19890 51718 19942 51770
rect 19994 51718 20046 51770
rect 20098 51718 48608 51770
rect 1344 51684 48608 51718
rect 5630 51602 5682 51614
rect 5630 51538 5682 51550
rect 5742 51602 5794 51614
rect 28030 51602 28082 51614
rect 11442 51550 11454 51602
rect 11506 51550 11518 51602
rect 14018 51550 14030 51602
rect 14082 51550 14094 51602
rect 25554 51550 25566 51602
rect 25618 51550 25630 51602
rect 5742 51538 5794 51550
rect 28030 51538 28082 51550
rect 35534 51602 35586 51614
rect 35534 51538 35586 51550
rect 35982 51602 36034 51614
rect 35982 51538 36034 51550
rect 36094 51602 36146 51614
rect 36094 51538 36146 51550
rect 37662 51602 37714 51614
rect 37662 51538 37714 51550
rect 39230 51602 39282 51614
rect 39230 51538 39282 51550
rect 39342 51602 39394 51614
rect 39342 51538 39394 51550
rect 40126 51602 40178 51614
rect 40126 51538 40178 51550
rect 44942 51602 44994 51614
rect 44942 51538 44994 51550
rect 28142 51490 28194 51502
rect 6850 51438 6862 51490
rect 6914 51438 6926 51490
rect 9874 51438 9886 51490
rect 9938 51438 9950 51490
rect 12114 51438 12126 51490
rect 12178 51438 12190 51490
rect 20850 51438 20862 51490
rect 20914 51438 20926 51490
rect 22194 51438 22206 51490
rect 22258 51438 22270 51490
rect 27010 51438 27022 51490
rect 27074 51438 27086 51490
rect 28142 51426 28194 51438
rect 29598 51490 29650 51502
rect 29598 51426 29650 51438
rect 31054 51490 31106 51502
rect 31054 51426 31106 51438
rect 34638 51490 34690 51502
rect 34638 51426 34690 51438
rect 36990 51490 37042 51502
rect 36990 51426 37042 51438
rect 37214 51490 37266 51502
rect 37214 51426 37266 51438
rect 38110 51490 38162 51502
rect 41234 51438 41246 51490
rect 41298 51438 41310 51490
rect 43026 51438 43038 51490
rect 43090 51438 43102 51490
rect 47394 51438 47406 51490
rect 47458 51438 47470 51490
rect 38110 51426 38162 51438
rect 5070 51378 5122 51390
rect 5070 51314 5122 51326
rect 5518 51378 5570 51390
rect 13694 51378 13746 51390
rect 15374 51378 15426 51390
rect 23774 51378 23826 51390
rect 30606 51378 30658 51390
rect 6066 51326 6078 51378
rect 6130 51326 6142 51378
rect 10322 51326 10334 51378
rect 10386 51326 10398 51378
rect 11106 51326 11118 51378
rect 11170 51326 11182 51378
rect 12338 51326 12350 51378
rect 12402 51326 12414 51378
rect 15026 51326 15038 51378
rect 15090 51326 15102 51378
rect 16034 51326 16046 51378
rect 16098 51326 16110 51378
rect 17490 51326 17502 51378
rect 17554 51326 17566 51378
rect 21970 51326 21982 51378
rect 22034 51326 22046 51378
rect 26002 51326 26014 51378
rect 26066 51326 26078 51378
rect 28914 51326 28926 51378
rect 28978 51326 28990 51378
rect 5518 51314 5570 51326
rect 13694 51314 13746 51326
rect 15374 51314 15426 51326
rect 23774 51314 23826 51326
rect 30606 51314 30658 51326
rect 31166 51378 31218 51390
rect 32510 51378 32562 51390
rect 39454 51378 39506 51390
rect 31490 51326 31502 51378
rect 31554 51326 31566 51378
rect 33954 51326 33966 51378
rect 34018 51326 34030 51378
rect 31166 51314 31218 51326
rect 32510 51314 32562 51326
rect 39454 51314 39506 51326
rect 39790 51378 39842 51390
rect 43486 51378 43538 51390
rect 41458 51326 41470 51378
rect 41522 51326 41534 51378
rect 42242 51326 42254 51378
rect 42306 51326 42318 51378
rect 42466 51326 42478 51378
rect 42530 51326 42542 51378
rect 39790 51314 39842 51326
rect 43486 51314 43538 51326
rect 44158 51378 44210 51390
rect 48178 51326 48190 51378
rect 48242 51326 48254 51378
rect 44158 51314 44210 51326
rect 1822 51266 1874 51278
rect 1822 51202 1874 51214
rect 4846 51266 4898 51278
rect 13358 51266 13410 51278
rect 20638 51266 20690 51278
rect 8978 51214 8990 51266
rect 9042 51214 9054 51266
rect 18162 51214 18174 51266
rect 18226 51214 18238 51266
rect 20290 51214 20302 51266
rect 20354 51214 20366 51266
rect 4846 51202 4898 51214
rect 13358 51202 13410 51214
rect 20638 51202 20690 51214
rect 23326 51266 23378 51278
rect 23326 51202 23378 51214
rect 27358 51266 27410 51278
rect 27358 51202 27410 51214
rect 27918 51266 27970 51278
rect 33182 51266 33234 51278
rect 37102 51266 37154 51278
rect 28690 51214 28702 51266
rect 28754 51214 28766 51266
rect 34290 51214 34302 51266
rect 34354 51214 34366 51266
rect 27918 51202 27970 51214
rect 33182 51202 33234 51214
rect 37102 51202 37154 51214
rect 38782 51266 38834 51278
rect 38782 51202 38834 51214
rect 40126 51266 40178 51278
rect 40126 51202 40178 51214
rect 40462 51266 40514 51278
rect 43934 51266 43986 51278
rect 42802 51214 42814 51266
rect 42866 51214 42878 51266
rect 45266 51214 45278 51266
rect 45330 51214 45342 51266
rect 40462 51202 40514 51214
rect 43934 51202 43986 51214
rect 23662 51154 23714 51166
rect 16482 51102 16494 51154
rect 16546 51102 16558 51154
rect 23662 51090 23714 51102
rect 35870 51154 35922 51166
rect 35870 51090 35922 51102
rect 38670 51154 38722 51166
rect 38670 51090 38722 51102
rect 44494 51154 44546 51166
rect 44494 51090 44546 51102
rect 1344 50986 48608 51020
rect 1344 50934 4478 50986
rect 4530 50934 4582 50986
rect 4634 50934 4686 50986
rect 4738 50934 35198 50986
rect 35250 50934 35302 50986
rect 35354 50934 35406 50986
rect 35458 50934 48608 50986
rect 1344 50900 48608 50934
rect 16494 50818 16546 50830
rect 16494 50754 16546 50766
rect 18398 50818 18450 50830
rect 18398 50754 18450 50766
rect 18734 50818 18786 50830
rect 18734 50754 18786 50766
rect 19294 50818 19346 50830
rect 19294 50754 19346 50766
rect 22094 50818 22146 50830
rect 22094 50754 22146 50766
rect 22430 50818 22482 50830
rect 22430 50754 22482 50766
rect 27470 50818 27522 50830
rect 29262 50818 29314 50830
rect 28578 50766 28590 50818
rect 28642 50766 28654 50818
rect 27470 50754 27522 50766
rect 29262 50754 29314 50766
rect 29598 50818 29650 50830
rect 29598 50754 29650 50766
rect 31614 50818 31666 50830
rect 31614 50754 31666 50766
rect 37102 50818 37154 50830
rect 43810 50766 43822 50818
rect 43874 50766 43886 50818
rect 47506 50766 47518 50818
rect 47570 50815 47582 50818
rect 48178 50815 48190 50818
rect 47570 50769 48190 50815
rect 47570 50766 47582 50769
rect 48178 50766 48190 50769
rect 48242 50766 48254 50818
rect 37102 50754 37154 50766
rect 5966 50706 6018 50718
rect 5966 50642 6018 50654
rect 6302 50706 6354 50718
rect 12910 50706 12962 50718
rect 7074 50654 7086 50706
rect 7138 50654 7150 50706
rect 9426 50654 9438 50706
rect 9490 50654 9502 50706
rect 10770 50654 10782 50706
rect 10834 50654 10846 50706
rect 6302 50642 6354 50654
rect 12910 50642 12962 50654
rect 14926 50706 14978 50718
rect 16606 50706 16658 50718
rect 16034 50654 16046 50706
rect 16098 50654 16110 50706
rect 14926 50642 14978 50654
rect 16606 50642 16658 50654
rect 19182 50706 19234 50718
rect 19182 50642 19234 50654
rect 21870 50706 21922 50718
rect 28030 50706 28082 50718
rect 37550 50706 37602 50718
rect 47070 50706 47122 50718
rect 24882 50654 24894 50706
rect 24946 50654 24958 50706
rect 27010 50654 27022 50706
rect 27074 50654 27086 50706
rect 30146 50654 30158 50706
rect 30210 50654 30222 50706
rect 36082 50654 36094 50706
rect 36146 50654 36158 50706
rect 38658 50654 38670 50706
rect 38722 50654 38734 50706
rect 40786 50654 40798 50706
rect 40850 50654 40862 50706
rect 42018 50654 42030 50706
rect 42082 50654 42094 50706
rect 21870 50642 21922 50654
rect 28030 50642 28082 50654
rect 37550 50642 37602 50654
rect 47070 50642 47122 50654
rect 47518 50706 47570 50718
rect 47518 50642 47570 50654
rect 48078 50706 48130 50718
rect 48078 50642 48130 50654
rect 2270 50594 2322 50606
rect 8318 50594 8370 50606
rect 5618 50542 5630 50594
rect 5682 50542 5694 50594
rect 6962 50542 6974 50594
rect 7026 50542 7038 50594
rect 2270 50530 2322 50542
rect 8318 50530 8370 50542
rect 8654 50594 8706 50606
rect 14814 50594 14866 50606
rect 21310 50594 21362 50606
rect 23662 50594 23714 50606
rect 8978 50542 8990 50594
rect 9042 50542 9054 50594
rect 9874 50542 9886 50594
rect 9938 50542 9950 50594
rect 14130 50542 14142 50594
rect 14194 50542 14206 50594
rect 15362 50542 15374 50594
rect 15426 50542 15438 50594
rect 16818 50542 16830 50594
rect 16882 50542 16894 50594
rect 19618 50542 19630 50594
rect 19682 50542 19694 50594
rect 20514 50542 20526 50594
rect 20578 50542 20590 50594
rect 23090 50542 23102 50594
rect 23154 50542 23166 50594
rect 8654 50530 8706 50542
rect 14814 50530 14866 50542
rect 21310 50530 21362 50542
rect 23662 50530 23714 50542
rect 23774 50594 23826 50606
rect 27582 50594 27634 50606
rect 24098 50542 24110 50594
rect 24162 50542 24174 50594
rect 23774 50530 23826 50542
rect 27582 50530 27634 50542
rect 28254 50594 28306 50606
rect 34078 50594 34130 50606
rect 30258 50542 30270 50594
rect 30322 50542 30334 50594
rect 32610 50542 32622 50594
rect 32674 50542 32686 50594
rect 33506 50542 33518 50594
rect 33570 50542 33582 50594
rect 28254 50530 28306 50542
rect 34078 50530 34130 50542
rect 34638 50594 34690 50606
rect 34638 50530 34690 50542
rect 35086 50594 35138 50606
rect 35086 50530 35138 50542
rect 35646 50594 35698 50606
rect 35970 50542 35982 50594
rect 36034 50542 36046 50594
rect 37874 50542 37886 50594
rect 37938 50542 37950 50594
rect 42354 50542 42366 50594
rect 42418 50542 42430 50594
rect 43586 50542 43598 50594
rect 43650 50542 43662 50594
rect 45490 50542 45502 50594
rect 45554 50542 45566 50594
rect 35646 50530 35698 50542
rect 1710 50482 1762 50494
rect 1710 50418 1762 50430
rect 4846 50482 4898 50494
rect 4846 50418 4898 50430
rect 8430 50482 8482 50494
rect 13582 50482 13634 50494
rect 17390 50482 17442 50494
rect 21422 50482 21474 50494
rect 9986 50430 9998 50482
rect 10050 50430 10062 50482
rect 10994 50430 11006 50482
rect 11058 50430 11070 50482
rect 12674 50430 12686 50482
rect 12738 50430 12750 50482
rect 15474 50430 15486 50482
rect 15538 50430 15550 50482
rect 20066 50430 20078 50482
rect 20130 50430 20142 50482
rect 8430 50418 8482 50430
rect 13582 50418 13634 50430
rect 17390 50418 17442 50430
rect 21422 50418 21474 50430
rect 21646 50482 21698 50494
rect 21646 50418 21698 50430
rect 27470 50482 27522 50494
rect 27470 50418 27522 50430
rect 29486 50482 29538 50494
rect 29486 50418 29538 50430
rect 29934 50482 29986 50494
rect 34414 50482 34466 50494
rect 31042 50430 31054 50482
rect 31106 50430 31118 50482
rect 32722 50430 32734 50482
rect 32786 50430 32798 50482
rect 29934 50418 29986 50430
rect 34414 50418 34466 50430
rect 35198 50482 35250 50494
rect 35198 50418 35250 50430
rect 36318 50482 36370 50494
rect 36318 50418 36370 50430
rect 36990 50482 37042 50494
rect 41458 50430 41470 50482
rect 41522 50430 41534 50482
rect 45154 50430 45166 50482
rect 45218 50430 45230 50482
rect 46834 50430 46846 50482
rect 46898 50430 46910 50482
rect 36990 50418 37042 50430
rect 5854 50370 5906 50382
rect 5854 50306 5906 50318
rect 18510 50370 18562 50382
rect 34190 50370 34242 50382
rect 20514 50318 20526 50370
rect 20578 50318 20590 50370
rect 33506 50318 33518 50370
rect 33570 50318 33582 50370
rect 18510 50306 18562 50318
rect 34190 50306 34242 50318
rect 34974 50370 35026 50382
rect 34974 50306 35026 50318
rect 41134 50370 41186 50382
rect 41134 50306 41186 50318
rect 1344 50202 48608 50236
rect 1344 50150 19838 50202
rect 19890 50150 19942 50202
rect 19994 50150 20046 50202
rect 20098 50150 48608 50202
rect 1344 50116 48608 50150
rect 11566 50034 11618 50046
rect 10882 49982 10894 50034
rect 10946 49982 10958 50034
rect 11566 49970 11618 49982
rect 11678 50034 11730 50046
rect 11678 49970 11730 49982
rect 13022 50034 13074 50046
rect 14814 50034 14866 50046
rect 13906 49982 13918 50034
rect 13970 49982 13982 50034
rect 14578 49982 14590 50034
rect 14642 49982 14654 50034
rect 13022 49970 13074 49982
rect 14814 49970 14866 49982
rect 15038 50034 15090 50046
rect 15038 49970 15090 49982
rect 32398 50034 32450 50046
rect 32398 49970 32450 49982
rect 36654 50034 36706 50046
rect 36654 49970 36706 49982
rect 37438 50034 37490 50046
rect 37438 49970 37490 49982
rect 38110 50034 38162 50046
rect 38110 49970 38162 49982
rect 39230 50034 39282 50046
rect 39230 49970 39282 49982
rect 39790 50034 39842 50046
rect 41570 49982 41582 50034
rect 41634 49982 41646 50034
rect 39790 49970 39842 49982
rect 12014 49922 12066 49934
rect 5618 49870 5630 49922
rect 5682 49870 5694 49922
rect 12014 49858 12066 49870
rect 13358 49922 13410 49934
rect 13358 49858 13410 49870
rect 15150 49922 15202 49934
rect 15150 49858 15202 49870
rect 22654 49922 22706 49934
rect 22654 49858 22706 49870
rect 22878 49922 22930 49934
rect 22878 49858 22930 49870
rect 23438 49922 23490 49934
rect 23438 49858 23490 49870
rect 23886 49922 23938 49934
rect 23886 49858 23938 49870
rect 23998 49922 24050 49934
rect 29374 49922 29426 49934
rect 26674 49870 26686 49922
rect 26738 49870 26750 49922
rect 28466 49870 28478 49922
rect 28530 49870 28542 49922
rect 23998 49858 24050 49870
rect 29374 49858 29426 49870
rect 32174 49922 32226 49934
rect 42142 49922 42194 49934
rect 33842 49870 33854 49922
rect 33906 49870 33918 49922
rect 32174 49858 32226 49870
rect 42142 49858 42194 49870
rect 46398 49922 46450 49934
rect 47842 49870 47854 49922
rect 47906 49870 47918 49922
rect 46398 49858 46450 49870
rect 11790 49810 11842 49822
rect 1810 49758 1822 49810
rect 1874 49758 1886 49810
rect 6514 49758 6526 49810
rect 6578 49758 6590 49810
rect 11106 49758 11118 49810
rect 11170 49758 11182 49810
rect 11790 49746 11842 49758
rect 14254 49810 14306 49822
rect 14254 49746 14306 49758
rect 22542 49810 22594 49822
rect 22542 49746 22594 49758
rect 23550 49810 23602 49822
rect 29710 49810 29762 49822
rect 36542 49810 36594 49822
rect 26786 49758 26798 49810
rect 26850 49758 26862 49810
rect 27346 49758 27358 49810
rect 27410 49758 27422 49810
rect 27570 49758 27582 49810
rect 27634 49758 27646 49810
rect 28690 49758 28702 49810
rect 28754 49758 28766 49810
rect 33170 49758 33182 49810
rect 33234 49758 33246 49810
rect 36306 49758 36318 49810
rect 36370 49758 36382 49810
rect 23550 49746 23602 49758
rect 29710 49746 29762 49758
rect 36542 49746 36594 49758
rect 36766 49810 36818 49822
rect 39118 49810 39170 49822
rect 40014 49810 40066 49822
rect 41918 49810 41970 49822
rect 36978 49758 36990 49810
rect 37042 49758 37054 49810
rect 39442 49758 39454 49810
rect 39506 49758 39518 49810
rect 39778 49758 39790 49810
rect 39842 49758 39854 49810
rect 41346 49758 41358 49810
rect 41410 49758 41422 49810
rect 36766 49746 36818 49758
rect 39118 49746 39170 49758
rect 40014 49746 40066 49758
rect 41918 49746 41970 49758
rect 42590 49810 42642 49822
rect 45826 49758 45838 49810
rect 45890 49758 45902 49810
rect 46722 49758 46734 49810
rect 46786 49758 46798 49810
rect 47730 49758 47742 49810
rect 47794 49758 47806 49810
rect 42590 49746 42642 49758
rect 7198 49698 7250 49710
rect 2482 49646 2494 49698
rect 2546 49646 2558 49698
rect 4610 49646 4622 49698
rect 4674 49646 4686 49698
rect 5058 49646 5070 49698
rect 5122 49646 5134 49698
rect 7198 49634 7250 49646
rect 7870 49698 7922 49710
rect 7870 49634 7922 49646
rect 10670 49698 10722 49710
rect 10670 49634 10722 49646
rect 25454 49698 25506 49710
rect 25454 49634 25506 49646
rect 25790 49698 25842 49710
rect 30158 49698 30210 49710
rect 38222 49698 38274 49710
rect 26562 49646 26574 49698
rect 26626 49646 26638 49698
rect 28242 49646 28254 49698
rect 28306 49646 28318 49698
rect 32498 49646 32510 49698
rect 32562 49646 32574 49698
rect 35970 49646 35982 49698
rect 36034 49646 36046 49698
rect 25790 49634 25842 49646
rect 30158 49634 30210 49646
rect 38222 49634 38274 49646
rect 38670 49698 38722 49710
rect 38670 49634 38722 49646
rect 40350 49698 40402 49710
rect 40350 49634 40402 49646
rect 42030 49698 42082 49710
rect 46286 49698 46338 49710
rect 42914 49646 42926 49698
rect 42978 49646 42990 49698
rect 45042 49646 45054 49698
rect 45106 49646 45118 49698
rect 47394 49646 47406 49698
rect 47458 49646 47470 49698
rect 42030 49634 42082 49646
rect 46286 49634 46338 49646
rect 13582 49586 13634 49598
rect 13582 49522 13634 49534
rect 23438 49586 23490 49598
rect 23438 49522 23490 49534
rect 23998 49586 24050 49598
rect 23998 49522 24050 49534
rect 25902 49586 25954 49598
rect 25902 49522 25954 49534
rect 1344 49418 48608 49452
rect 1344 49366 4478 49418
rect 4530 49366 4582 49418
rect 4634 49366 4686 49418
rect 4738 49366 35198 49418
rect 35250 49366 35302 49418
rect 35354 49366 35406 49418
rect 35458 49366 48608 49418
rect 1344 49332 48608 49366
rect 7310 49250 7362 49262
rect 26462 49250 26514 49262
rect 6402 49198 6414 49250
rect 6466 49198 6478 49250
rect 8754 49198 8766 49250
rect 8818 49198 8830 49250
rect 7310 49186 7362 49198
rect 26462 49186 26514 49198
rect 29598 49250 29650 49262
rect 29598 49186 29650 49198
rect 35982 49250 36034 49262
rect 35982 49186 36034 49198
rect 45054 49250 45106 49262
rect 45378 49198 45390 49250
rect 45442 49198 45454 49250
rect 45054 49186 45106 49198
rect 7422 49138 7474 49150
rect 6178 49086 6190 49138
rect 6242 49086 6254 49138
rect 7422 49074 7474 49086
rect 18510 49138 18562 49150
rect 25342 49138 25394 49150
rect 34638 49138 34690 49150
rect 19618 49086 19630 49138
rect 19682 49086 19694 49138
rect 30034 49086 30046 49138
rect 30098 49086 30110 49138
rect 32834 49086 32846 49138
rect 32898 49086 32910 49138
rect 33730 49086 33742 49138
rect 33794 49086 33806 49138
rect 18510 49074 18562 49086
rect 25342 49074 25394 49086
rect 34638 49074 34690 49086
rect 37102 49138 37154 49150
rect 37102 49074 37154 49086
rect 39006 49138 39058 49150
rect 39006 49074 39058 49086
rect 39454 49138 39506 49150
rect 39454 49074 39506 49086
rect 40126 49138 40178 49150
rect 42130 49086 42142 49138
rect 42194 49086 42206 49138
rect 44258 49086 44270 49138
rect 44322 49086 44334 49138
rect 40126 49074 40178 49086
rect 4734 49026 4786 49038
rect 9102 49026 9154 49038
rect 5506 48974 5518 49026
rect 5570 48974 5582 49026
rect 6290 48974 6302 49026
rect 6354 48974 6366 49026
rect 4734 48962 4786 48974
rect 9102 48962 9154 48974
rect 9326 49026 9378 49038
rect 14030 49026 14082 49038
rect 9762 48974 9774 49026
rect 9826 48974 9838 49026
rect 9326 48962 9378 48974
rect 14030 48962 14082 48974
rect 14366 49026 14418 49038
rect 18734 49026 18786 49038
rect 26350 49026 26402 49038
rect 29262 49026 29314 49038
rect 35198 49026 35250 49038
rect 44830 49026 44882 49038
rect 16370 48974 16382 49026
rect 16434 48974 16446 49026
rect 24546 48974 24558 49026
rect 24610 48974 24622 49026
rect 27346 48974 27358 49026
rect 27410 48974 27422 49026
rect 27906 48974 27918 49026
rect 27970 48974 27982 49026
rect 31490 48974 31502 49026
rect 31554 48974 31566 49026
rect 34178 48974 34190 49026
rect 34242 48974 34254 49026
rect 41346 48974 41358 49026
rect 41410 48974 41422 49026
rect 14366 48962 14418 48974
rect 18734 48962 18786 48974
rect 26350 48962 26402 48974
rect 29262 48962 29314 48974
rect 35198 48962 35250 48974
rect 44830 48962 44882 48974
rect 47630 49026 47682 49038
rect 47630 48962 47682 48974
rect 4958 48914 5010 48926
rect 4958 48850 5010 48862
rect 5070 48914 5122 48926
rect 5070 48850 5122 48862
rect 11566 48914 11618 48926
rect 11566 48850 11618 48862
rect 12238 48914 12290 48926
rect 12238 48850 12290 48862
rect 14142 48914 14194 48926
rect 18062 48914 18114 48926
rect 16034 48862 16046 48914
rect 16098 48862 16110 48914
rect 17490 48862 17502 48914
rect 17554 48862 17566 48914
rect 14142 48850 14194 48862
rect 18062 48850 18114 48862
rect 18286 48914 18338 48926
rect 18286 48850 18338 48862
rect 19966 48914 20018 48926
rect 19966 48850 20018 48862
rect 20302 48914 20354 48926
rect 35422 48914 35474 48926
rect 22530 48862 22542 48914
rect 22594 48862 22606 48914
rect 26002 48862 26014 48914
rect 26066 48862 26078 48914
rect 28578 48862 28590 48914
rect 28642 48862 28654 48914
rect 30258 48862 30270 48914
rect 30322 48862 30334 48914
rect 20302 48850 20354 48862
rect 35422 48850 35474 48862
rect 35534 48914 35586 48926
rect 35534 48850 35586 48862
rect 36094 48914 36146 48926
rect 36094 48850 36146 48862
rect 41022 48914 41074 48926
rect 41022 48850 41074 48862
rect 46734 48914 46786 48926
rect 46734 48850 46786 48862
rect 3726 48802 3778 48814
rect 3726 48738 3778 48750
rect 7534 48802 7586 48814
rect 7534 48738 7586 48750
rect 8430 48802 8482 48814
rect 10446 48802 10498 48814
rect 9986 48750 9998 48802
rect 10050 48750 10062 48802
rect 8430 48738 8482 48750
rect 10446 48738 10498 48750
rect 11678 48802 11730 48814
rect 11678 48738 11730 48750
rect 11902 48802 11954 48814
rect 19742 48802 19794 48814
rect 17378 48750 17390 48802
rect 17442 48750 17454 48802
rect 11902 48738 11954 48750
rect 19742 48738 19794 48750
rect 20414 48802 20466 48814
rect 20414 48738 20466 48750
rect 20638 48802 20690 48814
rect 20638 48738 20690 48750
rect 22878 48802 22930 48814
rect 22878 48738 22930 48750
rect 23438 48802 23490 48814
rect 23438 48738 23490 48750
rect 24110 48802 24162 48814
rect 25678 48802 25730 48814
rect 24322 48750 24334 48802
rect 24386 48750 24398 48802
rect 24110 48738 24162 48750
rect 25678 48738 25730 48750
rect 26462 48802 26514 48814
rect 26462 48738 26514 48750
rect 29486 48802 29538 48814
rect 29486 48738 29538 48750
rect 35982 48802 36034 48814
rect 35982 48738 36034 48750
rect 37774 48802 37826 48814
rect 37774 48738 37826 48750
rect 40574 48802 40626 48814
rect 40574 48738 40626 48750
rect 40910 48802 40962 48814
rect 40910 48738 40962 48750
rect 45838 48802 45890 48814
rect 45838 48738 45890 48750
rect 46510 48802 46562 48814
rect 46510 48738 46562 48750
rect 46622 48802 46674 48814
rect 46622 48738 46674 48750
rect 47406 48802 47458 48814
rect 47406 48738 47458 48750
rect 48190 48802 48242 48814
rect 48190 48738 48242 48750
rect 1344 48634 48608 48668
rect 1344 48582 19838 48634
rect 19890 48582 19942 48634
rect 19994 48582 20046 48634
rect 20098 48582 48608 48634
rect 1344 48548 48608 48582
rect 3054 48466 3106 48478
rect 3054 48402 3106 48414
rect 4398 48466 4450 48478
rect 4398 48402 4450 48414
rect 9438 48466 9490 48478
rect 12014 48466 12066 48478
rect 10658 48414 10670 48466
rect 10722 48414 10734 48466
rect 9438 48402 9490 48414
rect 12014 48402 12066 48414
rect 12574 48466 12626 48478
rect 12574 48402 12626 48414
rect 15822 48466 15874 48478
rect 15822 48402 15874 48414
rect 16718 48466 16770 48478
rect 16718 48402 16770 48414
rect 16830 48466 16882 48478
rect 16830 48402 16882 48414
rect 30382 48466 30434 48478
rect 30382 48402 30434 48414
rect 42478 48466 42530 48478
rect 42478 48402 42530 48414
rect 42590 48466 42642 48478
rect 42590 48402 42642 48414
rect 43374 48466 43426 48478
rect 43374 48402 43426 48414
rect 44046 48466 44098 48478
rect 44046 48402 44098 48414
rect 44494 48466 44546 48478
rect 44494 48402 44546 48414
rect 44942 48466 44994 48478
rect 44942 48402 44994 48414
rect 3390 48354 3442 48366
rect 3390 48290 3442 48302
rect 3950 48354 4002 48366
rect 3950 48290 4002 48302
rect 4846 48354 4898 48366
rect 4846 48290 4898 48302
rect 9662 48354 9714 48366
rect 9662 48290 9714 48302
rect 10110 48354 10162 48366
rect 11790 48354 11842 48366
rect 11666 48302 11678 48354
rect 11730 48302 11742 48354
rect 10110 48290 10162 48302
rect 11790 48290 11842 48302
rect 11902 48354 11954 48366
rect 11902 48290 11954 48302
rect 12910 48354 12962 48366
rect 12910 48290 12962 48302
rect 15710 48354 15762 48366
rect 24222 48354 24274 48366
rect 20850 48302 20862 48354
rect 20914 48302 20926 48354
rect 22194 48302 22206 48354
rect 22258 48302 22270 48354
rect 15710 48290 15762 48302
rect 24222 48290 24274 48302
rect 26238 48354 26290 48366
rect 41022 48354 41074 48366
rect 42366 48354 42418 48366
rect 27906 48302 27918 48354
rect 27970 48302 27982 48354
rect 40002 48302 40014 48354
rect 40066 48302 40078 48354
rect 41682 48302 41694 48354
rect 41746 48302 41758 48354
rect 26238 48290 26290 48302
rect 41022 48290 41074 48302
rect 42366 48290 42418 48302
rect 42926 48354 42978 48366
rect 47394 48302 47406 48354
rect 47458 48302 47470 48354
rect 42926 48290 42978 48302
rect 2158 48242 2210 48254
rect 2158 48178 2210 48190
rect 2382 48242 2434 48254
rect 2382 48178 2434 48190
rect 2718 48242 2770 48254
rect 2718 48178 2770 48190
rect 2942 48242 2994 48254
rect 2942 48178 2994 48190
rect 3166 48242 3218 48254
rect 3166 48178 3218 48190
rect 4174 48242 4226 48254
rect 4174 48178 4226 48190
rect 4958 48242 5010 48254
rect 9774 48242 9826 48254
rect 5842 48190 5854 48242
rect 5906 48190 5918 48242
rect 4958 48178 5010 48190
rect 9774 48178 9826 48190
rect 10334 48242 10386 48254
rect 10334 48178 10386 48190
rect 12126 48242 12178 48254
rect 12126 48178 12178 48190
rect 12462 48242 12514 48254
rect 12462 48178 12514 48190
rect 12686 48242 12738 48254
rect 12686 48178 12738 48190
rect 16158 48242 16210 48254
rect 16158 48178 16210 48190
rect 16606 48242 16658 48254
rect 26910 48242 26962 48254
rect 17490 48190 17502 48242
rect 17554 48190 17566 48242
rect 23762 48190 23774 48242
rect 23826 48190 23838 48242
rect 25554 48190 25566 48242
rect 25618 48190 25630 48242
rect 26562 48190 26574 48242
rect 26626 48190 26638 48242
rect 16606 48178 16658 48190
rect 26910 48178 26962 48190
rect 27134 48242 27186 48254
rect 30494 48242 30546 48254
rect 40350 48242 40402 48254
rect 42702 48242 42754 48254
rect 27346 48190 27358 48242
rect 27410 48239 27422 48242
rect 27570 48239 27582 48242
rect 27410 48193 27582 48239
rect 27410 48190 27422 48193
rect 27570 48190 27582 48193
rect 27634 48190 27646 48242
rect 28018 48190 28030 48242
rect 28082 48190 28094 48242
rect 29922 48190 29934 48242
rect 29986 48190 29998 48242
rect 31266 48190 31278 48242
rect 31330 48190 31342 48242
rect 35522 48190 35534 48242
rect 35586 48190 35598 48242
rect 39218 48190 39230 48242
rect 39282 48190 39294 48242
rect 41458 48190 41470 48242
rect 41522 48190 41534 48242
rect 48066 48190 48078 48242
rect 48130 48190 48142 48242
rect 27134 48178 27186 48190
rect 30494 48178 30546 48190
rect 40350 48178 40402 48190
rect 42702 48178 42754 48190
rect 2494 48130 2546 48142
rect 2494 48066 2546 48078
rect 4286 48130 4338 48142
rect 15374 48130 15426 48142
rect 20638 48130 20690 48142
rect 24670 48130 24722 48142
rect 27022 48130 27074 48142
rect 39678 48130 39730 48142
rect 6514 48078 6526 48130
rect 6578 48078 6590 48130
rect 8642 48078 8654 48130
rect 8706 48078 8718 48130
rect 18162 48078 18174 48130
rect 18226 48078 18238 48130
rect 20290 48078 20302 48130
rect 20354 48078 20366 48130
rect 22754 48078 22766 48130
rect 22818 48078 22830 48130
rect 23314 48078 23326 48130
rect 23378 48078 23390 48130
rect 25330 48078 25342 48130
rect 25394 48078 25406 48130
rect 35858 48078 35870 48130
rect 35922 48078 35934 48130
rect 36306 48078 36318 48130
rect 36370 48078 36382 48130
rect 38434 48078 38446 48130
rect 38498 48078 38510 48130
rect 45266 48078 45278 48130
rect 45330 48078 45342 48130
rect 4286 48066 4338 48078
rect 15374 48066 15426 48078
rect 20638 48066 20690 48078
rect 24670 48066 24722 48078
rect 27022 48066 27074 48078
rect 39678 48066 39730 48078
rect 4846 48018 4898 48030
rect 4846 47954 4898 47966
rect 15822 48018 15874 48030
rect 15822 47954 15874 47966
rect 39566 48018 39618 48030
rect 39566 47954 39618 47966
rect 1344 47850 48608 47884
rect 1344 47798 4478 47850
rect 4530 47798 4582 47850
rect 4634 47798 4686 47850
rect 4738 47798 35198 47850
rect 35250 47798 35302 47850
rect 35354 47798 35406 47850
rect 35458 47798 48608 47850
rect 1344 47764 48608 47798
rect 18286 47682 18338 47694
rect 12786 47630 12798 47682
rect 12850 47630 12862 47682
rect 18286 47618 18338 47630
rect 18622 47682 18674 47694
rect 18622 47618 18674 47630
rect 37550 47682 37602 47694
rect 46722 47630 46734 47682
rect 46786 47630 46798 47682
rect 37550 47618 37602 47630
rect 5070 47570 5122 47582
rect 9438 47570 9490 47582
rect 19630 47570 19682 47582
rect 35086 47570 35138 47582
rect 42142 47570 42194 47582
rect 2482 47518 2494 47570
rect 2546 47518 2558 47570
rect 4610 47518 4622 47570
rect 4674 47518 4686 47570
rect 8530 47518 8542 47570
rect 8594 47518 8606 47570
rect 12114 47518 12126 47570
rect 12178 47518 12190 47570
rect 16482 47518 16494 47570
rect 16546 47518 16558 47570
rect 23986 47518 23998 47570
rect 24050 47518 24062 47570
rect 27458 47518 27470 47570
rect 27522 47518 27534 47570
rect 29698 47518 29710 47570
rect 29762 47518 29774 47570
rect 30706 47518 30718 47570
rect 30770 47518 30782 47570
rect 38882 47518 38894 47570
rect 38946 47518 38958 47570
rect 41010 47518 41022 47570
rect 41074 47518 41086 47570
rect 46834 47518 46846 47570
rect 46898 47518 46910 47570
rect 5070 47506 5122 47518
rect 9438 47506 9490 47518
rect 19630 47506 19682 47518
rect 35086 47506 35138 47518
rect 42142 47506 42194 47518
rect 7086 47458 7138 47470
rect 8878 47458 8930 47470
rect 1810 47406 1822 47458
rect 1874 47406 1886 47458
rect 8306 47406 8318 47458
rect 8370 47406 8382 47458
rect 7086 47394 7138 47406
rect 8878 47394 8930 47406
rect 9326 47458 9378 47470
rect 9326 47394 9378 47406
rect 9550 47458 9602 47470
rect 9550 47394 9602 47406
rect 11230 47458 11282 47470
rect 11230 47394 11282 47406
rect 11566 47458 11618 47470
rect 21646 47458 21698 47470
rect 27694 47458 27746 47470
rect 12450 47406 12462 47458
rect 12514 47406 12526 47458
rect 13682 47406 13694 47458
rect 13746 47406 13758 47458
rect 18274 47406 18286 47458
rect 18338 47406 18350 47458
rect 20066 47406 20078 47458
rect 20130 47406 20142 47458
rect 20514 47406 20526 47458
rect 20578 47406 20590 47458
rect 23538 47406 23550 47458
rect 23602 47406 23614 47458
rect 24546 47406 24558 47458
rect 24610 47406 24622 47458
rect 11566 47394 11618 47406
rect 21646 47394 21698 47406
rect 27694 47394 27746 47406
rect 28030 47458 28082 47470
rect 28030 47394 28082 47406
rect 28366 47458 28418 47470
rect 31278 47458 31330 47470
rect 32174 47458 32226 47470
rect 29810 47406 29822 47458
rect 29874 47406 29886 47458
rect 31490 47406 31502 47458
rect 31554 47406 31566 47458
rect 28366 47394 28418 47406
rect 31278 47394 31330 47406
rect 32174 47394 32226 47406
rect 33406 47458 33458 47470
rect 33406 47394 33458 47406
rect 34974 47458 35026 47470
rect 34974 47394 35026 47406
rect 35422 47458 35474 47470
rect 35422 47394 35474 47406
rect 35646 47458 35698 47470
rect 44830 47458 44882 47470
rect 37538 47406 37550 47458
rect 37602 47406 37614 47458
rect 38210 47406 38222 47458
rect 38274 47406 38286 47458
rect 41570 47406 41582 47458
rect 41634 47406 41646 47458
rect 35646 47394 35698 47406
rect 44830 47394 44882 47406
rect 45054 47458 45106 47470
rect 47406 47458 47458 47470
rect 46610 47406 46622 47458
rect 46674 47406 46686 47458
rect 45054 47394 45106 47406
rect 47406 47394 47458 47406
rect 47966 47458 48018 47470
rect 47966 47394 48018 47406
rect 7310 47346 7362 47358
rect 7310 47282 7362 47294
rect 7646 47346 7698 47358
rect 7646 47282 7698 47294
rect 10222 47346 10274 47358
rect 10222 47282 10274 47294
rect 10558 47346 10610 47358
rect 21310 47346 21362 47358
rect 22766 47346 22818 47358
rect 27918 47346 27970 47358
rect 14354 47294 14366 47346
rect 14418 47294 14430 47346
rect 19394 47294 19406 47346
rect 19458 47294 19470 47346
rect 22082 47294 22094 47346
rect 22146 47294 22158 47346
rect 23426 47294 23438 47346
rect 23490 47294 23502 47346
rect 25330 47294 25342 47346
rect 25394 47294 25406 47346
rect 10558 47282 10610 47294
rect 21310 47282 21362 47294
rect 22766 47282 22818 47294
rect 27918 47282 27970 47294
rect 34526 47346 34578 47358
rect 34526 47282 34578 47294
rect 37214 47346 37266 47358
rect 37214 47282 37266 47294
rect 42478 47346 42530 47358
rect 42478 47282 42530 47294
rect 42702 47346 42754 47358
rect 42702 47282 42754 47294
rect 43038 47346 43090 47358
rect 43038 47282 43090 47294
rect 47630 47346 47682 47358
rect 47630 47282 47682 47294
rect 6862 47234 6914 47246
rect 6862 47170 6914 47182
rect 7198 47234 7250 47246
rect 7198 47170 7250 47182
rect 11342 47234 11394 47246
rect 11342 47170 11394 47182
rect 17054 47234 17106 47246
rect 17054 47170 17106 47182
rect 17390 47234 17442 47246
rect 17390 47170 17442 47182
rect 21422 47234 21474 47246
rect 21422 47170 21474 47182
rect 22430 47234 22482 47246
rect 22430 47170 22482 47182
rect 22878 47234 22930 47246
rect 22878 47170 22930 47182
rect 23102 47234 23154 47246
rect 23102 47170 23154 47182
rect 32734 47234 32786 47246
rect 32734 47170 32786 47182
rect 32846 47234 32898 47246
rect 32846 47170 32898 47182
rect 32958 47234 33010 47246
rect 32958 47170 33010 47182
rect 33742 47234 33794 47246
rect 33742 47170 33794 47182
rect 34414 47234 34466 47246
rect 34414 47170 34466 47182
rect 35198 47234 35250 47246
rect 35198 47170 35250 47182
rect 36206 47234 36258 47246
rect 42926 47234 42978 47246
rect 41346 47182 41358 47234
rect 41410 47182 41422 47234
rect 36206 47170 36258 47182
rect 42926 47170 42978 47182
rect 43486 47234 43538 47246
rect 43486 47170 43538 47182
rect 44270 47234 44322 47246
rect 47742 47234 47794 47246
rect 45378 47182 45390 47234
rect 45442 47182 45454 47234
rect 44270 47170 44322 47182
rect 47742 47170 47794 47182
rect 1344 47066 48608 47100
rect 1344 47014 19838 47066
rect 19890 47014 19942 47066
rect 19994 47014 20046 47066
rect 20098 47014 48608 47066
rect 1344 46980 48608 47014
rect 7758 46898 7810 46910
rect 5058 46846 5070 46898
rect 5122 46846 5134 46898
rect 7758 46834 7810 46846
rect 10446 46898 10498 46910
rect 10446 46834 10498 46846
rect 11678 46898 11730 46910
rect 11678 46834 11730 46846
rect 14926 46898 14978 46910
rect 14926 46834 14978 46846
rect 15934 46898 15986 46910
rect 15934 46834 15986 46846
rect 16718 46898 16770 46910
rect 25342 46898 25394 46910
rect 24658 46846 24670 46898
rect 24722 46846 24734 46898
rect 16718 46834 16770 46846
rect 25342 46834 25394 46846
rect 26462 46898 26514 46910
rect 34750 46898 34802 46910
rect 28690 46846 28702 46898
rect 28754 46846 28766 46898
rect 26462 46834 26514 46846
rect 34750 46834 34802 46846
rect 38782 46898 38834 46910
rect 38782 46834 38834 46846
rect 39678 46898 39730 46910
rect 39678 46834 39730 46846
rect 41022 46898 41074 46910
rect 41022 46834 41074 46846
rect 44718 46898 44770 46910
rect 44718 46834 44770 46846
rect 2830 46786 2882 46798
rect 2830 46722 2882 46734
rect 7310 46786 7362 46798
rect 7310 46722 7362 46734
rect 7534 46786 7586 46798
rect 7534 46722 7586 46734
rect 7870 46786 7922 46798
rect 7870 46722 7922 46734
rect 10222 46786 10274 46798
rect 10222 46722 10274 46734
rect 10782 46786 10834 46798
rect 10782 46722 10834 46734
rect 11006 46786 11058 46798
rect 11006 46722 11058 46734
rect 11342 46786 11394 46798
rect 11342 46722 11394 46734
rect 11454 46786 11506 46798
rect 11454 46722 11506 46734
rect 12238 46786 12290 46798
rect 12238 46722 12290 46734
rect 15822 46786 15874 46798
rect 15822 46722 15874 46734
rect 16046 46786 16098 46798
rect 16046 46722 16098 46734
rect 17726 46786 17778 46798
rect 17726 46722 17778 46734
rect 18398 46786 18450 46798
rect 18398 46722 18450 46734
rect 19182 46786 19234 46798
rect 19182 46722 19234 46734
rect 27806 46786 27858 46798
rect 27806 46722 27858 46734
rect 29934 46786 29986 46798
rect 29934 46722 29986 46734
rect 31950 46786 32002 46798
rect 31950 46722 32002 46734
rect 32510 46786 32562 46798
rect 32510 46722 32562 46734
rect 35310 46786 35362 46798
rect 35310 46722 35362 46734
rect 3726 46674 3778 46686
rect 3266 46622 3278 46674
rect 3330 46622 3342 46674
rect 3726 46610 3778 46622
rect 4510 46674 4562 46686
rect 4510 46610 4562 46622
rect 10110 46674 10162 46686
rect 10110 46610 10162 46622
rect 10670 46674 10722 46686
rect 10670 46610 10722 46622
rect 14702 46674 14754 46686
rect 14702 46610 14754 46622
rect 15150 46674 15202 46686
rect 15150 46610 15202 46622
rect 15374 46674 15426 46686
rect 15374 46610 15426 46622
rect 16494 46674 16546 46686
rect 16494 46610 16546 46622
rect 16830 46674 16882 46686
rect 16830 46610 16882 46622
rect 18510 46674 18562 46686
rect 18510 46610 18562 46622
rect 18958 46674 19010 46686
rect 24334 46674 24386 46686
rect 29150 46674 29202 46686
rect 20402 46622 20414 46674
rect 20466 46622 20478 46674
rect 23090 46622 23102 46674
rect 23154 46622 23166 46674
rect 27346 46622 27358 46674
rect 27410 46622 27422 46674
rect 18958 46610 19010 46622
rect 24334 46610 24386 46622
rect 29150 46610 29202 46622
rect 29374 46674 29426 46686
rect 29374 46610 29426 46622
rect 29486 46674 29538 46686
rect 29486 46610 29538 46622
rect 29710 46674 29762 46686
rect 29710 46610 29762 46622
rect 30270 46674 30322 46686
rect 30270 46610 30322 46622
rect 32286 46674 32338 46686
rect 32286 46610 32338 46622
rect 33294 46674 33346 46686
rect 34190 46674 34242 46686
rect 38894 46674 38946 46686
rect 33730 46622 33742 46674
rect 33794 46622 33806 46674
rect 36306 46622 36318 46674
rect 36370 46622 36382 46674
rect 33294 46610 33346 46622
rect 34190 46610 34242 46622
rect 38894 46610 38946 46622
rect 39230 46674 39282 46686
rect 39230 46610 39282 46622
rect 39342 46674 39394 46686
rect 39342 46610 39394 46622
rect 39902 46674 39954 46686
rect 44258 46622 44270 46674
rect 44322 46622 44334 46674
rect 48066 46622 48078 46674
rect 48130 46622 48142 46674
rect 39902 46610 39954 46622
rect 9774 46562 9826 46574
rect 9774 46498 9826 46510
rect 17838 46562 17890 46574
rect 23886 46562 23938 46574
rect 21074 46510 21086 46562
rect 21138 46510 21150 46562
rect 23202 46510 23214 46562
rect 23266 46510 23278 46562
rect 17838 46498 17890 46510
rect 23886 46498 23938 46510
rect 25790 46562 25842 46574
rect 28142 46562 28194 46574
rect 32062 46562 32114 46574
rect 39566 46562 39618 46574
rect 27010 46510 27022 46562
rect 27074 46510 27086 46562
rect 30370 46510 30382 46562
rect 30434 46510 30446 46562
rect 36978 46510 36990 46562
rect 37042 46510 37054 46562
rect 25790 46498 25842 46510
rect 28142 46498 28194 46510
rect 32062 46498 32114 46510
rect 39566 46498 39618 46510
rect 40350 46562 40402 46574
rect 41346 46510 41358 46562
rect 41410 46510 41422 46562
rect 43474 46510 43486 46562
rect 43538 46510 43550 46562
rect 45266 46510 45278 46562
rect 45330 46510 45342 46562
rect 47394 46510 47406 46562
rect 47458 46510 47470 46562
rect 40350 46498 40402 46510
rect 4734 46450 4786 46462
rect 4734 46386 4786 46398
rect 12350 46450 12402 46462
rect 12350 46386 12402 46398
rect 17950 46450 18002 46462
rect 17950 46386 18002 46398
rect 18622 46450 18674 46462
rect 18622 46386 18674 46398
rect 19294 46450 19346 46462
rect 19294 46386 19346 46398
rect 28366 46450 28418 46462
rect 28366 46386 28418 46398
rect 35086 46450 35138 46462
rect 35086 46386 35138 46398
rect 35422 46450 35474 46462
rect 35422 46386 35474 46398
rect 1344 46282 48608 46316
rect 1344 46230 4478 46282
rect 4530 46230 4582 46282
rect 4634 46230 4686 46282
rect 4738 46230 35198 46282
rect 35250 46230 35302 46282
rect 35354 46230 35406 46282
rect 35458 46230 48608 46282
rect 1344 46196 48608 46230
rect 25342 46114 25394 46126
rect 43150 46114 43202 46126
rect 27346 46062 27358 46114
rect 27410 46062 27422 46114
rect 25342 46050 25394 46062
rect 43150 46050 43202 46062
rect 43486 46114 43538 46126
rect 43486 46050 43538 46062
rect 45950 46114 46002 46126
rect 45950 46050 46002 46062
rect 46286 46114 46338 46126
rect 46286 46050 46338 46062
rect 47070 46114 47122 46126
rect 47070 46050 47122 46062
rect 10334 46002 10386 46014
rect 10334 45938 10386 45950
rect 12798 46002 12850 46014
rect 22542 46002 22594 46014
rect 15026 45950 15038 46002
rect 15090 45950 15102 46002
rect 17378 45950 17390 46002
rect 17442 45950 17454 46002
rect 20066 45950 20078 46002
rect 20130 45950 20142 46002
rect 22082 45950 22094 46002
rect 22146 45950 22158 46002
rect 12798 45938 12850 45950
rect 22542 45938 22594 45950
rect 27918 46002 27970 46014
rect 36430 46002 36482 46014
rect 46958 46002 47010 46014
rect 31602 45950 31614 46002
rect 31666 45950 31678 46002
rect 33730 45950 33742 46002
rect 33794 45950 33806 46002
rect 39890 45950 39902 46002
rect 39954 45950 39966 46002
rect 41906 45950 41918 46002
rect 41970 45950 41982 46002
rect 44818 45950 44830 46002
rect 44882 45950 44894 46002
rect 27918 45938 27970 45950
rect 36430 45938 36482 45950
rect 46958 45938 47010 45950
rect 4398 45890 4450 45902
rect 4398 45826 4450 45838
rect 6526 45890 6578 45902
rect 6526 45826 6578 45838
rect 6974 45890 7026 45902
rect 6974 45826 7026 45838
rect 7646 45890 7698 45902
rect 12350 45890 12402 45902
rect 10770 45838 10782 45890
rect 10834 45838 10846 45890
rect 7646 45826 7698 45838
rect 12350 45826 12402 45838
rect 12686 45890 12738 45902
rect 15598 45890 15650 45902
rect 13570 45838 13582 45890
rect 13634 45838 13646 45890
rect 13906 45838 13918 45890
rect 13970 45838 13982 45890
rect 12686 45826 12738 45838
rect 15598 45826 15650 45838
rect 16046 45890 16098 45902
rect 23214 45890 23266 45902
rect 19282 45838 19294 45890
rect 19346 45838 19358 45890
rect 19618 45838 19630 45890
rect 19682 45838 19694 45890
rect 20178 45838 20190 45890
rect 20242 45838 20254 45890
rect 21858 45838 21870 45890
rect 21922 45838 21934 45890
rect 16046 45826 16098 45838
rect 23214 45826 23266 45838
rect 25006 45890 25058 45902
rect 25006 45826 25058 45838
rect 27694 45890 27746 45902
rect 27694 45826 27746 45838
rect 29598 45890 29650 45902
rect 43262 45890 43314 45902
rect 30930 45838 30942 45890
rect 30994 45838 31006 45890
rect 34850 45838 34862 45890
rect 34914 45838 34926 45890
rect 35858 45838 35870 45890
rect 35922 45838 35934 45890
rect 37090 45838 37102 45890
rect 37154 45838 37166 45890
rect 40338 45838 40350 45890
rect 40402 45838 40414 45890
rect 29598 45826 29650 45838
rect 43262 45826 43314 45838
rect 43598 45890 43650 45902
rect 45838 45890 45890 45902
rect 45266 45838 45278 45890
rect 45330 45838 45342 45890
rect 43598 45826 43650 45838
rect 45838 45826 45890 45838
rect 46174 45890 46226 45902
rect 47630 45890 47682 45902
rect 46722 45838 46734 45890
rect 46786 45838 46798 45890
rect 46174 45826 46226 45838
rect 47630 45826 47682 45838
rect 2270 45778 2322 45790
rect 2270 45714 2322 45726
rect 2606 45778 2658 45790
rect 2606 45714 2658 45726
rect 2830 45778 2882 45790
rect 2830 45714 2882 45726
rect 3614 45778 3666 45790
rect 3614 45714 3666 45726
rect 4062 45778 4114 45790
rect 4062 45714 4114 45726
rect 4734 45778 4786 45790
rect 4734 45714 4786 45726
rect 4846 45778 4898 45790
rect 4846 45714 4898 45726
rect 5966 45778 6018 45790
rect 5966 45714 6018 45726
rect 6302 45778 6354 45790
rect 6302 45714 6354 45726
rect 7982 45778 8034 45790
rect 12910 45778 12962 45790
rect 23998 45778 24050 45790
rect 11218 45726 11230 45778
rect 11282 45726 11294 45778
rect 20290 45726 20302 45778
rect 20354 45726 20366 45778
rect 7982 45714 8034 45726
rect 12910 45714 12962 45726
rect 23998 45714 24050 45726
rect 25454 45778 25506 45790
rect 25454 45714 25506 45726
rect 25678 45778 25730 45790
rect 25678 45714 25730 45726
rect 26014 45778 26066 45790
rect 29922 45726 29934 45778
rect 29986 45726 29998 45778
rect 34514 45726 34526 45778
rect 34578 45726 34590 45778
rect 37762 45726 37774 45778
rect 37826 45726 37838 45778
rect 45154 45726 45166 45778
rect 45218 45726 45230 45778
rect 26014 45714 26066 45726
rect 2494 45666 2546 45678
rect 2494 45602 2546 45614
rect 3278 45666 3330 45678
rect 3278 45602 3330 45614
rect 3502 45666 3554 45678
rect 3502 45602 3554 45614
rect 3726 45666 3778 45678
rect 3726 45602 3778 45614
rect 4174 45666 4226 45678
rect 4174 45602 4226 45614
rect 4510 45666 4562 45678
rect 4510 45602 4562 45614
rect 6078 45666 6130 45678
rect 6078 45602 6130 45614
rect 6862 45666 6914 45678
rect 6862 45602 6914 45614
rect 7086 45666 7138 45678
rect 7086 45602 7138 45614
rect 7310 45666 7362 45678
rect 7310 45602 7362 45614
rect 7870 45666 7922 45678
rect 7870 45602 7922 45614
rect 11566 45666 11618 45678
rect 11566 45602 11618 45614
rect 16158 45666 16210 45678
rect 16158 45602 16210 45614
rect 16270 45666 16322 45678
rect 24334 45666 24386 45678
rect 22866 45614 22878 45666
rect 22930 45614 22942 45666
rect 16270 45602 16322 45614
rect 24334 45602 24386 45614
rect 24446 45666 24498 45678
rect 24446 45602 24498 45614
rect 24558 45666 24610 45678
rect 24558 45602 24610 45614
rect 25342 45666 25394 45678
rect 25342 45602 25394 45614
rect 25902 45666 25954 45678
rect 25902 45602 25954 45614
rect 44158 45666 44210 45678
rect 44158 45602 44210 45614
rect 48190 45666 48242 45678
rect 48190 45602 48242 45614
rect 1344 45498 48608 45532
rect 1344 45446 19838 45498
rect 19890 45446 19942 45498
rect 19994 45446 20046 45498
rect 20098 45446 48608 45498
rect 1344 45412 48608 45446
rect 3838 45330 3890 45342
rect 3838 45266 3890 45278
rect 8094 45330 8146 45342
rect 8094 45266 8146 45278
rect 21198 45330 21250 45342
rect 21198 45266 21250 45278
rect 33742 45330 33794 45342
rect 33742 45266 33794 45278
rect 34302 45330 34354 45342
rect 34302 45266 34354 45278
rect 34414 45330 34466 45342
rect 34414 45266 34466 45278
rect 34526 45330 34578 45342
rect 34526 45266 34578 45278
rect 38670 45330 38722 45342
rect 44830 45330 44882 45342
rect 40002 45278 40014 45330
rect 40066 45278 40078 45330
rect 40898 45278 40910 45330
rect 40962 45278 40974 45330
rect 45378 45278 45390 45330
rect 45442 45278 45454 45330
rect 47058 45278 47070 45330
rect 47122 45278 47134 45330
rect 38670 45266 38722 45278
rect 44830 45266 44882 45278
rect 2382 45218 2434 45230
rect 2382 45154 2434 45166
rect 3726 45218 3778 45230
rect 8430 45218 8482 45230
rect 5506 45166 5518 45218
rect 5570 45166 5582 45218
rect 3726 45154 3778 45166
rect 8430 45154 8482 45166
rect 11454 45218 11506 45230
rect 27582 45218 27634 45230
rect 13682 45166 13694 45218
rect 13746 45166 13758 45218
rect 18162 45166 18174 45218
rect 18226 45166 18238 45218
rect 26562 45166 26574 45218
rect 26626 45166 26638 45218
rect 11454 45154 11506 45166
rect 27582 45154 27634 45166
rect 29374 45218 29426 45230
rect 29374 45154 29426 45166
rect 33406 45218 33458 45230
rect 33406 45154 33458 45166
rect 33518 45218 33570 45230
rect 33518 45154 33570 45166
rect 38558 45218 38610 45230
rect 38558 45154 38610 45166
rect 3950 45106 4002 45118
rect 3042 45054 3054 45106
rect 3106 45054 3118 45106
rect 3950 45042 4002 45054
rect 4398 45106 4450 45118
rect 7982 45106 8034 45118
rect 4834 45054 4846 45106
rect 4898 45054 4910 45106
rect 4398 45042 4450 45054
rect 7982 45042 8034 45054
rect 8206 45106 8258 45118
rect 8206 45042 8258 45054
rect 8990 45106 9042 45118
rect 16270 45106 16322 45118
rect 27246 45106 27298 45118
rect 10770 45054 10782 45106
rect 10834 45054 10846 45106
rect 12898 45054 12910 45106
rect 12962 45054 12974 45106
rect 16818 45054 16830 45106
rect 16882 45054 16894 45106
rect 17490 45054 17502 45106
rect 17554 45054 17566 45106
rect 21746 45054 21758 45106
rect 21810 45054 21822 45106
rect 25442 45054 25454 45106
rect 25506 45054 25518 45106
rect 25890 45054 25902 45106
rect 25954 45054 25966 45106
rect 26786 45054 26798 45106
rect 26850 45054 26862 45106
rect 8990 45042 9042 45054
rect 16270 45042 16322 45054
rect 27246 45042 27298 45054
rect 29262 45106 29314 45118
rect 29262 45042 29314 45054
rect 29598 45106 29650 45118
rect 38782 45106 38834 45118
rect 30258 45054 30270 45106
rect 30322 45054 30334 45106
rect 31938 45054 31950 45106
rect 32002 45054 32014 45106
rect 34066 45054 34078 45106
rect 34130 45054 34142 45106
rect 34738 45054 34750 45106
rect 34802 45054 34814 45106
rect 35298 45054 35310 45106
rect 35362 45054 35374 45106
rect 29598 45042 29650 45054
rect 38782 45042 38834 45054
rect 39118 45106 39170 45118
rect 39118 45042 39170 45054
rect 39454 45106 39506 45118
rect 39454 45042 39506 45054
rect 39678 45106 39730 45118
rect 39678 45042 39730 45054
rect 40350 45106 40402 45118
rect 41582 45106 41634 45118
rect 41122 45054 41134 45106
rect 41186 45054 41198 45106
rect 40350 45042 40402 45054
rect 41582 45042 41634 45054
rect 42814 45106 42866 45118
rect 44494 45106 44546 45118
rect 43026 45054 43038 45106
rect 43090 45054 43102 45106
rect 43922 45054 43934 45106
rect 43986 45054 43998 45106
rect 42814 45042 42866 45054
rect 44494 45042 44546 45054
rect 44830 45106 44882 45118
rect 44830 45042 44882 45054
rect 45166 45106 45218 45118
rect 46510 45106 46562 45118
rect 45602 45054 45614 45106
rect 45666 45054 45678 45106
rect 46274 45054 46286 45106
rect 46338 45054 46350 45106
rect 45166 45042 45218 45054
rect 46510 45042 46562 45054
rect 46622 45106 46674 45118
rect 47954 45054 47966 45106
rect 48018 45054 48030 45106
rect 46622 45042 46674 45054
rect 9550 44994 9602 45006
rect 20750 44994 20802 45006
rect 25230 44994 25282 45006
rect 39566 44994 39618 45006
rect 43598 44994 43650 45006
rect 3154 44942 3166 44994
rect 3218 44942 3230 44994
rect 7634 44942 7646 44994
rect 7698 44942 7710 44994
rect 11106 44942 11118 44994
rect 11170 44942 11182 44994
rect 15810 44942 15822 44994
rect 15874 44942 15886 44994
rect 20290 44942 20302 44994
rect 20354 44942 20366 44994
rect 22530 44942 22542 44994
rect 22594 44942 22606 44994
rect 24658 44942 24670 44994
rect 24722 44942 24734 44994
rect 29810 44942 29822 44994
rect 29874 44942 29886 44994
rect 35970 44942 35982 44994
rect 36034 44942 36046 44994
rect 38098 44942 38110 44994
rect 38162 44942 38174 44994
rect 42018 44942 42030 44994
rect 42082 44942 42094 44994
rect 9550 44930 9602 44942
rect 20750 44930 20802 44942
rect 25230 44930 25282 44942
rect 39566 44930 39618 44942
rect 43598 44930 43650 44942
rect 47518 44994 47570 45006
rect 47518 44930 47570 44942
rect 9774 44882 9826 44894
rect 9774 44818 9826 44830
rect 10110 44882 10162 44894
rect 10110 44818 10162 44830
rect 16494 44882 16546 44894
rect 42702 44882 42754 44894
rect 47406 44882 47458 44894
rect 29922 44830 29934 44882
rect 29986 44830 29998 44882
rect 43474 44830 43486 44882
rect 43538 44830 43550 44882
rect 16494 44818 16546 44830
rect 42702 44818 42754 44830
rect 47406 44818 47458 44830
rect 47742 44882 47794 44894
rect 47742 44818 47794 44830
rect 1344 44714 48608 44748
rect 1344 44662 4478 44714
rect 4530 44662 4582 44714
rect 4634 44662 4686 44714
rect 4738 44662 35198 44714
rect 35250 44662 35302 44714
rect 35354 44662 35406 44714
rect 35458 44662 48608 44714
rect 1344 44628 48608 44662
rect 7758 44546 7810 44558
rect 26238 44546 26290 44558
rect 11330 44494 11342 44546
rect 11394 44494 11406 44546
rect 19842 44494 19854 44546
rect 19906 44543 19918 44546
rect 20738 44543 20750 44546
rect 19906 44497 20750 44543
rect 19906 44494 19918 44497
rect 20738 44494 20750 44497
rect 20802 44494 20814 44546
rect 24882 44494 24894 44546
rect 24946 44494 24958 44546
rect 7758 44482 7810 44494
rect 26238 44482 26290 44494
rect 34638 44546 34690 44558
rect 34638 44482 34690 44494
rect 35758 44546 35810 44558
rect 35758 44482 35810 44494
rect 38110 44546 38162 44558
rect 42926 44546 42978 44558
rect 41122 44494 41134 44546
rect 41186 44494 41198 44546
rect 38110 44482 38162 44494
rect 42926 44482 42978 44494
rect 6302 44434 6354 44446
rect 14478 44434 14530 44446
rect 2482 44382 2494 44434
rect 2546 44382 2558 44434
rect 4610 44382 4622 44434
rect 4674 44382 4686 44434
rect 6738 44382 6750 44434
rect 6802 44382 6814 44434
rect 6302 44370 6354 44382
rect 14478 44370 14530 44382
rect 14702 44434 14754 44446
rect 19854 44434 19906 44446
rect 15138 44382 15150 44434
rect 15202 44382 15214 44434
rect 14702 44370 14754 44382
rect 19854 44370 19906 44382
rect 20750 44434 20802 44446
rect 20750 44370 20802 44382
rect 23550 44434 23602 44446
rect 26014 44434 26066 44446
rect 31502 44434 31554 44446
rect 24658 44382 24670 44434
rect 24722 44382 24734 44434
rect 29362 44382 29374 44434
rect 29426 44382 29438 44434
rect 23550 44370 23602 44382
rect 26014 44370 26066 44382
rect 31502 44370 31554 44382
rect 32398 44434 32450 44446
rect 32398 44370 32450 44382
rect 34526 44434 34578 44446
rect 34526 44370 34578 44382
rect 35870 44434 35922 44446
rect 35870 44370 35922 44382
rect 37214 44434 37266 44446
rect 37214 44370 37266 44382
rect 38222 44434 38274 44446
rect 38222 44370 38274 44382
rect 38670 44434 38722 44446
rect 38670 44370 38722 44382
rect 43038 44434 43090 44446
rect 43038 44370 43090 44382
rect 44158 44434 44210 44446
rect 45266 44382 45278 44434
rect 45330 44382 45342 44434
rect 47394 44382 47406 44434
rect 47458 44382 47470 44434
rect 44158 44370 44210 44382
rect 10782 44322 10834 44334
rect 1810 44270 1822 44322
rect 1874 44270 1886 44322
rect 6850 44270 6862 44322
rect 6914 44270 6926 44322
rect 10546 44270 10558 44322
rect 10610 44270 10622 44322
rect 10782 44258 10834 44270
rect 12462 44322 12514 44334
rect 23438 44322 23490 44334
rect 15362 44270 15374 44322
rect 15426 44270 15438 44322
rect 18610 44270 18622 44322
rect 18674 44270 18686 44322
rect 12462 44258 12514 44270
rect 23438 44258 23490 44270
rect 23662 44322 23714 44334
rect 23662 44258 23714 44270
rect 23998 44322 24050 44334
rect 27918 44322 27970 44334
rect 30158 44322 30210 44334
rect 24882 44270 24894 44322
rect 24946 44270 24958 44322
rect 25330 44270 25342 44322
rect 25394 44270 25406 44322
rect 27234 44270 27246 44322
rect 27298 44270 27310 44322
rect 27682 44270 27694 44322
rect 27746 44270 27758 44322
rect 29586 44270 29598 44322
rect 29650 44270 29662 44322
rect 23998 44258 24050 44270
rect 27918 44258 27970 44270
rect 30158 44258 30210 44270
rect 30606 44322 30658 44334
rect 33854 44322 33906 44334
rect 41582 44322 41634 44334
rect 30818 44270 30830 44322
rect 30882 44270 30894 44322
rect 36082 44270 36094 44322
rect 36146 44270 36158 44322
rect 40786 44270 40798 44322
rect 40850 44270 40862 44322
rect 41122 44270 41134 44322
rect 41186 44270 41198 44322
rect 30606 44258 30658 44270
rect 33854 44258 33906 44270
rect 41582 44258 41634 44270
rect 41918 44322 41970 44334
rect 44270 44322 44322 44334
rect 42354 44270 42366 44322
rect 42418 44270 42430 44322
rect 48066 44270 48078 44322
rect 48130 44270 48142 44322
rect 41918 44258 41970 44270
rect 44270 44258 44322 44270
rect 7758 44210 7810 44222
rect 10894 44210 10946 44222
rect 7646 44154 7698 44166
rect 5070 44098 5122 44110
rect 5070 44034 5122 44046
rect 5742 44098 5794 44110
rect 8754 44158 8766 44210
rect 8818 44158 8830 44210
rect 7758 44146 7810 44158
rect 10894 44146 10946 44158
rect 12126 44210 12178 44222
rect 34190 44210 34242 44222
rect 43934 44210 43986 44222
rect 16818 44158 16830 44210
rect 16882 44158 16894 44210
rect 42578 44158 42590 44210
rect 42642 44158 42654 44210
rect 43810 44158 43822 44210
rect 43874 44158 43886 44210
rect 12126 44146 12178 44158
rect 34190 44146 34242 44158
rect 43934 44146 43986 44158
rect 44942 44210 44994 44222
rect 44942 44146 44994 44158
rect 7646 44090 7698 44102
rect 9102 44098 9154 44110
rect 9886 44098 9938 44110
rect 5742 44034 5794 44046
rect 9538 44046 9550 44098
rect 9602 44046 9614 44098
rect 9102 44034 9154 44046
rect 9886 44034 9938 44046
rect 12238 44098 12290 44110
rect 12238 44034 12290 44046
rect 19406 44098 19458 44110
rect 19406 44034 19458 44046
rect 20302 44098 20354 44110
rect 20302 44034 20354 44046
rect 22766 44098 22818 44110
rect 31838 44098 31890 44110
rect 26562 44046 26574 44098
rect 26626 44046 26638 44098
rect 22766 44034 22818 44046
rect 31838 44034 31890 44046
rect 34078 44098 34130 44110
rect 34078 44034 34130 44046
rect 40238 44098 40290 44110
rect 40238 44034 40290 44046
rect 41694 44098 41746 44110
rect 41694 44034 41746 44046
rect 44046 44098 44098 44110
rect 44046 44034 44098 44046
rect 1344 43930 48608 43964
rect 1344 43878 19838 43930
rect 19890 43878 19942 43930
rect 19994 43878 20046 43930
rect 20098 43878 48608 43930
rect 1344 43844 48608 43878
rect 10334 43762 10386 43774
rect 10334 43698 10386 43710
rect 12126 43762 12178 43774
rect 12126 43698 12178 43710
rect 25342 43762 25394 43774
rect 36430 43762 36482 43774
rect 28130 43710 28142 43762
rect 28194 43710 28206 43762
rect 25342 43698 25394 43710
rect 36430 43698 36482 43710
rect 38782 43762 38834 43774
rect 38782 43698 38834 43710
rect 41470 43762 41522 43774
rect 41470 43698 41522 43710
rect 47070 43762 47122 43774
rect 47070 43698 47122 43710
rect 5406 43650 5458 43662
rect 3826 43598 3838 43650
rect 3890 43598 3902 43650
rect 5406 43586 5458 43598
rect 8094 43650 8146 43662
rect 8094 43586 8146 43598
rect 11230 43650 11282 43662
rect 11230 43586 11282 43598
rect 11454 43650 11506 43662
rect 11454 43586 11506 43598
rect 15374 43650 15426 43662
rect 15374 43586 15426 43598
rect 15822 43650 15874 43662
rect 15822 43586 15874 43598
rect 16382 43650 16434 43662
rect 16382 43586 16434 43598
rect 16494 43650 16546 43662
rect 16494 43586 16546 43598
rect 20302 43650 20354 43662
rect 25230 43650 25282 43662
rect 21858 43598 21870 43650
rect 21922 43598 21934 43650
rect 20302 43586 20354 43598
rect 25230 43586 25282 43598
rect 26798 43650 26850 43662
rect 29710 43650 29762 43662
rect 27234 43598 27246 43650
rect 27298 43598 27310 43650
rect 26798 43586 26850 43598
rect 29710 43586 29762 43598
rect 31054 43650 31106 43662
rect 31054 43586 31106 43598
rect 36318 43650 36370 43662
rect 36318 43586 36370 43598
rect 37326 43650 37378 43662
rect 37326 43586 37378 43598
rect 37774 43650 37826 43662
rect 37774 43586 37826 43598
rect 40910 43650 40962 43662
rect 40910 43586 40962 43598
rect 41022 43650 41074 43662
rect 41022 43586 41074 43598
rect 43262 43650 43314 43662
rect 47182 43650 47234 43662
rect 44370 43598 44382 43650
rect 44434 43598 44446 43650
rect 43262 43586 43314 43598
rect 47182 43586 47234 43598
rect 48302 43650 48354 43662
rect 48302 43586 48354 43598
rect 5182 43538 5234 43550
rect 4274 43486 4286 43538
rect 4338 43486 4350 43538
rect 4946 43486 4958 43538
rect 5010 43486 5022 43538
rect 5182 43474 5234 43486
rect 5518 43538 5570 43550
rect 5518 43474 5570 43486
rect 7870 43538 7922 43550
rect 7870 43474 7922 43486
rect 8206 43538 8258 43550
rect 8206 43474 8258 43486
rect 10222 43538 10274 43550
rect 10222 43474 10274 43486
rect 10446 43538 10498 43550
rect 10446 43474 10498 43486
rect 10894 43538 10946 43550
rect 10894 43474 10946 43486
rect 11118 43538 11170 43550
rect 12014 43538 12066 43550
rect 11666 43486 11678 43538
rect 11730 43486 11742 43538
rect 11118 43474 11170 43486
rect 12014 43474 12066 43486
rect 12238 43538 12290 43550
rect 12238 43474 12290 43486
rect 12574 43538 12626 43550
rect 12574 43474 12626 43486
rect 15710 43538 15762 43550
rect 15710 43474 15762 43486
rect 16270 43538 16322 43550
rect 26686 43538 26738 43550
rect 36542 43538 36594 43550
rect 39006 43538 39058 43550
rect 46734 43538 46786 43550
rect 16818 43486 16830 43538
rect 16882 43486 16894 43538
rect 17938 43486 17950 43538
rect 18002 43486 18014 43538
rect 20738 43486 20750 43538
rect 20802 43486 20814 43538
rect 26338 43486 26350 43538
rect 26402 43486 26414 43538
rect 27682 43486 27694 43538
rect 27746 43486 27758 43538
rect 28018 43486 28030 43538
rect 28082 43486 28094 43538
rect 29138 43486 29150 43538
rect 29202 43486 29214 43538
rect 30370 43486 30382 43538
rect 30434 43486 30446 43538
rect 35858 43486 35870 43538
rect 35922 43486 35934 43538
rect 36866 43486 36878 43538
rect 36930 43486 36942 43538
rect 38546 43486 38558 43538
rect 38610 43486 38622 43538
rect 39218 43486 39230 43538
rect 39282 43486 39294 43538
rect 43586 43486 43598 43538
rect 43650 43486 43662 43538
rect 16270 43474 16322 43486
rect 26686 43474 26738 43486
rect 36542 43474 36594 43486
rect 39006 43474 39058 43486
rect 46734 43474 46786 43486
rect 47294 43538 47346 43550
rect 47294 43474 47346 43486
rect 14926 43426 14978 43438
rect 22318 43426 22370 43438
rect 39790 43426 39842 43438
rect 4386 43374 4398 43426
rect 4450 43374 4462 43426
rect 19618 43374 19630 43426
rect 19682 43374 19694 43426
rect 29362 43374 29374 43426
rect 29426 43374 29438 43426
rect 30706 43374 30718 43426
rect 30770 43374 30782 43426
rect 33058 43374 33070 43426
rect 33122 43374 33134 43426
rect 35186 43374 35198 43426
rect 35250 43374 35262 43426
rect 38770 43374 38782 43426
rect 38834 43374 38846 43426
rect 14926 43362 14978 43374
rect 22318 43362 22370 43374
rect 39790 43362 39842 43374
rect 40126 43426 40178 43438
rect 46498 43374 46510 43426
rect 46562 43374 46574 43426
rect 40126 43362 40178 43374
rect 12798 43314 12850 43326
rect 15822 43314 15874 43326
rect 13122 43262 13134 43314
rect 13186 43262 13198 43314
rect 12798 43250 12850 43262
rect 15822 43250 15874 43262
rect 1344 43146 48608 43180
rect 1344 43094 4478 43146
rect 4530 43094 4582 43146
rect 4634 43094 4686 43146
rect 4738 43094 35198 43146
rect 35250 43094 35302 43146
rect 35354 43094 35406 43146
rect 35458 43094 48608 43146
rect 1344 43060 48608 43094
rect 4734 42978 4786 42990
rect 12238 42978 12290 42990
rect 8306 42926 8318 42978
rect 8370 42926 8382 42978
rect 24546 42926 24558 42978
rect 24610 42975 24622 42978
rect 24770 42975 24782 42978
rect 24610 42929 24782 42975
rect 24610 42926 24622 42929
rect 24770 42926 24782 42929
rect 24834 42926 24846 42978
rect 4734 42914 4786 42926
rect 12238 42914 12290 42926
rect 11118 42866 11170 42878
rect 24558 42866 24610 42878
rect 30046 42866 30098 42878
rect 17154 42814 17166 42866
rect 17218 42814 17230 42866
rect 21746 42814 21758 42866
rect 21810 42814 21822 42866
rect 22642 42814 22654 42866
rect 22706 42814 22718 42866
rect 25890 42814 25902 42866
rect 25954 42814 25966 42866
rect 11118 42802 11170 42814
rect 24558 42802 24610 42814
rect 30046 42802 30098 42814
rect 34190 42866 34242 42878
rect 34190 42802 34242 42814
rect 36318 42866 36370 42878
rect 40014 42866 40066 42878
rect 38098 42814 38110 42866
rect 38162 42814 38174 42866
rect 36318 42802 36370 42814
rect 40014 42802 40066 42814
rect 40238 42866 40290 42878
rect 40238 42802 40290 42814
rect 40686 42866 40738 42878
rect 45054 42866 45106 42878
rect 42018 42814 42030 42866
rect 42082 42814 42094 42866
rect 44146 42814 44158 42866
rect 44210 42814 44222 42866
rect 40686 42802 40738 42814
rect 45054 42802 45106 42814
rect 3390 42754 3442 42766
rect 3390 42690 3442 42702
rect 3838 42754 3890 42766
rect 3838 42690 3890 42702
rect 4846 42754 4898 42766
rect 4846 42690 4898 42702
rect 5742 42754 5794 42766
rect 5742 42690 5794 42702
rect 5966 42754 6018 42766
rect 5966 42690 6018 42702
rect 6302 42754 6354 42766
rect 6302 42690 6354 42702
rect 7198 42754 7250 42766
rect 8990 42754 9042 42766
rect 7746 42702 7758 42754
rect 7810 42702 7822 42754
rect 8082 42702 8094 42754
rect 8146 42702 8158 42754
rect 8642 42702 8654 42754
rect 8706 42702 8718 42754
rect 7198 42690 7250 42702
rect 8990 42690 9042 42702
rect 9326 42754 9378 42766
rect 11790 42754 11842 42766
rect 10434 42702 10446 42754
rect 10498 42702 10510 42754
rect 10882 42702 10894 42754
rect 10946 42702 10958 42754
rect 9326 42690 9378 42702
rect 11790 42690 11842 42702
rect 12014 42754 12066 42766
rect 12014 42690 12066 42702
rect 14702 42754 14754 42766
rect 14702 42690 14754 42702
rect 15038 42754 15090 42766
rect 20862 42754 20914 42766
rect 26238 42754 26290 42766
rect 15586 42702 15598 42754
rect 15650 42702 15662 42754
rect 16258 42702 16270 42754
rect 16322 42702 16334 42754
rect 16482 42702 16494 42754
rect 16546 42702 16558 42754
rect 19954 42702 19966 42754
rect 20018 42702 20030 42754
rect 21970 42702 21982 42754
rect 22034 42702 22046 42754
rect 23090 42702 23102 42754
rect 23154 42702 23166 42754
rect 25666 42702 25678 42754
rect 25730 42702 25742 42754
rect 15038 42690 15090 42702
rect 20862 42690 20914 42702
rect 26238 42690 26290 42702
rect 27134 42754 27186 42766
rect 27134 42690 27186 42702
rect 27358 42754 27410 42766
rect 32062 42754 32114 42766
rect 31378 42702 31390 42754
rect 31442 42702 31454 42754
rect 27358 42690 27410 42702
rect 32062 42690 32114 42702
rect 32958 42754 33010 42766
rect 32958 42690 33010 42702
rect 33070 42754 33122 42766
rect 33070 42690 33122 42702
rect 33294 42754 33346 42766
rect 33294 42690 33346 42702
rect 33630 42754 33682 42766
rect 33630 42690 33682 42702
rect 34078 42754 34130 42766
rect 34078 42690 34130 42702
rect 34638 42754 34690 42766
rect 34638 42690 34690 42702
rect 36990 42754 37042 42766
rect 36990 42690 37042 42702
rect 37662 42754 37714 42766
rect 37662 42690 37714 42702
rect 38222 42754 38274 42766
rect 38222 42690 38274 42702
rect 38446 42754 38498 42766
rect 39230 42754 39282 42766
rect 38994 42702 39006 42754
rect 39058 42702 39070 42754
rect 38446 42690 38498 42702
rect 39230 42690 39282 42702
rect 39342 42754 39394 42766
rect 41234 42702 41246 42754
rect 41298 42702 41310 42754
rect 39342 42690 39394 42702
rect 2830 42642 2882 42654
rect 2830 42578 2882 42590
rect 3166 42642 3218 42654
rect 3166 42578 3218 42590
rect 6638 42642 6690 42654
rect 20526 42642 20578 42654
rect 16594 42590 16606 42642
rect 16658 42590 16670 42642
rect 19282 42590 19294 42642
rect 19346 42590 19358 42642
rect 6638 42578 6690 42590
rect 20526 42578 20578 42590
rect 21422 42642 21474 42654
rect 23774 42642 23826 42654
rect 23426 42590 23438 42642
rect 23490 42590 23502 42642
rect 21422 42578 21474 42590
rect 23774 42578 23826 42590
rect 23998 42642 24050 42654
rect 33406 42642 33458 42654
rect 30482 42590 30494 42642
rect 30546 42590 30558 42642
rect 23998 42578 24050 42590
rect 33406 42578 33458 42590
rect 38670 42642 38722 42654
rect 38670 42578 38722 42590
rect 39678 42642 39730 42654
rect 39678 42578 39730 42590
rect 2606 42530 2658 42542
rect 2606 42466 2658 42478
rect 2942 42530 2994 42542
rect 2942 42466 2994 42478
rect 3726 42530 3778 42542
rect 3726 42466 3778 42478
rect 3950 42530 4002 42542
rect 3950 42466 4002 42478
rect 4174 42530 4226 42542
rect 4174 42466 4226 42478
rect 4734 42530 4786 42542
rect 4734 42466 4786 42478
rect 6078 42530 6130 42542
rect 6078 42466 6130 42478
rect 6526 42530 6578 42542
rect 6526 42466 6578 42478
rect 6750 42530 6802 42542
rect 6750 42466 6802 42478
rect 9214 42530 9266 42542
rect 9214 42466 9266 42478
rect 12686 42530 12738 42542
rect 12686 42466 12738 42478
rect 14814 42530 14866 42542
rect 14814 42466 14866 42478
rect 20638 42530 20690 42542
rect 20638 42466 20690 42478
rect 21646 42530 21698 42542
rect 21646 42466 21698 42478
rect 23886 42530 23938 42542
rect 34302 42530 34354 42542
rect 27682 42478 27694 42530
rect 27746 42478 27758 42530
rect 23886 42466 23938 42478
rect 34302 42466 34354 42478
rect 34750 42530 34802 42542
rect 34750 42466 34802 42478
rect 34974 42530 35026 42542
rect 34974 42466 35026 42478
rect 37102 42530 37154 42542
rect 37102 42466 37154 42478
rect 37214 42530 37266 42542
rect 37214 42466 37266 42478
rect 38110 42530 38162 42542
rect 38110 42466 38162 42478
rect 40014 42530 40066 42542
rect 40014 42466 40066 42478
rect 46734 42530 46786 42542
rect 46734 42466 46786 42478
rect 47182 42530 47234 42542
rect 47182 42466 47234 42478
rect 48302 42530 48354 42542
rect 48302 42466 48354 42478
rect 1344 42362 48608 42396
rect 1344 42310 19838 42362
rect 19890 42310 19942 42362
rect 19994 42310 20046 42362
rect 20098 42310 48608 42362
rect 1344 42276 48608 42310
rect 18510 42194 18562 42206
rect 33182 42194 33234 42206
rect 29474 42142 29486 42194
rect 29538 42142 29550 42194
rect 18510 42130 18562 42142
rect 33182 42130 33234 42142
rect 34526 42194 34578 42206
rect 34526 42130 34578 42142
rect 34974 42194 35026 42206
rect 34974 42130 35026 42142
rect 41022 42194 41074 42206
rect 41022 42130 41074 42142
rect 9550 42082 9602 42094
rect 2482 42030 2494 42082
rect 2546 42030 2558 42082
rect 6066 42030 6078 42082
rect 6130 42030 6142 42082
rect 9550 42018 9602 42030
rect 12238 42082 12290 42094
rect 12238 42018 12290 42030
rect 17838 42082 17890 42094
rect 17838 42018 17890 42030
rect 19070 42082 19122 42094
rect 33294 42082 33346 42094
rect 30146 42030 30158 42082
rect 30210 42030 30222 42082
rect 19070 42018 19122 42030
rect 33294 42018 33346 42030
rect 34302 42082 34354 42094
rect 34302 42018 34354 42030
rect 34862 42082 34914 42094
rect 34862 42018 34914 42030
rect 40014 42082 40066 42094
rect 40014 42018 40066 42030
rect 47070 42082 47122 42094
rect 47070 42018 47122 42030
rect 8654 41970 8706 41982
rect 1810 41918 1822 41970
rect 1874 41918 1886 41970
rect 5394 41918 5406 41970
rect 5458 41918 5470 41970
rect 8654 41906 8706 41918
rect 9662 41970 9714 41982
rect 11902 41970 11954 41982
rect 19182 41970 19234 41982
rect 24670 41970 24722 41982
rect 48078 41970 48130 41982
rect 10434 41918 10446 41970
rect 10498 41918 10510 41970
rect 10994 41918 11006 41970
rect 11058 41918 11070 41970
rect 12562 41918 12574 41970
rect 12626 41918 12638 41970
rect 16370 41918 16382 41970
rect 16434 41918 16446 41970
rect 18274 41918 18286 41970
rect 18338 41918 18350 41970
rect 19730 41918 19742 41970
rect 19794 41918 19806 41970
rect 20514 41918 20526 41970
rect 20578 41918 20590 41970
rect 24210 41918 24222 41970
rect 24274 41918 24286 41970
rect 25330 41918 25342 41970
rect 25394 41918 25406 41970
rect 25554 41918 25566 41970
rect 25618 41918 25630 41970
rect 26226 41918 26238 41970
rect 26290 41918 26302 41970
rect 27346 41918 27358 41970
rect 27410 41918 27422 41970
rect 29250 41918 29262 41970
rect 29314 41918 29326 41970
rect 29810 41918 29822 41970
rect 29874 41918 29886 41970
rect 33954 41918 33966 41970
rect 34018 41918 34030 41970
rect 35186 41918 35198 41970
rect 35250 41918 35262 41970
rect 35522 41918 35534 41970
rect 35586 41918 35598 41970
rect 36306 41918 36318 41970
rect 36370 41918 36382 41970
rect 46498 41918 46510 41970
rect 46562 41918 46574 41970
rect 9662 41906 9714 41918
rect 11902 41906 11954 41918
rect 19182 41906 19234 41918
rect 24670 41906 24722 41918
rect 48078 41906 48130 41918
rect 11566 41858 11618 41870
rect 15822 41858 15874 41870
rect 17726 41858 17778 41870
rect 34414 41858 34466 41870
rect 38894 41858 38946 41870
rect 4610 41806 4622 41858
rect 4674 41806 4686 41858
rect 8194 41806 8206 41858
rect 8258 41806 8270 41858
rect 10322 41806 10334 41858
rect 10386 41806 10398 41858
rect 10882 41806 10894 41858
rect 10946 41806 10958 41858
rect 13346 41806 13358 41858
rect 13410 41806 13422 41858
rect 15474 41806 15486 41858
rect 15538 41806 15550 41858
rect 16706 41806 16718 41858
rect 16770 41806 16782 41858
rect 22642 41806 22654 41858
rect 22706 41806 22718 41858
rect 26450 41806 26462 41858
rect 26514 41806 26526 41858
rect 27458 41806 27470 41858
rect 27522 41806 27534 41858
rect 28578 41806 28590 41858
rect 28642 41806 28654 41858
rect 38434 41806 38446 41858
rect 38498 41806 38510 41858
rect 11566 41794 11618 41806
rect 15822 41794 15874 41806
rect 17726 41794 17778 41806
rect 34414 41794 34466 41806
rect 38894 41794 38946 41806
rect 39342 41858 39394 41870
rect 46386 41806 46398 41858
rect 46450 41806 46462 41858
rect 39342 41794 39394 41806
rect 10110 41746 10162 41758
rect 10110 41682 10162 41694
rect 17614 41746 17666 41758
rect 17614 41682 17666 41694
rect 18622 41746 18674 41758
rect 18622 41682 18674 41694
rect 19070 41746 19122 41758
rect 19070 41682 19122 41694
rect 33070 41746 33122 41758
rect 40126 41746 40178 41758
rect 47182 41746 47234 41758
rect 38882 41694 38894 41746
rect 38946 41743 38958 41746
rect 39554 41743 39566 41746
rect 38946 41697 39566 41743
rect 38946 41694 38958 41697
rect 39554 41694 39566 41697
rect 39618 41694 39630 41746
rect 45714 41694 45726 41746
rect 45778 41694 45790 41746
rect 33070 41682 33122 41694
rect 40126 41682 40178 41694
rect 47182 41682 47234 41694
rect 47406 41746 47458 41758
rect 47406 41682 47458 41694
rect 47518 41746 47570 41758
rect 47518 41682 47570 41694
rect 1344 41578 48608 41612
rect 1344 41526 4478 41578
rect 4530 41526 4582 41578
rect 4634 41526 4686 41578
rect 4738 41526 35198 41578
rect 35250 41526 35302 41578
rect 35354 41526 35406 41578
rect 35458 41526 48608 41578
rect 1344 41492 48608 41526
rect 12798 41410 12850 41422
rect 12798 41346 12850 41358
rect 25678 41410 25730 41422
rect 25678 41346 25730 41358
rect 26014 41410 26066 41422
rect 43486 41410 43538 41422
rect 30146 41358 30158 41410
rect 30210 41358 30222 41410
rect 26014 41346 26066 41358
rect 43486 41346 43538 41358
rect 3054 41298 3106 41310
rect 4958 41298 5010 41310
rect 3378 41246 3390 41298
rect 3442 41246 3454 41298
rect 3054 41234 3106 41246
rect 4958 41234 5010 41246
rect 6974 41298 7026 41310
rect 11566 41298 11618 41310
rect 14478 41298 14530 41310
rect 7298 41246 7310 41298
rect 7362 41246 7374 41298
rect 8530 41246 8542 41298
rect 8594 41246 8606 41298
rect 10770 41246 10782 41298
rect 10834 41246 10846 41298
rect 14018 41246 14030 41298
rect 14082 41246 14094 41298
rect 6974 41234 7026 41246
rect 11566 41234 11618 41246
rect 14478 41234 14530 41246
rect 15150 41298 15202 41310
rect 25454 41298 25506 41310
rect 21410 41246 21422 41298
rect 21474 41246 21486 41298
rect 24546 41246 24558 41298
rect 24610 41246 24622 41298
rect 15150 41234 15202 41246
rect 25454 41234 25506 41246
rect 27806 41298 27858 41310
rect 32510 41298 32562 41310
rect 29698 41246 29710 41298
rect 29762 41246 29774 41298
rect 27806 41234 27858 41246
rect 32510 41234 32562 41246
rect 33182 41298 33234 41310
rect 42814 41298 42866 41310
rect 35298 41246 35310 41298
rect 35362 41246 35374 41298
rect 39330 41246 39342 41298
rect 39394 41246 39406 41298
rect 41458 41246 41470 41298
rect 41522 41246 41534 41298
rect 46050 41246 46062 41298
rect 46114 41246 46126 41298
rect 48178 41246 48190 41298
rect 48242 41246 48254 41298
rect 33182 41234 33234 41246
rect 42814 41234 42866 41246
rect 4510 41186 4562 41198
rect 10222 41186 10274 41198
rect 15038 41186 15090 41198
rect 3490 41134 3502 41186
rect 3554 41134 3566 41186
rect 7634 41134 7646 41186
rect 7698 41134 7710 41186
rect 11218 41134 11230 41186
rect 11282 41134 11294 41186
rect 12114 41134 12126 41186
rect 12178 41134 12190 41186
rect 13794 41134 13806 41186
rect 13858 41134 13870 41186
rect 4510 41122 4562 41134
rect 10222 41122 10274 41134
rect 15038 41122 15090 41134
rect 15598 41186 15650 41198
rect 15598 41122 15650 41134
rect 16046 41186 16098 41198
rect 16046 41122 16098 41134
rect 16606 41186 16658 41198
rect 25118 41186 25170 41198
rect 17602 41134 17614 41186
rect 17666 41134 17678 41186
rect 18386 41134 18398 41186
rect 18450 41134 18462 41186
rect 19842 41134 19854 41186
rect 19906 41134 19918 41186
rect 24658 41134 24670 41186
rect 24722 41134 24734 41186
rect 16606 41122 16658 41134
rect 25118 41122 25170 41134
rect 27470 41186 27522 41198
rect 36990 41186 37042 41198
rect 29026 41134 29038 41186
rect 29090 41134 29102 41186
rect 29810 41134 29822 41186
rect 29874 41134 29886 41186
rect 32834 41134 32846 41186
rect 32898 41134 32910 41186
rect 33506 41134 33518 41186
rect 33570 41134 33582 41186
rect 33842 41134 33854 41186
rect 33906 41134 33918 41186
rect 38098 41134 38110 41186
rect 38162 41134 38174 41186
rect 38770 41134 38782 41186
rect 38834 41134 38846 41186
rect 42242 41134 42254 41186
rect 42306 41134 42318 41186
rect 43138 41134 43150 41186
rect 43202 41134 43214 41186
rect 45378 41134 45390 41186
rect 45442 41134 45454 41186
rect 27470 41122 27522 41134
rect 36990 41122 37042 41134
rect 12910 41074 12962 41086
rect 9874 41022 9886 41074
rect 9938 41022 9950 41074
rect 12910 41010 12962 41022
rect 15374 41074 15426 41086
rect 20526 41074 20578 41086
rect 17378 41022 17390 41074
rect 17442 41022 17454 41074
rect 15374 41010 15426 41022
rect 20526 41010 20578 41022
rect 20638 41074 20690 41086
rect 27246 41074 27298 41086
rect 21634 41022 21646 41074
rect 21698 41022 21710 41074
rect 23314 41022 23326 41074
rect 23378 41022 23390 41074
rect 20638 41010 20690 41022
rect 27246 41010 27298 41022
rect 33070 41074 33122 41086
rect 33070 41010 33122 41022
rect 37102 41074 37154 41086
rect 37102 41010 37154 41022
rect 37662 41074 37714 41086
rect 37662 41010 37714 41022
rect 38446 41074 38498 41086
rect 38446 41010 38498 41022
rect 4398 40962 4450 40974
rect 4398 40898 4450 40910
rect 8990 40962 9042 40974
rect 8990 40898 9042 40910
rect 12350 40962 12402 40974
rect 12350 40898 12402 40910
rect 12798 40962 12850 40974
rect 12798 40898 12850 40910
rect 15934 40962 15986 40974
rect 15934 40898 15986 40910
rect 16158 40962 16210 40974
rect 20862 40962 20914 40974
rect 33294 40962 33346 40974
rect 18722 40910 18734 40962
rect 18786 40910 18798 40962
rect 19618 40910 19630 40962
rect 19682 40910 19694 40962
rect 23426 40910 23438 40962
rect 23490 40910 23502 40962
rect 16158 40898 16210 40910
rect 20862 40898 20914 40910
rect 33294 40898 33346 40910
rect 37774 40962 37826 40974
rect 37774 40898 37826 40910
rect 38334 40962 38386 40974
rect 38334 40898 38386 40910
rect 38558 40962 38610 40974
rect 38558 40898 38610 40910
rect 43374 40962 43426 40974
rect 43374 40898 43426 40910
rect 1344 40794 48608 40828
rect 1344 40742 19838 40794
rect 19890 40742 19942 40794
rect 19994 40742 20046 40794
rect 20098 40742 48608 40794
rect 1344 40708 48608 40742
rect 8318 40626 8370 40638
rect 8318 40562 8370 40574
rect 11118 40626 11170 40638
rect 11118 40562 11170 40574
rect 16382 40626 16434 40638
rect 16382 40562 16434 40574
rect 20862 40626 20914 40638
rect 32174 40626 32226 40638
rect 21634 40574 21646 40626
rect 21698 40574 21710 40626
rect 34178 40574 34190 40626
rect 34242 40574 34254 40626
rect 47506 40574 47518 40626
rect 47570 40574 47582 40626
rect 20862 40562 20914 40574
rect 32174 40562 32226 40574
rect 4510 40514 4562 40526
rect 4510 40450 4562 40462
rect 8878 40514 8930 40526
rect 8878 40450 8930 40462
rect 8990 40514 9042 40526
rect 13358 40514 13410 40526
rect 10770 40462 10782 40514
rect 10834 40462 10846 40514
rect 12226 40462 12238 40514
rect 12290 40462 12302 40514
rect 12674 40462 12686 40514
rect 12738 40462 12750 40514
rect 8990 40450 9042 40462
rect 13358 40450 13410 40462
rect 14030 40514 14082 40526
rect 14030 40450 14082 40462
rect 14142 40514 14194 40526
rect 14142 40450 14194 40462
rect 16270 40514 16322 40526
rect 23886 40514 23938 40526
rect 17602 40462 17614 40514
rect 17666 40462 17678 40514
rect 16270 40450 16322 40462
rect 23886 40450 23938 40462
rect 30270 40514 30322 40526
rect 30270 40450 30322 40462
rect 33182 40514 33234 40526
rect 33182 40450 33234 40462
rect 33294 40514 33346 40526
rect 41918 40514 41970 40526
rect 45950 40514 46002 40526
rect 35746 40462 35758 40514
rect 35810 40462 35822 40514
rect 38210 40462 38222 40514
rect 38274 40462 38286 40514
rect 43362 40462 43374 40514
rect 43426 40462 43438 40514
rect 33294 40450 33346 40462
rect 41918 40450 41970 40462
rect 45950 40450 46002 40462
rect 48190 40514 48242 40526
rect 48190 40450 48242 40462
rect 4286 40402 4338 40414
rect 4286 40338 4338 40350
rect 4622 40402 4674 40414
rect 4622 40338 4674 40350
rect 7870 40402 7922 40414
rect 7870 40338 7922 40350
rect 8206 40402 8258 40414
rect 8206 40338 8258 40350
rect 9886 40402 9938 40414
rect 9886 40338 9938 40350
rect 10446 40402 10498 40414
rect 14366 40402 14418 40414
rect 11554 40350 11566 40402
rect 11618 40350 11630 40402
rect 11778 40350 11790 40402
rect 11842 40350 11854 40402
rect 12562 40350 12574 40402
rect 12626 40350 12638 40402
rect 13570 40350 13582 40402
rect 13634 40350 13646 40402
rect 10446 40338 10498 40350
rect 14366 40338 14418 40350
rect 15934 40402 15986 40414
rect 15934 40338 15986 40350
rect 16830 40402 16882 40414
rect 20414 40402 20466 40414
rect 17714 40350 17726 40402
rect 17778 40350 17790 40402
rect 17938 40350 17950 40402
rect 18002 40350 18014 40402
rect 19058 40350 19070 40402
rect 19122 40350 19134 40402
rect 19506 40350 19518 40402
rect 19570 40350 19582 40402
rect 16830 40338 16882 40350
rect 20414 40338 20466 40350
rect 21086 40402 21138 40414
rect 21086 40338 21138 40350
rect 21310 40402 21362 40414
rect 21310 40338 21362 40350
rect 21982 40402 22034 40414
rect 21982 40338 22034 40350
rect 22430 40402 22482 40414
rect 22430 40338 22482 40350
rect 24446 40402 24498 40414
rect 29822 40402 29874 40414
rect 27122 40350 27134 40402
rect 27186 40350 27198 40402
rect 28914 40350 28926 40402
rect 28978 40350 28990 40402
rect 24446 40338 24498 40350
rect 29822 40338 29874 40350
rect 30046 40402 30098 40414
rect 30046 40338 30098 40350
rect 30382 40402 30434 40414
rect 30382 40338 30434 40350
rect 31838 40402 31890 40414
rect 31838 40338 31890 40350
rect 32062 40402 32114 40414
rect 32062 40338 32114 40350
rect 32286 40402 32338 40414
rect 32286 40338 32338 40350
rect 33518 40402 33570 40414
rect 36542 40402 36594 40414
rect 40910 40402 40962 40414
rect 34514 40350 34526 40402
rect 34578 40350 34590 40402
rect 37426 40350 37438 40402
rect 37490 40350 37502 40402
rect 33518 40338 33570 40350
rect 36542 40338 36594 40350
rect 40910 40338 40962 40350
rect 41470 40402 41522 40414
rect 46958 40402 47010 40414
rect 42690 40350 42702 40402
rect 42754 40350 42766 40402
rect 46722 40350 46734 40402
rect 46786 40350 46798 40402
rect 41470 40338 41522 40350
rect 46958 40338 47010 40350
rect 47070 40402 47122 40414
rect 47070 40338 47122 40350
rect 15374 40290 15426 40302
rect 21198 40290 21250 40302
rect 27918 40290 27970 40302
rect 37102 40290 37154 40302
rect 46174 40290 46226 40302
rect 19730 40238 19742 40290
rect 19794 40238 19806 40290
rect 27458 40238 27470 40290
rect 27522 40238 27534 40290
rect 29026 40238 29038 40290
rect 29090 40238 29102 40290
rect 35970 40238 35982 40290
rect 36034 40238 36046 40290
rect 40338 40238 40350 40290
rect 40402 40238 40414 40290
rect 45490 40238 45502 40290
rect 45554 40238 45566 40290
rect 47842 40238 47854 40290
rect 47906 40238 47918 40290
rect 15374 40226 15426 40238
rect 21198 40226 21250 40238
rect 27918 40226 27970 40238
rect 37102 40226 37154 40238
rect 46174 40226 46226 40238
rect 8318 40178 8370 40190
rect 8318 40114 8370 40126
rect 8878 40178 8930 40190
rect 8878 40114 8930 40126
rect 45838 40178 45890 40190
rect 45838 40114 45890 40126
rect 1344 40010 48608 40044
rect 1344 39958 4478 40010
rect 4530 39958 4582 40010
rect 4634 39958 4686 40010
rect 4738 39958 35198 40010
rect 35250 39958 35302 40010
rect 35354 39958 35406 40010
rect 35458 39958 48608 40010
rect 1344 39924 48608 39958
rect 2830 39842 2882 39854
rect 35646 39842 35698 39854
rect 3938 39790 3950 39842
rect 4002 39790 4014 39842
rect 2830 39778 2882 39790
rect 35646 39778 35698 39790
rect 35982 39842 36034 39854
rect 45614 39842 45666 39854
rect 36194 39790 36206 39842
rect 36258 39839 36270 39842
rect 36530 39839 36542 39842
rect 36258 39793 36542 39839
rect 36258 39790 36270 39793
rect 36530 39790 36542 39793
rect 36594 39790 36606 39842
rect 35982 39778 36034 39790
rect 45614 39778 45666 39790
rect 10894 39730 10946 39742
rect 12910 39730 12962 39742
rect 3154 39678 3166 39730
rect 3218 39678 3230 39730
rect 8530 39678 8542 39730
rect 8594 39678 8606 39730
rect 12114 39678 12126 39730
rect 12178 39678 12190 39730
rect 10894 39666 10946 39678
rect 12910 39666 12962 39678
rect 13918 39730 13970 39742
rect 20078 39730 20130 39742
rect 17938 39678 17950 39730
rect 18002 39678 18014 39730
rect 13918 39666 13970 39678
rect 20078 39666 20130 39678
rect 20750 39730 20802 39742
rect 20750 39666 20802 39678
rect 22206 39730 22258 39742
rect 22206 39666 22258 39678
rect 24110 39730 24162 39742
rect 36990 39730 37042 39742
rect 42478 39730 42530 39742
rect 29250 39678 29262 39730
rect 29314 39678 29326 39730
rect 31714 39678 31726 39730
rect 31778 39678 31790 39730
rect 33170 39678 33182 39730
rect 33234 39678 33246 39730
rect 35298 39678 35310 39730
rect 35362 39678 35374 39730
rect 41122 39678 41134 39730
rect 41186 39678 41198 39730
rect 24110 39666 24162 39678
rect 36990 39666 37042 39678
rect 42478 39666 42530 39678
rect 43374 39730 43426 39742
rect 43374 39666 43426 39678
rect 47182 39730 47234 39742
rect 47182 39666 47234 39678
rect 13470 39618 13522 39630
rect 3602 39566 3614 39618
rect 3666 39566 3678 39618
rect 3826 39566 3838 39618
rect 3890 39566 3902 39618
rect 4498 39566 4510 39618
rect 4562 39566 4574 39618
rect 5730 39566 5742 39618
rect 5794 39566 5806 39618
rect 9538 39566 9550 39618
rect 9602 39566 9614 39618
rect 12226 39566 12238 39618
rect 12290 39566 12302 39618
rect 13470 39554 13522 39566
rect 13806 39618 13858 39630
rect 13806 39554 13858 39566
rect 14030 39618 14082 39630
rect 15374 39618 15426 39630
rect 21982 39618 22034 39630
rect 14802 39566 14814 39618
rect 14866 39566 14878 39618
rect 16034 39566 16046 39618
rect 16098 39566 16110 39618
rect 19506 39566 19518 39618
rect 19570 39566 19582 39618
rect 14030 39554 14082 39566
rect 15374 39554 15426 39566
rect 21982 39554 22034 39566
rect 22318 39618 22370 39630
rect 22318 39554 22370 39566
rect 23774 39618 23826 39630
rect 26014 39618 26066 39630
rect 24658 39566 24670 39618
rect 24722 39566 24734 39618
rect 24994 39566 25006 39618
rect 25058 39566 25070 39618
rect 23774 39554 23826 39566
rect 26014 39554 26066 39566
rect 26126 39618 26178 39630
rect 45838 39618 45890 39630
rect 28018 39566 28030 39618
rect 28082 39566 28094 39618
rect 28578 39566 28590 39618
rect 28642 39566 28654 39618
rect 30706 39566 30718 39618
rect 30770 39566 30782 39618
rect 32386 39566 32398 39618
rect 32450 39566 32462 39618
rect 39106 39566 39118 39618
rect 39170 39566 39182 39618
rect 42018 39566 42030 39618
rect 42082 39566 42094 39618
rect 26126 39554 26178 39566
rect 45838 39554 45890 39566
rect 47070 39618 47122 39630
rect 47070 39554 47122 39566
rect 47406 39618 47458 39630
rect 47406 39554 47458 39566
rect 47630 39618 47682 39630
rect 47630 39554 47682 39566
rect 3054 39506 3106 39518
rect 15486 39506 15538 39518
rect 6402 39454 6414 39506
rect 6466 39454 6478 39506
rect 10434 39454 10446 39506
rect 10498 39454 10510 39506
rect 3054 39442 3106 39454
rect 15486 39442 15538 39454
rect 15822 39506 15874 39518
rect 21422 39506 21474 39518
rect 18386 39454 18398 39506
rect 18450 39454 18462 39506
rect 15822 39442 15874 39454
rect 21422 39442 21474 39454
rect 21758 39506 21810 39518
rect 21758 39442 21810 39454
rect 22654 39506 22706 39518
rect 22654 39442 22706 39454
rect 23550 39506 23602 39518
rect 26462 39506 26514 39518
rect 37550 39506 37602 39518
rect 41694 39506 41746 39518
rect 25554 39454 25566 39506
rect 25618 39454 25630 39506
rect 27906 39454 27918 39506
rect 27970 39454 27982 39506
rect 29698 39454 29710 39506
rect 29762 39454 29774 39506
rect 37986 39454 37998 39506
rect 38050 39454 38062 39506
rect 23550 39442 23602 39454
rect 26462 39442 26514 39454
rect 37550 39442 37602 39454
rect 41694 39442 41746 39454
rect 42366 39506 42418 39518
rect 42366 39442 42418 39454
rect 42702 39506 42754 39518
rect 42702 39442 42754 39454
rect 42926 39506 42978 39518
rect 42926 39442 42978 39454
rect 46398 39506 46450 39518
rect 46398 39442 46450 39454
rect 46734 39506 46786 39518
rect 46734 39442 46786 39454
rect 17166 39394 17218 39406
rect 8978 39342 8990 39394
rect 9042 39342 9054 39394
rect 17166 39330 17218 39342
rect 17614 39394 17666 39406
rect 26350 39394 26402 39406
rect 35870 39394 35922 39406
rect 24546 39342 24558 39394
rect 24610 39342 24622 39394
rect 28466 39342 28478 39394
rect 28530 39342 28542 39394
rect 17614 39330 17666 39342
rect 26350 39330 26402 39342
rect 35870 39330 35922 39342
rect 36430 39394 36482 39406
rect 36430 39330 36482 39342
rect 38334 39394 38386 39406
rect 38334 39330 38386 39342
rect 41806 39394 41858 39406
rect 46062 39394 46114 39406
rect 45266 39342 45278 39394
rect 45330 39342 45342 39394
rect 41806 39330 41858 39342
rect 46062 39330 46114 39342
rect 46286 39394 46338 39406
rect 46286 39330 46338 39342
rect 48190 39394 48242 39406
rect 48190 39330 48242 39342
rect 1344 39226 48608 39260
rect 1344 39174 19838 39226
rect 19890 39174 19942 39226
rect 19994 39174 20046 39226
rect 20098 39174 48608 39226
rect 1344 39140 48608 39174
rect 6302 39058 6354 39070
rect 6302 38994 6354 39006
rect 6414 39058 6466 39070
rect 6414 38994 6466 39006
rect 6974 39058 7026 39070
rect 6974 38994 7026 39006
rect 7422 39058 7474 39070
rect 8318 39058 8370 39070
rect 11790 39058 11842 39070
rect 14030 39058 14082 39070
rect 7970 39006 7982 39058
rect 8034 39006 8046 39058
rect 8642 39006 8654 39058
rect 8706 39006 8718 39058
rect 12562 39006 12574 39058
rect 12626 39006 12638 39058
rect 7422 38994 7474 39006
rect 8318 38994 8370 39006
rect 11790 38994 11842 39006
rect 14030 38994 14082 39006
rect 17950 39058 18002 39070
rect 28926 39058 28978 39070
rect 18274 39006 18286 39058
rect 18338 39006 18350 39058
rect 22642 39006 22654 39058
rect 22706 39006 22718 39058
rect 17950 38994 18002 39006
rect 28926 38994 28978 39006
rect 30382 39058 30434 39070
rect 30382 38994 30434 39006
rect 33070 39058 33122 39070
rect 33070 38994 33122 39006
rect 33182 39058 33234 39070
rect 33182 38994 33234 39006
rect 33294 39058 33346 39070
rect 45378 39006 45390 39058
rect 45442 39006 45454 39058
rect 33294 38994 33346 39006
rect 6526 38946 6578 38958
rect 6526 38882 6578 38894
rect 7646 38946 7698 38958
rect 7646 38882 7698 38894
rect 8990 38946 9042 38958
rect 19070 38946 19122 38958
rect 10882 38894 10894 38946
rect 10946 38894 10958 38946
rect 12898 38894 12910 38946
rect 12962 38894 12974 38946
rect 16594 38894 16606 38946
rect 16658 38894 16670 38946
rect 8990 38882 9042 38894
rect 19070 38882 19122 38894
rect 24670 38946 24722 38958
rect 28814 38946 28866 38958
rect 27346 38894 27358 38946
rect 27410 38894 27422 38946
rect 24670 38882 24722 38894
rect 28814 38882 28866 38894
rect 32286 38946 32338 38958
rect 32286 38882 32338 38894
rect 33966 38946 34018 38958
rect 33966 38882 34018 38894
rect 34078 38946 34130 38958
rect 38446 38946 38498 38958
rect 36866 38894 36878 38946
rect 36930 38894 36942 38946
rect 34078 38882 34130 38894
rect 38446 38882 38498 38894
rect 39678 38946 39730 38958
rect 45502 38946 45554 38958
rect 41794 38894 41806 38946
rect 41858 38894 41870 38946
rect 39678 38882 39730 38894
rect 45502 38882 45554 38894
rect 47518 38946 47570 38958
rect 47518 38882 47570 38894
rect 13694 38834 13746 38846
rect 15374 38834 15426 38846
rect 17390 38834 17442 38846
rect 18846 38834 18898 38846
rect 4610 38782 4622 38834
rect 4674 38782 4686 38834
rect 5282 38782 5294 38834
rect 5346 38782 5358 38834
rect 9426 38782 9438 38834
rect 9490 38782 9502 38834
rect 10210 38782 10222 38834
rect 10274 38782 10286 38834
rect 11778 38782 11790 38834
rect 11842 38782 11854 38834
rect 12786 38782 12798 38834
rect 12850 38782 12862 38834
rect 14802 38782 14814 38834
rect 14866 38782 14878 38834
rect 16370 38782 16382 38834
rect 16434 38782 16446 38834
rect 18498 38782 18510 38834
rect 18562 38782 18574 38834
rect 13694 38770 13746 38782
rect 15374 38770 15426 38782
rect 17390 38770 17442 38782
rect 18846 38770 18898 38782
rect 19182 38834 19234 38846
rect 22990 38834 23042 38846
rect 20402 38782 20414 38834
rect 20466 38782 20478 38834
rect 21746 38782 21758 38834
rect 21810 38782 21822 38834
rect 19182 38770 19234 38782
rect 22990 38770 23042 38782
rect 23214 38834 23266 38846
rect 24558 38834 24610 38846
rect 30942 38834 30994 38846
rect 33742 38834 33794 38846
rect 23986 38782 23998 38834
rect 24050 38782 24062 38834
rect 28130 38782 28142 38834
rect 28194 38782 28206 38834
rect 29138 38782 29150 38834
rect 29202 38782 29214 38834
rect 31714 38782 31726 38834
rect 31778 38782 31790 38834
rect 23214 38770 23266 38782
rect 24558 38770 24610 38782
rect 30942 38770 30994 38782
rect 33742 38770 33794 38782
rect 34302 38834 34354 38846
rect 39006 38834 39058 38846
rect 48078 38834 48130 38846
rect 37538 38782 37550 38834
rect 37602 38782 37614 38834
rect 41122 38782 41134 38834
rect 41186 38782 41198 38834
rect 45938 38782 45950 38834
rect 46002 38782 46014 38834
rect 34302 38770 34354 38782
rect 39006 38770 39058 38782
rect 48078 38770 48130 38782
rect 5070 38722 5122 38734
rect 1698 38670 1710 38722
rect 1762 38670 1774 38722
rect 3826 38670 3838 38722
rect 3890 38670 3902 38722
rect 5070 38658 5122 38670
rect 5742 38722 5794 38734
rect 5742 38658 5794 38670
rect 7534 38722 7586 38734
rect 19630 38722 19682 38734
rect 21310 38722 21362 38734
rect 38110 38722 38162 38734
rect 10098 38670 10110 38722
rect 10162 38670 10174 38722
rect 13906 38670 13918 38722
rect 13970 38670 13982 38722
rect 19730 38670 19742 38722
rect 19794 38670 19806 38722
rect 22082 38670 22094 38722
rect 22146 38670 22158 38722
rect 25218 38670 25230 38722
rect 25282 38670 25294 38722
rect 31490 38670 31502 38722
rect 31554 38670 31566 38722
rect 34738 38670 34750 38722
rect 34802 38670 34814 38722
rect 7534 38658 7586 38670
rect 19630 38658 19682 38670
rect 21310 38658 21362 38670
rect 38110 38658 38162 38670
rect 40350 38722 40402 38734
rect 43922 38670 43934 38722
rect 43986 38670 43998 38722
rect 40350 38658 40402 38670
rect 4958 38610 5010 38622
rect 4958 38546 5010 38558
rect 39566 38610 39618 38622
rect 39566 38546 39618 38558
rect 39902 38610 39954 38622
rect 39902 38546 39954 38558
rect 1344 38442 48608 38476
rect 1344 38390 4478 38442
rect 4530 38390 4582 38442
rect 4634 38390 4686 38442
rect 4738 38390 35198 38442
rect 35250 38390 35302 38442
rect 35354 38390 35406 38442
rect 35458 38390 48608 38442
rect 1344 38356 48608 38390
rect 22430 38274 22482 38286
rect 8082 38222 8094 38274
rect 8146 38222 8158 38274
rect 12674 38222 12686 38274
rect 12738 38222 12750 38274
rect 17826 38222 17838 38274
rect 17890 38222 17902 38274
rect 22430 38210 22482 38222
rect 24558 38274 24610 38286
rect 36094 38274 36146 38286
rect 43822 38274 43874 38286
rect 24882 38222 24894 38274
rect 24946 38222 24958 38274
rect 42018 38222 42030 38274
rect 42082 38222 42094 38274
rect 24558 38210 24610 38222
rect 36094 38210 36146 38222
rect 43822 38210 43874 38222
rect 43934 38274 43986 38286
rect 43934 38210 43986 38222
rect 44158 38274 44210 38286
rect 44158 38210 44210 38222
rect 3950 38162 4002 38174
rect 3950 38098 4002 38110
rect 6414 38162 6466 38174
rect 6414 38098 6466 38110
rect 8654 38162 8706 38174
rect 11230 38162 11282 38174
rect 18398 38162 18450 38174
rect 9986 38110 9998 38162
rect 10050 38110 10062 38162
rect 15250 38110 15262 38162
rect 15314 38110 15326 38162
rect 16482 38110 16494 38162
rect 16546 38110 16558 38162
rect 8654 38098 8706 38110
rect 11230 38098 11282 38110
rect 18398 38098 18450 38110
rect 24334 38162 24386 38174
rect 24334 38098 24386 38110
rect 26014 38162 26066 38174
rect 26014 38098 26066 38110
rect 28366 38162 28418 38174
rect 31390 38162 31442 38174
rect 29250 38110 29262 38162
rect 29314 38110 29326 38162
rect 28366 38098 28418 38110
rect 31390 38098 31442 38110
rect 33070 38162 33122 38174
rect 34850 38110 34862 38162
rect 34914 38110 34926 38162
rect 39442 38110 39454 38162
rect 39506 38110 39518 38162
rect 41570 38110 41582 38162
rect 41634 38110 41646 38162
rect 42354 38110 42366 38162
rect 42418 38110 42430 38162
rect 33070 38098 33122 38110
rect 4510 38050 4562 38062
rect 2594 37998 2606 38050
rect 2658 37998 2670 38050
rect 3490 37998 3502 38050
rect 3554 37998 3566 38050
rect 4510 37986 4562 37998
rect 6190 38050 6242 38062
rect 6190 37986 6242 37998
rect 6526 38050 6578 38062
rect 6526 37986 6578 37998
rect 6862 38050 6914 38062
rect 6862 37986 6914 37998
rect 7310 38050 7362 38062
rect 7310 37986 7362 37998
rect 8430 38050 8482 38062
rect 12686 38050 12738 38062
rect 9090 37998 9102 38050
rect 9154 37998 9166 38050
rect 9874 37998 9886 38050
rect 9938 37998 9950 38050
rect 10770 37998 10782 38050
rect 10834 37998 10846 38050
rect 12002 37998 12014 38050
rect 12066 37998 12078 38050
rect 8430 37986 8482 37998
rect 12686 37986 12738 37998
rect 14254 38050 14306 38062
rect 18174 38050 18226 38062
rect 14354 37998 14366 38050
rect 14418 37998 14430 38050
rect 15138 37998 15150 38050
rect 15202 37998 15214 38050
rect 16146 37998 16158 38050
rect 16210 37998 16222 38050
rect 17154 37998 17166 38050
rect 17218 37998 17230 38050
rect 14254 37986 14306 37998
rect 18174 37986 18226 37998
rect 20078 38050 20130 38062
rect 21646 38050 21698 38062
rect 26126 38050 26178 38062
rect 32174 38050 32226 38062
rect 33630 38050 33682 38062
rect 36206 38050 36258 38062
rect 20514 37998 20526 38050
rect 20578 37998 20590 38050
rect 23090 37998 23102 38050
rect 23154 37998 23166 38050
rect 29138 37998 29150 38050
rect 29202 37998 29214 38050
rect 30146 37998 30158 38050
rect 30210 37998 30222 38050
rect 32386 37998 32398 38050
rect 32450 37998 32462 38050
rect 34738 37998 34750 38050
rect 34802 37998 34814 38050
rect 35522 37998 35534 38050
rect 35586 37998 35598 38050
rect 20078 37986 20130 37998
rect 21646 37986 21698 37998
rect 26126 37986 26178 37998
rect 32174 37986 32226 37998
rect 33630 37986 33682 37998
rect 36206 37986 36258 37998
rect 36990 38050 37042 38062
rect 46846 38050 46898 38062
rect 38770 37998 38782 38050
rect 38834 37998 38846 38050
rect 42802 37998 42814 38050
rect 42866 37998 42878 38050
rect 46050 37998 46062 38050
rect 46114 37998 46126 38050
rect 47618 37998 47630 38050
rect 47682 37998 47694 38050
rect 36990 37986 37042 37998
rect 46846 37986 46898 37998
rect 7422 37938 7474 37950
rect 13694 37938 13746 37950
rect 19182 37938 19234 37950
rect 2034 37886 2046 37938
rect 2098 37886 2110 37938
rect 9650 37886 9662 37938
rect 9714 37886 9726 37938
rect 15810 37886 15822 37938
rect 15874 37886 15886 37938
rect 16258 37886 16270 37938
rect 16322 37886 16334 37938
rect 7422 37874 7474 37886
rect 13694 37874 13746 37886
rect 19182 37874 19234 37886
rect 19294 37938 19346 37950
rect 22094 37938 22146 37950
rect 20738 37886 20750 37938
rect 20802 37886 20814 37938
rect 19294 37874 19346 37886
rect 22094 37874 22146 37886
rect 23326 37938 23378 37950
rect 23326 37874 23378 37886
rect 24110 37938 24162 37950
rect 30606 37938 30658 37950
rect 29250 37886 29262 37938
rect 29314 37886 29326 37938
rect 24110 37874 24162 37886
rect 30606 37874 30658 37886
rect 30942 37938 30994 37950
rect 36094 37938 36146 37950
rect 34290 37886 34302 37938
rect 34354 37886 34366 37938
rect 30942 37874 30994 37886
rect 36094 37874 36146 37886
rect 44270 37938 44322 37950
rect 45378 37886 45390 37938
rect 45442 37886 45454 37938
rect 44270 37874 44322 37886
rect 4174 37826 4226 37838
rect 4174 37762 4226 37774
rect 4398 37826 4450 37838
rect 4398 37762 4450 37774
rect 4958 37826 5010 37838
rect 4958 37762 5010 37774
rect 7198 37826 7250 37838
rect 7198 37762 7250 37774
rect 7646 37826 7698 37838
rect 7646 37762 7698 37774
rect 13918 37826 13970 37838
rect 13918 37762 13970 37774
rect 14142 37826 14194 37838
rect 14142 37762 14194 37774
rect 18846 37826 18898 37838
rect 18846 37762 18898 37774
rect 19518 37826 19570 37838
rect 21422 37826 21474 37838
rect 19730 37774 19742 37826
rect 19794 37774 19806 37826
rect 19518 37762 19570 37774
rect 21422 37762 21474 37774
rect 21534 37826 21586 37838
rect 21534 37762 21586 37774
rect 22318 37826 22370 37838
rect 22318 37762 22370 37774
rect 25678 37826 25730 37838
rect 25678 37762 25730 37774
rect 25902 37826 25954 37838
rect 25902 37762 25954 37774
rect 26574 37826 26626 37838
rect 26574 37762 26626 37774
rect 33406 37826 33458 37838
rect 33406 37762 33458 37774
rect 33518 37826 33570 37838
rect 33518 37762 33570 37774
rect 33854 37826 33906 37838
rect 33854 37762 33906 37774
rect 37550 37826 37602 37838
rect 37550 37762 37602 37774
rect 37886 37826 37938 37838
rect 38210 37774 38222 37826
rect 38274 37774 38286 37826
rect 46050 37774 46062 37826
rect 46114 37774 46126 37826
rect 37886 37762 37938 37774
rect 1344 37658 48608 37692
rect 1344 37606 19838 37658
rect 19890 37606 19942 37658
rect 19994 37606 20046 37658
rect 20098 37606 48608 37658
rect 1344 37572 48608 37606
rect 8766 37490 8818 37502
rect 8766 37426 8818 37438
rect 8878 37490 8930 37502
rect 8878 37426 8930 37438
rect 10222 37490 10274 37502
rect 10222 37426 10274 37438
rect 19854 37490 19906 37502
rect 19854 37426 19906 37438
rect 20190 37490 20242 37502
rect 20190 37426 20242 37438
rect 21198 37490 21250 37502
rect 21198 37426 21250 37438
rect 21646 37490 21698 37502
rect 21646 37426 21698 37438
rect 22990 37490 23042 37502
rect 22990 37426 23042 37438
rect 23550 37490 23602 37502
rect 23550 37426 23602 37438
rect 24782 37490 24834 37502
rect 24782 37426 24834 37438
rect 25454 37490 25506 37502
rect 25454 37426 25506 37438
rect 26014 37490 26066 37502
rect 26014 37426 26066 37438
rect 28030 37490 28082 37502
rect 37886 37490 37938 37502
rect 36082 37438 36094 37490
rect 36146 37438 36158 37490
rect 28030 37426 28082 37438
rect 37886 37426 37938 37438
rect 38222 37490 38274 37502
rect 38222 37426 38274 37438
rect 38558 37490 38610 37502
rect 38558 37426 38610 37438
rect 39230 37490 39282 37502
rect 39230 37426 39282 37438
rect 41918 37490 41970 37502
rect 41918 37426 41970 37438
rect 2830 37378 2882 37390
rect 2830 37314 2882 37326
rect 2942 37378 2994 37390
rect 10334 37378 10386 37390
rect 3378 37326 3390 37378
rect 3442 37326 3454 37378
rect 5842 37326 5854 37378
rect 5906 37326 5918 37378
rect 2942 37314 2994 37326
rect 10334 37314 10386 37326
rect 10782 37378 10834 37390
rect 10782 37314 10834 37326
rect 11902 37378 11954 37390
rect 11902 37314 11954 37326
rect 12574 37378 12626 37390
rect 12574 37314 12626 37326
rect 14478 37378 14530 37390
rect 14478 37314 14530 37326
rect 15150 37378 15202 37390
rect 15150 37314 15202 37326
rect 20862 37378 20914 37390
rect 20862 37314 20914 37326
rect 21086 37378 21138 37390
rect 21086 37314 21138 37326
rect 25342 37378 25394 37390
rect 25342 37314 25394 37326
rect 27806 37378 27858 37390
rect 33630 37378 33682 37390
rect 41470 37378 41522 37390
rect 28802 37326 28814 37378
rect 28866 37326 28878 37378
rect 34626 37326 34638 37378
rect 34690 37326 34702 37378
rect 27806 37314 27858 37326
rect 33630 37314 33682 37326
rect 41470 37314 41522 37326
rect 42366 37378 42418 37390
rect 42366 37314 42418 37326
rect 43598 37378 43650 37390
rect 44594 37326 44606 37378
rect 44658 37326 44670 37378
rect 47170 37326 47182 37378
rect 47234 37326 47246 37378
rect 43598 37314 43650 37326
rect 8206 37266 8258 37278
rect 3714 37214 3726 37266
rect 3778 37214 3790 37266
rect 4386 37214 4398 37266
rect 4450 37214 4462 37266
rect 5170 37214 5182 37266
rect 5234 37214 5246 37266
rect 8206 37202 8258 37214
rect 8654 37266 8706 37278
rect 8654 37202 8706 37214
rect 9662 37266 9714 37278
rect 11566 37266 11618 37278
rect 16270 37266 16322 37278
rect 18286 37266 18338 37278
rect 10994 37214 11006 37266
rect 11058 37214 11070 37266
rect 12338 37214 12350 37266
rect 12402 37214 12414 37266
rect 14690 37214 14702 37266
rect 14754 37214 14766 37266
rect 15362 37214 15374 37266
rect 15426 37214 15438 37266
rect 17938 37214 17950 37266
rect 18002 37214 18014 37266
rect 9662 37202 9714 37214
rect 11566 37202 11618 37214
rect 16270 37202 16322 37214
rect 18286 37202 18338 37214
rect 18398 37266 18450 37278
rect 18398 37202 18450 37214
rect 18734 37266 18786 37278
rect 18734 37202 18786 37214
rect 19182 37266 19234 37278
rect 19182 37202 19234 37214
rect 19294 37266 19346 37278
rect 19294 37202 19346 37214
rect 19742 37266 19794 37278
rect 19742 37202 19794 37214
rect 19966 37266 20018 37278
rect 19966 37202 20018 37214
rect 20526 37266 20578 37278
rect 20526 37202 20578 37214
rect 21870 37266 21922 37278
rect 21870 37202 21922 37214
rect 22318 37266 22370 37278
rect 22318 37202 22370 37214
rect 23438 37266 23490 37278
rect 23438 37202 23490 37214
rect 23662 37266 23714 37278
rect 25230 37266 25282 37278
rect 23986 37214 23998 37266
rect 24050 37214 24062 37266
rect 23662 37202 23714 37214
rect 25230 37202 25282 37214
rect 26462 37266 26514 37278
rect 26462 37202 26514 37214
rect 27694 37266 27746 37278
rect 32510 37266 32562 37278
rect 29362 37214 29374 37266
rect 29426 37214 29438 37266
rect 30034 37214 30046 37266
rect 30098 37214 30110 37266
rect 27694 37202 27746 37214
rect 32510 37202 32562 37214
rect 32958 37266 33010 37278
rect 32958 37202 33010 37214
rect 33294 37266 33346 37278
rect 38894 37266 38946 37278
rect 34738 37214 34750 37266
rect 34802 37214 34814 37266
rect 35634 37214 35646 37266
rect 35698 37214 35710 37266
rect 33294 37202 33346 37214
rect 38894 37202 38946 37214
rect 39790 37266 39842 37278
rect 39790 37202 39842 37214
rect 41582 37266 41634 37278
rect 42702 37266 42754 37278
rect 42130 37214 42142 37266
rect 42194 37214 42206 37266
rect 43810 37214 43822 37266
rect 43874 37214 43886 37266
rect 47058 37214 47070 37266
rect 47122 37214 47134 37266
rect 47954 37214 47966 37266
rect 48018 37214 48030 37266
rect 41582 37202 41634 37214
rect 42702 37202 42754 37214
rect 16046 37154 16098 37166
rect 18958 37154 19010 37166
rect 3490 37102 3502 37154
rect 3554 37102 3566 37154
rect 7970 37102 7982 37154
rect 8034 37102 8046 37154
rect 16706 37102 16718 37154
rect 16770 37102 16782 37154
rect 16046 37090 16098 37102
rect 18958 37090 19010 37102
rect 21758 37154 21810 37166
rect 21758 37090 21810 37102
rect 27470 37154 27522 37166
rect 27470 37090 27522 37102
rect 30718 37154 30770 37166
rect 30718 37090 30770 37102
rect 33182 37154 33234 37166
rect 33182 37090 33234 37102
rect 40238 37154 40290 37166
rect 40238 37090 40290 37102
rect 42926 37154 42978 37166
rect 46722 37102 46734 37154
rect 46786 37102 46798 37154
rect 47170 37102 47182 37154
rect 47234 37102 47246 37154
rect 42926 37090 42978 37102
rect 2830 37042 2882 37054
rect 2830 36978 2882 36990
rect 10110 37042 10162 37054
rect 10110 36978 10162 36990
rect 22654 37042 22706 37054
rect 22654 36978 22706 36990
rect 22878 37042 22930 37054
rect 22878 36978 22930 36990
rect 22990 37042 23042 37054
rect 41470 37042 41522 37054
rect 25778 36990 25790 37042
rect 25842 37039 25854 37042
rect 26562 37039 26574 37042
rect 25842 36993 26574 37039
rect 25842 36990 25854 36993
rect 26562 36990 26574 36993
rect 26626 36990 26638 37042
rect 22990 36978 23042 36990
rect 41470 36978 41522 36990
rect 42254 37042 42306 37054
rect 42254 36978 42306 36990
rect 43150 37042 43202 37054
rect 43150 36978 43202 36990
rect 1344 36874 48608 36908
rect 1344 36822 4478 36874
rect 4530 36822 4582 36874
rect 4634 36822 4686 36874
rect 4738 36822 35198 36874
rect 35250 36822 35302 36874
rect 35354 36822 35406 36874
rect 35458 36822 48608 36874
rect 1344 36788 48608 36822
rect 4958 36706 5010 36718
rect 4958 36642 5010 36654
rect 20302 36706 20354 36718
rect 20302 36642 20354 36654
rect 24670 36706 24722 36718
rect 26798 36706 26850 36718
rect 34526 36706 34578 36718
rect 25666 36654 25678 36706
rect 25730 36654 25742 36706
rect 30146 36654 30158 36706
rect 30210 36654 30222 36706
rect 24670 36642 24722 36654
rect 26798 36642 26850 36654
rect 34526 36642 34578 36654
rect 34862 36706 34914 36718
rect 34862 36642 34914 36654
rect 36094 36706 36146 36718
rect 36094 36642 36146 36654
rect 5070 36594 5122 36606
rect 4610 36542 4622 36594
rect 4674 36542 4686 36594
rect 5070 36530 5122 36542
rect 5742 36594 5794 36606
rect 5742 36530 5794 36542
rect 6190 36594 6242 36606
rect 18398 36594 18450 36606
rect 7074 36542 7086 36594
rect 7138 36542 7150 36594
rect 10994 36542 11006 36594
rect 11058 36542 11070 36594
rect 12450 36542 12462 36594
rect 12514 36542 12526 36594
rect 6190 36530 6242 36542
rect 18398 36530 18450 36542
rect 18846 36594 18898 36606
rect 18846 36530 18898 36542
rect 21982 36594 22034 36606
rect 24222 36594 24274 36606
rect 28366 36594 28418 36606
rect 38558 36594 38610 36606
rect 47742 36594 47794 36606
rect 23314 36542 23326 36594
rect 23378 36542 23390 36594
rect 25554 36542 25566 36594
rect 25618 36542 25630 36594
rect 27570 36542 27582 36594
rect 27634 36542 27646 36594
rect 29474 36542 29486 36594
rect 29538 36542 29550 36594
rect 34178 36542 34190 36594
rect 34242 36542 34254 36594
rect 41794 36542 41806 36594
rect 41858 36542 41870 36594
rect 21982 36530 22034 36542
rect 24222 36530 24274 36542
rect 28366 36530 28418 36542
rect 38558 36530 38610 36542
rect 47742 36530 47794 36542
rect 10670 36482 10722 36494
rect 18286 36482 18338 36494
rect 1810 36430 1822 36482
rect 1874 36430 1886 36482
rect 6626 36430 6638 36482
rect 6690 36430 6702 36482
rect 8530 36430 8542 36482
rect 8594 36430 8606 36482
rect 13570 36430 13582 36482
rect 13634 36430 13646 36482
rect 15250 36430 15262 36482
rect 15314 36430 15326 36482
rect 17266 36430 17278 36482
rect 17330 36430 17342 36482
rect 10670 36418 10722 36430
rect 18286 36418 18338 36430
rect 18510 36482 18562 36494
rect 18510 36418 18562 36430
rect 19406 36482 19458 36494
rect 19406 36418 19458 36430
rect 20078 36482 20130 36494
rect 27022 36482 27074 36494
rect 35198 36482 35250 36494
rect 21410 36430 21422 36482
rect 21474 36430 21486 36482
rect 22306 36430 22318 36482
rect 22370 36430 22382 36482
rect 22866 36430 22878 36482
rect 22930 36430 22942 36482
rect 23538 36430 23550 36482
rect 23602 36430 23614 36482
rect 27794 36430 27806 36482
rect 27858 36430 27870 36482
rect 29586 36430 29598 36482
rect 29650 36430 29662 36482
rect 31266 36430 31278 36482
rect 31330 36430 31342 36482
rect 32050 36430 32062 36482
rect 32114 36430 32126 36482
rect 20078 36418 20130 36430
rect 27022 36418 27074 36430
rect 35198 36418 35250 36430
rect 35534 36482 35586 36494
rect 42254 36482 42306 36494
rect 47294 36482 47346 36494
rect 38882 36430 38894 36482
rect 38946 36430 38958 36482
rect 42802 36430 42814 36482
rect 42866 36430 42878 36482
rect 35534 36418 35586 36430
rect 42254 36418 42306 36430
rect 47294 36418 47346 36430
rect 47630 36482 47682 36494
rect 47630 36418 47682 36430
rect 47854 36482 47906 36494
rect 47854 36418 47906 36430
rect 18062 36370 18114 36382
rect 24670 36370 24722 36382
rect 2482 36318 2494 36370
rect 2546 36318 2558 36370
rect 10434 36318 10446 36370
rect 10498 36318 10510 36370
rect 11666 36318 11678 36370
rect 11730 36318 11742 36370
rect 13458 36318 13470 36370
rect 13522 36318 13534 36370
rect 17602 36318 17614 36370
rect 17666 36318 17678 36370
rect 21522 36318 21534 36370
rect 21586 36318 21598 36370
rect 18062 36306 18114 36318
rect 24670 36306 24722 36318
rect 24782 36370 24834 36382
rect 34750 36370 34802 36382
rect 25218 36318 25230 36370
rect 25282 36318 25294 36370
rect 24782 36306 24834 36318
rect 34750 36306 34802 36318
rect 35310 36370 35362 36382
rect 35310 36306 35362 36318
rect 36318 36370 36370 36382
rect 42142 36370 42194 36382
rect 39666 36318 39678 36370
rect 39730 36318 39742 36370
rect 46610 36318 46622 36370
rect 46674 36318 46686 36370
rect 36318 36306 36370 36318
rect 42142 36306 42194 36318
rect 8318 36258 8370 36270
rect 8318 36194 8370 36206
rect 9886 36258 9938 36270
rect 9886 36194 9938 36206
rect 11006 36258 11058 36270
rect 11006 36194 11058 36206
rect 11230 36258 11282 36270
rect 30718 36258 30770 36270
rect 13682 36206 13694 36258
rect 13746 36206 13758 36258
rect 20626 36206 20638 36258
rect 20690 36206 20702 36258
rect 11230 36194 11282 36206
rect 30718 36194 30770 36206
rect 36206 36258 36258 36270
rect 36206 36194 36258 36206
rect 37102 36258 37154 36270
rect 37102 36194 37154 36206
rect 45726 36258 45778 36270
rect 45726 36194 45778 36206
rect 46958 36258 47010 36270
rect 46958 36194 47010 36206
rect 1344 36090 48608 36124
rect 1344 36038 19838 36090
rect 19890 36038 19942 36090
rect 19994 36038 20046 36090
rect 20098 36038 48608 36090
rect 1344 36004 48608 36038
rect 4734 35922 4786 35934
rect 3714 35870 3726 35922
rect 3778 35870 3790 35922
rect 4734 35858 4786 35870
rect 8206 35922 8258 35934
rect 12574 35922 12626 35934
rect 8978 35870 8990 35922
rect 9042 35870 9054 35922
rect 8206 35858 8258 35870
rect 12574 35858 12626 35870
rect 16494 35922 16546 35934
rect 16494 35858 16546 35870
rect 19406 35922 19458 35934
rect 47406 35922 47458 35934
rect 22418 35870 22430 35922
rect 22482 35870 22494 35922
rect 19406 35858 19458 35870
rect 47406 35858 47458 35870
rect 4286 35810 4338 35822
rect 10110 35810 10162 35822
rect 16718 35810 16770 35822
rect 21534 35810 21586 35822
rect 39902 35810 39954 35822
rect 7074 35758 7086 35810
rect 7138 35758 7150 35810
rect 13010 35758 13022 35810
rect 13074 35758 13086 35810
rect 17490 35758 17502 35810
rect 17554 35758 17566 35810
rect 22530 35758 22542 35810
rect 22594 35758 22606 35810
rect 26002 35758 26014 35810
rect 26066 35758 26078 35810
rect 27122 35758 27134 35810
rect 27186 35758 27198 35810
rect 29586 35758 29598 35810
rect 29650 35758 29662 35810
rect 37762 35758 37774 35810
rect 37826 35758 37838 35810
rect 4286 35746 4338 35758
rect 10110 35746 10162 35758
rect 16718 35746 16770 35758
rect 21534 35746 21586 35758
rect 39902 35746 39954 35758
rect 40126 35810 40178 35822
rect 40126 35746 40178 35758
rect 47630 35810 47682 35822
rect 47630 35746 47682 35758
rect 4062 35698 4114 35710
rect 9886 35698 9938 35710
rect 2930 35646 2942 35698
rect 2994 35646 3006 35698
rect 6178 35646 6190 35698
rect 6242 35646 6254 35698
rect 8754 35646 8766 35698
rect 8818 35646 8830 35698
rect 4062 35634 4114 35646
rect 9886 35634 9938 35646
rect 10334 35698 10386 35710
rect 16830 35698 16882 35710
rect 21086 35698 21138 35710
rect 31502 35698 31554 35710
rect 10994 35646 11006 35698
rect 11058 35646 11070 35698
rect 11666 35646 11678 35698
rect 11730 35646 11742 35698
rect 12002 35646 12014 35698
rect 12066 35646 12078 35698
rect 13346 35646 13358 35698
rect 13410 35646 13422 35698
rect 14242 35646 14254 35698
rect 14306 35646 14318 35698
rect 15810 35646 15822 35698
rect 15874 35646 15886 35698
rect 17378 35646 17390 35698
rect 17442 35646 17454 35698
rect 18610 35646 18622 35698
rect 18674 35646 18686 35698
rect 20402 35646 20414 35698
rect 20466 35646 20478 35698
rect 20626 35646 20638 35698
rect 20690 35646 20702 35698
rect 21858 35646 21870 35698
rect 21922 35646 21934 35698
rect 22194 35646 22206 35698
rect 22258 35646 22270 35698
rect 22978 35646 22990 35698
rect 23042 35646 23054 35698
rect 24098 35646 24110 35698
rect 24162 35646 24174 35698
rect 25778 35646 25790 35698
rect 25842 35646 25854 35698
rect 28578 35646 28590 35698
rect 28642 35646 28654 35698
rect 28914 35646 28926 35698
rect 28978 35646 28990 35698
rect 29474 35646 29486 35698
rect 29538 35646 29550 35698
rect 31154 35646 31166 35698
rect 31218 35646 31230 35698
rect 10334 35634 10386 35646
rect 16830 35634 16882 35646
rect 21086 35634 21138 35646
rect 31502 35634 31554 35646
rect 31726 35698 31778 35710
rect 38894 35698 38946 35710
rect 38546 35646 38558 35698
rect 38610 35646 38622 35698
rect 42690 35646 42702 35698
rect 42754 35646 42766 35698
rect 46274 35646 46286 35698
rect 46338 35646 46350 35698
rect 31726 35634 31778 35646
rect 38894 35634 38946 35646
rect 2270 35586 2322 35598
rect 5518 35586 5570 35598
rect 18174 35586 18226 35598
rect 30830 35586 30882 35598
rect 3042 35534 3054 35586
rect 3106 35534 3118 35586
rect 7634 35534 7646 35586
rect 7698 35534 7710 35586
rect 10882 35534 10894 35586
rect 10946 35534 10958 35586
rect 17490 35534 17502 35586
rect 17554 35534 17566 35586
rect 20738 35534 20750 35586
rect 20802 35534 20814 35586
rect 23650 35534 23662 35586
rect 23714 35534 23726 35586
rect 28354 35534 28366 35586
rect 28418 35534 28430 35586
rect 29698 35534 29710 35586
rect 29762 35534 29774 35586
rect 2270 35522 2322 35534
rect 5518 35522 5570 35534
rect 18174 35522 18226 35534
rect 30830 35522 30882 35534
rect 31614 35586 31666 35598
rect 31614 35522 31666 35534
rect 34414 35586 34466 35598
rect 46062 35586 46114 35598
rect 35634 35534 35646 35586
rect 35698 35534 35710 35586
rect 39330 35534 39342 35586
rect 39394 35534 39406 35586
rect 39778 35534 39790 35586
rect 39842 35534 39854 35586
rect 43362 35534 43374 35586
rect 43426 35534 43438 35586
rect 45490 35534 45502 35586
rect 45554 35534 45566 35586
rect 47282 35534 47294 35586
rect 47346 35534 47358 35586
rect 34414 35522 34466 35534
rect 46062 35522 46114 35534
rect 9662 35474 9714 35486
rect 9662 35410 9714 35422
rect 10446 35474 10498 35486
rect 45950 35474 46002 35486
rect 24098 35422 24110 35474
rect 24162 35422 24174 35474
rect 10446 35410 10498 35422
rect 45950 35410 46002 35422
rect 1344 35306 48608 35340
rect 1344 35254 4478 35306
rect 4530 35254 4582 35306
rect 4634 35254 4686 35306
rect 4738 35254 35198 35306
rect 35250 35254 35302 35306
rect 35354 35254 35406 35306
rect 35458 35254 48608 35306
rect 1344 35220 48608 35254
rect 2606 35138 2658 35150
rect 2606 35074 2658 35086
rect 4398 35138 4450 35150
rect 11006 35138 11058 35150
rect 6514 35086 6526 35138
rect 6578 35086 6590 35138
rect 4398 35074 4450 35086
rect 11006 35074 11058 35086
rect 11342 35138 11394 35150
rect 29374 35138 29426 35150
rect 18834 35086 18846 35138
rect 18898 35086 18910 35138
rect 11342 35074 11394 35086
rect 29374 35074 29426 35086
rect 20526 35026 20578 35038
rect 2818 34974 2830 35026
rect 2882 34974 2894 35026
rect 14466 34974 14478 35026
rect 14530 34974 14542 35026
rect 16370 34974 16382 35026
rect 16434 34974 16446 35026
rect 18498 34974 18510 35026
rect 18562 34974 18574 35026
rect 20526 34962 20578 34974
rect 21422 35026 21474 35038
rect 25118 35026 25170 35038
rect 23538 34974 23550 35026
rect 23602 34974 23614 35026
rect 21422 34962 21474 34974
rect 25118 34962 25170 34974
rect 28030 35026 28082 35038
rect 28030 34962 28082 34974
rect 29150 35026 29202 35038
rect 33630 35026 33682 35038
rect 33170 34974 33182 35026
rect 33234 34974 33246 35026
rect 29150 34962 29202 34974
rect 33630 34962 33682 34974
rect 43822 35026 43874 35038
rect 46050 34974 46062 35026
rect 46114 34974 46126 35026
rect 48178 34974 48190 35026
rect 48242 34974 48254 35026
rect 43822 34962 43874 34974
rect 4958 34914 5010 34926
rect 7758 34914 7810 34926
rect 19406 34914 19458 34926
rect 23214 34914 23266 34926
rect 27918 34914 27970 34926
rect 36990 34914 37042 34926
rect 38446 34914 38498 34926
rect 2930 34862 2942 34914
rect 2994 34862 3006 34914
rect 5842 34862 5854 34914
rect 5906 34862 5918 34914
rect 6402 34862 6414 34914
rect 6466 34862 6478 34914
rect 7186 34862 7198 34914
rect 7250 34862 7262 34914
rect 8754 34862 8766 34914
rect 8818 34862 8830 34914
rect 9986 34862 9998 34914
rect 10050 34862 10062 34914
rect 11666 34862 11678 34914
rect 11730 34862 11742 34914
rect 12114 34862 12126 34914
rect 12178 34862 12190 34914
rect 12898 34862 12910 34914
rect 12962 34862 12974 34914
rect 13794 34862 13806 34914
rect 13858 34862 13870 34914
rect 14130 34862 14142 34914
rect 14194 34862 14206 34914
rect 15698 34862 15710 34914
rect 15762 34862 15774 34914
rect 19618 34862 19630 34914
rect 19682 34862 19694 34914
rect 22754 34862 22766 34914
rect 22818 34862 22830 34914
rect 25330 34862 25342 34914
rect 25394 34862 25406 34914
rect 27570 34862 27582 34914
rect 27634 34862 27646 34914
rect 29698 34862 29710 34914
rect 29762 34862 29774 34914
rect 30370 34862 30382 34914
rect 30434 34862 30446 34914
rect 37426 34862 37438 34914
rect 37490 34862 37502 34914
rect 4958 34850 5010 34862
rect 7758 34850 7810 34862
rect 19406 34850 19458 34862
rect 23214 34850 23266 34862
rect 27918 34850 27970 34862
rect 36990 34850 37042 34862
rect 38446 34850 38498 34862
rect 44046 34914 44098 34926
rect 44046 34850 44098 34862
rect 44270 34914 44322 34926
rect 45378 34862 45390 34914
rect 45442 34862 45454 34914
rect 44270 34850 44322 34862
rect 3614 34802 3666 34814
rect 3614 34738 3666 34750
rect 4174 34802 4226 34814
rect 4174 34738 4226 34750
rect 5070 34802 5122 34814
rect 5070 34738 5122 34750
rect 7422 34802 7474 34814
rect 15038 34802 15090 34814
rect 8642 34750 8654 34802
rect 8706 34750 8718 34802
rect 12786 34750 12798 34802
rect 12850 34750 12862 34802
rect 7422 34738 7474 34750
rect 15038 34738 15090 34750
rect 15374 34802 15426 34814
rect 15374 34738 15426 34750
rect 19294 34802 19346 34814
rect 19294 34738 19346 34750
rect 21310 34802 21362 34814
rect 38782 34802 38834 34814
rect 31042 34750 31054 34802
rect 31106 34750 31118 34802
rect 21310 34738 21362 34750
rect 38782 34738 38834 34750
rect 39118 34802 39170 34814
rect 39118 34738 39170 34750
rect 43150 34802 43202 34814
rect 43150 34738 43202 34750
rect 43710 34802 43762 34814
rect 43710 34738 43762 34750
rect 2382 34690 2434 34702
rect 2382 34626 2434 34638
rect 3278 34690 3330 34702
rect 3278 34626 3330 34638
rect 3502 34690 3554 34702
rect 3502 34626 3554 34638
rect 4286 34690 4338 34702
rect 4286 34626 4338 34638
rect 4846 34690 4898 34702
rect 15150 34690 15202 34702
rect 13794 34638 13806 34690
rect 13858 34638 13870 34690
rect 4846 34626 4898 34638
rect 15150 34626 15202 34638
rect 19966 34690 20018 34702
rect 19966 34626 20018 34638
rect 21534 34690 21586 34702
rect 21534 34626 21586 34638
rect 21758 34690 21810 34702
rect 21758 34626 21810 34638
rect 28702 34690 28754 34702
rect 28702 34626 28754 34638
rect 37886 34690 37938 34702
rect 37886 34626 37938 34638
rect 39566 34690 39618 34702
rect 39566 34626 39618 34638
rect 43262 34690 43314 34702
rect 43262 34626 43314 34638
rect 43486 34690 43538 34702
rect 43486 34626 43538 34638
rect 1344 34522 48608 34556
rect 1344 34470 19838 34522
rect 19890 34470 19942 34522
rect 19994 34470 20046 34522
rect 20098 34470 48608 34522
rect 1344 34436 48608 34470
rect 7198 34354 7250 34366
rect 7198 34290 7250 34302
rect 7422 34354 7474 34366
rect 10782 34354 10834 34366
rect 8866 34302 8878 34354
rect 8930 34302 8942 34354
rect 7422 34290 7474 34302
rect 10782 34290 10834 34302
rect 13694 34354 13746 34366
rect 24222 34354 24274 34366
rect 21858 34302 21870 34354
rect 21922 34302 21934 34354
rect 13694 34290 13746 34302
rect 24222 34290 24274 34302
rect 25454 34354 25506 34366
rect 25454 34290 25506 34302
rect 25566 34354 25618 34366
rect 25566 34290 25618 34302
rect 25678 34354 25730 34366
rect 25678 34290 25730 34302
rect 25790 34354 25842 34366
rect 25790 34290 25842 34302
rect 29374 34354 29426 34366
rect 29374 34290 29426 34302
rect 31054 34354 31106 34366
rect 31054 34290 31106 34302
rect 31950 34354 32002 34366
rect 31950 34290 32002 34302
rect 36094 34354 36146 34366
rect 36094 34290 36146 34302
rect 3390 34242 3442 34254
rect 7534 34242 7586 34254
rect 11342 34242 11394 34254
rect 4834 34190 4846 34242
rect 4898 34190 4910 34242
rect 8306 34190 8318 34242
rect 8370 34190 8382 34242
rect 3390 34178 3442 34190
rect 7534 34178 7586 34190
rect 11342 34178 11394 34190
rect 14254 34242 14306 34254
rect 14254 34178 14306 34190
rect 15598 34242 15650 34254
rect 17278 34242 17330 34254
rect 19966 34242 20018 34254
rect 26014 34242 26066 34254
rect 15922 34190 15934 34242
rect 15986 34190 15998 34242
rect 16706 34190 16718 34242
rect 16770 34190 16782 34242
rect 17826 34190 17838 34242
rect 17890 34190 17902 34242
rect 18162 34190 18174 34242
rect 18226 34190 18238 34242
rect 20626 34190 20638 34242
rect 20690 34190 20702 34242
rect 15598 34178 15650 34190
rect 17278 34178 17330 34190
rect 19966 34178 20018 34190
rect 26014 34178 26066 34190
rect 30046 34242 30098 34254
rect 30046 34178 30098 34190
rect 31278 34242 31330 34254
rect 31278 34178 31330 34190
rect 31502 34242 31554 34254
rect 31502 34178 31554 34190
rect 31838 34242 31890 34254
rect 34862 34242 34914 34254
rect 33058 34190 33070 34242
rect 33122 34190 33134 34242
rect 31838 34178 31890 34190
rect 34862 34178 34914 34190
rect 37326 34242 37378 34254
rect 37326 34178 37378 34190
rect 10558 34130 10610 34142
rect 3602 34078 3614 34130
rect 3666 34078 3678 34130
rect 4050 34078 4062 34130
rect 4114 34078 4126 34130
rect 8194 34078 8206 34130
rect 8258 34078 8270 34130
rect 8978 34078 8990 34130
rect 9042 34078 9054 34130
rect 10558 34066 10610 34078
rect 12238 34130 12290 34142
rect 15710 34130 15762 34142
rect 15250 34078 15262 34130
rect 15314 34078 15326 34130
rect 12238 34066 12290 34078
rect 15710 34066 15762 34078
rect 17502 34130 17554 34142
rect 17502 34066 17554 34078
rect 19406 34130 19458 34142
rect 24110 34130 24162 34142
rect 20514 34078 20526 34130
rect 20578 34078 20590 34130
rect 22306 34078 22318 34130
rect 22370 34078 22382 34130
rect 23090 34078 23102 34130
rect 23154 34078 23166 34130
rect 19406 34066 19458 34078
rect 24110 34066 24162 34078
rect 24334 34130 24386 34142
rect 26574 34130 26626 34142
rect 29262 34130 29314 34142
rect 24658 34078 24670 34130
rect 24722 34078 24734 34130
rect 28354 34078 28366 34130
rect 28418 34078 28430 34130
rect 24334 34066 24386 34078
rect 26574 34066 26626 34078
rect 29262 34066 29314 34078
rect 29598 34130 29650 34142
rect 29598 34066 29650 34078
rect 30830 34130 30882 34142
rect 34750 34130 34802 34142
rect 33730 34078 33742 34130
rect 33794 34078 33806 34130
rect 34514 34078 34526 34130
rect 34578 34078 34590 34130
rect 30830 34066 30882 34078
rect 34750 34066 34802 34078
rect 35086 34130 35138 34142
rect 35086 34066 35138 34078
rect 37214 34130 37266 34142
rect 44046 34130 44098 34142
rect 41010 34078 41022 34130
rect 41074 34078 41086 34130
rect 37214 34066 37266 34078
rect 44046 34066 44098 34078
rect 44382 34130 44434 34142
rect 44382 34066 44434 34078
rect 44606 34130 44658 34142
rect 45378 34078 45390 34130
rect 45442 34078 45454 34130
rect 44606 34066 44658 34078
rect 13470 34018 13522 34030
rect 6962 33966 6974 34018
rect 7026 33966 7038 34018
rect 13470 33954 13522 33966
rect 19182 34018 19234 34030
rect 21310 34018 21362 34030
rect 26350 34018 26402 34030
rect 28814 34018 28866 34030
rect 35534 34018 35586 34030
rect 44270 34018 44322 34030
rect 20850 33966 20862 34018
rect 20914 33966 20926 34018
rect 22530 33966 22542 34018
rect 22594 33966 22606 34018
rect 23202 33966 23214 34018
rect 23266 33966 23278 34018
rect 28466 33966 28478 34018
rect 28530 33966 28542 34018
rect 33842 33966 33854 34018
rect 33906 33966 33918 34018
rect 41682 33966 41694 34018
rect 41746 33966 41758 34018
rect 43810 33966 43822 34018
rect 43874 33966 43886 34018
rect 46050 33966 46062 34018
rect 46114 33966 46126 34018
rect 48178 33966 48190 34018
rect 48242 33966 48254 34018
rect 19182 33954 19234 33966
rect 21310 33954 21362 33966
rect 26350 33954 26402 33966
rect 28814 33954 28866 33966
rect 35534 33954 35586 33966
rect 44270 33954 44322 33966
rect 21534 33906 21586 33918
rect 29822 33906 29874 33918
rect 26898 33854 26910 33906
rect 26962 33854 26974 33906
rect 21534 33842 21586 33854
rect 29822 33842 29874 33854
rect 30158 33906 30210 33918
rect 30158 33842 30210 33854
rect 31950 33906 32002 33918
rect 31950 33842 32002 33854
rect 37326 33906 37378 33918
rect 37326 33842 37378 33854
rect 1344 33738 48608 33772
rect 1344 33686 4478 33738
rect 4530 33686 4582 33738
rect 4634 33686 4686 33738
rect 4738 33686 35198 33738
rect 35250 33686 35302 33738
rect 35354 33686 35406 33738
rect 35458 33686 48608 33738
rect 1344 33652 48608 33686
rect 2718 33570 2770 33582
rect 2718 33506 2770 33518
rect 3502 33570 3554 33582
rect 3502 33506 3554 33518
rect 14030 33570 14082 33582
rect 28702 33570 28754 33582
rect 44942 33570 44994 33582
rect 26562 33518 26574 33570
rect 26626 33518 26638 33570
rect 30818 33518 30830 33570
rect 30882 33518 30894 33570
rect 14030 33506 14082 33518
rect 28702 33506 28754 33518
rect 44942 33506 44994 33518
rect 2606 33458 2658 33470
rect 5742 33458 5794 33470
rect 9998 33458 10050 33470
rect 33182 33458 33234 33470
rect 3602 33406 3614 33458
rect 3666 33406 3678 33458
rect 6626 33406 6638 33458
rect 6690 33406 6702 33458
rect 12338 33406 12350 33458
rect 12402 33406 12414 33458
rect 18050 33406 18062 33458
rect 18114 33406 18126 33458
rect 20290 33406 20302 33458
rect 20354 33406 20366 33458
rect 26786 33406 26798 33458
rect 26850 33406 26862 33458
rect 30594 33406 30606 33458
rect 30658 33406 30670 33458
rect 36418 33406 36430 33458
rect 36482 33406 36494 33458
rect 36978 33406 36990 33458
rect 37042 33406 37054 33458
rect 43138 33406 43150 33458
rect 43202 33406 43214 33458
rect 2606 33394 2658 33406
rect 5742 33394 5794 33406
rect 9998 33394 10050 33406
rect 33182 33394 33234 33406
rect 13918 33346 13970 33358
rect 3266 33294 3278 33346
rect 3330 33294 3342 33346
rect 3714 33294 3726 33346
rect 3778 33294 3790 33346
rect 5058 33294 5070 33346
rect 5122 33294 5134 33346
rect 9090 33294 9102 33346
rect 9154 33294 9166 33346
rect 10770 33294 10782 33346
rect 10834 33294 10846 33346
rect 12450 33294 12462 33346
rect 12514 33294 12526 33346
rect 13918 33282 13970 33294
rect 15262 33346 15314 33358
rect 22094 33346 22146 33358
rect 24782 33346 24834 33358
rect 25678 33346 25730 33358
rect 27806 33346 27858 33358
rect 32286 33346 32338 33358
rect 43934 33346 43986 33358
rect 17042 33294 17054 33346
rect 17106 33294 17118 33346
rect 17378 33294 17390 33346
rect 17442 33294 17454 33346
rect 19058 33294 19070 33346
rect 19122 33294 19134 33346
rect 22306 33294 22318 33346
rect 22370 33294 22382 33346
rect 25218 33294 25230 33346
rect 25282 33294 25294 33346
rect 26338 33294 26350 33346
rect 26402 33294 26414 33346
rect 27458 33294 27470 33346
rect 27522 33294 27534 33346
rect 28242 33294 28254 33346
rect 28306 33294 28318 33346
rect 29922 33294 29934 33346
rect 29986 33294 29998 33346
rect 31042 33294 31054 33346
rect 31106 33294 31118 33346
rect 32722 33294 32734 33346
rect 32786 33294 32798 33346
rect 33618 33294 33630 33346
rect 33682 33294 33694 33346
rect 39890 33294 39902 33346
rect 39954 33294 39966 33346
rect 40338 33294 40350 33346
rect 40402 33294 40414 33346
rect 15262 33282 15314 33294
rect 22094 33282 22146 33294
rect 24782 33282 24834 33294
rect 25678 33282 25730 33294
rect 27806 33282 27858 33294
rect 32286 33282 32338 33294
rect 43934 33282 43986 33294
rect 45726 33346 45778 33358
rect 45726 33282 45778 33294
rect 46174 33346 46226 33358
rect 46174 33282 46226 33294
rect 46622 33346 46674 33358
rect 46622 33282 46674 33294
rect 2494 33234 2546 33246
rect 2494 33170 2546 33182
rect 4734 33234 4786 33246
rect 8878 33234 8930 33246
rect 16046 33234 16098 33246
rect 20302 33234 20354 33246
rect 7410 33182 7422 33234
rect 7474 33182 7486 33234
rect 10658 33182 10670 33234
rect 10722 33182 10734 33234
rect 12898 33182 12910 33234
rect 12962 33182 12974 33234
rect 17938 33182 17950 33234
rect 18002 33182 18014 33234
rect 4734 33170 4786 33182
rect 8878 33170 8930 33182
rect 16046 33170 16098 33182
rect 20302 33170 20354 33182
rect 20750 33234 20802 33246
rect 20750 33170 20802 33182
rect 22878 33234 22930 33246
rect 22878 33170 22930 33182
rect 27918 33234 27970 33246
rect 29150 33234 29202 33246
rect 43598 33234 43650 33246
rect 28130 33182 28142 33234
rect 28194 33182 28206 33234
rect 34290 33182 34302 33234
rect 34354 33182 34366 33234
rect 39106 33182 39118 33234
rect 39170 33182 39182 33234
rect 41010 33182 41022 33234
rect 41074 33182 41086 33234
rect 27918 33170 27970 33182
rect 29150 33170 29202 33182
rect 43598 33170 43650 33182
rect 44830 33234 44882 33246
rect 44830 33170 44882 33182
rect 44942 33234 44994 33246
rect 44942 33170 44994 33182
rect 46398 33234 46450 33246
rect 46398 33170 46450 33182
rect 46846 33234 46898 33246
rect 46846 33170 46898 33182
rect 46958 33234 47010 33246
rect 46958 33170 47010 33182
rect 4846 33122 4898 33134
rect 4846 33058 4898 33070
rect 6302 33122 6354 33134
rect 6302 33058 6354 33070
rect 7086 33122 7138 33134
rect 7086 33058 7138 33070
rect 7758 33122 7810 33134
rect 7758 33058 7810 33070
rect 8318 33122 8370 33134
rect 8318 33058 8370 33070
rect 9662 33122 9714 33134
rect 9662 33058 9714 33070
rect 13694 33122 13746 33134
rect 13694 33058 13746 33070
rect 14030 33122 14082 33134
rect 20526 33122 20578 33134
rect 15138 33070 15150 33122
rect 15202 33070 15214 33122
rect 14030 33058 14082 33070
rect 20526 33058 20578 33070
rect 23774 33122 23826 33134
rect 23774 33058 23826 33070
rect 24446 33122 24498 33134
rect 24446 33058 24498 33070
rect 29486 33122 29538 33134
rect 29486 33058 29538 33070
rect 31838 33122 31890 33134
rect 31838 33058 31890 33070
rect 43710 33122 43762 33134
rect 43710 33058 43762 33070
rect 46062 33122 46114 33134
rect 46062 33058 46114 33070
rect 47630 33122 47682 33134
rect 48190 33122 48242 33134
rect 47842 33070 47854 33122
rect 47906 33070 47918 33122
rect 47630 33058 47682 33070
rect 48190 33058 48242 33070
rect 1344 32954 48608 32988
rect 1344 32902 19838 32954
rect 19890 32902 19942 32954
rect 19994 32902 20046 32954
rect 20098 32902 48608 32954
rect 1344 32868 48608 32902
rect 5070 32786 5122 32798
rect 5070 32722 5122 32734
rect 6974 32786 7026 32798
rect 6974 32722 7026 32734
rect 8878 32786 8930 32798
rect 20862 32786 20914 32798
rect 17714 32734 17726 32786
rect 17778 32734 17790 32786
rect 8878 32722 8930 32734
rect 20862 32722 20914 32734
rect 20974 32786 21026 32798
rect 20974 32722 21026 32734
rect 33406 32786 33458 32798
rect 33406 32722 33458 32734
rect 34638 32786 34690 32798
rect 34638 32722 34690 32734
rect 35758 32786 35810 32798
rect 35758 32722 35810 32734
rect 37550 32786 37602 32798
rect 37550 32722 37602 32734
rect 40014 32786 40066 32798
rect 40014 32722 40066 32734
rect 43822 32786 43874 32798
rect 43822 32722 43874 32734
rect 45390 32786 45442 32798
rect 45390 32722 45442 32734
rect 45614 32786 45666 32798
rect 45614 32722 45666 32734
rect 46958 32786 47010 32798
rect 46958 32722 47010 32734
rect 9774 32674 9826 32686
rect 13134 32674 13186 32686
rect 10882 32622 10894 32674
rect 10946 32622 10958 32674
rect 9774 32610 9826 32622
rect 13134 32610 13186 32622
rect 19182 32674 19234 32686
rect 19182 32610 19234 32622
rect 21198 32674 21250 32686
rect 21198 32610 21250 32622
rect 21310 32674 21362 32686
rect 33294 32674 33346 32686
rect 30146 32622 30158 32674
rect 30210 32622 30222 32674
rect 21310 32610 21362 32622
rect 33294 32610 33346 32622
rect 33854 32674 33906 32686
rect 33854 32610 33906 32622
rect 34078 32674 34130 32686
rect 34078 32610 34130 32622
rect 34750 32674 34802 32686
rect 34750 32610 34802 32622
rect 35870 32674 35922 32686
rect 35870 32610 35922 32622
rect 37438 32674 37490 32686
rect 37438 32610 37490 32622
rect 41246 32674 41298 32686
rect 41246 32610 41298 32622
rect 43486 32674 43538 32686
rect 43486 32610 43538 32622
rect 43598 32674 43650 32686
rect 43598 32610 43650 32622
rect 44046 32674 44098 32686
rect 44046 32610 44098 32622
rect 44830 32674 44882 32686
rect 44830 32610 44882 32622
rect 44942 32674 44994 32686
rect 44942 32610 44994 32622
rect 45278 32674 45330 32686
rect 45278 32610 45330 32622
rect 47406 32674 47458 32686
rect 47406 32610 47458 32622
rect 47518 32674 47570 32686
rect 47518 32610 47570 32622
rect 6078 32562 6130 32574
rect 3826 32510 3838 32562
rect 3890 32510 3902 32562
rect 4610 32510 4622 32562
rect 4674 32510 4686 32562
rect 6078 32498 6130 32510
rect 6190 32562 6242 32574
rect 6190 32498 6242 32510
rect 6526 32562 6578 32574
rect 6526 32498 6578 32510
rect 8990 32562 9042 32574
rect 18622 32562 18674 32574
rect 22990 32562 23042 32574
rect 26574 32562 26626 32574
rect 9986 32510 9998 32562
rect 10050 32510 10062 32562
rect 10994 32510 11006 32562
rect 11058 32510 11070 32562
rect 11330 32510 11342 32562
rect 11394 32510 11406 32562
rect 12338 32510 12350 32562
rect 12402 32510 12414 32562
rect 13570 32510 13582 32562
rect 13634 32510 13646 32562
rect 14914 32510 14926 32562
rect 14978 32510 14990 32562
rect 16594 32510 16606 32562
rect 16658 32510 16670 32562
rect 19618 32510 19630 32562
rect 19682 32510 19694 32562
rect 20178 32510 20190 32562
rect 20242 32510 20254 32562
rect 20402 32510 20414 32562
rect 20466 32510 20478 32562
rect 22082 32510 22094 32562
rect 22146 32510 22158 32562
rect 22642 32510 22654 32562
rect 22706 32510 22718 32562
rect 23202 32510 23214 32562
rect 23266 32510 23278 32562
rect 24546 32510 24558 32562
rect 24610 32510 24622 32562
rect 25554 32510 25566 32562
rect 25618 32510 25630 32562
rect 8990 32498 9042 32510
rect 18622 32498 18674 32510
rect 22990 32498 23042 32510
rect 26574 32498 26626 32510
rect 28366 32562 28418 32574
rect 39678 32562 39730 32574
rect 44606 32562 44658 32574
rect 29026 32510 29038 32562
rect 29090 32510 29102 32562
rect 31042 32510 31054 32562
rect 31106 32510 31118 32562
rect 32386 32510 32398 32562
rect 32450 32510 32462 32562
rect 37762 32510 37774 32562
rect 37826 32510 37838 32562
rect 40226 32510 40238 32562
rect 40290 32510 40302 32562
rect 44258 32510 44270 32562
rect 44322 32510 44334 32562
rect 28366 32498 28418 32510
rect 39678 32498 39730 32510
rect 44606 32498 44658 32510
rect 46734 32562 46786 32574
rect 46734 32498 46786 32510
rect 47070 32562 47122 32574
rect 47070 32498 47122 32510
rect 6414 32450 6466 32462
rect 1698 32398 1710 32450
rect 1762 32398 1774 32450
rect 6414 32386 6466 32398
rect 7758 32450 7810 32462
rect 7758 32386 7810 32398
rect 7982 32450 8034 32462
rect 7982 32386 8034 32398
rect 8430 32450 8482 32462
rect 18286 32450 18338 32462
rect 31726 32450 31778 32462
rect 10882 32398 10894 32450
rect 10946 32398 10958 32450
rect 11666 32398 11678 32450
rect 11730 32398 11742 32450
rect 12002 32398 12014 32450
rect 12066 32398 12078 32450
rect 16482 32398 16494 32450
rect 16546 32398 16558 32450
rect 21970 32398 21982 32450
rect 22034 32398 22046 32450
rect 25890 32398 25902 32450
rect 25954 32398 25966 32450
rect 29586 32398 29598 32450
rect 29650 32398 29662 32450
rect 8430 32386 8482 32398
rect 18286 32386 18338 32398
rect 31726 32386 31778 32398
rect 32062 32450 32114 32462
rect 36654 32450 36706 32462
rect 32274 32398 32286 32450
rect 32338 32398 32350 32450
rect 34178 32398 34190 32450
rect 34242 32398 34254 32450
rect 32062 32386 32114 32398
rect 36654 32386 36706 32398
rect 8878 32338 8930 32350
rect 18062 32338 18114 32350
rect 24222 32338 24274 32350
rect 7410 32286 7422 32338
rect 7474 32286 7486 32338
rect 15362 32286 15374 32338
rect 15426 32286 15438 32338
rect 23426 32286 23438 32338
rect 23490 32286 23502 32338
rect 8878 32274 8930 32286
rect 18062 32274 18114 32286
rect 24222 32274 24274 32286
rect 24558 32338 24610 32350
rect 24558 32274 24610 32286
rect 33406 32338 33458 32350
rect 33406 32274 33458 32286
rect 34526 32338 34578 32350
rect 34526 32274 34578 32286
rect 39902 32338 39954 32350
rect 39902 32274 39954 32286
rect 41470 32338 41522 32350
rect 41470 32274 41522 32286
rect 41806 32338 41858 32350
rect 41806 32274 41858 32286
rect 47518 32338 47570 32350
rect 47518 32274 47570 32286
rect 1344 32170 48608 32204
rect 1344 32118 4478 32170
rect 4530 32118 4582 32170
rect 4634 32118 4686 32170
rect 4738 32118 35198 32170
rect 35250 32118 35302 32170
rect 35354 32118 35406 32170
rect 35458 32118 48608 32170
rect 1344 32084 48608 32118
rect 19966 32002 20018 32014
rect 8866 31950 8878 32002
rect 8930 31950 8942 32002
rect 19966 31938 20018 31950
rect 20190 32002 20242 32014
rect 20190 31938 20242 31950
rect 23998 32002 24050 32014
rect 28478 32002 28530 32014
rect 25442 31950 25454 32002
rect 25506 31950 25518 32002
rect 23998 31938 24050 31950
rect 28478 31938 28530 31950
rect 33406 32002 33458 32014
rect 33406 31938 33458 31950
rect 34862 32002 34914 32014
rect 34862 31938 34914 31950
rect 4958 31890 5010 31902
rect 4958 31826 5010 31838
rect 7310 31890 7362 31902
rect 7310 31826 7362 31838
rect 7870 31890 7922 31902
rect 16158 31890 16210 31902
rect 20750 31890 20802 31902
rect 29150 31890 29202 31902
rect 35758 31890 35810 31902
rect 10994 31838 11006 31890
rect 11058 31838 11070 31890
rect 14354 31838 14366 31890
rect 14418 31838 14430 31890
rect 16930 31838 16942 31890
rect 16994 31838 17006 31890
rect 20402 31838 20414 31890
rect 20466 31838 20478 31890
rect 21522 31838 21534 31890
rect 21586 31838 21598 31890
rect 25218 31838 25230 31890
rect 25282 31838 25294 31890
rect 30146 31838 30158 31890
rect 30210 31838 30222 31890
rect 32274 31838 32286 31890
rect 32338 31838 32350 31890
rect 7870 31826 7922 31838
rect 16158 31826 16210 31838
rect 20750 31826 20802 31838
rect 29150 31826 29202 31838
rect 35758 31826 35810 31838
rect 38222 31890 38274 31902
rect 44146 31838 44158 31890
rect 44210 31838 44222 31890
rect 48178 31838 48190 31890
rect 48242 31838 48254 31890
rect 38222 31826 38274 31838
rect 4174 31778 4226 31790
rect 2594 31726 2606 31778
rect 2658 31726 2670 31778
rect 4174 31714 4226 31726
rect 5742 31778 5794 31790
rect 5742 31714 5794 31726
rect 6190 31778 6242 31790
rect 6190 31714 6242 31726
rect 6414 31778 6466 31790
rect 9774 31778 9826 31790
rect 6850 31726 6862 31778
rect 6914 31726 6926 31778
rect 8306 31726 8318 31778
rect 8370 31726 8382 31778
rect 9202 31726 9214 31778
rect 9266 31726 9278 31778
rect 6414 31714 6466 31726
rect 9774 31714 9826 31726
rect 9886 31778 9938 31790
rect 20638 31778 20690 31790
rect 23774 31778 23826 31790
rect 36094 31778 36146 31790
rect 12450 31726 12462 31778
rect 12514 31726 12526 31778
rect 14242 31726 14254 31778
rect 14306 31726 14318 31778
rect 15026 31726 15038 31778
rect 15090 31726 15102 31778
rect 16818 31726 16830 31778
rect 16882 31726 16894 31778
rect 18274 31726 18286 31778
rect 18338 31726 18350 31778
rect 21970 31726 21982 31778
rect 22034 31726 22046 31778
rect 22978 31726 22990 31778
rect 23042 31726 23054 31778
rect 23426 31726 23438 31778
rect 23490 31726 23502 31778
rect 26786 31726 26798 31778
rect 26850 31726 26862 31778
rect 28242 31726 28254 31778
rect 28306 31726 28318 31778
rect 29586 31726 29598 31778
rect 29650 31726 29662 31778
rect 33058 31726 33070 31778
rect 33122 31726 33134 31778
rect 9886 31714 9938 31726
rect 20638 31714 20690 31726
rect 23774 31714 23826 31726
rect 36094 31714 36146 31726
rect 38110 31778 38162 31790
rect 41346 31726 41358 31778
rect 41410 31726 41422 31778
rect 45378 31726 45390 31778
rect 45442 31726 45454 31778
rect 38110 31714 38162 31726
rect 4510 31666 4562 31678
rect 2034 31614 2046 31666
rect 2098 31614 2110 31666
rect 3714 31614 3726 31666
rect 3778 31614 3790 31666
rect 4510 31602 4562 31614
rect 9438 31666 9490 31678
rect 16270 31666 16322 31678
rect 21310 31666 21362 31678
rect 25678 31666 25730 31678
rect 33742 31666 33794 31678
rect 13570 31614 13582 31666
rect 13634 31614 13646 31666
rect 17490 31614 17502 31666
rect 17554 31614 17566 31666
rect 22418 31614 22430 31666
rect 22482 31614 22494 31666
rect 22754 31614 22766 31666
rect 22818 31614 22830 31666
rect 28018 31614 28030 31666
rect 28082 31614 28094 31666
rect 9438 31602 9490 31614
rect 16270 31602 16322 31614
rect 21310 31602 21362 31614
rect 25678 31602 25730 31614
rect 33742 31602 33794 31614
rect 34302 31666 34354 31678
rect 34302 31602 34354 31614
rect 35198 31666 35250 31678
rect 35198 31602 35250 31614
rect 37774 31666 37826 31678
rect 37774 31602 37826 31614
rect 38334 31666 38386 31678
rect 38334 31602 38386 31614
rect 38670 31666 38722 31678
rect 42018 31614 42030 31666
rect 42082 31614 42094 31666
rect 46050 31614 46062 31666
rect 46114 31614 46126 31666
rect 38670 31602 38722 31614
rect 4398 31554 4450 31566
rect 3602 31502 3614 31554
rect 3666 31502 3678 31554
rect 4398 31490 4450 31502
rect 6302 31554 6354 31566
rect 6302 31490 6354 31502
rect 15710 31554 15762 31566
rect 15710 31490 15762 31502
rect 16046 31554 16098 31566
rect 16046 31490 16098 31502
rect 33518 31554 33570 31566
rect 33518 31490 33570 31502
rect 33966 31554 34018 31566
rect 33966 31490 34018 31502
rect 34190 31554 34242 31566
rect 34190 31490 34242 31502
rect 34974 31554 35026 31566
rect 34974 31490 35026 31502
rect 37438 31554 37490 31566
rect 37438 31490 37490 31502
rect 39006 31554 39058 31566
rect 39006 31490 39058 31502
rect 1344 31386 48608 31420
rect 1344 31334 19838 31386
rect 19890 31334 19942 31386
rect 19994 31334 20046 31386
rect 20098 31334 48608 31386
rect 1344 31300 48608 31334
rect 3390 31218 3442 31230
rect 3390 31154 3442 31166
rect 7310 31218 7362 31230
rect 7310 31154 7362 31166
rect 7534 31218 7586 31230
rect 8990 31218 9042 31230
rect 7970 31166 7982 31218
rect 8034 31166 8046 31218
rect 7534 31154 7586 31166
rect 8990 31154 9042 31166
rect 9886 31218 9938 31230
rect 15374 31218 15426 31230
rect 11218 31166 11230 31218
rect 11282 31166 11294 31218
rect 9886 31154 9938 31166
rect 15374 31154 15426 31166
rect 18510 31218 18562 31230
rect 36990 31218 37042 31230
rect 30930 31166 30942 31218
rect 30994 31166 31006 31218
rect 18510 31154 18562 31166
rect 36990 31154 37042 31166
rect 37214 31218 37266 31230
rect 37214 31154 37266 31166
rect 38110 31218 38162 31230
rect 38110 31154 38162 31166
rect 39678 31218 39730 31230
rect 39678 31154 39730 31166
rect 42478 31218 42530 31230
rect 42478 31154 42530 31166
rect 43822 31218 43874 31230
rect 43822 31154 43874 31166
rect 44494 31218 44546 31230
rect 44494 31154 44546 31166
rect 44718 31218 44770 31230
rect 44718 31154 44770 31166
rect 45278 31218 45330 31230
rect 45278 31154 45330 31166
rect 46958 31218 47010 31230
rect 46958 31154 47010 31166
rect 47854 31218 47906 31230
rect 47854 31154 47906 31166
rect 2718 31106 2770 31118
rect 2718 31042 2770 31054
rect 2942 31106 2994 31118
rect 7646 31106 7698 31118
rect 11790 31106 11842 31118
rect 15038 31106 15090 31118
rect 4946 31054 4958 31106
rect 5010 31054 5022 31106
rect 10210 31054 10222 31106
rect 10274 31054 10286 31106
rect 14578 31054 14590 31106
rect 14642 31054 14654 31106
rect 2942 31042 2994 31054
rect 7646 31042 7698 31054
rect 11790 31042 11842 31054
rect 15038 31042 15090 31054
rect 15150 31106 15202 31118
rect 15150 31042 15202 31054
rect 20974 31106 21026 31118
rect 20974 31042 21026 31054
rect 24558 31106 24610 31118
rect 32398 31106 32450 31118
rect 28578 31054 28590 31106
rect 28642 31054 28654 31106
rect 31266 31054 31278 31106
rect 31330 31054 31342 31106
rect 31602 31054 31614 31106
rect 31666 31054 31678 31106
rect 24558 31042 24610 31054
rect 32398 31042 32450 31054
rect 32510 31106 32562 31118
rect 32510 31042 32562 31054
rect 39230 31106 39282 31118
rect 39230 31042 39282 31054
rect 41358 31106 41410 31118
rect 43710 31106 43762 31118
rect 42802 31054 42814 31106
rect 42866 31054 42878 31106
rect 41358 31042 41410 31054
rect 43710 31042 43762 31054
rect 44046 31106 44098 31118
rect 44046 31042 44098 31054
rect 44830 31106 44882 31118
rect 44830 31042 44882 31054
rect 46398 31106 46450 31118
rect 46398 31042 46450 31054
rect 47182 31106 47234 31118
rect 47182 31042 47234 31054
rect 2382 30994 2434 31006
rect 2382 30930 2434 30942
rect 3278 30994 3330 31006
rect 3278 30930 3330 30942
rect 3502 30994 3554 31006
rect 3502 30930 3554 30942
rect 3950 30994 4002 31006
rect 9550 30994 9602 31006
rect 12798 30994 12850 31006
rect 4274 30942 4286 30994
rect 4338 30942 4350 30994
rect 10770 30942 10782 30994
rect 10834 30942 10846 30994
rect 11106 30942 11118 30994
rect 11170 30942 11182 30994
rect 12338 30942 12350 30994
rect 12402 30942 12414 30994
rect 3950 30930 4002 30942
rect 9550 30930 9602 30942
rect 12798 30930 12850 30942
rect 13470 30994 13522 31006
rect 13470 30930 13522 30942
rect 13582 30994 13634 31006
rect 17390 30994 17442 31006
rect 16594 30942 16606 30994
rect 16658 30942 16670 30994
rect 13582 30930 13634 30942
rect 17390 30930 17442 30942
rect 17950 30994 18002 31006
rect 17950 30930 18002 30942
rect 18846 30994 18898 31006
rect 18846 30930 18898 30942
rect 20078 30994 20130 31006
rect 20078 30930 20130 30942
rect 20526 30994 20578 31006
rect 20526 30930 20578 30942
rect 20638 30994 20690 31006
rect 37662 30994 37714 31006
rect 21522 30942 21534 30994
rect 21586 30942 21598 30994
rect 23874 30942 23886 30994
rect 23938 30942 23950 30994
rect 25218 30942 25230 30994
rect 25282 30942 25294 30994
rect 31826 30942 31838 30994
rect 31890 30942 31902 30994
rect 33170 30942 33182 30994
rect 33234 30942 33246 30994
rect 33842 30942 33854 30994
rect 33906 30942 33918 30994
rect 37426 30942 37438 30994
rect 37490 30942 37502 30994
rect 20638 30930 20690 30942
rect 37662 30930 37714 30942
rect 38222 30994 38274 31006
rect 38222 30930 38274 30942
rect 38334 30994 38386 31006
rect 38334 30930 38386 30942
rect 38670 30994 38722 31006
rect 38670 30930 38722 30942
rect 39006 30994 39058 31006
rect 44270 30994 44322 31006
rect 46062 30994 46114 31006
rect 41682 30942 41694 30994
rect 41746 30942 41758 30994
rect 45490 30942 45502 30994
rect 45554 30942 45566 30994
rect 39006 30930 39058 30942
rect 44270 30930 44322 30942
rect 46062 30930 46114 30942
rect 46734 30994 46786 31006
rect 46734 30930 46786 30942
rect 47294 30994 47346 31006
rect 47294 30930 47346 30942
rect 47742 30994 47794 31006
rect 47742 30930 47794 30942
rect 2494 30882 2546 30894
rect 8542 30882 8594 30894
rect 20862 30882 20914 30894
rect 36542 30882 36594 30894
rect 39118 30882 39170 30894
rect 7074 30830 7086 30882
rect 7138 30830 7150 30882
rect 12450 30830 12462 30882
rect 12514 30830 12526 30882
rect 18610 30830 18622 30882
rect 18674 30830 18686 30882
rect 19618 30830 19630 30882
rect 19682 30830 19694 30882
rect 21858 30830 21870 30882
rect 21922 30830 21934 30882
rect 24658 30830 24670 30882
rect 24722 30830 24734 30882
rect 35970 30830 35982 30882
rect 36034 30830 36046 30882
rect 37090 30830 37102 30882
rect 37154 30830 37166 30882
rect 2494 30818 2546 30830
rect 8542 30818 8594 30830
rect 20862 30818 20914 30830
rect 36542 30818 36594 30830
rect 39118 30818 39170 30830
rect 39566 30882 39618 30894
rect 41570 30830 41582 30882
rect 41634 30830 41646 30882
rect 39566 30818 39618 30830
rect 8318 30770 8370 30782
rect 8318 30706 8370 30718
rect 13022 30770 13074 30782
rect 13022 30706 13074 30718
rect 15822 30770 15874 30782
rect 24334 30770 24386 30782
rect 22306 30718 22318 30770
rect 22370 30718 22382 30770
rect 15822 30706 15874 30718
rect 24334 30706 24386 30718
rect 32398 30770 32450 30782
rect 32398 30706 32450 30718
rect 47854 30770 47906 30782
rect 47854 30706 47906 30718
rect 1344 30602 48608 30636
rect 1344 30550 4478 30602
rect 4530 30550 4582 30602
rect 4634 30550 4686 30602
rect 4738 30550 35198 30602
rect 35250 30550 35302 30602
rect 35354 30550 35406 30602
rect 35458 30550 48608 30602
rect 1344 30516 48608 30550
rect 9550 30434 9602 30446
rect 9550 30370 9602 30382
rect 22206 30434 22258 30446
rect 22206 30370 22258 30382
rect 7198 30322 7250 30334
rect 2482 30270 2494 30322
rect 2546 30270 2558 30322
rect 4610 30270 4622 30322
rect 4674 30270 4686 30322
rect 7198 30258 7250 30270
rect 9214 30322 9266 30334
rect 27022 30322 27074 30334
rect 10546 30270 10558 30322
rect 10610 30270 10622 30322
rect 11106 30270 11118 30322
rect 11170 30270 11182 30322
rect 12674 30270 12686 30322
rect 12738 30270 12750 30322
rect 13906 30270 13918 30322
rect 13970 30270 13982 30322
rect 18946 30270 18958 30322
rect 19010 30270 19022 30322
rect 9214 30258 9266 30270
rect 27022 30258 27074 30270
rect 29038 30322 29090 30334
rect 29038 30258 29090 30270
rect 33630 30322 33682 30334
rect 33630 30258 33682 30270
rect 34862 30322 34914 30334
rect 40798 30322 40850 30334
rect 35746 30270 35758 30322
rect 35810 30270 35822 30322
rect 37538 30270 37550 30322
rect 37602 30270 37614 30322
rect 39666 30270 39678 30322
rect 39730 30270 39742 30322
rect 34862 30258 34914 30270
rect 40798 30258 40850 30270
rect 5182 30210 5234 30222
rect 1810 30158 1822 30210
rect 1874 30158 1886 30210
rect 5182 30146 5234 30158
rect 7646 30210 7698 30222
rect 12014 30210 12066 30222
rect 15486 30210 15538 30222
rect 20414 30210 20466 30222
rect 30494 30210 30546 30222
rect 11442 30158 11454 30210
rect 11506 30158 11518 30210
rect 12562 30158 12574 30210
rect 12626 30158 12638 30210
rect 13682 30158 13694 30210
rect 13746 30158 13758 30210
rect 14578 30158 14590 30210
rect 14642 30158 14654 30210
rect 16034 30158 16046 30210
rect 16098 30158 16110 30210
rect 19618 30158 19630 30210
rect 19682 30158 19694 30210
rect 20738 30158 20750 30210
rect 20802 30158 20814 30210
rect 21410 30158 21422 30210
rect 21474 30158 21486 30210
rect 21858 30158 21870 30210
rect 21922 30158 21934 30210
rect 22306 30158 22318 30210
rect 22370 30158 22382 30210
rect 22978 30158 22990 30210
rect 23042 30158 23054 30210
rect 23538 30158 23550 30210
rect 23602 30158 23614 30210
rect 24770 30158 24782 30210
rect 24834 30158 24846 30210
rect 26674 30158 26686 30210
rect 26738 30158 26750 30210
rect 28578 30158 28590 30210
rect 28642 30158 28654 30210
rect 30146 30158 30158 30210
rect 30210 30158 30222 30210
rect 7646 30146 7698 30158
rect 12014 30146 12066 30158
rect 15486 30146 15538 30158
rect 20414 30146 20466 30158
rect 30494 30146 30546 30158
rect 31502 30210 31554 30222
rect 32398 30210 32450 30222
rect 41022 30210 41074 30222
rect 42702 30210 42754 30222
rect 31938 30158 31950 30210
rect 32002 30158 32014 30210
rect 32834 30158 32846 30210
rect 32898 30158 32910 30210
rect 35522 30158 35534 30210
rect 35586 30158 35598 30210
rect 40450 30158 40462 30210
rect 40514 30158 40526 30210
rect 42242 30158 42254 30210
rect 42306 30158 42318 30210
rect 31502 30146 31554 30158
rect 32398 30146 32450 30158
rect 41022 30146 41074 30158
rect 42702 30146 42754 30158
rect 43822 30210 43874 30222
rect 43822 30146 43874 30158
rect 47070 30210 47122 30222
rect 47070 30146 47122 30158
rect 47406 30210 47458 30222
rect 47406 30146 47458 30158
rect 7310 30098 7362 30110
rect 14926 30098 14978 30110
rect 20078 30098 20130 30110
rect 34526 30098 34578 30110
rect 8418 30046 8430 30098
rect 8482 30046 8494 30098
rect 8978 30046 8990 30098
rect 9042 30046 9054 30098
rect 14242 30046 14254 30098
rect 14306 30046 14318 30098
rect 16818 30046 16830 30098
rect 16882 30046 16894 30098
rect 23650 30046 23662 30098
rect 23714 30046 23726 30098
rect 25106 30046 25118 30098
rect 25170 30046 25182 30098
rect 28466 30046 28478 30098
rect 28530 30046 28542 30098
rect 29474 30046 29486 30098
rect 29538 30046 29550 30098
rect 29922 30046 29934 30098
rect 29986 30046 29998 30098
rect 7310 30034 7362 30046
rect 14926 30034 14978 30046
rect 20078 30034 20130 30046
rect 34526 30034 34578 30046
rect 46734 30098 46786 30110
rect 46734 30034 46786 30046
rect 7086 29986 7138 29998
rect 7086 29922 7138 29934
rect 7758 29986 7810 29998
rect 7758 29922 7810 29934
rect 7982 29986 8034 29998
rect 30942 29986 30994 29998
rect 23090 29934 23102 29986
rect 23154 29934 23166 29986
rect 7982 29922 8034 29934
rect 30942 29922 30994 29934
rect 31054 29986 31106 29998
rect 31054 29922 31106 29934
rect 31166 29986 31218 29998
rect 31166 29922 31218 29934
rect 33518 29986 33570 29998
rect 33518 29922 33570 29934
rect 33742 29986 33794 29998
rect 33742 29922 33794 29934
rect 33966 29986 34018 29998
rect 33966 29922 34018 29934
rect 36430 29986 36482 29998
rect 42030 29986 42082 29998
rect 41346 29934 41358 29986
rect 41410 29934 41422 29986
rect 36430 29922 36482 29934
rect 42030 29922 42082 29934
rect 43038 29986 43090 29998
rect 43038 29922 43090 29934
rect 43486 29986 43538 29998
rect 43486 29922 43538 29934
rect 43710 29986 43762 29998
rect 43710 29922 43762 29934
rect 47182 29986 47234 29998
rect 47182 29922 47234 29934
rect 1344 29818 48608 29852
rect 1344 29766 19838 29818
rect 19890 29766 19942 29818
rect 19994 29766 20046 29818
rect 20098 29766 48608 29818
rect 1344 29732 48608 29766
rect 1710 29650 1762 29662
rect 1710 29586 1762 29598
rect 8766 29650 8818 29662
rect 8766 29586 8818 29598
rect 14590 29650 14642 29662
rect 14590 29586 14642 29598
rect 16830 29650 16882 29662
rect 16830 29586 16882 29598
rect 17502 29650 17554 29662
rect 17502 29586 17554 29598
rect 18734 29650 18786 29662
rect 18734 29586 18786 29598
rect 20750 29650 20802 29662
rect 20750 29586 20802 29598
rect 24558 29650 24610 29662
rect 24558 29586 24610 29598
rect 26686 29650 26738 29662
rect 26686 29586 26738 29598
rect 33182 29650 33234 29662
rect 36082 29598 36094 29650
rect 36146 29598 36158 29650
rect 33182 29586 33234 29598
rect 9662 29538 9714 29550
rect 7746 29486 7758 29538
rect 7810 29486 7822 29538
rect 9662 29474 9714 29486
rect 10110 29538 10162 29550
rect 10110 29474 10162 29486
rect 11566 29538 11618 29550
rect 11566 29474 11618 29486
rect 12798 29538 12850 29550
rect 12798 29474 12850 29486
rect 13694 29538 13746 29550
rect 13694 29474 13746 29486
rect 18846 29538 18898 29550
rect 18846 29474 18898 29486
rect 19742 29538 19794 29550
rect 19742 29474 19794 29486
rect 24110 29538 24162 29550
rect 24110 29474 24162 29486
rect 25790 29538 25842 29550
rect 25790 29474 25842 29486
rect 29710 29538 29762 29550
rect 31278 29538 31330 29550
rect 30370 29486 30382 29538
rect 30434 29486 30446 29538
rect 30594 29486 30606 29538
rect 30658 29486 30670 29538
rect 29710 29474 29762 29486
rect 31278 29474 31330 29486
rect 33630 29538 33682 29550
rect 33630 29474 33682 29486
rect 35086 29538 35138 29550
rect 35086 29474 35138 29486
rect 42814 29538 42866 29550
rect 42814 29474 42866 29486
rect 43150 29538 43202 29550
rect 45602 29486 45614 29538
rect 45666 29486 45678 29538
rect 43150 29474 43202 29486
rect 6302 29426 6354 29438
rect 5506 29374 5518 29426
rect 5570 29374 5582 29426
rect 6302 29362 6354 29374
rect 6862 29426 6914 29438
rect 9774 29426 9826 29438
rect 12014 29426 12066 29438
rect 16046 29426 16098 29438
rect 18398 29426 18450 29438
rect 7970 29374 7982 29426
rect 8034 29374 8046 29426
rect 11106 29374 11118 29426
rect 11170 29374 11182 29426
rect 12562 29374 12574 29426
rect 12626 29374 12638 29426
rect 14690 29374 14702 29426
rect 14754 29374 14766 29426
rect 17378 29374 17390 29426
rect 17442 29374 17454 29426
rect 6862 29362 6914 29374
rect 9774 29362 9826 29374
rect 12014 29362 12066 29374
rect 16046 29362 16098 29374
rect 18398 29362 18450 29374
rect 18622 29426 18674 29438
rect 20974 29426 21026 29438
rect 27022 29426 27074 29438
rect 29934 29426 29986 29438
rect 19170 29374 19182 29426
rect 19234 29374 19246 29426
rect 24658 29374 24670 29426
rect 24722 29374 24734 29426
rect 26786 29374 26798 29426
rect 26850 29374 26862 29426
rect 28578 29374 28590 29426
rect 28642 29374 28654 29426
rect 29138 29374 29150 29426
rect 29202 29374 29214 29426
rect 18622 29362 18674 29374
rect 20974 29362 21026 29374
rect 27022 29362 27074 29374
rect 29934 29362 29986 29374
rect 31614 29426 31666 29438
rect 31614 29362 31666 29374
rect 32510 29426 32562 29438
rect 32510 29362 32562 29374
rect 32958 29426 33010 29438
rect 32958 29362 33010 29374
rect 33294 29426 33346 29438
rect 34526 29426 34578 29438
rect 36766 29426 36818 29438
rect 43262 29426 43314 29438
rect 34066 29374 34078 29426
rect 34130 29374 34142 29426
rect 35410 29374 35422 29426
rect 35474 29374 35486 29426
rect 35858 29374 35870 29426
rect 35922 29374 35934 29426
rect 37090 29374 37102 29426
rect 37154 29374 37166 29426
rect 38098 29374 38110 29426
rect 38162 29374 38174 29426
rect 44818 29374 44830 29426
rect 44882 29374 44894 29426
rect 33294 29362 33346 29374
rect 34526 29362 34578 29374
rect 36766 29362 36818 29374
rect 43262 29362 43314 29374
rect 2270 29314 2322 29326
rect 2270 29250 2322 29262
rect 5966 29314 6018 29326
rect 5966 29250 6018 29262
rect 8430 29314 8482 29326
rect 8430 29250 8482 29262
rect 14926 29314 14978 29326
rect 14926 29250 14978 29262
rect 22878 29314 22930 29326
rect 31502 29314 31554 29326
rect 28802 29262 28814 29314
rect 28866 29262 28878 29314
rect 29250 29262 29262 29314
rect 29314 29262 29326 29314
rect 22878 29250 22930 29262
rect 31502 29250 31554 29262
rect 41022 29314 41074 29326
rect 41022 29250 41074 29262
rect 42926 29314 42978 29326
rect 42926 29250 42978 29262
rect 44494 29314 44546 29326
rect 47730 29262 47742 29314
rect 47794 29262 47806 29314
rect 44494 29250 44546 29262
rect 9662 29202 9714 29214
rect 10322 29150 10334 29202
rect 10386 29150 10398 29202
rect 40786 29150 40798 29202
rect 40850 29199 40862 29202
rect 41010 29199 41022 29202
rect 40850 29153 41022 29199
rect 40850 29150 40862 29153
rect 41010 29150 41022 29153
rect 41074 29150 41086 29202
rect 9662 29138 9714 29150
rect 1344 29034 48608 29068
rect 1344 28982 4478 29034
rect 4530 28982 4582 29034
rect 4634 28982 4686 29034
rect 4738 28982 35198 29034
rect 35250 28982 35302 29034
rect 35354 28982 35406 29034
rect 35458 28982 48608 29034
rect 1344 28948 48608 28982
rect 35646 28866 35698 28878
rect 47070 28866 47122 28878
rect 6962 28814 6974 28866
rect 7026 28814 7038 28866
rect 9538 28814 9550 28866
rect 9602 28814 9614 28866
rect 23426 28814 23438 28866
rect 23490 28814 23502 28866
rect 35970 28814 35982 28866
rect 36034 28814 36046 28866
rect 37538 28814 37550 28866
rect 37602 28814 37614 28866
rect 35646 28802 35698 28814
rect 47070 28802 47122 28814
rect 1822 28754 1874 28766
rect 1822 28690 1874 28702
rect 4958 28754 5010 28766
rect 4958 28690 5010 28702
rect 7198 28754 7250 28766
rect 19854 28754 19906 28766
rect 22990 28754 23042 28766
rect 12450 28702 12462 28754
rect 12514 28702 12526 28754
rect 14130 28702 14142 28754
rect 14194 28702 14206 28754
rect 16370 28702 16382 28754
rect 16434 28702 16446 28754
rect 20290 28702 20302 28754
rect 20354 28702 20366 28754
rect 21410 28702 21422 28754
rect 21474 28702 21486 28754
rect 7198 28690 7250 28702
rect 19854 28690 19906 28702
rect 22990 28690 23042 28702
rect 23998 28754 24050 28766
rect 23998 28690 24050 28702
rect 26910 28754 26962 28766
rect 35422 28754 35474 28766
rect 32050 28702 32062 28754
rect 32114 28702 32126 28754
rect 34178 28702 34190 28754
rect 34242 28702 34254 28754
rect 34962 28702 34974 28754
rect 35026 28702 35038 28754
rect 26910 28690 26962 28702
rect 35422 28690 35474 28702
rect 36430 28754 36482 28766
rect 44942 28754 44994 28766
rect 42130 28702 42142 28754
rect 42194 28702 42206 28754
rect 44258 28702 44270 28754
rect 44322 28702 44334 28754
rect 36430 28690 36482 28702
rect 44942 28690 44994 28702
rect 4622 28642 4674 28654
rect 4622 28578 4674 28590
rect 4846 28642 4898 28654
rect 4846 28578 4898 28590
rect 5182 28642 5234 28654
rect 17726 28642 17778 28654
rect 5954 28590 5966 28642
rect 6018 28590 6030 28642
rect 6738 28590 6750 28642
rect 6802 28590 6814 28642
rect 8418 28590 8430 28642
rect 8482 28590 8494 28642
rect 9426 28590 9438 28642
rect 9490 28590 9502 28642
rect 9762 28590 9774 28642
rect 9826 28590 9838 28642
rect 10434 28590 10446 28642
rect 10498 28590 10510 28642
rect 11218 28590 11230 28642
rect 11282 28590 11294 28642
rect 12898 28590 12910 28642
rect 12962 28590 12974 28642
rect 17042 28590 17054 28642
rect 17106 28590 17118 28642
rect 5182 28578 5234 28590
rect 17726 28578 17778 28590
rect 17950 28642 18002 28654
rect 17950 28578 18002 28590
rect 18174 28642 18226 28654
rect 18174 28578 18226 28590
rect 18958 28642 19010 28654
rect 18958 28578 19010 28590
rect 20750 28642 20802 28654
rect 22430 28642 22482 28654
rect 21746 28590 21758 28642
rect 21810 28590 21822 28642
rect 20750 28578 20802 28590
rect 22430 28578 22482 28590
rect 23774 28642 23826 28654
rect 27022 28642 27074 28654
rect 29486 28642 29538 28654
rect 24434 28590 24446 28642
rect 24498 28590 24510 28642
rect 26002 28590 26014 28642
rect 26066 28590 26078 28642
rect 27794 28590 27806 28642
rect 27858 28590 27870 28642
rect 23774 28578 23826 28590
rect 27022 28578 27074 28590
rect 29486 28578 29538 28590
rect 30606 28642 30658 28654
rect 36990 28642 37042 28654
rect 31378 28590 31390 28642
rect 31442 28590 31454 28642
rect 34626 28590 34638 28642
rect 34690 28590 34702 28642
rect 30606 28578 30658 28590
rect 36990 28578 37042 28590
rect 37214 28642 37266 28654
rect 37214 28578 37266 28590
rect 37886 28642 37938 28654
rect 37886 28578 37938 28590
rect 39006 28642 39058 28654
rect 46398 28642 46450 28654
rect 39218 28590 39230 28642
rect 39282 28590 39294 28642
rect 41346 28590 41358 28642
rect 41410 28590 41422 28642
rect 45714 28590 45726 28642
rect 45778 28590 45790 28642
rect 39006 28578 39058 28590
rect 46398 28578 46450 28590
rect 17502 28530 17554 28542
rect 11330 28478 11342 28530
rect 11394 28478 11406 28530
rect 17502 28466 17554 28478
rect 22878 28530 22930 28542
rect 22878 28466 22930 28478
rect 23102 28530 23154 28542
rect 29150 28530 29202 28542
rect 24322 28478 24334 28530
rect 24386 28478 24398 28530
rect 23102 28466 23154 28478
rect 29150 28466 29202 28478
rect 29822 28530 29874 28542
rect 29822 28466 29874 28478
rect 30158 28530 30210 28542
rect 30158 28466 30210 28478
rect 30942 28530 30994 28542
rect 30942 28466 30994 28478
rect 39902 28530 39954 28542
rect 47070 28530 47122 28542
rect 45938 28478 45950 28530
rect 46002 28478 46014 28530
rect 47630 28530 47682 28542
rect 39902 28466 39954 28478
rect 47070 28466 47122 28478
rect 47182 28474 47234 28486
rect 18398 28418 18450 28430
rect 10434 28366 10446 28418
rect 10498 28366 10510 28418
rect 11442 28366 11454 28418
rect 11506 28366 11518 28418
rect 18398 28354 18450 28366
rect 19294 28418 19346 28430
rect 46510 28418 46562 28430
rect 38210 28366 38222 28418
rect 38274 28366 38286 28418
rect 19294 28354 19346 28366
rect 46510 28354 46562 28366
rect 46734 28418 46786 28430
rect 47630 28466 47682 28478
rect 47742 28530 47794 28542
rect 47742 28466 47794 28478
rect 47182 28410 47234 28422
rect 47406 28418 47458 28430
rect 46734 28354 46786 28366
rect 47406 28354 47458 28366
rect 1344 28250 48608 28284
rect 1344 28198 19838 28250
rect 19890 28198 19942 28250
rect 19994 28198 20046 28250
rect 20098 28198 48608 28250
rect 1344 28164 48608 28198
rect 15038 28082 15090 28094
rect 15038 28018 15090 28030
rect 17390 28082 17442 28094
rect 17390 28018 17442 28030
rect 21982 28082 22034 28094
rect 21982 28018 22034 28030
rect 22206 28082 22258 28094
rect 22766 28082 22818 28094
rect 22418 28030 22430 28082
rect 22482 28030 22494 28082
rect 22206 28018 22258 28030
rect 22766 28018 22818 28030
rect 23662 28082 23714 28094
rect 23662 28018 23714 28030
rect 32958 28082 33010 28094
rect 32958 28018 33010 28030
rect 33070 28082 33122 28094
rect 33070 28018 33122 28030
rect 34078 28082 34130 28094
rect 34078 28018 34130 28030
rect 35646 28082 35698 28094
rect 35646 28018 35698 28030
rect 40910 28082 40962 28094
rect 40910 28018 40962 28030
rect 41918 28082 41970 28094
rect 41918 28018 41970 28030
rect 44606 28082 44658 28094
rect 44606 28018 44658 28030
rect 4510 27970 4562 27982
rect 12910 27970 12962 27982
rect 10658 27918 10670 27970
rect 10722 27918 10734 27970
rect 11218 27918 11230 27970
rect 11282 27918 11294 27970
rect 12002 27918 12014 27970
rect 12066 27918 12078 27970
rect 12226 27918 12238 27970
rect 12290 27918 12302 27970
rect 4510 27906 4562 27918
rect 12910 27906 12962 27918
rect 14030 27970 14082 27982
rect 23326 27970 23378 27982
rect 16818 27918 16830 27970
rect 16882 27918 16894 27970
rect 14030 27906 14082 27918
rect 23326 27906 23378 27918
rect 23438 27970 23490 27982
rect 23438 27906 23490 27918
rect 25566 27970 25618 27982
rect 25566 27906 25618 27918
rect 31838 27970 31890 27982
rect 31838 27906 31890 27918
rect 32174 27970 32226 27982
rect 32174 27906 32226 27918
rect 42142 27970 42194 27982
rect 42142 27906 42194 27918
rect 42814 27970 42866 27982
rect 42814 27906 42866 27918
rect 42926 27970 42978 27982
rect 44930 27918 44942 27970
rect 44994 27918 45006 27970
rect 42926 27906 42978 27918
rect 6414 27858 6466 27870
rect 14926 27858 14978 27870
rect 4274 27806 4286 27858
rect 4338 27806 4350 27858
rect 7186 27806 7198 27858
rect 7250 27806 7262 27858
rect 9762 27806 9774 27858
rect 9826 27806 9838 27858
rect 10098 27806 10110 27858
rect 10162 27806 10174 27858
rect 10882 27806 10894 27858
rect 10946 27806 10958 27858
rect 11778 27806 11790 27858
rect 11842 27806 11854 27858
rect 6414 27794 6466 27806
rect 14926 27794 14978 27806
rect 15262 27858 15314 27870
rect 15262 27794 15314 27806
rect 16494 27858 16546 27870
rect 21870 27858 21922 27870
rect 32510 27858 32562 27870
rect 41134 27858 41186 27870
rect 18610 27806 18622 27858
rect 18674 27806 18686 27858
rect 19394 27806 19406 27858
rect 19458 27806 19470 27858
rect 24322 27806 24334 27858
rect 24386 27806 24398 27858
rect 26114 27806 26126 27858
rect 26178 27806 26190 27858
rect 27346 27806 27358 27858
rect 27410 27806 27422 27858
rect 27794 27806 27806 27858
rect 27858 27806 27870 27858
rect 29698 27806 29710 27858
rect 29762 27806 29774 27858
rect 33282 27806 33294 27858
rect 33346 27806 33358 27858
rect 33506 27806 33518 27858
rect 33570 27806 33582 27858
rect 34738 27806 34750 27858
rect 34802 27806 34814 27858
rect 39106 27806 39118 27858
rect 39170 27806 39182 27858
rect 16494 27794 16546 27806
rect 21870 27794 21922 27806
rect 32510 27794 32562 27806
rect 41134 27794 41186 27806
rect 41582 27858 41634 27870
rect 41582 27794 41634 27806
rect 41694 27858 41746 27870
rect 41694 27794 41746 27806
rect 42254 27858 42306 27870
rect 48066 27806 48078 27858
rect 48130 27806 48142 27858
rect 42254 27794 42306 27806
rect 6302 27746 6354 27758
rect 23886 27746 23938 27758
rect 26910 27746 26962 27758
rect 29374 27746 29426 27758
rect 31278 27746 31330 27758
rect 17826 27694 17838 27746
rect 17890 27694 17902 27746
rect 21522 27694 21534 27746
rect 21586 27694 21598 27746
rect 26226 27694 26238 27746
rect 26290 27694 26302 27746
rect 27906 27694 27918 27746
rect 27970 27694 27982 27746
rect 30370 27694 30382 27746
rect 30434 27694 30446 27746
rect 6302 27682 6354 27694
rect 23886 27682 23938 27694
rect 26910 27682 26962 27694
rect 29374 27682 29426 27694
rect 31278 27682 31330 27694
rect 34414 27746 34466 27758
rect 39566 27746 39618 27758
rect 36194 27694 36206 27746
rect 36258 27694 36270 27746
rect 38322 27694 38334 27746
rect 38386 27694 38398 27746
rect 34414 27682 34466 27694
rect 39566 27682 39618 27694
rect 41022 27746 41074 27758
rect 41022 27682 41074 27694
rect 44270 27746 44322 27758
rect 45266 27694 45278 27746
rect 45330 27694 45342 27746
rect 47394 27694 47406 27746
rect 47458 27694 47470 27746
rect 44270 27682 44322 27694
rect 34750 27634 34802 27646
rect 34750 27570 34802 27582
rect 35086 27634 35138 27646
rect 35086 27570 35138 27582
rect 42814 27634 42866 27646
rect 42814 27570 42866 27582
rect 1344 27466 48608 27500
rect 1344 27414 4478 27466
rect 4530 27414 4582 27466
rect 4634 27414 4686 27466
rect 4738 27414 35198 27466
rect 35250 27414 35302 27466
rect 35354 27414 35406 27466
rect 35458 27414 48608 27466
rect 1344 27380 48608 27414
rect 29710 27298 29762 27310
rect 6402 27246 6414 27298
rect 6466 27246 6478 27298
rect 8978 27246 8990 27298
rect 9042 27246 9054 27298
rect 13794 27246 13806 27298
rect 13858 27246 13870 27298
rect 5070 27186 5122 27198
rect 5070 27122 5122 27134
rect 8654 27186 8706 27198
rect 19170 27190 19182 27242
rect 19234 27190 19246 27242
rect 29710 27234 29762 27246
rect 38222 27298 38274 27310
rect 38222 27234 38274 27246
rect 31278 27186 31330 27198
rect 35870 27186 35922 27198
rect 43598 27186 43650 27198
rect 11106 27134 11118 27186
rect 11170 27134 11182 27186
rect 13906 27134 13918 27186
rect 13970 27134 13982 27186
rect 24322 27134 24334 27186
rect 24386 27134 24398 27186
rect 31714 27134 31726 27186
rect 31778 27134 31790 27186
rect 33282 27134 33294 27186
rect 33346 27134 33358 27186
rect 35410 27134 35422 27186
rect 35474 27134 35486 27186
rect 40226 27134 40238 27186
rect 40290 27134 40302 27186
rect 42354 27134 42366 27186
rect 42418 27134 42430 27186
rect 8654 27122 8706 27134
rect 31278 27122 31330 27134
rect 35870 27122 35922 27134
rect 43598 27122 43650 27134
rect 47294 27186 47346 27198
rect 47294 27122 47346 27134
rect 7086 27074 7138 27086
rect 4610 27022 4622 27074
rect 4674 27022 4686 27074
rect 6738 27022 6750 27074
rect 6802 27022 6814 27074
rect 7086 27010 7138 27022
rect 9774 27074 9826 27086
rect 14478 27074 14530 27086
rect 19518 27074 19570 27086
rect 10546 27022 10558 27074
rect 10610 27022 10622 27074
rect 12114 27022 12126 27074
rect 12178 27022 12190 27074
rect 13682 27022 13694 27074
rect 13746 27022 13758 27074
rect 14690 27022 14702 27074
rect 14754 27022 14766 27074
rect 16258 27022 16270 27074
rect 16322 27022 16334 27074
rect 9774 27010 9826 27022
rect 14478 27010 14530 27022
rect 19518 27010 19570 27022
rect 20190 27074 20242 27086
rect 26798 27074 26850 27086
rect 30718 27074 30770 27086
rect 36990 27074 37042 27086
rect 21410 27022 21422 27074
rect 21474 27022 21486 27074
rect 26562 27022 26574 27074
rect 26626 27022 26638 27074
rect 28130 27022 28142 27074
rect 28194 27022 28206 27074
rect 29138 27022 29150 27074
rect 29202 27022 29214 27074
rect 32610 27022 32622 27074
rect 32674 27022 32686 27074
rect 20190 27010 20242 27022
rect 26798 27010 26850 27022
rect 30718 27010 30770 27022
rect 36990 27010 37042 27022
rect 37102 27074 37154 27086
rect 37102 27010 37154 27022
rect 37886 27074 37938 27086
rect 44830 27074 44882 27086
rect 39554 27022 39566 27074
rect 39618 27022 39630 27074
rect 37886 27010 37938 27022
rect 44830 27010 44882 27022
rect 46286 27074 46338 27086
rect 46286 27010 46338 27022
rect 47070 27074 47122 27086
rect 47070 27010 47122 27022
rect 47518 27074 47570 27086
rect 47518 27010 47570 27022
rect 9326 26962 9378 26974
rect 9326 26898 9378 26910
rect 9550 26962 9602 26974
rect 12910 26962 12962 26974
rect 12450 26910 12462 26962
rect 12514 26910 12526 26962
rect 9550 26898 9602 26910
rect 12910 26898 12962 26910
rect 15486 26962 15538 26974
rect 15486 26898 15538 26910
rect 15598 26962 15650 26974
rect 15598 26898 15650 26910
rect 15822 26962 15874 26974
rect 26014 26962 26066 26974
rect 32174 26962 32226 26974
rect 17042 26910 17054 26962
rect 17106 26910 17118 26962
rect 19842 26910 19854 26962
rect 19906 26910 19918 26962
rect 20514 26910 20526 26962
rect 20578 26910 20590 26962
rect 22082 26910 22094 26962
rect 22146 26910 22158 26962
rect 27906 26910 27918 26962
rect 27970 26910 27982 26962
rect 15822 26898 15874 26910
rect 26014 26898 26066 26910
rect 32174 26898 32226 26910
rect 38110 26962 38162 26974
rect 38110 26898 38162 26910
rect 42926 26962 42978 26974
rect 42926 26898 42978 26910
rect 46398 26962 46450 26974
rect 46398 26898 46450 26910
rect 46846 26962 46898 26974
rect 46846 26898 46898 26910
rect 47854 26962 47906 26974
rect 47854 26898 47906 26910
rect 48190 26962 48242 26974
rect 48190 26898 48242 26910
rect 25118 26850 25170 26862
rect 25118 26786 25170 26798
rect 35758 26850 35810 26862
rect 35758 26786 35810 26798
rect 35982 26850 36034 26862
rect 35982 26786 36034 26798
rect 36206 26850 36258 26862
rect 36206 26786 36258 26798
rect 37214 26850 37266 26862
rect 37214 26786 37266 26798
rect 37438 26850 37490 26862
rect 37438 26786 37490 26798
rect 43038 26850 43090 26862
rect 43038 26786 43090 26798
rect 43262 26850 43314 26862
rect 46622 26850 46674 26862
rect 45154 26798 45166 26850
rect 45218 26798 45230 26850
rect 43262 26786 43314 26798
rect 46622 26786 46674 26798
rect 1344 26682 48608 26716
rect 1344 26630 19838 26682
rect 19890 26630 19942 26682
rect 19994 26630 20046 26682
rect 20098 26630 48608 26682
rect 1344 26596 48608 26630
rect 8094 26514 8146 26526
rect 8094 26450 8146 26462
rect 9102 26514 9154 26526
rect 9102 26450 9154 26462
rect 10110 26514 10162 26526
rect 10110 26450 10162 26462
rect 10894 26514 10946 26526
rect 10894 26450 10946 26462
rect 15598 26514 15650 26526
rect 15598 26450 15650 26462
rect 15822 26514 15874 26526
rect 18286 26514 18338 26526
rect 17938 26462 17950 26514
rect 18002 26462 18014 26514
rect 15822 26450 15874 26462
rect 18286 26450 18338 26462
rect 19070 26514 19122 26526
rect 19070 26450 19122 26462
rect 19518 26514 19570 26526
rect 19518 26450 19570 26462
rect 20302 26514 20354 26526
rect 23886 26514 23938 26526
rect 23538 26462 23550 26514
rect 23602 26462 23614 26514
rect 20302 26450 20354 26462
rect 23886 26450 23938 26462
rect 26014 26514 26066 26526
rect 26014 26450 26066 26462
rect 27470 26514 27522 26526
rect 33070 26514 33122 26526
rect 28466 26462 28478 26514
rect 28530 26462 28542 26514
rect 27470 26450 27522 26462
rect 33070 26450 33122 26462
rect 34862 26514 34914 26526
rect 37102 26514 37154 26526
rect 35186 26462 35198 26514
rect 35250 26462 35262 26514
rect 34862 26450 34914 26462
rect 37102 26450 37154 26462
rect 37998 26514 38050 26526
rect 37998 26450 38050 26462
rect 39118 26514 39170 26526
rect 45614 26514 45666 26526
rect 42354 26462 42366 26514
rect 42418 26462 42430 26514
rect 39118 26450 39170 26462
rect 45614 26450 45666 26462
rect 48302 26514 48354 26526
rect 48302 26450 48354 26462
rect 7198 26402 7250 26414
rect 7198 26338 7250 26350
rect 8990 26402 9042 26414
rect 8990 26338 9042 26350
rect 18622 26402 18674 26414
rect 18622 26338 18674 26350
rect 18958 26402 19010 26414
rect 18958 26338 19010 26350
rect 20190 26402 20242 26414
rect 20190 26338 20242 26350
rect 20862 26402 20914 26414
rect 32510 26402 32562 26414
rect 25554 26350 25566 26402
rect 25618 26350 25630 26402
rect 20862 26338 20914 26350
rect 32510 26338 32562 26350
rect 39342 26402 39394 26414
rect 39342 26338 39394 26350
rect 41022 26402 41074 26414
rect 43374 26402 43426 26414
rect 41234 26350 41246 26402
rect 41298 26350 41310 26402
rect 41022 26338 41074 26350
rect 43374 26338 43426 26350
rect 43710 26402 43762 26414
rect 45266 26350 45278 26402
rect 45330 26350 45342 26402
rect 43710 26338 43762 26350
rect 8430 26290 8482 26302
rect 9550 26290 9602 26302
rect 15150 26290 15202 26302
rect 8194 26238 8206 26290
rect 8258 26238 8270 26290
rect 8754 26238 8766 26290
rect 8818 26238 8830 26290
rect 14690 26238 14702 26290
rect 14754 26238 14766 26290
rect 8430 26226 8482 26238
rect 9550 26226 9602 26238
rect 15150 26226 15202 26238
rect 15710 26290 15762 26302
rect 19630 26290 19682 26302
rect 16594 26238 16606 26290
rect 16658 26238 16670 26290
rect 17378 26238 17390 26290
rect 17442 26238 17454 26290
rect 15710 26226 15762 26238
rect 19630 26226 19682 26238
rect 20974 26290 21026 26302
rect 27022 26290 27074 26302
rect 28142 26290 28194 26302
rect 35758 26290 35810 26302
rect 25330 26238 25342 26290
rect 25394 26238 25406 26290
rect 27346 26238 27358 26290
rect 27410 26238 27422 26290
rect 29250 26238 29262 26290
rect 29314 26238 29326 26290
rect 20974 26226 21026 26238
rect 27022 26226 27074 26238
rect 28142 26226 28194 26238
rect 35758 26226 35810 26238
rect 39454 26290 39506 26302
rect 46622 26290 46674 26302
rect 41794 26238 41806 26290
rect 41858 26238 41870 26290
rect 42578 26238 42590 26290
rect 42642 26238 42654 26290
rect 39454 26226 39506 26238
rect 46622 26226 46674 26238
rect 46958 26290 47010 26302
rect 46958 26226 47010 26238
rect 47182 26290 47234 26302
rect 47182 26226 47234 26238
rect 6414 26178 6466 26190
rect 16158 26178 16210 26190
rect 11666 26126 11678 26178
rect 11730 26126 11742 26178
rect 14018 26126 14030 26178
rect 14082 26126 14094 26178
rect 6414 26114 6466 26126
rect 16158 26114 16210 26126
rect 21758 26178 21810 26190
rect 21758 26114 21810 26126
rect 22318 26178 22370 26190
rect 22318 26114 22370 26126
rect 22654 26178 22706 26190
rect 22654 26114 22706 26126
rect 23102 26178 23154 26190
rect 23102 26114 23154 26126
rect 24670 26178 24722 26190
rect 24670 26114 24722 26126
rect 27918 26178 27970 26190
rect 34078 26178 34130 26190
rect 29922 26126 29934 26178
rect 29986 26126 29998 26178
rect 32050 26126 32062 26178
rect 32114 26126 32126 26178
rect 33506 26126 33518 26178
rect 33570 26126 33582 26178
rect 27918 26114 27970 26126
rect 34078 26114 34130 26126
rect 36206 26178 36258 26190
rect 36206 26114 36258 26126
rect 36654 26178 36706 26190
rect 36654 26114 36706 26126
rect 37550 26178 37602 26190
rect 37550 26114 37602 26126
rect 41134 26178 41186 26190
rect 41134 26114 41186 26126
rect 46846 26178 46898 26190
rect 46846 26114 46898 26126
rect 19518 26066 19570 26078
rect 19518 26002 19570 26014
rect 20302 26066 20354 26078
rect 20302 26002 20354 26014
rect 20862 26066 20914 26078
rect 32398 26066 32450 26078
rect 21746 26014 21758 26066
rect 21810 26063 21822 26066
rect 23090 26063 23102 26066
rect 21810 26017 23102 26063
rect 21810 26014 21822 26017
rect 23090 26014 23102 26017
rect 23154 26014 23166 26066
rect 20862 26002 20914 26014
rect 32398 26002 32450 26014
rect 35534 26066 35586 26078
rect 36418 26014 36430 26066
rect 36482 26063 36494 26066
rect 37538 26063 37550 26066
rect 36482 26017 37550 26063
rect 36482 26014 36494 26017
rect 37538 26014 37550 26017
rect 37602 26014 37614 26066
rect 41570 26014 41582 26066
rect 41634 26014 41646 26066
rect 35534 26002 35586 26014
rect 1344 25898 48608 25932
rect 1344 25846 4478 25898
rect 4530 25846 4582 25898
rect 4634 25846 4686 25898
rect 4738 25846 35198 25898
rect 35250 25846 35302 25898
rect 35354 25846 35406 25898
rect 35458 25846 48608 25898
rect 1344 25812 48608 25846
rect 18622 25730 18674 25742
rect 18622 25666 18674 25678
rect 37438 25730 37490 25742
rect 37438 25666 37490 25678
rect 41918 25730 41970 25742
rect 41918 25666 41970 25678
rect 42254 25730 42306 25742
rect 42254 25666 42306 25678
rect 28590 25618 28642 25630
rect 34078 25618 34130 25630
rect 10770 25566 10782 25618
rect 10834 25566 10846 25618
rect 18274 25566 18286 25618
rect 18338 25566 18350 25618
rect 19282 25566 19294 25618
rect 19346 25566 19358 25618
rect 21858 25566 21870 25618
rect 21922 25566 21934 25618
rect 23314 25566 23326 25618
rect 23378 25566 23390 25618
rect 26114 25566 26126 25618
rect 26178 25566 26190 25618
rect 27122 25566 27134 25618
rect 27186 25566 27198 25618
rect 27458 25566 27470 25618
rect 27522 25566 27534 25618
rect 28242 25566 28254 25618
rect 28306 25566 28318 25618
rect 29922 25566 29934 25618
rect 29986 25566 29998 25618
rect 33618 25566 33630 25618
rect 33682 25566 33694 25618
rect 34514 25566 34526 25618
rect 34578 25566 34590 25618
rect 38210 25566 38222 25618
rect 38274 25566 38286 25618
rect 40338 25566 40350 25618
rect 40402 25566 40414 25618
rect 46050 25566 46062 25618
rect 46114 25566 46126 25618
rect 48178 25566 48190 25618
rect 48242 25566 48254 25618
rect 28590 25554 28642 25566
rect 34078 25554 34130 25566
rect 4846 25506 4898 25518
rect 13694 25506 13746 25518
rect 9650 25454 9662 25506
rect 9714 25454 9726 25506
rect 10546 25454 10558 25506
rect 10610 25454 10622 25506
rect 11778 25454 11790 25506
rect 11842 25454 11854 25506
rect 12786 25454 12798 25506
rect 12850 25454 12862 25506
rect 4846 25442 4898 25454
rect 13694 25442 13746 25454
rect 14030 25506 14082 25518
rect 25678 25506 25730 25518
rect 35534 25506 35586 25518
rect 37214 25506 37266 25518
rect 43374 25506 43426 25518
rect 15362 25454 15374 25506
rect 15426 25454 15438 25506
rect 25778 25454 25790 25506
rect 25842 25454 25854 25506
rect 26898 25454 26910 25506
rect 26962 25454 26974 25506
rect 27682 25454 27694 25506
rect 27746 25454 27758 25506
rect 30706 25454 30718 25506
rect 30770 25454 30782 25506
rect 36978 25454 36990 25506
rect 37042 25454 37054 25506
rect 41122 25454 41134 25506
rect 41186 25454 41198 25506
rect 41906 25454 41918 25506
rect 41970 25454 41982 25506
rect 14030 25442 14082 25454
rect 25678 25442 25730 25454
rect 35534 25442 35586 25454
rect 37214 25442 37266 25454
rect 43374 25442 43426 25454
rect 43486 25506 43538 25518
rect 43486 25442 43538 25454
rect 43934 25506 43986 25518
rect 45378 25454 45390 25506
rect 45442 25454 45454 25506
rect 43934 25442 43986 25454
rect 4510 25394 4562 25406
rect 4510 25330 4562 25342
rect 5070 25394 5122 25406
rect 5070 25330 5122 25342
rect 8430 25394 8482 25406
rect 8430 25330 8482 25342
rect 13806 25394 13858 25406
rect 18734 25394 18786 25406
rect 14354 25342 14366 25394
rect 14418 25342 14430 25394
rect 14914 25342 14926 25394
rect 14978 25342 14990 25394
rect 16146 25342 16158 25394
rect 16210 25342 16222 25394
rect 13806 25330 13858 25342
rect 18734 25330 18786 25342
rect 19294 25394 19346 25406
rect 19294 25330 19346 25342
rect 19406 25394 19458 25406
rect 20302 25394 20354 25406
rect 19506 25342 19518 25394
rect 19570 25342 19582 25394
rect 19406 25330 19458 25342
rect 20302 25330 20354 25342
rect 20414 25394 20466 25406
rect 21870 25394 21922 25406
rect 21634 25342 21646 25394
rect 21698 25342 21710 25394
rect 20414 25330 20466 25342
rect 21870 25330 21922 25342
rect 21982 25394 22034 25406
rect 21982 25330 22034 25342
rect 22766 25394 22818 25406
rect 22766 25330 22818 25342
rect 22878 25394 22930 25406
rect 23550 25394 23602 25406
rect 22978 25342 22990 25394
rect 23042 25342 23054 25394
rect 22878 25330 22930 25342
rect 23550 25330 23602 25342
rect 23774 25394 23826 25406
rect 23774 25330 23826 25342
rect 23886 25394 23938 25406
rect 23886 25330 23938 25342
rect 24446 25394 24498 25406
rect 24446 25330 24498 25342
rect 24558 25394 24610 25406
rect 29934 25394 29986 25406
rect 29810 25342 29822 25394
rect 29874 25342 29886 25394
rect 24558 25330 24610 25342
rect 29934 25330 29986 25342
rect 30046 25394 30098 25406
rect 34638 25394 34690 25406
rect 31490 25342 31502 25394
rect 31554 25342 31566 25394
rect 30046 25330 30098 25342
rect 34638 25330 34690 25342
rect 34862 25394 34914 25406
rect 34862 25330 34914 25342
rect 35646 25394 35698 25406
rect 35646 25330 35698 25342
rect 35870 25394 35922 25406
rect 35870 25330 35922 25342
rect 35982 25394 36034 25406
rect 35982 25330 36034 25342
rect 36430 25394 36482 25406
rect 36430 25330 36482 25342
rect 37550 25394 37602 25406
rect 37550 25330 37602 25342
rect 4734 25282 4786 25294
rect 4734 25218 4786 25230
rect 6302 25282 6354 25294
rect 6302 25218 6354 25230
rect 19070 25282 19122 25294
rect 19070 25218 19122 25230
rect 20078 25282 20130 25294
rect 20078 25218 20130 25230
rect 22206 25282 22258 25294
rect 22206 25218 22258 25230
rect 22542 25282 22594 25294
rect 22542 25218 22594 25230
rect 24782 25282 24834 25294
rect 30270 25282 30322 25294
rect 25554 25230 25566 25282
rect 25618 25230 25630 25282
rect 24782 25218 24834 25230
rect 30270 25218 30322 25230
rect 36206 25282 36258 25294
rect 36206 25218 36258 25230
rect 41582 25282 41634 25294
rect 41582 25218 41634 25230
rect 43598 25282 43650 25294
rect 43598 25218 43650 25230
rect 44942 25282 44994 25294
rect 44942 25218 44994 25230
rect 1344 25114 48608 25148
rect 1344 25062 19838 25114
rect 19890 25062 19942 25114
rect 19994 25062 20046 25114
rect 20098 25062 48608 25114
rect 1344 25028 48608 25062
rect 6526 24946 6578 24958
rect 6526 24882 6578 24894
rect 9438 24946 9490 24958
rect 19406 24946 19458 24958
rect 26798 24946 26850 24958
rect 16034 24894 16046 24946
rect 16098 24894 16110 24946
rect 26002 24894 26014 24946
rect 26066 24894 26078 24946
rect 9438 24882 9490 24894
rect 19406 24882 19458 24894
rect 26798 24882 26850 24894
rect 28590 24946 28642 24958
rect 28590 24882 28642 24894
rect 29934 24946 29986 24958
rect 29934 24882 29986 24894
rect 30718 24946 30770 24958
rect 30718 24882 30770 24894
rect 31502 24946 31554 24958
rect 31502 24882 31554 24894
rect 31614 24946 31666 24958
rect 31614 24882 31666 24894
rect 44830 24946 44882 24958
rect 44830 24882 44882 24894
rect 47294 24946 47346 24958
rect 47294 24882 47346 24894
rect 47630 24946 47682 24958
rect 47630 24882 47682 24894
rect 6974 24834 7026 24846
rect 6974 24770 7026 24782
rect 9662 24834 9714 24846
rect 9662 24770 9714 24782
rect 9774 24834 9826 24846
rect 18174 24834 18226 24846
rect 10994 24782 11006 24834
rect 11058 24782 11070 24834
rect 9774 24770 9826 24782
rect 18174 24770 18226 24782
rect 18286 24834 18338 24846
rect 18286 24770 18338 24782
rect 19518 24834 19570 24846
rect 19518 24770 19570 24782
rect 19630 24834 19682 24846
rect 19630 24770 19682 24782
rect 20526 24834 20578 24846
rect 24446 24834 24498 24846
rect 23314 24782 23326 24834
rect 23378 24782 23390 24834
rect 20526 24770 20578 24782
rect 24446 24770 24498 24782
rect 24558 24834 24610 24846
rect 24558 24770 24610 24782
rect 29710 24834 29762 24846
rect 29710 24770 29762 24782
rect 31054 24834 31106 24846
rect 31054 24770 31106 24782
rect 31838 24834 31890 24846
rect 45054 24834 45106 24846
rect 33842 24782 33854 24834
rect 33906 24782 33918 24834
rect 38434 24782 38446 24834
rect 38498 24782 38510 24834
rect 43474 24782 43486 24834
rect 43538 24782 43550 24834
rect 31838 24770 31890 24782
rect 45054 24770 45106 24782
rect 45166 24834 45218 24846
rect 45166 24770 45218 24782
rect 45614 24834 45666 24846
rect 45614 24770 45666 24782
rect 47070 24834 47122 24846
rect 47070 24770 47122 24782
rect 7870 24722 7922 24734
rect 18510 24722 18562 24734
rect 6066 24670 6078 24722
rect 6130 24670 6142 24722
rect 11442 24670 11454 24722
rect 11506 24670 11518 24722
rect 12114 24670 12126 24722
rect 12178 24670 12190 24722
rect 13122 24670 13134 24722
rect 13186 24670 13198 24722
rect 17714 24670 17726 24722
rect 17778 24670 17790 24722
rect 7870 24658 7922 24670
rect 18510 24658 18562 24670
rect 18958 24722 19010 24734
rect 18958 24658 19010 24670
rect 19294 24722 19346 24734
rect 20302 24722 20354 24734
rect 20066 24670 20078 24722
rect 20130 24670 20142 24722
rect 19294 24658 19346 24670
rect 20302 24658 20354 24670
rect 20638 24722 20690 24734
rect 29598 24722 29650 24734
rect 24098 24670 24110 24722
rect 24162 24670 24174 24722
rect 25778 24670 25790 24722
rect 25842 24670 25854 24722
rect 26114 24670 26126 24722
rect 26178 24670 26190 24722
rect 28130 24670 28142 24722
rect 28194 24670 28206 24722
rect 20638 24658 20690 24670
rect 29598 24658 29650 24670
rect 30494 24722 30546 24734
rect 30494 24658 30546 24670
rect 30830 24722 30882 24734
rect 30830 24658 30882 24670
rect 31390 24722 31442 24734
rect 45726 24722 45778 24734
rect 33170 24670 33182 24722
rect 33234 24670 33246 24722
rect 39218 24670 39230 24722
rect 39282 24670 39294 24722
rect 44258 24670 44270 24722
rect 44322 24670 44334 24722
rect 31390 24658 31442 24670
rect 45726 24658 45778 24670
rect 46958 24722 47010 24734
rect 46958 24658 47010 24670
rect 47518 24722 47570 24734
rect 47518 24658 47570 24670
rect 8206 24610 8258 24622
rect 16718 24610 16770 24622
rect 27694 24610 27746 24622
rect 32398 24610 32450 24622
rect 39678 24610 39730 24622
rect 46174 24610 46226 24622
rect 3154 24558 3166 24610
rect 3218 24558 3230 24610
rect 5282 24558 5294 24610
rect 5346 24558 5358 24610
rect 10546 24558 10558 24610
rect 10610 24558 10622 24610
rect 13794 24558 13806 24610
rect 13858 24558 13870 24610
rect 18162 24558 18174 24610
rect 18226 24558 18238 24610
rect 21186 24558 21198 24610
rect 21250 24558 21262 24610
rect 26226 24558 26238 24610
rect 26290 24558 26302 24610
rect 27234 24558 27246 24610
rect 27298 24558 27310 24610
rect 29026 24558 29038 24610
rect 29090 24558 29102 24610
rect 35970 24558 35982 24610
rect 36034 24558 36046 24610
rect 36306 24558 36318 24610
rect 36370 24558 36382 24610
rect 41346 24558 41358 24610
rect 41410 24558 41422 24610
rect 8206 24546 8258 24558
rect 16718 24546 16770 24558
rect 27694 24546 27746 24558
rect 32398 24546 32450 24558
rect 39678 24546 39730 24558
rect 46174 24546 46226 24558
rect 16830 24498 16882 24510
rect 16830 24434 16882 24446
rect 24558 24498 24610 24510
rect 24558 24434 24610 24446
rect 45614 24498 45666 24510
rect 45614 24434 45666 24446
rect 47630 24498 47682 24510
rect 47630 24434 47682 24446
rect 1344 24330 48608 24364
rect 1344 24278 4478 24330
rect 4530 24278 4582 24330
rect 4634 24278 4686 24330
rect 4738 24278 35198 24330
rect 35250 24278 35302 24330
rect 35354 24278 35406 24330
rect 35458 24278 48608 24330
rect 1344 24244 48608 24278
rect 12798 24162 12850 24174
rect 8642 24110 8654 24162
rect 8706 24110 8718 24162
rect 31042 24159 31054 24162
rect 12798 24098 12850 24110
rect 30609 24113 31054 24159
rect 14142 24050 14194 24062
rect 22318 24050 22370 24062
rect 29710 24050 29762 24062
rect 7186 23998 7198 24050
rect 7250 23998 7262 24050
rect 8418 23998 8430 24050
rect 8482 23998 8494 24050
rect 14802 23998 14814 24050
rect 14866 23998 14878 24050
rect 15922 23998 15934 24050
rect 15986 23998 15998 24050
rect 24546 23998 24558 24050
rect 24610 23998 24622 24050
rect 27794 23998 27806 24050
rect 27858 23998 27870 24050
rect 14142 23986 14194 23998
rect 22318 23986 22370 23998
rect 29710 23986 29762 23998
rect 12350 23938 12402 23950
rect 7522 23886 7534 23938
rect 7586 23886 7598 23938
rect 8642 23886 8654 23938
rect 8706 23886 8718 23938
rect 10882 23886 10894 23938
rect 10946 23886 10958 23938
rect 12350 23874 12402 23886
rect 12686 23938 12738 23950
rect 21646 23938 21698 23950
rect 29262 23938 29314 23950
rect 18834 23886 18846 23938
rect 18898 23886 18910 23938
rect 19282 23886 19294 23938
rect 19346 23886 19358 23938
rect 20178 23886 20190 23938
rect 20242 23886 20254 23938
rect 22642 23886 22654 23938
rect 22706 23886 22718 23938
rect 24882 23886 24894 23938
rect 24946 23886 24958 23938
rect 12686 23874 12738 23886
rect 21646 23874 21698 23886
rect 29262 23874 29314 23886
rect 30382 23938 30434 23950
rect 30609 23938 30655 24113
rect 31042 24110 31054 24113
rect 31106 24110 31118 24162
rect 35086 24050 35138 24062
rect 35086 23986 35138 23998
rect 35982 24050 36034 24062
rect 40674 23998 40686 24050
rect 40738 23998 40750 24050
rect 44818 23998 44830 24050
rect 44882 23998 44894 24050
rect 35982 23986 36034 23998
rect 31614 23938 31666 23950
rect 34974 23938 35026 23950
rect 30594 23886 30606 23938
rect 30658 23886 30670 23938
rect 34626 23886 34638 23938
rect 34690 23886 34702 23938
rect 30382 23874 30434 23886
rect 31614 23874 31666 23886
rect 34974 23874 35026 23886
rect 35758 23938 35810 23950
rect 35758 23874 35810 23886
rect 36094 23938 36146 23950
rect 36094 23874 36146 23886
rect 36318 23938 36370 23950
rect 37874 23886 37886 23938
rect 37938 23886 37950 23938
rect 47730 23886 47742 23938
rect 47794 23886 47806 23938
rect 36318 23874 36370 23886
rect 6526 23826 6578 23838
rect 12798 23826 12850 23838
rect 13918 23826 13970 23838
rect 11554 23774 11566 23826
rect 11618 23774 11630 23826
rect 12114 23774 12126 23826
rect 12178 23774 12190 23826
rect 13682 23774 13694 23826
rect 13746 23774 13758 23826
rect 6526 23762 6578 23774
rect 12798 23762 12850 23774
rect 13918 23762 13970 23774
rect 14254 23826 14306 23838
rect 14254 23762 14306 23774
rect 14926 23826 14978 23838
rect 19518 23826 19570 23838
rect 23102 23826 23154 23838
rect 15138 23774 15150 23826
rect 15202 23774 15214 23826
rect 18050 23774 18062 23826
rect 18114 23774 18126 23826
rect 21298 23774 21310 23826
rect 21362 23774 21374 23826
rect 14926 23762 14978 23774
rect 19518 23762 19570 23774
rect 23102 23762 23154 23774
rect 23214 23826 23266 23838
rect 23214 23762 23266 23774
rect 23998 23826 24050 23838
rect 23998 23762 24050 23774
rect 24110 23826 24162 23838
rect 31278 23826 31330 23838
rect 24210 23774 24222 23826
rect 24274 23774 24286 23826
rect 25666 23774 25678 23826
rect 25730 23774 25742 23826
rect 28466 23774 28478 23826
rect 28530 23774 28542 23826
rect 24110 23762 24162 23774
rect 31278 23762 31330 23774
rect 32062 23826 32114 23838
rect 32062 23762 32114 23774
rect 35646 23826 35698 23838
rect 38546 23774 38558 23826
rect 38610 23774 38622 23826
rect 46946 23774 46958 23826
rect 47010 23774 47022 23826
rect 35646 23762 35698 23774
rect 5070 23714 5122 23726
rect 5070 23650 5122 23662
rect 5966 23714 6018 23726
rect 14030 23714 14082 23726
rect 12002 23662 12014 23714
rect 12066 23662 12078 23714
rect 5966 23650 6018 23662
rect 14030 23650 14082 23662
rect 14590 23714 14642 23726
rect 14590 23650 14642 23662
rect 14814 23714 14866 23726
rect 20750 23714 20802 23726
rect 19954 23662 19966 23714
rect 20018 23662 20030 23714
rect 14814 23650 14866 23662
rect 20750 23650 20802 23662
rect 23326 23714 23378 23726
rect 23326 23650 23378 23662
rect 23438 23714 23490 23726
rect 23438 23650 23490 23662
rect 23774 23714 23826 23726
rect 23774 23650 23826 23662
rect 28142 23714 28194 23726
rect 28142 23650 28194 23662
rect 29150 23714 29202 23726
rect 30830 23714 30882 23726
rect 30034 23662 30046 23714
rect 30098 23662 30110 23714
rect 29150 23650 29202 23662
rect 30830 23650 30882 23662
rect 37102 23714 37154 23726
rect 37102 23650 37154 23662
rect 41134 23714 41186 23726
rect 41134 23650 41186 23662
rect 44270 23714 44322 23726
rect 44270 23650 44322 23662
rect 1344 23546 48608 23580
rect 1344 23494 19838 23546
rect 19890 23494 19942 23546
rect 19994 23494 20046 23546
rect 20098 23494 48608 23546
rect 1344 23460 48608 23494
rect 18286 23378 18338 23390
rect 10210 23326 10222 23378
rect 10274 23326 10286 23378
rect 18286 23314 18338 23326
rect 18398 23378 18450 23390
rect 22990 23378 23042 23390
rect 19058 23326 19070 23378
rect 19122 23326 19134 23378
rect 21522 23326 21534 23378
rect 21586 23326 21598 23378
rect 22194 23326 22206 23378
rect 22258 23326 22270 23378
rect 18398 23314 18450 23326
rect 22990 23314 23042 23326
rect 23214 23378 23266 23390
rect 23214 23314 23266 23326
rect 27918 23378 27970 23390
rect 27918 23314 27970 23326
rect 39566 23378 39618 23390
rect 39566 23314 39618 23326
rect 44942 23378 44994 23390
rect 44942 23314 44994 23326
rect 45614 23378 45666 23390
rect 45614 23314 45666 23326
rect 11230 23266 11282 23278
rect 18174 23266 18226 23278
rect 12674 23214 12686 23266
rect 12738 23214 12750 23266
rect 11230 23202 11282 23214
rect 18174 23202 18226 23214
rect 44606 23266 44658 23278
rect 44606 23202 44658 23214
rect 44718 23266 44770 23278
rect 44718 23202 44770 23214
rect 45166 23266 45218 23278
rect 45166 23202 45218 23214
rect 45950 23266 46002 23278
rect 45950 23202 46002 23214
rect 46174 23266 46226 23278
rect 46174 23202 46226 23214
rect 46286 23266 46338 23278
rect 46286 23202 46338 23214
rect 46622 23266 46674 23278
rect 46622 23202 46674 23214
rect 48078 23266 48130 23278
rect 48078 23202 48130 23214
rect 12126 23154 12178 23166
rect 19406 23154 19458 23166
rect 6290 23102 6302 23154
rect 6354 23102 6366 23154
rect 7970 23102 7982 23154
rect 8034 23102 8046 23154
rect 8418 23102 8430 23154
rect 8482 23102 8494 23154
rect 12562 23102 12574 23154
rect 12626 23102 12638 23154
rect 13458 23102 13470 23154
rect 13522 23102 13534 23154
rect 13906 23102 13918 23154
rect 13970 23102 13982 23154
rect 16370 23102 16382 23154
rect 16434 23102 16446 23154
rect 17602 23102 17614 23154
rect 17666 23102 17678 23154
rect 17938 23102 17950 23154
rect 18002 23102 18014 23154
rect 12126 23090 12178 23102
rect 19406 23090 19458 23102
rect 19742 23154 19794 23166
rect 21870 23154 21922 23166
rect 21298 23102 21310 23154
rect 21362 23102 21374 23154
rect 19742 23090 19794 23102
rect 21870 23090 21922 23102
rect 23326 23154 23378 23166
rect 45502 23154 45554 23166
rect 28242 23102 28254 23154
rect 28306 23102 28318 23154
rect 40898 23102 40910 23154
rect 40962 23102 40974 23154
rect 23326 23090 23378 23102
rect 45502 23090 45554 23102
rect 45838 23154 45890 23166
rect 45838 23090 45890 23102
rect 46958 23154 47010 23166
rect 46958 23090 47010 23102
rect 47294 23154 47346 23166
rect 47294 23090 47346 23102
rect 47406 23154 47458 23166
rect 47406 23090 47458 23102
rect 47742 23154 47794 23166
rect 47742 23090 47794 23102
rect 8878 23042 8930 23054
rect 3490 22990 3502 23042
rect 3554 22990 3566 23042
rect 5618 22990 5630 23042
rect 5682 22990 5694 23042
rect 8878 22978 8930 22990
rect 10446 23042 10498 23054
rect 20302 23042 20354 23054
rect 15810 22990 15822 23042
rect 15874 22990 15886 23042
rect 10446 22978 10498 22990
rect 20302 22978 20354 22990
rect 20750 23042 20802 23054
rect 20750 22978 20802 22990
rect 22654 23042 22706 23054
rect 22654 22978 22706 22990
rect 23886 23042 23938 23054
rect 23886 22978 23938 22990
rect 24334 23042 24386 23054
rect 24334 22978 24386 22990
rect 25342 23042 25394 23054
rect 31614 23042 31666 23054
rect 29026 22990 29038 23042
rect 29090 22990 29102 23042
rect 31154 22990 31166 23042
rect 31218 22990 31230 23042
rect 25342 22978 25394 22990
rect 31614 22978 31666 22990
rect 36766 23042 36818 23054
rect 36766 22978 36818 22990
rect 39118 23042 39170 23054
rect 39118 22978 39170 22990
rect 40462 23042 40514 23054
rect 44270 23042 44322 23054
rect 41682 22990 41694 23042
rect 41746 22990 41758 23042
rect 43810 22990 43822 23042
rect 43874 22990 43886 23042
rect 40462 22978 40514 22990
rect 44270 22978 44322 22990
rect 47070 23042 47122 23054
rect 47070 22978 47122 22990
rect 47630 23042 47682 23054
rect 47630 22978 47682 22990
rect 7422 22930 7474 22942
rect 7422 22866 7474 22878
rect 19854 22930 19906 22942
rect 19854 22866 19906 22878
rect 1344 22762 48608 22796
rect 1344 22710 4478 22762
rect 4530 22710 4582 22762
rect 4634 22710 4686 22762
rect 4738 22710 35198 22762
rect 35250 22710 35302 22762
rect 35354 22710 35406 22762
rect 35458 22710 48608 22762
rect 1344 22676 48608 22710
rect 35198 22594 35250 22606
rect 44706 22542 44718 22594
rect 44770 22591 44782 22594
rect 45042 22591 45054 22594
rect 44770 22545 45054 22591
rect 44770 22542 44782 22545
rect 45042 22542 45054 22545
rect 45106 22542 45118 22594
rect 35198 22530 35250 22542
rect 7086 22482 7138 22494
rect 4722 22430 4734 22482
rect 4786 22430 4798 22482
rect 6066 22430 6078 22482
rect 6130 22430 6142 22482
rect 7086 22418 7138 22430
rect 7198 22482 7250 22494
rect 7198 22418 7250 22430
rect 11118 22482 11170 22494
rect 21422 22482 21474 22494
rect 16370 22430 16382 22482
rect 16434 22430 16446 22482
rect 16930 22430 16942 22482
rect 16994 22430 17006 22482
rect 11118 22418 11170 22430
rect 21422 22418 21474 22430
rect 22430 22482 22482 22494
rect 29486 22482 29538 22494
rect 36318 22482 36370 22494
rect 40910 22482 40962 22494
rect 23650 22430 23662 22482
rect 23714 22430 23726 22482
rect 25778 22430 25790 22482
rect 25842 22430 25854 22482
rect 28466 22430 28478 22482
rect 28530 22430 28542 22482
rect 34178 22430 34190 22482
rect 34242 22430 34254 22482
rect 40450 22430 40462 22482
rect 40514 22430 40526 22482
rect 22430 22418 22482 22430
rect 29486 22418 29538 22430
rect 36318 22418 36370 22430
rect 40910 22418 40962 22430
rect 43150 22482 43202 22494
rect 45266 22430 45278 22482
rect 45330 22430 45342 22482
rect 47394 22430 47406 22482
rect 47458 22430 47470 22482
rect 43150 22418 43202 22430
rect 12686 22370 12738 22382
rect 17614 22370 17666 22382
rect 4946 22318 4958 22370
rect 5010 22318 5022 22370
rect 5842 22318 5854 22370
rect 5906 22318 5918 22370
rect 8978 22318 8990 22370
rect 9042 22318 9054 22370
rect 9314 22318 9326 22370
rect 9378 22318 9390 22370
rect 13570 22318 13582 22370
rect 13634 22318 13646 22370
rect 16706 22318 16718 22370
rect 16770 22318 16782 22370
rect 12686 22306 12738 22318
rect 17614 22306 17666 22318
rect 18174 22370 18226 22382
rect 19630 22370 19682 22382
rect 18610 22318 18622 22370
rect 18674 22318 18686 22370
rect 18174 22306 18226 22318
rect 19630 22306 19682 22318
rect 19966 22370 20018 22382
rect 19966 22306 20018 22318
rect 20190 22370 20242 22382
rect 27022 22370 27074 22382
rect 22978 22318 22990 22370
rect 23042 22318 23054 22370
rect 20190 22306 20242 22318
rect 27022 22306 27074 22318
rect 27582 22370 27634 22382
rect 27582 22306 27634 22318
rect 28030 22370 28082 22382
rect 28030 22306 28082 22318
rect 30382 22370 30434 22382
rect 30382 22306 30434 22318
rect 30606 22370 30658 22382
rect 30606 22306 30658 22318
rect 31726 22370 31778 22382
rect 31726 22306 31778 22318
rect 32286 22370 32338 22382
rect 32286 22306 32338 22318
rect 32622 22370 32674 22382
rect 34862 22370 34914 22382
rect 33842 22318 33854 22370
rect 33906 22318 33918 22370
rect 34626 22318 34638 22370
rect 34690 22318 34702 22370
rect 32622 22306 32674 22318
rect 34862 22306 34914 22318
rect 35086 22370 35138 22382
rect 42254 22370 42306 22382
rect 37538 22318 37550 22370
rect 37602 22318 37614 22370
rect 48178 22318 48190 22370
rect 48242 22318 48254 22370
rect 35086 22306 35138 22318
rect 42254 22306 42306 22318
rect 7982 22258 8034 22270
rect 7982 22194 8034 22206
rect 10334 22258 10386 22270
rect 10334 22194 10386 22206
rect 12350 22258 12402 22270
rect 12350 22194 12402 22206
rect 12798 22258 12850 22270
rect 20526 22258 20578 22270
rect 14242 22206 14254 22258
rect 14306 22206 14318 22258
rect 18498 22206 18510 22258
rect 18562 22206 18574 22258
rect 19170 22206 19182 22258
rect 19234 22206 19246 22258
rect 12798 22194 12850 22206
rect 20526 22194 20578 22206
rect 27694 22258 27746 22270
rect 27694 22194 27746 22206
rect 29374 22258 29426 22270
rect 29374 22194 29426 22206
rect 29710 22258 29762 22270
rect 29710 22194 29762 22206
rect 29934 22258 29986 22270
rect 42478 22258 42530 22270
rect 35522 22206 35534 22258
rect 35586 22206 35598 22258
rect 38322 22206 38334 22258
rect 38386 22206 38398 22258
rect 29934 22194 29986 22206
rect 42478 22194 42530 22206
rect 43598 22258 43650 22270
rect 43598 22194 43650 22206
rect 9438 22146 9490 22158
rect 9438 22082 9490 22094
rect 13022 22146 13074 22158
rect 13022 22082 13074 22094
rect 19854 22146 19906 22158
rect 19854 22082 19906 22094
rect 20414 22146 20466 22158
rect 20414 22082 20466 22094
rect 21982 22146 22034 22158
rect 21982 22082 22034 22094
rect 26238 22146 26290 22158
rect 26238 22082 26290 22094
rect 27134 22146 27186 22158
rect 27134 22082 27186 22094
rect 27358 22146 27410 22158
rect 27358 22082 27410 22094
rect 30494 22146 30546 22158
rect 30494 22082 30546 22094
rect 30830 22146 30882 22158
rect 30830 22082 30882 22094
rect 31390 22146 31442 22158
rect 33406 22146 33458 22158
rect 32946 22094 32958 22146
rect 33010 22094 33022 22146
rect 31390 22082 31442 22094
rect 33406 22082 33458 22094
rect 35870 22146 35922 22158
rect 35870 22082 35922 22094
rect 37102 22146 37154 22158
rect 37102 22082 37154 22094
rect 41582 22146 41634 22158
rect 41582 22082 41634 22094
rect 41694 22146 41746 22158
rect 41694 22082 41746 22094
rect 41806 22146 41858 22158
rect 41806 22082 41858 22094
rect 42590 22146 42642 22158
rect 42590 22082 42642 22094
rect 42814 22146 42866 22158
rect 42814 22082 42866 22094
rect 43486 22146 43538 22158
rect 43486 22082 43538 22094
rect 44158 22146 44210 22158
rect 44158 22082 44210 22094
rect 44942 22146 44994 22158
rect 44942 22082 44994 22094
rect 1344 21978 48608 22012
rect 1344 21926 19838 21978
rect 19890 21926 19942 21978
rect 19994 21926 20046 21978
rect 20098 21926 48608 21978
rect 1344 21892 48608 21926
rect 10894 21810 10946 21822
rect 8194 21758 8206 21810
rect 8258 21758 8270 21810
rect 10894 21746 10946 21758
rect 12910 21810 12962 21822
rect 12910 21746 12962 21758
rect 13918 21810 13970 21822
rect 13918 21746 13970 21758
rect 14590 21810 14642 21822
rect 14590 21746 14642 21758
rect 15150 21810 15202 21822
rect 15934 21810 15986 21822
rect 15586 21758 15598 21810
rect 15650 21758 15662 21810
rect 15150 21746 15202 21758
rect 15934 21746 15986 21758
rect 18286 21810 18338 21822
rect 18286 21746 18338 21758
rect 18734 21810 18786 21822
rect 18734 21746 18786 21758
rect 20078 21810 20130 21822
rect 20078 21746 20130 21758
rect 21310 21810 21362 21822
rect 21310 21746 21362 21758
rect 21646 21810 21698 21822
rect 21646 21746 21698 21758
rect 22206 21810 22258 21822
rect 22206 21746 22258 21758
rect 22878 21810 22930 21822
rect 22878 21746 22930 21758
rect 23438 21810 23490 21822
rect 29150 21810 29202 21822
rect 24322 21758 24334 21810
rect 24386 21758 24398 21810
rect 26338 21758 26350 21810
rect 26402 21758 26414 21810
rect 23438 21746 23490 21758
rect 29150 21746 29202 21758
rect 40350 21810 40402 21822
rect 40350 21746 40402 21758
rect 41134 21810 41186 21822
rect 41134 21746 41186 21758
rect 46622 21810 46674 21822
rect 46622 21746 46674 21758
rect 46846 21810 46898 21822
rect 46846 21746 46898 21758
rect 47182 21810 47234 21822
rect 47182 21746 47234 21758
rect 10782 21698 10834 21710
rect 9538 21646 9550 21698
rect 9602 21646 9614 21698
rect 10658 21646 10670 21698
rect 10722 21646 10734 21698
rect 10782 21634 10834 21646
rect 11678 21698 11730 21710
rect 14142 21698 14194 21710
rect 12562 21646 12574 21698
rect 12626 21646 12638 21698
rect 11678 21634 11730 21646
rect 14142 21634 14194 21646
rect 21086 21698 21138 21710
rect 21086 21634 21138 21646
rect 23102 21698 23154 21710
rect 23102 21634 23154 21646
rect 23886 21698 23938 21710
rect 23886 21634 23938 21646
rect 31054 21698 31106 21710
rect 31054 21634 31106 21646
rect 31390 21698 31442 21710
rect 31390 21634 31442 21646
rect 31614 21698 31666 21710
rect 31614 21634 31666 21646
rect 39566 21698 39618 21710
rect 39566 21634 39618 21646
rect 41470 21698 41522 21710
rect 41470 21634 41522 21646
rect 46510 21698 46562 21710
rect 46510 21634 46562 21646
rect 47070 21698 47122 21710
rect 47070 21634 47122 21646
rect 47854 21698 47906 21710
rect 47854 21634 47906 21646
rect 9886 21586 9938 21598
rect 4834 21534 4846 21586
rect 4898 21534 4910 21586
rect 9886 21522 9938 21534
rect 11118 21586 11170 21598
rect 11118 21522 11170 21534
rect 11454 21586 11506 21598
rect 14702 21586 14754 21598
rect 11890 21534 11902 21586
rect 11954 21534 11966 21586
rect 12226 21534 12238 21586
rect 12290 21534 12302 21586
rect 13346 21534 13358 21586
rect 13410 21534 13422 21586
rect 13682 21534 13694 21586
rect 13746 21534 13758 21586
rect 11454 21522 11506 21534
rect 14702 21522 14754 21534
rect 14926 21586 14978 21598
rect 14926 21522 14978 21534
rect 15262 21586 15314 21598
rect 15262 21522 15314 21534
rect 16270 21586 16322 21598
rect 17950 21586 18002 21598
rect 17714 21534 17726 21586
rect 17778 21534 17790 21586
rect 16270 21522 16322 21534
rect 17950 21522 18002 21534
rect 19966 21586 20018 21598
rect 19966 21522 20018 21534
rect 20190 21586 20242 21598
rect 20190 21522 20242 21534
rect 20974 21586 21026 21598
rect 20974 21522 21026 21534
rect 21758 21586 21810 21598
rect 21758 21522 21810 21534
rect 22766 21586 22818 21598
rect 22766 21522 22818 21534
rect 23662 21586 23714 21598
rect 23662 21522 23714 21534
rect 23998 21586 24050 21598
rect 23998 21522 24050 21534
rect 24670 21586 24722 21598
rect 26686 21586 26738 21598
rect 39342 21586 39394 21598
rect 25330 21534 25342 21586
rect 25394 21534 25406 21586
rect 27346 21534 27358 21586
rect 27410 21534 27422 21586
rect 27570 21534 27582 21586
rect 27634 21534 27646 21586
rect 32050 21534 32062 21586
rect 32114 21534 32126 21586
rect 35186 21534 35198 21586
rect 35250 21534 35262 21586
rect 38546 21534 38558 21586
rect 38610 21534 38622 21586
rect 24670 21522 24722 21534
rect 26686 21522 26738 21534
rect 39342 21522 39394 21534
rect 39790 21586 39842 21598
rect 39790 21522 39842 21534
rect 40014 21586 40066 21598
rect 40014 21522 40066 21534
rect 40798 21586 40850 21598
rect 40798 21522 40850 21534
rect 41134 21586 41186 21598
rect 48190 21586 48242 21598
rect 41906 21534 41918 21586
rect 41970 21534 41982 21586
rect 41134 21522 41186 21534
rect 48190 21522 48242 21534
rect 9102 21474 9154 21486
rect 14030 21474 14082 21486
rect 19294 21474 19346 21486
rect 5506 21422 5518 21474
rect 5570 21422 5582 21474
rect 10322 21422 10334 21474
rect 10386 21422 10398 21474
rect 11778 21422 11790 21474
rect 11842 21422 11854 21474
rect 16706 21422 16718 21474
rect 16770 21422 16782 21474
rect 9102 21410 9154 21422
rect 14030 21410 14082 21422
rect 19294 21410 19346 21422
rect 20414 21474 20466 21486
rect 28702 21474 28754 21486
rect 25666 21422 25678 21474
rect 25730 21422 25742 21474
rect 28018 21422 28030 21474
rect 28082 21422 28094 21474
rect 20414 21410 20466 21422
rect 28702 21410 28754 21422
rect 29598 21474 29650 21486
rect 32286 21474 32338 21486
rect 46286 21474 46338 21486
rect 31266 21422 31278 21474
rect 31330 21422 31342 21474
rect 35970 21422 35982 21474
rect 36034 21422 36046 21474
rect 38098 21422 38110 21474
rect 38162 21422 38174 21474
rect 38882 21422 38894 21474
rect 38946 21422 38958 21474
rect 42578 21422 42590 21474
rect 42642 21422 42654 21474
rect 44706 21422 44718 21474
rect 44770 21422 44782 21474
rect 29598 21410 29650 21422
rect 32286 21410 32338 21422
rect 46286 21410 46338 21422
rect 14590 21362 14642 21374
rect 14590 21298 14642 21310
rect 20638 21362 20690 21374
rect 20638 21298 20690 21310
rect 21646 21362 21698 21374
rect 32398 21362 32450 21374
rect 28130 21310 28142 21362
rect 28194 21310 28206 21362
rect 21646 21298 21698 21310
rect 32398 21298 32450 21310
rect 47182 21362 47234 21374
rect 47182 21298 47234 21310
rect 1344 21194 48608 21228
rect 1344 21142 4478 21194
rect 4530 21142 4582 21194
rect 4634 21142 4686 21194
rect 4738 21142 35198 21194
rect 35250 21142 35302 21194
rect 35354 21142 35406 21194
rect 35458 21142 48608 21194
rect 1344 21108 48608 21142
rect 6862 21026 6914 21038
rect 4946 20974 4958 21026
rect 5010 20974 5022 21026
rect 6862 20962 6914 20974
rect 19966 21026 20018 21038
rect 19966 20962 20018 20974
rect 21422 21026 21474 21038
rect 21422 20962 21474 20974
rect 26462 21026 26514 21038
rect 26462 20962 26514 20974
rect 27134 21026 27186 21038
rect 35758 21026 35810 21038
rect 28018 20974 28030 21026
rect 28082 21023 28094 21026
rect 28690 21023 28702 21026
rect 28082 20977 28702 21023
rect 28082 20974 28094 20977
rect 28690 20974 28702 20977
rect 28754 20974 28766 21026
rect 27134 20962 27186 20974
rect 35758 20962 35810 20974
rect 4846 20914 4898 20926
rect 17950 20914 18002 20926
rect 9650 20862 9662 20914
rect 9714 20862 9726 20914
rect 10658 20862 10670 20914
rect 10722 20862 10734 20914
rect 14130 20862 14142 20914
rect 14194 20862 14206 20914
rect 4846 20850 4898 20862
rect 17950 20850 18002 20862
rect 19406 20914 19458 20926
rect 19406 20850 19458 20862
rect 20526 20914 20578 20926
rect 20526 20850 20578 20862
rect 22542 20914 22594 20926
rect 22542 20850 22594 20862
rect 22654 20914 22706 20926
rect 22654 20850 22706 20862
rect 27358 20914 27410 20926
rect 27358 20850 27410 20862
rect 28030 20914 28082 20926
rect 28030 20850 28082 20862
rect 29822 20914 29874 20926
rect 36094 20914 36146 20926
rect 32274 20862 32286 20914
rect 32338 20862 32350 20914
rect 34402 20862 34414 20914
rect 34466 20862 34478 20914
rect 29822 20850 29874 20862
rect 36094 20850 36146 20862
rect 37662 20914 37714 20926
rect 37662 20850 37714 20862
rect 39342 20914 39394 20926
rect 42814 20914 42866 20926
rect 41906 20862 41918 20914
rect 41970 20862 41982 20914
rect 39342 20850 39394 20862
rect 42814 20850 42866 20862
rect 44942 20914 44994 20926
rect 45266 20862 45278 20914
rect 45330 20862 45342 20914
rect 47394 20862 47406 20914
rect 47458 20862 47470 20914
rect 44942 20850 44994 20862
rect 4734 20802 4786 20814
rect 11902 20802 11954 20814
rect 17726 20802 17778 20814
rect 8754 20750 8766 20802
rect 8818 20750 8830 20802
rect 10994 20750 11006 20802
rect 11058 20750 11070 20802
rect 17042 20750 17054 20802
rect 17106 20750 17118 20802
rect 4734 20738 4786 20750
rect 11902 20738 11954 20750
rect 17726 20738 17778 20750
rect 19630 20802 19682 20814
rect 19630 20738 19682 20750
rect 20190 20802 20242 20814
rect 20190 20738 20242 20750
rect 20414 20802 20466 20814
rect 20414 20738 20466 20750
rect 20638 20802 20690 20814
rect 20638 20738 20690 20750
rect 21534 20802 21586 20814
rect 21534 20738 21586 20750
rect 23998 20802 24050 20814
rect 26126 20802 26178 20814
rect 35982 20802 36034 20814
rect 25106 20750 25118 20802
rect 25170 20750 25182 20802
rect 26898 20750 26910 20802
rect 26962 20750 26974 20802
rect 31490 20750 31502 20802
rect 31554 20750 31566 20802
rect 23998 20738 24050 20750
rect 26126 20738 26178 20750
rect 35982 20738 36034 20750
rect 38222 20802 38274 20814
rect 40002 20750 40014 20802
rect 40066 20750 40078 20802
rect 48066 20750 48078 20802
rect 48130 20750 48142 20802
rect 38222 20738 38274 20750
rect 11566 20690 11618 20702
rect 11566 20626 11618 20638
rect 11678 20690 11730 20702
rect 12574 20690 12626 20702
rect 21422 20690 21474 20702
rect 12450 20638 12462 20690
rect 12514 20638 12526 20690
rect 13458 20638 13470 20690
rect 13522 20638 13534 20690
rect 16258 20638 16270 20690
rect 16322 20638 16334 20690
rect 11678 20626 11730 20638
rect 12574 20626 12626 20638
rect 21422 20626 21474 20638
rect 22094 20690 22146 20702
rect 22094 20626 22146 20638
rect 22206 20690 22258 20702
rect 22206 20626 22258 20638
rect 23438 20690 23490 20702
rect 23438 20626 23490 20638
rect 23886 20690 23938 20702
rect 23886 20626 23938 20638
rect 24334 20690 24386 20702
rect 24334 20626 24386 20638
rect 24446 20690 24498 20702
rect 26574 20690 26626 20702
rect 24882 20638 24894 20690
rect 24946 20638 24958 20690
rect 24446 20626 24498 20638
rect 26574 20626 26626 20638
rect 27470 20690 27522 20702
rect 27470 20626 27522 20638
rect 34862 20690 34914 20702
rect 34862 20626 34914 20638
rect 35310 20690 35362 20702
rect 36206 20690 36258 20702
rect 35522 20638 35534 20690
rect 35586 20638 35598 20690
rect 35310 20626 35362 20638
rect 36206 20626 36258 20638
rect 36990 20690 37042 20702
rect 36990 20626 37042 20638
rect 37102 20690 37154 20702
rect 39006 20690 39058 20702
rect 38546 20638 38558 20690
rect 38610 20638 38622 20690
rect 37102 20626 37154 20638
rect 39006 20626 39058 20638
rect 42702 20690 42754 20702
rect 42702 20626 42754 20638
rect 43038 20690 43090 20702
rect 43934 20690 43986 20702
rect 43138 20638 43150 20690
rect 43202 20638 43214 20690
rect 43038 20626 43090 20638
rect 43934 20626 43986 20638
rect 6302 20578 6354 20590
rect 6302 20514 6354 20526
rect 12686 20578 12738 20590
rect 12686 20514 12738 20526
rect 12798 20578 12850 20590
rect 12798 20514 12850 20526
rect 12910 20578 12962 20590
rect 12910 20514 12962 20526
rect 13806 20578 13858 20590
rect 13806 20514 13858 20526
rect 18286 20578 18338 20590
rect 18286 20514 18338 20526
rect 18958 20578 19010 20590
rect 18958 20514 19010 20526
rect 19070 20578 19122 20590
rect 19070 20514 19122 20526
rect 19182 20578 19234 20590
rect 19182 20514 19234 20526
rect 21870 20578 21922 20590
rect 23662 20578 23714 20590
rect 28366 20578 28418 20590
rect 23090 20526 23102 20578
rect 23154 20526 23166 20578
rect 25778 20526 25790 20578
rect 25842 20526 25854 20578
rect 21870 20514 21922 20526
rect 23662 20514 23714 20526
rect 28366 20514 28418 20526
rect 39230 20578 39282 20590
rect 39230 20514 39282 20526
rect 39454 20578 39506 20590
rect 39454 20514 39506 20526
rect 42926 20578 42978 20590
rect 42926 20514 42978 20526
rect 1344 20410 48608 20444
rect 1344 20358 19838 20410
rect 19890 20358 19942 20410
rect 19994 20358 20046 20410
rect 20098 20358 48608 20410
rect 1344 20324 48608 20358
rect 15822 20242 15874 20254
rect 14466 20190 14478 20242
rect 14530 20190 14542 20242
rect 15822 20178 15874 20190
rect 16830 20242 16882 20254
rect 16830 20178 16882 20190
rect 17614 20242 17666 20254
rect 17614 20178 17666 20190
rect 20414 20242 20466 20254
rect 23326 20242 23378 20254
rect 21298 20190 21310 20242
rect 21362 20190 21374 20242
rect 20414 20178 20466 20190
rect 23326 20178 23378 20190
rect 24782 20242 24834 20254
rect 39566 20242 39618 20254
rect 39106 20190 39118 20242
rect 39170 20190 39182 20242
rect 24782 20178 24834 20190
rect 39566 20178 39618 20190
rect 5406 20130 5458 20142
rect 5406 20066 5458 20078
rect 9662 20130 9714 20142
rect 9662 20066 9714 20078
rect 9774 20130 9826 20142
rect 11902 20130 11954 20142
rect 10434 20078 10446 20130
rect 10498 20078 10510 20130
rect 9774 20066 9826 20078
rect 11902 20066 11954 20078
rect 12014 20130 12066 20142
rect 12014 20066 12066 20078
rect 12462 20130 12514 20142
rect 12462 20066 12514 20078
rect 13246 20130 13298 20142
rect 13246 20066 13298 20078
rect 15262 20130 15314 20142
rect 15262 20066 15314 20078
rect 15374 20130 15426 20142
rect 17390 20130 17442 20142
rect 16482 20078 16494 20130
rect 16546 20078 16558 20130
rect 15374 20066 15426 20078
rect 17390 20066 17442 20078
rect 20526 20130 20578 20142
rect 20526 20066 20578 20078
rect 22094 20130 22146 20142
rect 22094 20066 22146 20078
rect 22318 20130 22370 20142
rect 22318 20066 22370 20078
rect 22654 20130 22706 20142
rect 22654 20066 22706 20078
rect 22766 20130 22818 20142
rect 25566 20130 25618 20142
rect 23874 20078 23886 20130
rect 23938 20078 23950 20130
rect 22766 20066 22818 20078
rect 25566 20066 25618 20078
rect 30718 20130 30770 20142
rect 30718 20066 30770 20078
rect 31166 20130 31218 20142
rect 31166 20066 31218 20078
rect 32174 20130 32226 20142
rect 32174 20066 32226 20078
rect 32510 20130 32562 20142
rect 32510 20066 32562 20078
rect 33742 20130 33794 20142
rect 33742 20066 33794 20078
rect 33966 20130 34018 20142
rect 35086 20130 35138 20142
rect 34738 20078 34750 20130
rect 34802 20078 34814 20130
rect 33966 20066 34018 20078
rect 35086 20066 35138 20078
rect 35646 20130 35698 20142
rect 35646 20066 35698 20078
rect 38782 20130 38834 20142
rect 38782 20066 38834 20078
rect 41806 20130 41858 20142
rect 41806 20066 41858 20078
rect 42254 20130 42306 20142
rect 42254 20066 42306 20078
rect 43262 20130 43314 20142
rect 47854 20130 47906 20142
rect 47506 20078 47518 20130
rect 47570 20078 47582 20130
rect 43262 20066 43314 20078
rect 47854 20066 47906 20078
rect 5070 20018 5122 20030
rect 12126 20018 12178 20030
rect 8642 19966 8654 20018
rect 8706 19966 8718 20018
rect 10658 19966 10670 20018
rect 10722 19966 10734 20018
rect 11442 19966 11454 20018
rect 11506 19966 11518 20018
rect 11666 19966 11678 20018
rect 11730 19966 11742 20018
rect 5070 19954 5122 19966
rect 12126 19954 12178 19966
rect 13582 20018 13634 20030
rect 19182 20018 19234 20030
rect 14690 19966 14702 20018
rect 14754 19966 14766 20018
rect 17826 19966 17838 20018
rect 17890 19966 17902 20018
rect 18050 19966 18062 20018
rect 18114 19966 18126 20018
rect 13582 19954 13634 19966
rect 19182 19954 19234 19966
rect 19966 20018 20018 20030
rect 19966 19954 20018 19966
rect 20190 20018 20242 20030
rect 20190 19954 20242 19966
rect 20638 20018 20690 20030
rect 21982 20018 22034 20030
rect 21522 19966 21534 20018
rect 21586 19966 21598 20018
rect 20638 19954 20690 19966
rect 21982 19954 22034 19966
rect 23550 20018 23602 20030
rect 30158 20018 30210 20030
rect 26898 19966 26910 20018
rect 26962 19966 26974 20018
rect 23550 19954 23602 19966
rect 30158 19954 30210 19966
rect 30382 20018 30434 20030
rect 30382 19954 30434 19966
rect 31054 20018 31106 20030
rect 31054 19954 31106 19966
rect 31278 20018 31330 20030
rect 31278 19954 31330 19966
rect 31726 20018 31778 20030
rect 40798 20018 40850 20030
rect 35858 19966 35870 20018
rect 35922 19966 35934 20018
rect 31726 19954 31778 19966
rect 40798 19954 40850 19966
rect 41134 20018 41186 20030
rect 41134 19954 41186 19966
rect 41358 20018 41410 20030
rect 41358 19954 41410 19966
rect 41918 20018 41970 20030
rect 41918 19954 41970 19966
rect 42030 20018 42082 20030
rect 42030 19954 42082 19966
rect 43710 20018 43762 20030
rect 45726 20018 45778 20030
rect 45042 19966 45054 20018
rect 45106 19966 45118 20018
rect 43710 19954 43762 19966
rect 45726 19954 45778 19966
rect 46174 20018 46226 20030
rect 46174 19954 46226 19966
rect 15710 19906 15762 19918
rect 4946 19854 4958 19906
rect 5010 19854 5022 19906
rect 5730 19854 5742 19906
rect 5794 19854 5806 19906
rect 7858 19854 7870 19906
rect 7922 19854 7934 19906
rect 14018 19854 14030 19906
rect 14082 19854 14094 19906
rect 15710 19842 15762 19854
rect 17502 19906 17554 19918
rect 17502 19842 17554 19854
rect 18622 19906 18674 19918
rect 18622 19842 18674 19854
rect 19630 19906 19682 19918
rect 19630 19842 19682 19854
rect 26574 19906 26626 19918
rect 30270 19906 30322 19918
rect 27682 19854 27694 19906
rect 27746 19854 27758 19906
rect 29810 19854 29822 19906
rect 29874 19854 29886 19906
rect 26574 19842 26626 19854
rect 30270 19842 30322 19854
rect 33854 19906 33906 19918
rect 33854 19842 33906 19854
rect 34414 19906 34466 19918
rect 40014 19906 40066 19918
rect 37090 19854 37102 19906
rect 37154 19854 37166 19906
rect 34414 19842 34466 19854
rect 40014 19842 40066 19854
rect 41022 19906 41074 19918
rect 42814 19906 42866 19918
rect 42354 19854 42366 19906
rect 42418 19903 42430 19906
rect 42418 19857 42527 19903
rect 42418 19854 42430 19857
rect 41022 19842 41074 19854
rect 9774 19794 9826 19806
rect 9774 19730 9826 19742
rect 15262 19794 15314 19806
rect 15262 19730 15314 19742
rect 22654 19794 22706 19806
rect 42481 19791 42527 19857
rect 42814 19842 42866 19854
rect 44270 19906 44322 19918
rect 44270 19842 44322 19854
rect 44606 19906 44658 19918
rect 44606 19842 44658 19854
rect 43250 19791 43262 19794
rect 42481 19745 43262 19791
rect 43250 19742 43262 19745
rect 43314 19742 43326 19794
rect 22654 19730 22706 19742
rect 1344 19626 48608 19660
rect 1344 19574 4478 19626
rect 4530 19574 4582 19626
rect 4634 19574 4686 19626
rect 4738 19574 35198 19626
rect 35250 19574 35302 19626
rect 35354 19574 35406 19626
rect 35458 19574 48608 19626
rect 1344 19540 48608 19574
rect 6738 19406 6750 19458
rect 6802 19406 6814 19458
rect 12910 19346 12962 19358
rect 8306 19294 8318 19346
rect 8370 19294 8382 19346
rect 12114 19294 12126 19346
rect 12178 19294 12190 19346
rect 12910 19282 12962 19294
rect 16046 19346 16098 19358
rect 28142 19346 28194 19358
rect 34526 19346 34578 19358
rect 17826 19294 17838 19346
rect 17890 19343 17902 19346
rect 18162 19343 18174 19346
rect 17890 19297 18174 19343
rect 17890 19294 17902 19297
rect 18162 19294 18174 19297
rect 18226 19294 18238 19346
rect 20290 19294 20302 19346
rect 20354 19294 20366 19346
rect 23650 19294 23662 19346
rect 23714 19294 23726 19346
rect 29922 19294 29934 19346
rect 29986 19294 29998 19346
rect 32050 19294 32062 19346
rect 32114 19294 32126 19346
rect 33170 19294 33182 19346
rect 33234 19294 33246 19346
rect 16046 19282 16098 19294
rect 28142 19282 28194 19294
rect 34526 19282 34578 19294
rect 35310 19346 35362 19358
rect 35310 19282 35362 19294
rect 36206 19346 36258 19358
rect 36206 19282 36258 19294
rect 39118 19346 39170 19358
rect 46846 19346 46898 19358
rect 40226 19294 40238 19346
rect 40290 19294 40302 19346
rect 42354 19294 42366 19346
rect 42418 19294 42430 19346
rect 45154 19294 45166 19346
rect 45218 19294 45230 19346
rect 39118 19282 39170 19294
rect 46846 19282 46898 19294
rect 12462 19234 12514 19246
rect 7298 19182 7310 19234
rect 7362 19182 7374 19234
rect 11442 19182 11454 19234
rect 11506 19182 11518 19234
rect 11666 19182 11678 19234
rect 11730 19182 11742 19234
rect 12002 19182 12014 19234
rect 12066 19182 12078 19234
rect 12462 19170 12514 19182
rect 14142 19234 14194 19246
rect 14142 19170 14194 19182
rect 14254 19234 14306 19246
rect 14254 19170 14306 19182
rect 14590 19234 14642 19246
rect 14590 19170 14642 19182
rect 16382 19234 16434 19246
rect 16382 19170 16434 19182
rect 16718 19234 16770 19246
rect 16718 19170 16770 19182
rect 17278 19234 17330 19246
rect 25118 19234 25170 19246
rect 17826 19182 17838 19234
rect 17890 19182 17902 19234
rect 18722 19182 18734 19234
rect 18786 19182 18798 19234
rect 21522 19182 21534 19234
rect 21586 19182 21598 19234
rect 22082 19182 22094 19234
rect 22146 19182 22158 19234
rect 17278 19170 17330 19182
rect 25118 19170 25170 19182
rect 25454 19234 25506 19246
rect 25454 19170 25506 19182
rect 26238 19234 26290 19246
rect 26238 19170 26290 19182
rect 27918 19234 27970 19246
rect 27918 19170 27970 19182
rect 28254 19234 28306 19246
rect 32398 19234 32450 19246
rect 34750 19234 34802 19246
rect 29250 19182 29262 19234
rect 29314 19182 29326 19234
rect 33282 19182 33294 19234
rect 33346 19182 33358 19234
rect 28254 19170 28306 19182
rect 32398 19170 32450 19182
rect 34750 19170 34802 19182
rect 35198 19234 35250 19246
rect 36878 19234 36930 19246
rect 35746 19182 35758 19234
rect 35810 19182 35822 19234
rect 35198 19170 35250 19182
rect 36878 19170 36930 19182
rect 37214 19234 37266 19246
rect 43598 19234 43650 19246
rect 39554 19182 39566 19234
rect 39618 19182 39630 19234
rect 37214 19170 37266 19182
rect 43598 19170 43650 19182
rect 43822 19234 43874 19246
rect 44818 19182 44830 19234
rect 44882 19182 44894 19234
rect 45938 19182 45950 19234
rect 46002 19182 46014 19234
rect 43822 19170 43874 19182
rect 13694 19122 13746 19134
rect 10546 19070 10558 19122
rect 10610 19070 10622 19122
rect 13694 19058 13746 19070
rect 14478 19122 14530 19134
rect 14478 19058 14530 19070
rect 15150 19122 15202 19134
rect 15150 19058 15202 19070
rect 16942 19122 16994 19134
rect 25790 19122 25842 19134
rect 21746 19070 21758 19122
rect 21810 19070 21822 19122
rect 16942 19058 16994 19070
rect 25790 19058 25842 19070
rect 28590 19122 28642 19134
rect 28590 19058 28642 19070
rect 34414 19122 34466 19134
rect 34414 19058 34466 19070
rect 35422 19122 35474 19134
rect 35422 19058 35474 19070
rect 36094 19122 36146 19134
rect 36094 19058 36146 19070
rect 36318 19122 36370 19134
rect 36318 19058 36370 19070
rect 37550 19122 37602 19134
rect 37550 19058 37602 19070
rect 38222 19122 38274 19134
rect 38222 19058 38274 19070
rect 43374 19122 43426 19134
rect 46398 19122 46450 19134
rect 44930 19070 44942 19122
rect 44994 19070 45006 19122
rect 46498 19070 46510 19122
rect 46562 19119 46574 19122
rect 46722 19119 46734 19122
rect 46562 19073 46734 19119
rect 46562 19070 46574 19073
rect 46722 19070 46734 19073
rect 46786 19070 46798 19122
rect 43374 19058 43426 19070
rect 46398 19058 46450 19070
rect 12238 19010 12290 19022
rect 12238 18946 12290 18958
rect 13470 19010 13522 19022
rect 13470 18946 13522 18958
rect 13582 19010 13634 19022
rect 13582 18946 13634 18958
rect 15710 19010 15762 19022
rect 15710 18946 15762 18958
rect 16494 19010 16546 19022
rect 16494 18946 16546 18958
rect 17390 19010 17442 19022
rect 17390 18946 17442 18958
rect 17502 19010 17554 19022
rect 17502 18946 17554 18958
rect 25454 19010 25506 19022
rect 25454 18946 25506 18958
rect 27806 19010 27858 19022
rect 27806 18946 27858 18958
rect 34190 19010 34242 19022
rect 34190 18946 34242 18958
rect 37102 19010 37154 19022
rect 37102 18946 37154 18958
rect 37886 19010 37938 19022
rect 37886 18946 37938 18958
rect 38670 19010 38722 19022
rect 38670 18946 38722 18958
rect 42926 19010 42978 19022
rect 42926 18946 42978 18958
rect 43486 19010 43538 19022
rect 43486 18946 43538 18958
rect 46286 19010 46338 19022
rect 46286 18946 46338 18958
rect 1344 18842 48608 18876
rect 1344 18790 19838 18842
rect 19890 18790 19942 18842
rect 19994 18790 20046 18842
rect 20098 18790 48608 18842
rect 1344 18756 48608 18790
rect 8878 18674 8930 18686
rect 17614 18674 17666 18686
rect 24110 18674 24162 18686
rect 14578 18622 14590 18674
rect 14642 18622 14654 18674
rect 18722 18622 18734 18674
rect 18786 18622 18798 18674
rect 8878 18610 8930 18622
rect 17614 18610 17666 18622
rect 24110 18610 24162 18622
rect 24670 18674 24722 18686
rect 24670 18610 24722 18622
rect 28814 18674 28866 18686
rect 28814 18610 28866 18622
rect 33182 18674 33234 18686
rect 33182 18610 33234 18622
rect 35870 18674 35922 18686
rect 35870 18610 35922 18622
rect 16270 18562 16322 18574
rect 16270 18498 16322 18510
rect 16830 18562 16882 18574
rect 16830 18498 16882 18510
rect 19070 18562 19122 18574
rect 19070 18498 19122 18510
rect 21646 18562 21698 18574
rect 21646 18498 21698 18510
rect 28926 18562 28978 18574
rect 41246 18562 41298 18574
rect 40002 18510 40014 18562
rect 40066 18510 40078 18562
rect 28926 18498 28978 18510
rect 41246 18498 41298 18510
rect 42478 18562 42530 18574
rect 42478 18498 42530 18510
rect 44270 18562 44322 18574
rect 46050 18510 46062 18562
rect 46114 18510 46126 18562
rect 44270 18498 44322 18510
rect 10894 18450 10946 18462
rect 15150 18450 15202 18462
rect 10210 18398 10222 18450
rect 10274 18398 10286 18450
rect 11666 18398 11678 18450
rect 11730 18398 11742 18450
rect 12338 18398 12350 18450
rect 12402 18398 12414 18450
rect 10894 18386 10946 18398
rect 15150 18386 15202 18398
rect 15598 18450 15650 18462
rect 15598 18386 15650 18398
rect 16606 18450 16658 18462
rect 16606 18386 16658 18398
rect 17726 18450 17778 18462
rect 17726 18386 17778 18398
rect 17838 18450 17890 18462
rect 17838 18386 17890 18398
rect 18286 18450 18338 18462
rect 22206 18450 22258 18462
rect 20066 18398 20078 18450
rect 20130 18398 20142 18450
rect 18286 18386 18338 18398
rect 22206 18386 22258 18398
rect 22654 18450 22706 18462
rect 22654 18386 22706 18398
rect 22990 18450 23042 18462
rect 22990 18386 23042 18398
rect 23214 18450 23266 18462
rect 23214 18386 23266 18398
rect 23438 18450 23490 18462
rect 23438 18386 23490 18398
rect 23886 18450 23938 18462
rect 23886 18386 23938 18398
rect 23998 18450 24050 18462
rect 28702 18450 28754 18462
rect 32958 18450 33010 18462
rect 25218 18398 25230 18450
rect 25282 18398 25294 18450
rect 26002 18398 26014 18450
rect 26066 18398 26078 18450
rect 29250 18398 29262 18450
rect 29314 18398 29326 18450
rect 31938 18398 31950 18450
rect 32002 18398 32014 18450
rect 23998 18386 24050 18398
rect 28702 18386 28754 18398
rect 32958 18386 33010 18398
rect 33294 18450 33346 18462
rect 33294 18386 33346 18398
rect 33630 18450 33682 18462
rect 35534 18450 35586 18462
rect 40350 18450 40402 18462
rect 35074 18398 35086 18450
rect 35138 18398 35150 18450
rect 36082 18398 36094 18450
rect 36146 18398 36158 18450
rect 36866 18398 36878 18450
rect 36930 18398 36942 18450
rect 33630 18386 33682 18398
rect 35534 18386 35586 18398
rect 40350 18386 40402 18398
rect 40910 18450 40962 18462
rect 40910 18386 40962 18398
rect 41470 18450 41522 18462
rect 42702 18450 42754 18462
rect 42130 18398 42142 18450
rect 42194 18398 42206 18450
rect 41470 18386 41522 18398
rect 42702 18386 42754 18398
rect 42926 18450 42978 18462
rect 42926 18386 42978 18398
rect 43262 18450 43314 18462
rect 43262 18386 43314 18398
rect 43598 18450 43650 18462
rect 44830 18450 44882 18462
rect 44594 18398 44606 18450
rect 44658 18398 44670 18450
rect 45378 18398 45390 18450
rect 45442 18398 45454 18450
rect 43598 18386 43650 18398
rect 44830 18386 44882 18398
rect 16382 18338 16434 18350
rect 16382 18274 16434 18286
rect 22766 18338 22818 18350
rect 29710 18338 29762 18350
rect 28130 18286 28142 18338
rect 28194 18286 28206 18338
rect 29362 18286 29374 18338
rect 29426 18286 29438 18338
rect 22766 18274 22818 18286
rect 29377 18223 29423 18286
rect 29710 18274 29762 18286
rect 32510 18338 32562 18350
rect 39454 18338 39506 18350
rect 34626 18286 34638 18338
rect 34690 18286 34702 18338
rect 38994 18286 39006 18338
rect 39058 18286 39070 18338
rect 32510 18274 32562 18286
rect 39454 18274 39506 18286
rect 41022 18338 41074 18350
rect 41022 18274 41074 18286
rect 42590 18338 42642 18350
rect 42590 18274 42642 18286
rect 43150 18338 43202 18350
rect 43150 18274 43202 18286
rect 43934 18338 43986 18350
rect 44930 18286 44942 18338
rect 44994 18286 45006 18338
rect 48178 18286 48190 18338
rect 48242 18286 48254 18338
rect 43934 18274 43986 18286
rect 32286 18226 32338 18238
rect 29698 18223 29710 18226
rect 29377 18177 29710 18223
rect 29698 18174 29710 18177
rect 29762 18174 29774 18226
rect 32286 18162 32338 18174
rect 44046 18226 44098 18238
rect 44046 18162 44098 18174
rect 1344 18058 48608 18092
rect 1344 18006 4478 18058
rect 4530 18006 4582 18058
rect 4634 18006 4686 18058
rect 4738 18006 35198 18058
rect 35250 18006 35302 18058
rect 35354 18006 35406 18058
rect 35458 18006 48608 18058
rect 1344 17972 48608 18006
rect 33182 17890 33234 17902
rect 35086 17890 35138 17902
rect 19058 17838 19070 17890
rect 19122 17887 19134 17890
rect 19282 17887 19294 17890
rect 19122 17841 19294 17887
rect 19122 17838 19134 17841
rect 19282 17838 19294 17841
rect 19346 17887 19358 17890
rect 20066 17887 20078 17890
rect 19346 17841 20078 17887
rect 19346 17838 19358 17841
rect 20066 17838 20078 17841
rect 20130 17838 20142 17890
rect 33506 17838 33518 17890
rect 33570 17838 33582 17890
rect 33182 17826 33234 17838
rect 35086 17826 35138 17838
rect 35310 17890 35362 17902
rect 35310 17826 35362 17838
rect 37214 17890 37266 17902
rect 37214 17826 37266 17838
rect 10670 17778 10722 17790
rect 9986 17726 9998 17778
rect 10050 17726 10062 17778
rect 10670 17714 10722 17726
rect 11566 17778 11618 17790
rect 11566 17714 11618 17726
rect 12462 17778 12514 17790
rect 12462 17714 12514 17726
rect 13582 17778 13634 17790
rect 17390 17778 17442 17790
rect 14802 17726 14814 17778
rect 14866 17726 14878 17778
rect 16930 17726 16942 17778
rect 16994 17726 17006 17778
rect 13582 17714 13634 17726
rect 17390 17714 17442 17726
rect 17950 17778 18002 17790
rect 17950 17714 18002 17726
rect 19742 17778 19794 17790
rect 19742 17714 19794 17726
rect 20190 17778 20242 17790
rect 20190 17714 20242 17726
rect 20526 17778 20578 17790
rect 20526 17714 20578 17726
rect 21422 17778 21474 17790
rect 26126 17778 26178 17790
rect 22530 17726 22542 17778
rect 22594 17726 22606 17778
rect 24658 17726 24670 17778
rect 24722 17726 24734 17778
rect 21422 17714 21474 17726
rect 26126 17714 26178 17726
rect 31054 17778 31106 17790
rect 31054 17714 31106 17726
rect 32958 17778 33010 17790
rect 32958 17714 33010 17726
rect 36206 17778 36258 17790
rect 36206 17714 36258 17726
rect 37774 17778 37826 17790
rect 44830 17778 44882 17790
rect 40338 17726 40350 17778
rect 40402 17726 40414 17778
rect 44258 17726 44270 17778
rect 44322 17726 44334 17778
rect 48178 17726 48190 17778
rect 48242 17726 48254 17778
rect 37774 17714 37826 17726
rect 44830 17714 44882 17726
rect 9550 17666 9602 17678
rect 9550 17602 9602 17614
rect 10894 17666 10946 17678
rect 10894 17602 10946 17614
rect 11118 17666 11170 17678
rect 25006 17666 25058 17678
rect 14018 17614 14030 17666
rect 14082 17614 14094 17666
rect 21858 17614 21870 17666
rect 21922 17614 21934 17666
rect 11118 17602 11170 17614
rect 25006 17602 25058 17614
rect 26014 17666 26066 17678
rect 26014 17602 26066 17614
rect 26238 17666 26290 17678
rect 28590 17666 28642 17678
rect 27122 17614 27134 17666
rect 27186 17614 27198 17666
rect 26238 17602 26290 17614
rect 28590 17602 28642 17614
rect 29374 17666 29426 17678
rect 29374 17602 29426 17614
rect 29710 17666 29762 17678
rect 29710 17602 29762 17614
rect 29934 17666 29986 17678
rect 29934 17602 29986 17614
rect 30382 17666 30434 17678
rect 30382 17602 30434 17614
rect 30606 17666 30658 17678
rect 30606 17602 30658 17614
rect 33966 17666 34018 17678
rect 36094 17666 36146 17678
rect 34850 17614 34862 17666
rect 34914 17614 34926 17666
rect 33966 17602 34018 17614
rect 36094 17602 36146 17614
rect 36318 17666 36370 17678
rect 36318 17602 36370 17614
rect 37998 17666 38050 17678
rect 37998 17602 38050 17614
rect 38222 17666 38274 17678
rect 38222 17602 38274 17614
rect 38446 17666 38498 17678
rect 43262 17666 43314 17678
rect 39106 17614 39118 17666
rect 39170 17614 39182 17666
rect 42914 17614 42926 17666
rect 42978 17614 42990 17666
rect 38446 17602 38498 17614
rect 43262 17602 43314 17614
rect 43374 17666 43426 17678
rect 44158 17666 44210 17678
rect 43922 17614 43934 17666
rect 43986 17614 43998 17666
rect 45378 17614 45390 17666
rect 45442 17614 45454 17666
rect 43374 17602 43426 17614
rect 44158 17602 44210 17614
rect 10558 17554 10610 17566
rect 10558 17490 10610 17502
rect 18734 17554 18786 17566
rect 28478 17554 28530 17566
rect 25330 17502 25342 17554
rect 25394 17502 25406 17554
rect 18734 17490 18786 17502
rect 28478 17490 28530 17502
rect 29150 17554 29202 17566
rect 29150 17490 29202 17502
rect 31390 17554 31442 17566
rect 31390 17490 31442 17502
rect 34302 17554 34354 17566
rect 34302 17490 34354 17502
rect 34526 17554 34578 17566
rect 34526 17490 34578 17502
rect 35422 17554 35474 17566
rect 35422 17490 35474 17502
rect 35758 17554 35810 17566
rect 35758 17490 35810 17502
rect 37102 17554 37154 17566
rect 37102 17490 37154 17502
rect 38894 17554 38946 17566
rect 41806 17554 41858 17566
rect 39218 17502 39230 17554
rect 39282 17502 39294 17554
rect 38894 17490 38946 17502
rect 41806 17490 41858 17502
rect 43710 17554 43762 17566
rect 43710 17490 43762 17502
rect 44942 17554 44994 17566
rect 46050 17502 46062 17554
rect 46114 17502 46126 17554
rect 44942 17490 44994 17502
rect 13022 17442 13074 17454
rect 13022 17378 13074 17390
rect 18174 17442 18226 17454
rect 18174 17378 18226 17390
rect 19182 17442 19234 17454
rect 19182 17378 19234 17390
rect 26462 17442 26514 17454
rect 27694 17442 27746 17454
rect 26898 17390 26910 17442
rect 26962 17390 26974 17442
rect 26462 17378 26514 17390
rect 27694 17378 27746 17390
rect 28142 17442 28194 17454
rect 28142 17378 28194 17390
rect 28366 17442 28418 17454
rect 28366 17378 28418 17390
rect 29598 17442 29650 17454
rect 29598 17378 29650 17390
rect 30158 17442 30210 17454
rect 30158 17378 30210 17390
rect 30942 17442 30994 17454
rect 30942 17378 30994 17390
rect 31166 17442 31218 17454
rect 31166 17378 31218 17390
rect 34190 17442 34242 17454
rect 34190 17378 34242 17390
rect 37214 17442 37266 17454
rect 37214 17378 37266 17390
rect 1344 17274 48608 17308
rect 1344 17222 19838 17274
rect 19890 17222 19942 17274
rect 19994 17222 20046 17274
rect 20098 17222 48608 17274
rect 1344 17188 48608 17222
rect 12014 17106 12066 17118
rect 12014 17042 12066 17054
rect 12798 17106 12850 17118
rect 12798 17042 12850 17054
rect 13582 17106 13634 17118
rect 13582 17042 13634 17054
rect 17502 17106 17554 17118
rect 17502 17042 17554 17054
rect 18062 17106 18114 17118
rect 18062 17042 18114 17054
rect 21534 17106 21586 17118
rect 21534 17042 21586 17054
rect 25342 17106 25394 17118
rect 25342 17042 25394 17054
rect 30830 17106 30882 17118
rect 30830 17042 30882 17054
rect 31726 17106 31778 17118
rect 31726 17042 31778 17054
rect 34190 17106 34242 17118
rect 34190 17042 34242 17054
rect 34414 17106 34466 17118
rect 34414 17042 34466 17054
rect 35422 17106 35474 17118
rect 35422 17042 35474 17054
rect 36318 17106 36370 17118
rect 36318 17042 36370 17054
rect 43598 17106 43650 17118
rect 43598 17042 43650 17054
rect 43822 17106 43874 17118
rect 45614 17106 45666 17118
rect 45042 17054 45054 17106
rect 45106 17054 45118 17106
rect 43822 17042 43874 17054
rect 45614 17042 45666 17054
rect 47854 17106 47906 17118
rect 47854 17042 47906 17054
rect 18622 16994 18674 17006
rect 14690 16942 14702 16994
rect 14754 16942 14766 16994
rect 18622 16930 18674 16942
rect 19630 16994 19682 17006
rect 19630 16930 19682 16942
rect 21646 16994 21698 17006
rect 21646 16930 21698 16942
rect 26910 16994 26962 17006
rect 33294 16994 33346 17006
rect 29362 16942 29374 16994
rect 29426 16942 29438 16994
rect 26910 16930 26962 16942
rect 33294 16930 33346 16942
rect 36094 16994 36146 17006
rect 36094 16930 36146 16942
rect 36430 16994 36482 17006
rect 36430 16930 36482 16942
rect 37438 16994 37490 17006
rect 37438 16930 37490 16942
rect 38334 16994 38386 17006
rect 38334 16930 38386 16942
rect 38894 16994 38946 17006
rect 38894 16930 38946 16942
rect 41134 16994 41186 17006
rect 41134 16930 41186 16942
rect 42366 16994 42418 17006
rect 42366 16930 42418 16942
rect 11566 16882 11618 16894
rect 18734 16882 18786 16894
rect 22766 16882 22818 16894
rect 14018 16830 14030 16882
rect 14082 16830 14094 16882
rect 19058 16830 19070 16882
rect 19122 16830 19134 16882
rect 11566 16818 11618 16830
rect 18734 16818 18786 16830
rect 22766 16818 22818 16830
rect 26574 16882 26626 16894
rect 31390 16882 31442 16894
rect 34974 16882 35026 16894
rect 30146 16830 30158 16882
rect 30210 16830 30222 16882
rect 33506 16830 33518 16882
rect 33570 16830 33582 16882
rect 26574 16818 26626 16830
rect 31390 16818 31442 16830
rect 34974 16818 35026 16830
rect 36654 16882 36706 16894
rect 37886 16882 37938 16894
rect 37650 16830 37662 16882
rect 37714 16830 37726 16882
rect 36654 16818 36706 16830
rect 37886 16818 37938 16830
rect 38558 16882 38610 16894
rect 38558 16818 38610 16830
rect 38782 16882 38834 16894
rect 38782 16818 38834 16830
rect 39566 16882 39618 16894
rect 39566 16818 39618 16830
rect 39790 16882 39842 16894
rect 39790 16818 39842 16830
rect 40910 16882 40962 16894
rect 40910 16818 40962 16830
rect 41582 16882 41634 16894
rect 41582 16818 41634 16830
rect 41694 16882 41746 16894
rect 41694 16818 41746 16830
rect 42030 16882 42082 16894
rect 42030 16818 42082 16830
rect 42702 16882 42754 16894
rect 42702 16818 42754 16830
rect 42926 16882 42978 16894
rect 44494 16882 44546 16894
rect 44146 16830 44158 16882
rect 44210 16830 44222 16882
rect 42926 16818 42978 16830
rect 44494 16818 44546 16830
rect 45390 16882 45442 16894
rect 45390 16818 45442 16830
rect 46062 16882 46114 16894
rect 46062 16818 46114 16830
rect 46286 16882 46338 16894
rect 46286 16818 46338 16830
rect 47182 16882 47234 16894
rect 47182 16818 47234 16830
rect 47406 16882 47458 16894
rect 47406 16818 47458 16830
rect 40238 16770 40290 16782
rect 16818 16718 16830 16770
rect 16882 16718 16894 16770
rect 27234 16718 27246 16770
rect 27298 16718 27310 16770
rect 37986 16718 37998 16770
rect 38050 16718 38062 16770
rect 40238 16706 40290 16718
rect 41022 16770 41074 16782
rect 41022 16706 41074 16718
rect 41918 16770 41970 16782
rect 41918 16706 41970 16718
rect 43710 16770 43762 16782
rect 43710 16706 43762 16718
rect 44718 16770 44770 16782
rect 44718 16706 44770 16718
rect 45502 16770 45554 16782
rect 45502 16706 45554 16718
rect 46734 16770 46786 16782
rect 46734 16706 46786 16718
rect 46958 16770 47010 16782
rect 46958 16706 47010 16718
rect 36990 16658 37042 16670
rect 30818 16606 30830 16658
rect 30882 16655 30894 16658
rect 31602 16655 31614 16658
rect 30882 16609 31614 16655
rect 30882 16606 30894 16609
rect 31602 16606 31614 16609
rect 31666 16606 31678 16658
rect 36990 16594 37042 16606
rect 37102 16658 37154 16670
rect 39218 16606 39230 16658
rect 39282 16606 39294 16658
rect 43250 16606 43262 16658
rect 43314 16606 43326 16658
rect 37102 16594 37154 16606
rect 1344 16490 48608 16524
rect 1344 16438 4478 16490
rect 4530 16438 4582 16490
rect 4634 16438 4686 16490
rect 4738 16438 35198 16490
rect 35250 16438 35302 16490
rect 35354 16438 35406 16490
rect 35458 16438 48608 16490
rect 1344 16404 48608 16438
rect 19742 16322 19794 16334
rect 19742 16258 19794 16270
rect 36094 16322 36146 16334
rect 36094 16258 36146 16270
rect 36430 16322 36482 16334
rect 36430 16258 36482 16270
rect 43822 16322 43874 16334
rect 43822 16258 43874 16270
rect 45950 16322 46002 16334
rect 46274 16270 46286 16322
rect 46338 16270 46350 16322
rect 45950 16258 46002 16270
rect 14590 16210 14642 16222
rect 14590 16146 14642 16158
rect 14926 16210 14978 16222
rect 14926 16146 14978 16158
rect 16270 16210 16322 16222
rect 16270 16146 16322 16158
rect 16830 16210 16882 16222
rect 16830 16146 16882 16158
rect 23102 16210 23154 16222
rect 35198 16210 35250 16222
rect 44270 16210 44322 16222
rect 26450 16158 26462 16210
rect 26514 16158 26526 16210
rect 30146 16158 30158 16210
rect 30210 16158 30222 16210
rect 32274 16158 32286 16210
rect 32338 16158 32350 16210
rect 39218 16158 39230 16210
rect 39282 16158 39294 16210
rect 41794 16158 41806 16210
rect 41858 16158 41870 16210
rect 23102 16146 23154 16158
rect 35198 16146 35250 16158
rect 44270 16146 44322 16158
rect 46734 16210 46786 16222
rect 46734 16146 46786 16158
rect 17502 16098 17554 16110
rect 17502 16034 17554 16046
rect 21646 16098 21698 16110
rect 21646 16034 21698 16046
rect 22206 16098 22258 16110
rect 33966 16098 34018 16110
rect 23650 16046 23662 16098
rect 23714 16046 23726 16098
rect 29362 16046 29374 16098
rect 29426 16046 29438 16098
rect 33506 16046 33518 16098
rect 33570 16046 33582 16098
rect 22206 16034 22258 16046
rect 33966 16034 34018 16046
rect 35534 16098 35586 16110
rect 35534 16034 35586 16046
rect 35870 16098 35922 16110
rect 42926 16098 42978 16110
rect 43710 16098 43762 16110
rect 37538 16046 37550 16098
rect 37602 16046 37614 16098
rect 39890 16046 39902 16098
rect 39954 16046 39966 16098
rect 43138 16046 43150 16098
rect 43202 16046 43214 16098
rect 35870 16034 35922 16046
rect 42926 16034 42978 16046
rect 43710 16034 43762 16046
rect 45054 16098 45106 16110
rect 45726 16098 45778 16110
rect 45378 16046 45390 16098
rect 45442 16046 45454 16098
rect 45054 16034 45106 16046
rect 45726 16034 45778 16046
rect 17166 15986 17218 15998
rect 17166 15922 17218 15934
rect 17726 15986 17778 15998
rect 17726 15922 17778 15934
rect 18510 15986 18562 15998
rect 19742 15986 19794 15998
rect 18510 15922 18562 15934
rect 19630 15930 19682 15942
rect 17278 15874 17330 15886
rect 19182 15874 19234 15886
rect 18834 15822 18846 15874
rect 18898 15822 18910 15874
rect 19742 15922 19794 15934
rect 20414 15986 20466 15998
rect 20414 15922 20466 15934
rect 20750 15986 20802 15998
rect 20750 15922 20802 15934
rect 21310 15986 21362 15998
rect 21310 15922 21362 15934
rect 21870 15986 21922 15998
rect 34302 15986 34354 15998
rect 36318 15986 36370 15998
rect 22530 15934 22542 15986
rect 22594 15934 22606 15986
rect 24322 15934 24334 15986
rect 24386 15934 24398 15986
rect 34626 15934 34638 15986
rect 34690 15934 34702 15986
rect 21870 15922 21922 15934
rect 34302 15922 34354 15934
rect 36318 15922 36370 15934
rect 44942 15986 44994 15998
rect 44942 15922 44994 15934
rect 47854 15986 47906 15998
rect 47854 15922 47906 15934
rect 48190 15986 48242 15998
rect 48190 15922 48242 15934
rect 19630 15866 19682 15878
rect 21422 15874 21474 15886
rect 17278 15810 17330 15822
rect 19182 15810 19234 15822
rect 21422 15810 21474 15822
rect 35646 15874 35698 15886
rect 35646 15810 35698 15822
rect 43038 15874 43090 15886
rect 43038 15810 43090 15822
rect 43374 15874 43426 15886
rect 43374 15810 43426 15822
rect 44830 15874 44882 15886
rect 44830 15810 44882 15822
rect 47630 15874 47682 15886
rect 47630 15810 47682 15822
rect 1344 15706 48608 15740
rect 1344 15654 19838 15706
rect 19890 15654 19942 15706
rect 19994 15654 20046 15706
rect 20098 15654 48608 15706
rect 1344 15620 48608 15654
rect 17614 15538 17666 15550
rect 17614 15474 17666 15486
rect 18062 15538 18114 15550
rect 26574 15538 26626 15550
rect 20514 15486 20526 15538
rect 20578 15486 20590 15538
rect 25218 15486 25230 15538
rect 25282 15486 25294 15538
rect 18062 15474 18114 15486
rect 26574 15474 26626 15486
rect 27134 15538 27186 15550
rect 27134 15474 27186 15486
rect 29598 15538 29650 15550
rect 33294 15538 33346 15550
rect 31602 15486 31614 15538
rect 31666 15486 31678 15538
rect 29598 15474 29650 15486
rect 33294 15474 33346 15486
rect 33854 15538 33906 15550
rect 33854 15474 33906 15486
rect 40238 15538 40290 15550
rect 40238 15474 40290 15486
rect 41582 15538 41634 15550
rect 41582 15474 41634 15486
rect 16606 15426 16658 15438
rect 22206 15426 22258 15438
rect 19170 15374 19182 15426
rect 19234 15374 19246 15426
rect 16606 15362 16658 15374
rect 22206 15362 22258 15374
rect 30718 15426 30770 15438
rect 30718 15362 30770 15374
rect 38446 15426 38498 15438
rect 38446 15362 38498 15374
rect 38894 15426 38946 15438
rect 38894 15362 38946 15374
rect 39454 15426 39506 15438
rect 39454 15362 39506 15374
rect 41470 15426 41522 15438
rect 42030 15426 42082 15438
rect 41682 15374 41694 15426
rect 41746 15374 41758 15426
rect 41470 15362 41522 15374
rect 42030 15362 42082 15374
rect 43598 15426 43650 15438
rect 43598 15362 43650 15374
rect 16270 15314 16322 15326
rect 16270 15250 16322 15262
rect 16830 15314 16882 15326
rect 16830 15250 16882 15262
rect 17950 15314 18002 15326
rect 17950 15250 18002 15262
rect 18174 15314 18226 15326
rect 18174 15250 18226 15262
rect 18622 15314 18674 15326
rect 22766 15314 22818 15326
rect 25790 15314 25842 15326
rect 19058 15262 19070 15314
rect 19122 15262 19134 15314
rect 24098 15262 24110 15314
rect 24162 15262 24174 15314
rect 18622 15250 18674 15262
rect 22766 15250 22818 15262
rect 25790 15250 25842 15262
rect 26014 15314 26066 15326
rect 26798 15314 26850 15326
rect 26338 15262 26350 15314
rect 26402 15262 26414 15314
rect 26014 15250 26066 15262
rect 26798 15250 26850 15262
rect 27246 15314 27298 15326
rect 27246 15250 27298 15262
rect 27470 15314 27522 15326
rect 27470 15250 27522 15262
rect 30158 15314 30210 15326
rect 30158 15250 30210 15262
rect 30942 15314 30994 15326
rect 30942 15250 30994 15262
rect 31278 15314 31330 15326
rect 31278 15250 31330 15262
rect 32174 15314 32226 15326
rect 39006 15314 39058 15326
rect 39678 15314 39730 15326
rect 35074 15262 35086 15314
rect 35138 15262 35150 15314
rect 39106 15262 39118 15314
rect 39170 15262 39182 15314
rect 32174 15250 32226 15262
rect 39006 15250 39058 15262
rect 39678 15250 39730 15262
rect 39790 15314 39842 15326
rect 39790 15250 39842 15262
rect 42254 15314 42306 15326
rect 42254 15250 42306 15262
rect 42366 15314 42418 15326
rect 43038 15314 43090 15326
rect 42690 15262 42702 15314
rect 42754 15262 42766 15314
rect 42366 15250 42418 15262
rect 43038 15250 43090 15262
rect 43262 15314 43314 15326
rect 43262 15250 43314 15262
rect 43710 15314 43762 15326
rect 44146 15262 44158 15314
rect 44210 15262 44222 15314
rect 44818 15262 44830 15314
rect 44882 15262 44894 15314
rect 43710 15250 43762 15262
rect 16382 15202 16434 15214
rect 25566 15202 25618 15214
rect 23874 15150 23886 15202
rect 23938 15150 23950 15202
rect 16382 15138 16434 15150
rect 25566 15138 25618 15150
rect 26238 15202 26290 15214
rect 26238 15138 26290 15150
rect 27918 15202 27970 15214
rect 27918 15138 27970 15150
rect 30830 15202 30882 15214
rect 38334 15202 38386 15214
rect 35858 15150 35870 15202
rect 35922 15150 35934 15202
rect 37986 15150 37998 15202
rect 38050 15150 38062 15202
rect 46946 15150 46958 15202
rect 47010 15150 47022 15202
rect 30830 15138 30882 15150
rect 38334 15138 38386 15150
rect 31950 15090 32002 15102
rect 17266 15038 17278 15090
rect 17330 15087 17342 15090
rect 17602 15087 17614 15090
rect 17330 15041 17614 15087
rect 17330 15038 17342 15041
rect 17602 15038 17614 15041
rect 17666 15038 17678 15090
rect 24546 15038 24558 15090
rect 24610 15038 24622 15090
rect 31950 15026 32002 15038
rect 33070 15090 33122 15102
rect 33070 15026 33122 15038
rect 33406 15090 33458 15102
rect 33406 15026 33458 15038
rect 1344 14922 48608 14956
rect 1344 14870 4478 14922
rect 4530 14870 4582 14922
rect 4634 14870 4686 14922
rect 4738 14870 35198 14922
rect 35250 14870 35302 14922
rect 35354 14870 35406 14922
rect 35458 14870 48608 14922
rect 1344 14836 48608 14870
rect 30258 14702 30270 14754
rect 30322 14751 30334 14754
rect 31042 14751 31054 14754
rect 30322 14705 31054 14751
rect 30322 14702 30334 14705
rect 31042 14702 31054 14705
rect 31106 14702 31118 14754
rect 18846 14642 18898 14654
rect 16034 14590 16046 14642
rect 16098 14590 16110 14642
rect 18162 14590 18174 14642
rect 18226 14590 18238 14642
rect 18846 14578 18898 14590
rect 20638 14642 20690 14654
rect 30494 14642 30546 14654
rect 35534 14642 35586 14654
rect 25666 14590 25678 14642
rect 25730 14590 25742 14642
rect 27794 14590 27806 14642
rect 27858 14590 27870 14642
rect 29586 14590 29598 14642
rect 29650 14590 29662 14642
rect 31378 14590 31390 14642
rect 31442 14590 31454 14642
rect 33506 14590 33518 14642
rect 33570 14590 33582 14642
rect 20638 14578 20690 14590
rect 30494 14578 30546 14590
rect 35534 14578 35586 14590
rect 36430 14642 36482 14654
rect 44942 14642 44994 14654
rect 38098 14590 38110 14642
rect 38162 14590 38174 14642
rect 41346 14590 41358 14642
rect 41410 14590 41422 14642
rect 36430 14578 36482 14590
rect 44942 14578 44994 14590
rect 19182 14530 19234 14542
rect 15250 14478 15262 14530
rect 15314 14478 15326 14530
rect 19182 14466 19234 14478
rect 19294 14530 19346 14542
rect 19294 14466 19346 14478
rect 19742 14530 19794 14542
rect 24782 14530 24834 14542
rect 23874 14478 23886 14530
rect 23938 14478 23950 14530
rect 19742 14466 19794 14478
rect 24782 14466 24834 14478
rect 25006 14530 25058 14542
rect 34526 14530 34578 14542
rect 28578 14478 28590 14530
rect 28642 14478 28654 14530
rect 34290 14478 34302 14530
rect 34354 14478 34366 14530
rect 25006 14466 25058 14478
rect 34526 14466 34578 14478
rect 37326 14530 37378 14542
rect 41010 14478 41022 14530
rect 41074 14478 41086 14530
rect 44146 14478 44158 14530
rect 44210 14478 44222 14530
rect 37326 14466 37378 14478
rect 20526 14418 20578 14430
rect 25342 14418 25394 14430
rect 22082 14366 22094 14418
rect 22146 14366 22158 14418
rect 20526 14354 20578 14366
rect 25342 14354 25394 14366
rect 35086 14418 35138 14430
rect 37650 14366 37662 14418
rect 37714 14366 37726 14418
rect 40226 14366 40238 14418
rect 40290 14366 40302 14418
rect 43474 14366 43486 14418
rect 43538 14366 43550 14418
rect 35086 14354 35138 14366
rect 19518 14306 19570 14318
rect 19518 14242 19570 14254
rect 20302 14306 20354 14318
rect 20302 14242 20354 14254
rect 20750 14306 20802 14318
rect 20750 14242 20802 14254
rect 24334 14306 24386 14318
rect 24334 14242 24386 14254
rect 25006 14306 25058 14318
rect 25006 14242 25058 14254
rect 30046 14306 30098 14318
rect 30046 14242 30098 14254
rect 31054 14306 31106 14318
rect 31054 14242 31106 14254
rect 34862 14306 34914 14318
rect 34862 14242 34914 14254
rect 35198 14306 35250 14318
rect 35198 14242 35250 14254
rect 1344 14138 48608 14172
rect 1344 14086 19838 14138
rect 19890 14086 19942 14138
rect 19994 14086 20046 14138
rect 20098 14086 48608 14138
rect 1344 14052 48608 14086
rect 17726 13970 17778 13982
rect 17726 13906 17778 13918
rect 19518 13970 19570 13982
rect 19518 13906 19570 13918
rect 23550 13970 23602 13982
rect 23550 13906 23602 13918
rect 26798 13970 26850 13982
rect 26798 13906 26850 13918
rect 27694 13970 27746 13982
rect 27694 13906 27746 13918
rect 30830 13970 30882 13982
rect 30830 13906 30882 13918
rect 33630 13970 33682 13982
rect 33630 13906 33682 13918
rect 35422 13970 35474 13982
rect 35422 13906 35474 13918
rect 36206 13970 36258 13982
rect 36206 13906 36258 13918
rect 36990 13970 37042 13982
rect 36990 13906 37042 13918
rect 39230 13970 39282 13982
rect 41918 13970 41970 13982
rect 41458 13918 41470 13970
rect 41522 13918 41534 13970
rect 39230 13906 39282 13918
rect 41918 13906 41970 13918
rect 43038 13970 43090 13982
rect 43038 13906 43090 13918
rect 43374 13970 43426 13982
rect 43374 13906 43426 13918
rect 43822 13970 43874 13982
rect 43822 13906 43874 13918
rect 46174 13970 46226 13982
rect 46174 13906 46226 13918
rect 17838 13858 17890 13870
rect 23886 13858 23938 13870
rect 14690 13806 14702 13858
rect 14754 13806 14766 13858
rect 20738 13806 20750 13858
rect 20802 13806 20814 13858
rect 17838 13794 17890 13806
rect 23886 13794 23938 13806
rect 27246 13858 27298 13870
rect 27246 13794 27298 13806
rect 32510 13858 32562 13870
rect 32510 13794 32562 13806
rect 33406 13858 33458 13870
rect 33406 13794 33458 13806
rect 33742 13858 33794 13870
rect 33742 13794 33794 13806
rect 35534 13858 35586 13870
rect 35534 13794 35586 13806
rect 35758 13858 35810 13870
rect 35758 13794 35810 13806
rect 39118 13858 39170 13870
rect 39118 13794 39170 13806
rect 42366 13858 42418 13870
rect 42366 13794 42418 13806
rect 45614 13858 45666 13870
rect 45614 13794 45666 13806
rect 45726 13858 45778 13870
rect 45726 13794 45778 13806
rect 17950 13746 18002 13758
rect 14018 13694 14030 13746
rect 14082 13694 14094 13746
rect 17950 13682 18002 13694
rect 18398 13746 18450 13758
rect 18398 13682 18450 13694
rect 18958 13746 19010 13758
rect 18958 13682 19010 13694
rect 19406 13746 19458 13758
rect 19406 13682 19458 13694
rect 19630 13746 19682 13758
rect 23662 13746 23714 13758
rect 20066 13694 20078 13746
rect 20130 13694 20142 13746
rect 19630 13682 19682 13694
rect 23662 13682 23714 13694
rect 23998 13746 24050 13758
rect 23998 13682 24050 13694
rect 24334 13746 24386 13758
rect 24334 13682 24386 13694
rect 25230 13746 25282 13758
rect 25230 13682 25282 13694
rect 25454 13746 25506 13758
rect 25454 13682 25506 13694
rect 25902 13746 25954 13758
rect 25902 13682 25954 13694
rect 26686 13746 26738 13758
rect 26686 13682 26738 13694
rect 27022 13746 27074 13758
rect 33966 13746 34018 13758
rect 29922 13694 29934 13746
rect 29986 13694 29998 13746
rect 31826 13694 31838 13746
rect 31890 13694 31902 13746
rect 27022 13682 27074 13694
rect 33966 13682 34018 13694
rect 34414 13746 34466 13758
rect 34414 13682 34466 13694
rect 35086 13746 35138 13758
rect 35086 13682 35138 13694
rect 41134 13746 41186 13758
rect 41134 13682 41186 13694
rect 44494 13746 44546 13758
rect 44494 13682 44546 13694
rect 44942 13746 44994 13758
rect 44942 13682 44994 13694
rect 45054 13746 45106 13758
rect 45054 13682 45106 13694
rect 45390 13746 45442 13758
rect 45390 13682 45442 13694
rect 18734 13634 18786 13646
rect 25342 13634 25394 13646
rect 16818 13582 16830 13634
rect 16882 13582 16894 13634
rect 22866 13582 22878 13634
rect 22930 13582 22942 13634
rect 18734 13570 18786 13582
rect 25342 13570 25394 13582
rect 26126 13634 26178 13646
rect 26126 13570 26178 13582
rect 27694 13634 27746 13646
rect 44270 13634 44322 13646
rect 30258 13582 30270 13634
rect 30322 13582 30334 13634
rect 31938 13582 31950 13634
rect 32002 13582 32014 13634
rect 27694 13570 27746 13582
rect 44270 13570 44322 13582
rect 44718 13634 44770 13646
rect 44718 13570 44770 13582
rect 26238 13522 26290 13534
rect 26238 13458 26290 13470
rect 27806 13522 27858 13534
rect 27806 13458 27858 13470
rect 28030 13522 28082 13534
rect 28030 13458 28082 13470
rect 34526 13522 34578 13534
rect 34526 13458 34578 13470
rect 34750 13522 34802 13534
rect 34750 13458 34802 13470
rect 34862 13522 34914 13534
rect 34862 13458 34914 13470
rect 42478 13522 42530 13534
rect 42690 13470 42702 13522
rect 42754 13519 42766 13522
rect 43474 13519 43486 13522
rect 42754 13473 43486 13519
rect 42754 13470 42766 13473
rect 43474 13470 43486 13473
rect 43538 13470 43550 13522
rect 42478 13458 42530 13470
rect 1344 13354 48608 13388
rect 1344 13302 4478 13354
rect 4530 13302 4582 13354
rect 4634 13302 4686 13354
rect 4738 13302 35198 13354
rect 35250 13302 35302 13354
rect 35354 13302 35406 13354
rect 35458 13302 48608 13354
rect 1344 13268 48608 13302
rect 17054 13074 17106 13086
rect 27694 13074 27746 13086
rect 34190 13074 34242 13086
rect 24210 13022 24222 13074
rect 24274 13022 24286 13074
rect 25666 13022 25678 13074
rect 25730 13022 25742 13074
rect 32162 13022 32174 13074
rect 32226 13022 32238 13074
rect 45602 13022 45614 13074
rect 45666 13022 45678 13074
rect 47730 13022 47742 13074
rect 47794 13022 47806 13074
rect 17054 13010 17106 13022
rect 27694 13010 27746 13022
rect 34190 13010 34242 13022
rect 34414 12962 34466 12974
rect 18722 12910 18734 12962
rect 18786 12910 18798 12962
rect 21298 12910 21310 12962
rect 21362 12910 21374 12962
rect 25106 12910 25118 12962
rect 25170 12910 25182 12962
rect 29362 12910 29374 12962
rect 29426 12910 29438 12962
rect 34414 12898 34466 12910
rect 34638 12962 34690 12974
rect 34638 12898 34690 12910
rect 43934 12962 43986 12974
rect 43934 12898 43986 12910
rect 44270 12962 44322 12974
rect 44818 12910 44830 12962
rect 44882 12910 44894 12962
rect 44270 12898 44322 12910
rect 18174 12850 18226 12862
rect 34078 12850 34130 12862
rect 22082 12798 22094 12850
rect 22146 12798 22158 12850
rect 30034 12798 30046 12850
rect 30098 12798 30110 12850
rect 18174 12786 18226 12798
rect 34078 12786 34130 12798
rect 35086 12850 35138 12862
rect 35086 12786 35138 12798
rect 41918 12738 41970 12750
rect 17826 12686 17838 12738
rect 17890 12686 17902 12738
rect 18946 12686 18958 12738
rect 19010 12686 19022 12738
rect 41918 12674 41970 12686
rect 42366 12738 42418 12750
rect 42366 12674 42418 12686
rect 43710 12738 43762 12750
rect 43710 12674 43762 12686
rect 44046 12738 44098 12750
rect 44046 12674 44098 12686
rect 1344 12570 48608 12604
rect 1344 12518 19838 12570
rect 19890 12518 19942 12570
rect 19994 12518 20046 12570
rect 20098 12518 48608 12570
rect 1344 12484 48608 12518
rect 17502 12402 17554 12414
rect 17502 12338 17554 12350
rect 17838 12402 17890 12414
rect 19070 12402 19122 12414
rect 26574 12402 26626 12414
rect 18722 12350 18734 12402
rect 18786 12350 18798 12402
rect 20514 12350 20526 12402
rect 20578 12350 20590 12402
rect 17838 12338 17890 12350
rect 19070 12338 19122 12350
rect 26574 12338 26626 12350
rect 29598 12402 29650 12414
rect 39790 12402 39842 12414
rect 38098 12350 38110 12402
rect 38162 12350 38174 12402
rect 29598 12338 29650 12350
rect 39790 12338 39842 12350
rect 44494 12402 44546 12414
rect 44494 12338 44546 12350
rect 16270 12290 16322 12302
rect 16270 12226 16322 12238
rect 16606 12290 16658 12302
rect 16606 12226 16658 12238
rect 16830 12290 16882 12302
rect 16830 12226 16882 12238
rect 19742 12290 19794 12302
rect 19742 12226 19794 12238
rect 27134 12290 27186 12302
rect 28478 12290 28530 12302
rect 30382 12290 30434 12302
rect 28130 12238 28142 12290
rect 28194 12238 28206 12290
rect 28802 12238 28814 12290
rect 28866 12238 28878 12290
rect 30146 12238 30158 12290
rect 30210 12238 30222 12290
rect 31166 12290 31218 12302
rect 27134 12226 27186 12238
rect 28478 12226 28530 12238
rect 30382 12226 30434 12238
rect 30494 12234 30546 12246
rect 17950 12178 18002 12190
rect 17950 12114 18002 12126
rect 18062 12178 18114 12190
rect 31166 12226 31218 12238
rect 31614 12290 31666 12302
rect 31614 12226 31666 12238
rect 31726 12290 31778 12302
rect 31726 12226 31778 12238
rect 32174 12290 32226 12302
rect 35298 12238 35310 12290
rect 35362 12238 35374 12290
rect 38770 12238 38782 12290
rect 38834 12238 38846 12290
rect 39106 12238 39118 12290
rect 39170 12238 39182 12290
rect 40114 12238 40126 12290
rect 40178 12238 40190 12290
rect 32174 12226 32226 12238
rect 18386 12126 18398 12178
rect 18450 12126 18462 12178
rect 20290 12126 20302 12178
rect 20354 12126 20366 12178
rect 24546 12126 24558 12178
rect 24610 12126 24622 12178
rect 25778 12126 25790 12178
rect 25842 12126 25854 12178
rect 26114 12126 26126 12178
rect 26178 12126 26190 12178
rect 26786 12126 26798 12178
rect 26850 12126 26862 12178
rect 27906 12126 27918 12178
rect 27970 12126 27982 12178
rect 30494 12170 30546 12182
rect 30718 12178 30770 12190
rect 18062 12114 18114 12126
rect 30718 12114 30770 12126
rect 30942 12178 30994 12190
rect 30942 12114 30994 12126
rect 31278 12178 31330 12190
rect 37774 12178 37826 12190
rect 33842 12126 33854 12178
rect 33906 12126 33918 12178
rect 34514 12126 34526 12178
rect 34578 12126 34590 12178
rect 38546 12126 38558 12178
rect 38610 12126 38622 12178
rect 39330 12126 39342 12178
rect 39394 12126 39406 12178
rect 40898 12126 40910 12178
rect 40962 12126 40974 12178
rect 31278 12114 31330 12126
rect 37774 12114 37826 12126
rect 16382 12066 16434 12078
rect 34078 12066 34130 12078
rect 21746 12014 21758 12066
rect 21810 12014 21822 12066
rect 23874 12014 23886 12066
rect 23938 12014 23950 12066
rect 25330 12014 25342 12066
rect 25394 12014 25406 12066
rect 30370 12014 30382 12066
rect 30434 12014 30446 12066
rect 37426 12014 37438 12066
rect 37490 12014 37502 12066
rect 41682 12014 41694 12066
rect 41746 12014 41758 12066
rect 43810 12014 43822 12066
rect 43874 12014 43886 12066
rect 16382 12002 16434 12014
rect 34078 12002 34130 12014
rect 26798 11954 26850 11966
rect 26798 11890 26850 11902
rect 34190 11954 34242 11966
rect 34190 11890 34242 11902
rect 1344 11786 48608 11820
rect 1344 11734 4478 11786
rect 4530 11734 4582 11786
rect 4634 11734 4686 11786
rect 4738 11734 35198 11786
rect 35250 11734 35302 11786
rect 35354 11734 35406 11786
rect 35458 11734 48608 11786
rect 1344 11700 48608 11734
rect 23438 11618 23490 11630
rect 24446 11618 24498 11630
rect 32734 11618 32786 11630
rect 23762 11566 23774 11618
rect 23826 11566 23838 11618
rect 27010 11566 27022 11618
rect 27074 11615 27086 11618
rect 27794 11615 27806 11618
rect 27074 11569 27806 11615
rect 27074 11566 27086 11569
rect 27794 11566 27806 11569
rect 27858 11566 27870 11618
rect 34178 11566 34190 11618
rect 34242 11566 34254 11618
rect 23438 11554 23490 11566
rect 24446 11554 24498 11566
rect 32734 11554 32786 11566
rect 23214 11506 23266 11518
rect 41246 11506 41298 11518
rect 15586 11454 15598 11506
rect 15650 11454 15662 11506
rect 17714 11454 17726 11506
rect 17778 11454 17790 11506
rect 34290 11454 34302 11506
rect 34354 11454 34366 11506
rect 43026 11454 43038 11506
rect 43090 11454 43102 11506
rect 23214 11442 23266 11454
rect 41246 11442 41298 11454
rect 19966 11394 20018 11406
rect 14914 11342 14926 11394
rect 14978 11342 14990 11394
rect 18274 11342 18286 11394
rect 18338 11342 18350 11394
rect 18834 11342 18846 11394
rect 18898 11342 18910 11394
rect 19966 11330 20018 11342
rect 20414 11394 20466 11406
rect 22990 11394 23042 11406
rect 21858 11342 21870 11394
rect 21922 11342 21934 11394
rect 20414 11330 20466 11342
rect 22990 11330 23042 11342
rect 24334 11394 24386 11406
rect 24334 11330 24386 11342
rect 25230 11394 25282 11406
rect 25230 11330 25282 11342
rect 25678 11394 25730 11406
rect 25678 11330 25730 11342
rect 25790 11394 25842 11406
rect 25790 11330 25842 11342
rect 26014 11394 26066 11406
rect 26014 11330 26066 11342
rect 26238 11394 26290 11406
rect 26238 11330 26290 11342
rect 26686 11394 26738 11406
rect 26686 11330 26738 11342
rect 27806 11394 27858 11406
rect 27806 11330 27858 11342
rect 28366 11394 28418 11406
rect 28366 11330 28418 11342
rect 31166 11394 31218 11406
rect 31166 11330 31218 11342
rect 32510 11394 32562 11406
rect 33406 11394 33458 11406
rect 35646 11394 35698 11406
rect 33058 11342 33070 11394
rect 33122 11342 33134 11394
rect 34626 11342 34638 11394
rect 34690 11342 34702 11394
rect 34962 11342 34974 11394
rect 35026 11342 35038 11394
rect 32510 11330 32562 11342
rect 33406 11330 33458 11342
rect 35646 11330 35698 11342
rect 38110 11394 38162 11406
rect 38110 11330 38162 11342
rect 38894 11394 38946 11406
rect 38894 11330 38946 11342
rect 39118 11394 39170 11406
rect 39118 11330 39170 11342
rect 39902 11394 39954 11406
rect 39902 11330 39954 11342
rect 40014 11394 40066 11406
rect 40014 11330 40066 11342
rect 41134 11394 41186 11406
rect 41134 11330 41186 11342
rect 41358 11394 41410 11406
rect 41358 11330 41410 11342
rect 42254 11394 42306 11406
rect 42254 11330 42306 11342
rect 43374 11394 43426 11406
rect 43374 11330 43426 11342
rect 20638 11282 20690 11294
rect 20638 11218 20690 11230
rect 21422 11282 21474 11294
rect 21422 11218 21474 11230
rect 24222 11282 24274 11294
rect 24222 11218 24274 11230
rect 28030 11282 28082 11294
rect 28030 11218 28082 11230
rect 28590 11282 28642 11294
rect 28590 11218 28642 11230
rect 36094 11282 36146 11294
rect 36094 11218 36146 11230
rect 37102 11282 37154 11294
rect 37102 11218 37154 11230
rect 38558 11282 38610 11294
rect 38558 11218 38610 11230
rect 41694 11282 41746 11294
rect 41694 11218 41746 11230
rect 42590 11282 42642 11294
rect 43486 11282 43538 11294
rect 42690 11230 42702 11282
rect 42754 11230 42766 11282
rect 42590 11218 42642 11230
rect 43486 11218 43538 11230
rect 44942 11282 44994 11294
rect 44942 11218 44994 11230
rect 19406 11170 19458 11182
rect 20190 11170 20242 11182
rect 18050 11118 18062 11170
rect 18114 11118 18126 11170
rect 19058 11118 19070 11170
rect 19122 11118 19134 11170
rect 19730 11118 19742 11170
rect 19794 11118 19806 11170
rect 19406 11106 19458 11118
rect 20190 11106 20242 11118
rect 21310 11170 21362 11182
rect 21310 11106 21362 11118
rect 21534 11170 21586 11182
rect 21534 11106 21586 11118
rect 24894 11170 24946 11182
rect 27134 11170 27186 11182
rect 25666 11118 25678 11170
rect 25730 11118 25742 11170
rect 24894 11106 24946 11118
rect 27134 11106 27186 11118
rect 28142 11170 28194 11182
rect 28142 11106 28194 11118
rect 29150 11170 29202 11182
rect 29150 11106 29202 11118
rect 29262 11170 29314 11182
rect 29262 11106 29314 11118
rect 29374 11170 29426 11182
rect 29374 11106 29426 11118
rect 29598 11170 29650 11182
rect 29598 11106 29650 11118
rect 30718 11170 30770 11182
rect 30718 11106 30770 11118
rect 30942 11170 30994 11182
rect 30942 11106 30994 11118
rect 31054 11170 31106 11182
rect 35758 11170 35810 11182
rect 33730 11118 33742 11170
rect 33794 11118 33806 11170
rect 31054 11106 31106 11118
rect 35758 11106 35810 11118
rect 35870 11170 35922 11182
rect 35870 11106 35922 11118
rect 36990 11170 37042 11182
rect 36990 11106 37042 11118
rect 37662 11170 37714 11182
rect 37662 11106 37714 11118
rect 38670 11170 38722 11182
rect 38670 11106 38722 11118
rect 39566 11170 39618 11182
rect 39566 11106 39618 11118
rect 39790 11170 39842 11182
rect 39790 11106 39842 11118
rect 40574 11170 40626 11182
rect 40574 11106 40626 11118
rect 42478 11170 42530 11182
rect 42478 11106 42530 11118
rect 43598 11170 43650 11182
rect 43598 11106 43650 11118
rect 43822 11170 43874 11182
rect 43822 11106 43874 11118
rect 44830 11170 44882 11182
rect 44830 11106 44882 11118
rect 1344 11002 48608 11036
rect 1344 10950 19838 11002
rect 19890 10950 19942 11002
rect 19994 10950 20046 11002
rect 20098 10950 48608 11002
rect 1344 10916 48608 10950
rect 16046 10834 16098 10846
rect 16046 10770 16098 10782
rect 17614 10834 17666 10846
rect 17614 10770 17666 10782
rect 17950 10834 18002 10846
rect 17950 10770 18002 10782
rect 23662 10834 23714 10846
rect 23662 10770 23714 10782
rect 25342 10834 25394 10846
rect 25342 10770 25394 10782
rect 30158 10834 30210 10846
rect 30158 10770 30210 10782
rect 37998 10834 38050 10846
rect 37998 10770 38050 10782
rect 38446 10834 38498 10846
rect 38446 10770 38498 10782
rect 38894 10834 38946 10846
rect 38894 10770 38946 10782
rect 39454 10834 39506 10846
rect 39454 10770 39506 10782
rect 41470 10834 41522 10846
rect 41470 10770 41522 10782
rect 42254 10834 42306 10846
rect 42254 10770 42306 10782
rect 47518 10834 47570 10846
rect 47518 10770 47570 10782
rect 16270 10722 16322 10734
rect 16270 10658 16322 10670
rect 16606 10722 16658 10734
rect 16606 10658 16658 10670
rect 16830 10722 16882 10734
rect 24334 10722 24386 10734
rect 29486 10722 29538 10734
rect 19954 10670 19966 10722
rect 20018 10670 20030 10722
rect 26674 10670 26686 10722
rect 26738 10670 26750 10722
rect 16830 10658 16882 10670
rect 24334 10658 24386 10670
rect 29486 10658 29538 10670
rect 33182 10722 33234 10734
rect 33182 10658 33234 10670
rect 33518 10722 33570 10734
rect 39678 10722 39730 10734
rect 37650 10670 37662 10722
rect 37714 10670 37726 10722
rect 33518 10658 33570 10670
rect 39678 10658 39730 10670
rect 41918 10722 41970 10734
rect 41918 10658 41970 10670
rect 42030 10722 42082 10734
rect 43250 10670 43262 10722
rect 43314 10670 43326 10722
rect 42030 10658 42082 10670
rect 18062 10610 18114 10622
rect 18062 10546 18114 10558
rect 18174 10610 18226 10622
rect 23550 10610 23602 10622
rect 18498 10558 18510 10610
rect 18562 10558 18574 10610
rect 19170 10558 19182 10610
rect 19234 10558 19246 10610
rect 18174 10546 18226 10558
rect 23550 10546 23602 10558
rect 23886 10610 23938 10622
rect 23886 10546 23938 10558
rect 25454 10610 25506 10622
rect 29150 10610 29202 10622
rect 25890 10558 25902 10610
rect 25954 10558 25966 10610
rect 25454 10546 25506 10558
rect 29150 10546 29202 10558
rect 29710 10610 29762 10622
rect 29710 10546 29762 10558
rect 30046 10610 30098 10622
rect 30046 10546 30098 10558
rect 30270 10610 30322 10622
rect 30270 10546 30322 10558
rect 30718 10610 30770 10622
rect 30718 10546 30770 10558
rect 30830 10610 30882 10622
rect 30830 10546 30882 10558
rect 31278 10610 31330 10622
rect 31278 10546 31330 10558
rect 31390 10610 31442 10622
rect 31390 10546 31442 10558
rect 31950 10610 32002 10622
rect 40014 10610 40066 10622
rect 34402 10558 34414 10610
rect 34466 10558 34478 10610
rect 31950 10546 32002 10558
rect 40014 10546 40066 10558
rect 40238 10610 40290 10622
rect 40238 10546 40290 10558
rect 40798 10610 40850 10622
rect 40798 10546 40850 10558
rect 41246 10610 41298 10622
rect 41246 10546 41298 10558
rect 41358 10610 41410 10622
rect 42466 10558 42478 10610
rect 42530 10558 42542 10610
rect 41358 10546 41410 10558
rect 16382 10498 16434 10510
rect 22654 10498 22706 10510
rect 22082 10446 22094 10498
rect 22146 10446 22158 10498
rect 16382 10434 16434 10446
rect 22654 10434 22706 10446
rect 23102 10498 23154 10510
rect 29262 10498 29314 10510
rect 28802 10446 28814 10498
rect 28866 10446 28878 10498
rect 23102 10434 23154 10446
rect 29262 10434 29314 10446
rect 31054 10498 31106 10510
rect 39790 10498 39842 10510
rect 47630 10498 47682 10510
rect 35186 10446 35198 10498
rect 35250 10446 35262 10498
rect 37314 10446 37326 10498
rect 37378 10446 37390 10498
rect 45378 10446 45390 10498
rect 45442 10446 45454 10498
rect 31054 10434 31106 10446
rect 39790 10434 39842 10446
rect 47630 10434 47682 10446
rect 22542 10386 22594 10398
rect 22542 10322 22594 10334
rect 24110 10386 24162 10398
rect 24110 10322 24162 10334
rect 24446 10386 24498 10398
rect 24446 10322 24498 10334
rect 25342 10386 25394 10398
rect 25342 10322 25394 10334
rect 1344 10218 48608 10252
rect 1344 10166 4478 10218
rect 4530 10166 4582 10218
rect 4634 10166 4686 10218
rect 4738 10166 35198 10218
rect 35250 10166 35302 10218
rect 35354 10166 35406 10218
rect 35458 10166 48608 10218
rect 1344 10132 48608 10166
rect 25454 10050 25506 10062
rect 25454 9986 25506 9998
rect 25566 10050 25618 10062
rect 25566 9986 25618 9998
rect 18286 9938 18338 9950
rect 26126 9938 26178 9950
rect 15698 9886 15710 9938
rect 15762 9886 15774 9938
rect 17826 9886 17838 9938
rect 17890 9886 17902 9938
rect 22082 9886 22094 9938
rect 22146 9886 22158 9938
rect 24210 9886 24222 9938
rect 24274 9886 24286 9938
rect 24658 9886 24670 9938
rect 24722 9886 24734 9938
rect 18286 9874 18338 9886
rect 26126 9874 26178 9886
rect 27358 9938 27410 9950
rect 27358 9874 27410 9886
rect 28702 9938 28754 9950
rect 35310 9938 35362 9950
rect 32386 9886 32398 9938
rect 32450 9886 32462 9938
rect 28702 9874 28754 9886
rect 35310 9874 35362 9886
rect 36094 9938 36146 9950
rect 36094 9874 36146 9886
rect 36542 9938 36594 9950
rect 41246 9938 41298 9950
rect 37986 9886 37998 9938
rect 38050 9886 38062 9938
rect 40114 9886 40126 9938
rect 40178 9886 40190 9938
rect 36542 9874 36594 9886
rect 41246 9874 41298 9886
rect 41806 9938 41858 9950
rect 41806 9874 41858 9886
rect 45838 9938 45890 9950
rect 45838 9874 45890 9886
rect 26910 9826 26962 9838
rect 35086 9826 35138 9838
rect 15026 9774 15038 9826
rect 15090 9774 15102 9826
rect 21298 9774 21310 9826
rect 21362 9774 21374 9826
rect 29586 9774 29598 9826
rect 29650 9774 29662 9826
rect 34626 9774 34638 9826
rect 34690 9774 34702 9826
rect 34850 9774 34862 9826
rect 34914 9774 34926 9826
rect 26910 9762 26962 9774
rect 35086 9762 35138 9774
rect 35534 9826 35586 9838
rect 44830 9826 44882 9838
rect 37202 9774 37214 9826
rect 37266 9774 37278 9826
rect 42690 9774 42702 9826
rect 42754 9774 42766 9826
rect 43362 9774 43374 9826
rect 43426 9774 43438 9826
rect 43922 9774 43934 9826
rect 43986 9774 43998 9826
rect 35534 9762 35586 9774
rect 44830 9762 44882 9774
rect 45166 9826 45218 9838
rect 45166 9762 45218 9774
rect 24670 9714 24722 9726
rect 25230 9714 25282 9726
rect 40910 9714 40962 9726
rect 45390 9714 45442 9726
rect 24882 9662 24894 9714
rect 24946 9662 24958 9714
rect 26562 9662 26574 9714
rect 26626 9662 26638 9714
rect 30258 9662 30270 9714
rect 30322 9662 30334 9714
rect 44258 9662 44270 9714
rect 44322 9662 44334 9714
rect 24670 9650 24722 9662
rect 25230 9650 25282 9662
rect 40910 9650 40962 9662
rect 45390 9650 45442 9662
rect 47854 9714 47906 9726
rect 47854 9650 47906 9662
rect 48190 9714 48242 9726
rect 48190 9650 48242 9662
rect 42142 9602 42194 9614
rect 34962 9550 34974 9602
rect 35026 9550 35038 9602
rect 42142 9538 42194 9550
rect 42254 9602 42306 9614
rect 42254 9538 42306 9550
rect 42366 9602 42418 9614
rect 45278 9602 45330 9614
rect 43250 9550 43262 9602
rect 43314 9550 43326 9602
rect 42366 9538 42418 9550
rect 45278 9538 45330 9550
rect 47630 9602 47682 9614
rect 47630 9538 47682 9550
rect 1344 9434 48608 9468
rect 1344 9382 19838 9434
rect 19890 9382 19942 9434
rect 19994 9382 20046 9434
rect 20098 9382 48608 9434
rect 1344 9348 48608 9382
rect 18286 9266 18338 9278
rect 18286 9202 18338 9214
rect 19070 9266 19122 9278
rect 19070 9202 19122 9214
rect 19854 9266 19906 9278
rect 19854 9202 19906 9214
rect 21198 9266 21250 9278
rect 23662 9266 23714 9278
rect 23202 9214 23214 9266
rect 23266 9214 23278 9266
rect 21198 9202 21250 9214
rect 23662 9202 23714 9214
rect 24558 9266 24610 9278
rect 24558 9202 24610 9214
rect 35086 9266 35138 9278
rect 37326 9266 37378 9278
rect 35634 9214 35646 9266
rect 35698 9214 35710 9266
rect 35086 9202 35138 9214
rect 37326 9202 37378 9214
rect 39566 9266 39618 9278
rect 39566 9202 39618 9214
rect 18398 9154 18450 9166
rect 18398 9090 18450 9102
rect 20078 9154 20130 9166
rect 20078 9090 20130 9102
rect 20414 9154 20466 9166
rect 20414 9090 20466 9102
rect 20638 9154 20690 9166
rect 20638 9090 20690 9102
rect 21310 9154 21362 9166
rect 34078 9154 34130 9166
rect 27458 9102 27470 9154
rect 27522 9102 27534 9154
rect 21310 9090 21362 9102
rect 34078 9090 34130 9102
rect 34190 9154 34242 9166
rect 34190 9090 34242 9102
rect 38670 9154 38722 9166
rect 41682 9102 41694 9154
rect 41746 9102 41758 9154
rect 46610 9102 46622 9154
rect 46674 9102 46686 9154
rect 38670 9090 38722 9102
rect 17950 9042 18002 9054
rect 17950 8978 18002 8990
rect 18622 9042 18674 9054
rect 18622 8978 18674 8990
rect 21086 9042 21138 9054
rect 23438 9042 23490 9054
rect 21634 8990 21646 9042
rect 21698 8990 21710 9042
rect 22978 8990 22990 9042
rect 23042 8990 23054 9042
rect 21086 8978 21138 8990
rect 23438 8978 23490 8990
rect 23774 9042 23826 9054
rect 23774 8978 23826 8990
rect 24110 9042 24162 9054
rect 33182 9042 33234 9054
rect 26674 8990 26686 9042
rect 26738 8990 26750 9042
rect 24110 8978 24162 8990
rect 33182 8978 33234 8990
rect 33406 9042 33458 9054
rect 33406 8978 33458 8990
rect 33742 9042 33794 9054
rect 33742 8978 33794 8990
rect 33854 9042 33906 9054
rect 33854 8978 33906 8990
rect 34750 9042 34802 9054
rect 39006 9042 39058 9054
rect 35858 8990 35870 9042
rect 35922 8990 35934 9042
rect 41010 8990 41022 9042
rect 41074 8990 41086 9042
rect 47282 8990 47294 9042
rect 47346 8990 47358 9042
rect 34750 8978 34802 8990
rect 39006 8978 39058 8990
rect 20190 8930 20242 8942
rect 20190 8866 20242 8878
rect 25790 8930 25842 8942
rect 33518 8930 33570 8942
rect 29586 8878 29598 8930
rect 29650 8878 29662 8930
rect 37762 8878 37774 8930
rect 37826 8878 37838 8930
rect 43810 8878 43822 8930
rect 43874 8878 43886 8930
rect 44482 8878 44494 8930
rect 44546 8878 44558 8930
rect 25790 8866 25842 8878
rect 33518 8866 33570 8878
rect 24210 8766 24222 8818
rect 24274 8815 24286 8818
rect 24770 8815 24782 8818
rect 24274 8769 24782 8815
rect 24274 8766 24286 8769
rect 24770 8766 24782 8769
rect 24834 8766 24846 8818
rect 1344 8650 48608 8684
rect 1344 8598 4478 8650
rect 4530 8598 4582 8650
rect 4634 8598 4686 8650
rect 4738 8598 35198 8650
rect 35250 8598 35302 8650
rect 35354 8598 35406 8650
rect 35458 8598 48608 8650
rect 1344 8564 48608 8598
rect 25006 8482 25058 8494
rect 25006 8418 25058 8430
rect 43598 8482 43650 8494
rect 43598 8418 43650 8430
rect 44942 8482 44994 8494
rect 44942 8418 44994 8430
rect 45502 8482 45554 8494
rect 45502 8418 45554 8430
rect 18846 8370 18898 8382
rect 18162 8318 18174 8370
rect 18226 8318 18238 8370
rect 18846 8306 18898 8318
rect 19742 8370 19794 8382
rect 46062 8370 46114 8382
rect 31490 8318 31502 8370
rect 31554 8318 31566 8370
rect 33618 8318 33630 8370
rect 33682 8318 33694 8370
rect 19742 8306 19794 8318
rect 46062 8306 46114 8318
rect 18734 8258 18786 8270
rect 15362 8206 15374 8258
rect 15426 8206 15438 8258
rect 18734 8194 18786 8206
rect 18958 8258 19010 8270
rect 18958 8194 19010 8206
rect 23774 8258 23826 8270
rect 23774 8194 23826 8206
rect 23998 8258 24050 8270
rect 23998 8194 24050 8206
rect 24334 8258 24386 8270
rect 24334 8194 24386 8206
rect 24782 8258 24834 8270
rect 24782 8194 24834 8206
rect 25230 8258 25282 8270
rect 25230 8194 25282 8206
rect 25454 8258 25506 8270
rect 34638 8258 34690 8270
rect 39678 8258 39730 8270
rect 30258 8206 30270 8258
rect 30322 8206 30334 8258
rect 31154 8206 31166 8258
rect 31218 8206 31230 8258
rect 34402 8206 34414 8258
rect 34466 8206 34478 8258
rect 37538 8206 37550 8258
rect 37602 8206 37614 8258
rect 25454 8194 25506 8206
rect 34638 8194 34690 8206
rect 39678 8194 39730 8206
rect 42478 8258 42530 8270
rect 42478 8194 42530 8206
rect 43150 8258 43202 8270
rect 43150 8194 43202 8206
rect 43822 8258 43874 8270
rect 43822 8194 43874 8206
rect 44046 8258 44098 8270
rect 44046 8194 44098 8206
rect 44830 8258 44882 8270
rect 44830 8194 44882 8206
rect 45614 8258 45666 8270
rect 45614 8194 45666 8206
rect 19182 8146 19234 8158
rect 35086 8146 35138 8158
rect 16034 8094 16046 8146
rect 16098 8094 16110 8146
rect 26674 8094 26686 8146
rect 26738 8094 26750 8146
rect 30482 8094 30494 8146
rect 30546 8094 30558 8146
rect 19182 8082 19234 8094
rect 35086 8082 35138 8094
rect 35310 8146 35362 8158
rect 40238 8146 40290 8158
rect 35634 8094 35646 8146
rect 35698 8094 35710 8146
rect 37650 8094 37662 8146
rect 37714 8094 37726 8146
rect 35310 8082 35362 8094
rect 40238 8082 40290 8094
rect 42142 8146 42194 8158
rect 42142 8082 42194 8094
rect 42702 8146 42754 8158
rect 42702 8082 42754 8094
rect 44270 8146 44322 8158
rect 44270 8082 44322 8094
rect 44942 8146 44994 8158
rect 44942 8082 44994 8094
rect 23886 8034 23938 8046
rect 23886 7970 23938 7982
rect 25902 8034 25954 8046
rect 25902 7970 25954 7982
rect 27022 8034 27074 8046
rect 34862 8034 34914 8046
rect 31042 7982 31054 8034
rect 31106 7982 31118 8034
rect 27022 7970 27074 7982
rect 34862 7970 34914 7982
rect 35982 8034 36034 8046
rect 35982 7970 36034 7982
rect 36430 8034 36482 8046
rect 42254 8034 42306 8046
rect 41234 7982 41246 8034
rect 41298 7982 41310 8034
rect 36430 7970 36482 7982
rect 42254 7970 42306 7982
rect 45502 8034 45554 8046
rect 45502 7970 45554 7982
rect 1344 7866 48608 7900
rect 1344 7814 19838 7866
rect 19890 7814 19942 7866
rect 19994 7814 20046 7866
rect 20098 7814 48608 7866
rect 1344 7780 48608 7814
rect 16382 7698 16434 7710
rect 16382 7634 16434 7646
rect 17950 7698 18002 7710
rect 17950 7634 18002 7646
rect 18062 7698 18114 7710
rect 18062 7634 18114 7646
rect 27022 7698 27074 7710
rect 27022 7634 27074 7646
rect 33406 7698 33458 7710
rect 33406 7634 33458 7646
rect 35646 7698 35698 7710
rect 35646 7634 35698 7646
rect 37550 7698 37602 7710
rect 37550 7634 37602 7646
rect 38558 7698 38610 7710
rect 39902 7698 39954 7710
rect 38882 7646 38894 7698
rect 38946 7646 38958 7698
rect 38558 7634 38610 7646
rect 39902 7634 39954 7646
rect 45390 7698 45442 7710
rect 45390 7634 45442 7646
rect 16830 7586 16882 7598
rect 23662 7586 23714 7598
rect 19954 7534 19966 7586
rect 20018 7534 20030 7586
rect 16830 7522 16882 7534
rect 23662 7522 23714 7534
rect 27470 7586 27522 7598
rect 27470 7522 27522 7534
rect 28926 7586 28978 7598
rect 28926 7522 28978 7534
rect 33182 7586 33234 7598
rect 33182 7522 33234 7534
rect 33742 7586 33794 7598
rect 33742 7522 33794 7534
rect 34078 7586 34130 7598
rect 34078 7522 34130 7534
rect 34190 7586 34242 7598
rect 34190 7522 34242 7534
rect 34750 7586 34802 7598
rect 34750 7522 34802 7534
rect 34862 7586 34914 7598
rect 34862 7522 34914 7534
rect 35422 7586 35474 7598
rect 35422 7522 35474 7534
rect 36430 7586 36482 7598
rect 40014 7586 40066 7598
rect 37874 7534 37886 7586
rect 37938 7534 37950 7586
rect 36430 7522 36482 7534
rect 40014 7522 40066 7534
rect 42590 7586 42642 7598
rect 43486 7586 43538 7598
rect 42802 7534 42814 7586
rect 42866 7534 42878 7586
rect 42590 7522 42642 7534
rect 43486 7522 43538 7534
rect 16270 7474 16322 7486
rect 16270 7410 16322 7422
rect 16606 7474 16658 7486
rect 16606 7410 16658 7422
rect 18174 7474 18226 7486
rect 23886 7474 23938 7486
rect 18498 7422 18510 7474
rect 18562 7422 18574 7474
rect 19282 7422 19294 7474
rect 19346 7422 19358 7474
rect 18174 7410 18226 7422
rect 23886 7410 23938 7422
rect 24222 7474 24274 7486
rect 24222 7410 24274 7422
rect 25454 7474 25506 7486
rect 25454 7410 25506 7422
rect 27918 7474 27970 7486
rect 31054 7474 31106 7486
rect 30034 7422 30046 7474
rect 30098 7422 30110 7474
rect 27918 7410 27970 7422
rect 31054 7410 31106 7422
rect 31502 7474 31554 7486
rect 31502 7410 31554 7422
rect 31614 7474 31666 7486
rect 31614 7410 31666 7422
rect 31950 7474 32002 7486
rect 31950 7410 32002 7422
rect 32174 7474 32226 7486
rect 32174 7410 32226 7422
rect 33070 7474 33122 7486
rect 33070 7410 33122 7422
rect 34414 7474 34466 7486
rect 34414 7410 34466 7422
rect 34526 7474 34578 7486
rect 34526 7410 34578 7422
rect 35758 7474 35810 7486
rect 35758 7410 35810 7422
rect 35982 7474 36034 7486
rect 35982 7410 36034 7422
rect 36654 7474 36706 7486
rect 39566 7474 39618 7486
rect 38098 7422 38110 7474
rect 38162 7422 38174 7474
rect 36654 7410 36706 7422
rect 39566 7410 39618 7422
rect 40238 7474 40290 7486
rect 40238 7410 40290 7422
rect 41582 7474 41634 7486
rect 41582 7410 41634 7422
rect 41806 7474 41858 7486
rect 41806 7410 41858 7422
rect 42926 7474 42978 7486
rect 43710 7474 43762 7486
rect 43138 7422 43150 7474
rect 43202 7422 43214 7474
rect 42926 7410 42978 7422
rect 43710 7410 43762 7422
rect 44046 7474 44098 7486
rect 44046 7410 44098 7422
rect 17502 7362 17554 7374
rect 22542 7362 22594 7374
rect 22082 7310 22094 7362
rect 22146 7310 22158 7362
rect 17502 7298 17554 7310
rect 22542 7298 22594 7310
rect 23774 7362 23826 7374
rect 23774 7298 23826 7310
rect 30382 7362 30434 7374
rect 30382 7298 30434 7310
rect 31838 7362 31890 7374
rect 31838 7298 31890 7310
rect 43598 7362 43650 7374
rect 43598 7298 43650 7310
rect 44494 7362 44546 7374
rect 44494 7298 44546 7310
rect 44942 7362 44994 7374
rect 44942 7298 44994 7310
rect 30606 7250 30658 7262
rect 30606 7186 30658 7198
rect 30830 7250 30882 7262
rect 30830 7186 30882 7198
rect 36878 7250 36930 7262
rect 36878 7186 36930 7198
rect 37102 7250 37154 7262
rect 42142 7250 42194 7262
rect 41234 7198 41246 7250
rect 41298 7198 41310 7250
rect 37102 7186 37154 7198
rect 42142 7186 42194 7198
rect 42254 7250 42306 7262
rect 42254 7186 42306 7198
rect 1344 7082 48608 7116
rect 1344 7030 4478 7082
rect 4530 7030 4582 7082
rect 4634 7030 4686 7082
rect 4738 7030 35198 7082
rect 35250 7030 35302 7082
rect 35354 7030 35406 7082
rect 35458 7030 48608 7082
rect 1344 6996 48608 7030
rect 22766 6914 22818 6926
rect 22766 6850 22818 6862
rect 25790 6914 25842 6926
rect 25790 6850 25842 6862
rect 31390 6914 31442 6926
rect 31390 6850 31442 6862
rect 34638 6914 34690 6926
rect 34638 6850 34690 6862
rect 42366 6914 42418 6926
rect 42366 6850 42418 6862
rect 42478 6914 42530 6926
rect 42478 6850 42530 6862
rect 24334 6802 24386 6814
rect 34414 6802 34466 6814
rect 19282 6750 19294 6802
rect 19346 6750 19358 6802
rect 25106 6750 25118 6802
rect 25170 6750 25182 6802
rect 24334 6738 24386 6750
rect 34414 6738 34466 6750
rect 35646 6802 35698 6814
rect 35646 6738 35698 6750
rect 40686 6802 40738 6814
rect 40686 6738 40738 6750
rect 41918 6802 41970 6814
rect 43362 6750 43374 6802
rect 43426 6750 43438 6802
rect 44818 6750 44830 6802
rect 44882 6750 44894 6802
rect 41918 6738 41970 6750
rect 19742 6690 19794 6702
rect 16482 6638 16494 6690
rect 16546 6638 16558 6690
rect 17154 6638 17166 6690
rect 17218 6638 17230 6690
rect 19742 6626 19794 6638
rect 20302 6690 20354 6702
rect 20302 6626 20354 6638
rect 21982 6690 22034 6702
rect 21982 6626 22034 6638
rect 22990 6690 23042 6702
rect 22990 6626 23042 6638
rect 23886 6690 23938 6702
rect 23886 6626 23938 6638
rect 24222 6690 24274 6702
rect 25566 6690 25618 6702
rect 27022 6690 27074 6702
rect 24882 6638 24894 6690
rect 24946 6638 24958 6690
rect 25218 6638 25230 6690
rect 25282 6638 25294 6690
rect 26114 6638 26126 6690
rect 26178 6638 26190 6690
rect 24222 6626 24274 6638
rect 25566 6626 25618 6638
rect 27022 6626 27074 6638
rect 27470 6690 27522 6702
rect 27470 6626 27522 6638
rect 27694 6690 27746 6702
rect 27694 6626 27746 6638
rect 28366 6690 28418 6702
rect 28366 6626 28418 6638
rect 28590 6690 28642 6702
rect 28590 6626 28642 6638
rect 29038 6690 29090 6702
rect 29038 6626 29090 6638
rect 29262 6690 29314 6702
rect 29262 6626 29314 6638
rect 29486 6690 29538 6702
rect 29486 6626 29538 6638
rect 30046 6690 30098 6702
rect 30046 6626 30098 6638
rect 31614 6690 31666 6702
rect 31614 6626 31666 6638
rect 31950 6690 32002 6702
rect 31950 6626 32002 6638
rect 32174 6690 32226 6702
rect 32174 6626 32226 6638
rect 33182 6690 33234 6702
rect 35870 6690 35922 6702
rect 35298 6638 35310 6690
rect 35362 6638 35374 6690
rect 33182 6626 33234 6638
rect 35870 6626 35922 6638
rect 37326 6690 37378 6702
rect 37326 6626 37378 6638
rect 37998 6690 38050 6702
rect 37998 6626 38050 6638
rect 40126 6690 40178 6702
rect 40126 6626 40178 6638
rect 40462 6690 40514 6702
rect 41806 6690 41858 6702
rect 41458 6638 41470 6690
rect 41522 6638 41534 6690
rect 40462 6626 40514 6638
rect 41806 6626 41858 6638
rect 42030 6690 42082 6702
rect 43262 6690 43314 6702
rect 43026 6638 43038 6690
rect 43090 6638 43102 6690
rect 42030 6626 42082 6638
rect 43262 6626 43314 6638
rect 43822 6690 43874 6702
rect 47618 6638 47630 6690
rect 47682 6638 47694 6690
rect 43822 6626 43874 6638
rect 24670 6578 24722 6590
rect 24670 6514 24722 6526
rect 29710 6578 29762 6590
rect 29710 6514 29762 6526
rect 30270 6578 30322 6590
rect 34862 6578 34914 6590
rect 31042 6526 31054 6578
rect 31106 6526 31118 6578
rect 30270 6514 30322 6526
rect 34862 6514 34914 6526
rect 37550 6578 37602 6590
rect 37550 6514 37602 6526
rect 37774 6578 37826 6590
rect 37774 6514 37826 6526
rect 38782 6578 38834 6590
rect 38782 6514 38834 6526
rect 44158 6578 44210 6590
rect 44158 6514 44210 6526
rect 44270 6578 44322 6590
rect 46946 6526 46958 6578
rect 47010 6526 47022 6578
rect 44270 6514 44322 6526
rect 21534 6466 21586 6478
rect 21534 6402 21586 6414
rect 22094 6466 22146 6478
rect 23438 6466 23490 6478
rect 22418 6414 22430 6466
rect 22482 6414 22494 6466
rect 22094 6402 22146 6414
rect 23438 6402 23490 6414
rect 23662 6466 23714 6478
rect 23662 6402 23714 6414
rect 23774 6466 23826 6478
rect 23774 6402 23826 6414
rect 27358 6466 27410 6478
rect 30158 6466 30210 6478
rect 28018 6414 28030 6466
rect 28082 6414 28094 6466
rect 27358 6402 27410 6414
rect 30158 6402 30210 6414
rect 30494 6466 30546 6478
rect 30494 6402 30546 6414
rect 32062 6466 32114 6478
rect 32062 6402 32114 6414
rect 32398 6466 32450 6478
rect 34750 6466 34802 6478
rect 32834 6414 32846 6466
rect 32898 6414 32910 6466
rect 32398 6402 32450 6414
rect 34750 6402 34802 6414
rect 36542 6466 36594 6478
rect 36542 6402 36594 6414
rect 38334 6466 38386 6478
rect 38334 6402 38386 6414
rect 38558 6466 38610 6478
rect 38558 6402 38610 6414
rect 38670 6466 38722 6478
rect 38670 6402 38722 6414
rect 39678 6466 39730 6478
rect 39678 6402 39730 6414
rect 39902 6466 39954 6478
rect 39902 6402 39954 6414
rect 40014 6466 40066 6478
rect 42814 6466 42866 6478
rect 41010 6414 41022 6466
rect 41074 6414 41086 6466
rect 40014 6402 40066 6414
rect 42814 6402 42866 6414
rect 1344 6298 48608 6332
rect 1344 6246 19838 6298
rect 19890 6246 19942 6298
rect 19994 6246 20046 6298
rect 20098 6246 48608 6298
rect 1344 6212 48608 6246
rect 18398 6130 18450 6142
rect 18398 6066 18450 6078
rect 20638 6130 20690 6142
rect 20638 6066 20690 6078
rect 24670 6130 24722 6142
rect 24670 6066 24722 6078
rect 27918 6130 27970 6142
rect 27918 6066 27970 6078
rect 32622 6130 32674 6142
rect 33058 6078 33070 6130
rect 33122 6078 33134 6130
rect 42242 6078 42254 6130
rect 42306 6078 42318 6130
rect 32622 6066 32674 6078
rect 19518 6018 19570 6030
rect 19518 5954 19570 5966
rect 19854 6018 19906 6030
rect 26686 6018 26738 6030
rect 27246 6018 27298 6030
rect 29598 6018 29650 6030
rect 31502 6018 31554 6030
rect 22082 5966 22094 6018
rect 22146 5966 22158 6018
rect 27010 5966 27022 6018
rect 27074 5966 27086 6018
rect 29250 5966 29262 6018
rect 29314 5966 29326 6018
rect 31266 5966 31278 6018
rect 31330 5966 31342 6018
rect 19854 5954 19906 5966
rect 26686 5954 26738 5966
rect 27246 5954 27298 5966
rect 29598 5954 29650 5966
rect 31502 5954 31554 5966
rect 33742 6018 33794 6030
rect 33742 5954 33794 5966
rect 34078 6018 34130 6030
rect 34078 5954 34130 5966
rect 34974 6018 35026 6030
rect 34974 5954 35026 5966
rect 35534 6018 35586 6030
rect 35534 5954 35586 5966
rect 36318 6018 36370 6030
rect 36318 5954 36370 5966
rect 37438 6018 37490 6030
rect 37438 5954 37490 5966
rect 37774 6018 37826 6030
rect 37774 5954 37826 5966
rect 38222 6018 38274 6030
rect 38222 5954 38274 5966
rect 38670 6018 38722 6030
rect 38670 5954 38722 5966
rect 41246 6018 41298 6030
rect 41570 5966 41582 6018
rect 41634 5966 41646 6018
rect 41246 5954 41298 5966
rect 18622 5906 18674 5918
rect 18622 5842 18674 5854
rect 18846 5906 18898 5918
rect 18846 5842 18898 5854
rect 19294 5906 19346 5918
rect 19294 5842 19346 5854
rect 19966 5906 20018 5918
rect 19966 5842 20018 5854
rect 20414 5906 20466 5918
rect 20414 5842 20466 5854
rect 20526 5906 20578 5918
rect 26014 5906 26066 5918
rect 20962 5854 20974 5906
rect 21026 5854 21038 5906
rect 21298 5854 21310 5906
rect 21362 5854 21374 5906
rect 20526 5842 20578 5854
rect 26014 5842 26066 5854
rect 27134 5906 27186 5918
rect 27134 5842 27186 5854
rect 27694 5906 27746 5918
rect 27694 5842 27746 5854
rect 28366 5906 28418 5918
rect 28366 5842 28418 5854
rect 29038 5906 29090 5918
rect 29038 5842 29090 5854
rect 29150 5906 29202 5918
rect 29150 5842 29202 5854
rect 29822 5906 29874 5918
rect 29822 5842 29874 5854
rect 29934 5906 29986 5918
rect 29934 5842 29986 5854
rect 31054 5906 31106 5918
rect 31054 5842 31106 5854
rect 31166 5906 31218 5918
rect 31166 5842 31218 5854
rect 31838 5906 31890 5918
rect 31838 5842 31890 5854
rect 31950 5906 32002 5918
rect 31950 5842 32002 5854
rect 33406 5906 33458 5918
rect 33406 5842 33458 5854
rect 34638 5906 34690 5918
rect 34638 5842 34690 5854
rect 34750 5906 34802 5918
rect 35422 5906 35474 5918
rect 35298 5854 35310 5906
rect 35362 5854 35374 5906
rect 34750 5842 34802 5854
rect 35422 5842 35474 5854
rect 36094 5906 36146 5918
rect 36766 5906 36818 5918
rect 39006 5906 39058 5918
rect 36642 5854 36654 5906
rect 36706 5854 36718 5906
rect 36978 5854 36990 5906
rect 37042 5854 37054 5906
rect 38434 5854 38446 5906
rect 38498 5854 38510 5906
rect 36094 5842 36146 5854
rect 36766 5842 36818 5854
rect 39006 5842 39058 5854
rect 39118 5906 39170 5918
rect 39790 5906 39842 5918
rect 39442 5854 39454 5906
rect 39506 5854 39518 5906
rect 39118 5842 39170 5854
rect 39790 5842 39842 5854
rect 40014 5906 40066 5918
rect 40014 5842 40066 5854
rect 40910 5906 40962 5918
rect 40910 5842 40962 5854
rect 41022 5906 41074 5918
rect 41022 5842 41074 5854
rect 41806 5906 41858 5918
rect 41806 5842 41858 5854
rect 42590 5906 42642 5918
rect 42590 5842 42642 5854
rect 42814 5906 42866 5918
rect 42814 5842 42866 5854
rect 19070 5794 19122 5806
rect 19070 5730 19122 5742
rect 19630 5794 19682 5806
rect 26350 5794 26402 5806
rect 24210 5742 24222 5794
rect 24274 5742 24286 5794
rect 25442 5742 25454 5794
rect 25506 5742 25518 5794
rect 19630 5730 19682 5742
rect 26350 5730 26402 5742
rect 27806 5794 27858 5806
rect 38098 5742 38110 5794
rect 38162 5742 38174 5794
rect 41906 5742 41918 5794
rect 41970 5742 41982 5794
rect 27806 5730 27858 5742
rect 25790 5682 25842 5694
rect 25790 5618 25842 5630
rect 26462 5682 26514 5694
rect 26462 5618 26514 5630
rect 35982 5682 36034 5694
rect 35982 5618 36034 5630
rect 1344 5514 48608 5548
rect 1344 5462 4478 5514
rect 4530 5462 4582 5514
rect 4634 5462 4686 5514
rect 4738 5462 35198 5514
rect 35250 5462 35302 5514
rect 35354 5462 35406 5514
rect 35458 5462 48608 5514
rect 1344 5428 48608 5462
rect 24222 5346 24274 5358
rect 41458 5294 41470 5346
rect 41522 5343 41534 5346
rect 41794 5343 41806 5346
rect 41522 5297 41806 5343
rect 41522 5294 41534 5297
rect 41794 5294 41806 5297
rect 41858 5294 41870 5346
rect 24222 5282 24274 5294
rect 21422 5234 21474 5246
rect 18610 5182 18622 5234
rect 18674 5182 18686 5234
rect 20738 5182 20750 5234
rect 20802 5182 20814 5234
rect 21422 5170 21474 5182
rect 22318 5234 22370 5246
rect 29262 5234 29314 5246
rect 33518 5234 33570 5246
rect 24994 5182 25006 5234
rect 25058 5182 25070 5234
rect 28354 5182 28366 5234
rect 28418 5182 28430 5234
rect 32722 5182 32734 5234
rect 32786 5182 32798 5234
rect 22318 5170 22370 5182
rect 29262 5170 29314 5182
rect 33518 5170 33570 5182
rect 36318 5234 36370 5246
rect 36318 5170 36370 5182
rect 37214 5234 37266 5246
rect 37214 5170 37266 5182
rect 37438 5234 37490 5246
rect 41134 5234 41186 5246
rect 37874 5182 37886 5234
rect 37938 5182 37950 5234
rect 37438 5170 37490 5182
rect 41134 5170 41186 5182
rect 41694 5234 41746 5246
rect 41694 5170 41746 5182
rect 42814 5234 42866 5246
rect 42814 5170 42866 5182
rect 44046 5234 44098 5246
rect 44046 5170 44098 5182
rect 23326 5122 23378 5134
rect 17938 5070 17950 5122
rect 18002 5070 18014 5122
rect 21858 5070 21870 5122
rect 21922 5070 21934 5122
rect 23326 5058 23378 5070
rect 23438 5122 23490 5134
rect 24110 5122 24162 5134
rect 33182 5122 33234 5134
rect 23762 5070 23774 5122
rect 23826 5070 23838 5122
rect 25106 5070 25118 5122
rect 25170 5070 25182 5122
rect 25554 5070 25566 5122
rect 25618 5070 25630 5122
rect 29922 5070 29934 5122
rect 29986 5070 29998 5122
rect 23438 5058 23490 5070
rect 24110 5058 24162 5070
rect 33182 5058 33234 5070
rect 35422 5122 35474 5134
rect 35422 5058 35474 5070
rect 35534 5122 35586 5134
rect 35534 5058 35586 5070
rect 37550 5122 37602 5134
rect 40002 5070 40014 5122
rect 40066 5070 40078 5122
rect 40786 5070 40798 5122
rect 40850 5070 40862 5122
rect 37550 5058 37602 5070
rect 21310 5010 21362 5022
rect 21310 4946 21362 4958
rect 21534 5010 21586 5022
rect 21534 4946 21586 4958
rect 23214 5010 23266 5022
rect 23214 4946 23266 4958
rect 24558 5010 24610 5022
rect 29150 5010 29202 5022
rect 35646 5010 35698 5022
rect 24770 4958 24782 5010
rect 24834 4958 24846 5010
rect 26226 4958 26238 5010
rect 26290 4958 26302 5010
rect 30594 4958 30606 5010
rect 30658 4958 30670 5010
rect 24558 4946 24610 4958
rect 29150 4946 29202 4958
rect 35646 4946 35698 4958
rect 33630 4898 33682 4910
rect 33630 4834 33682 4846
rect 35870 4898 35922 4910
rect 35870 4834 35922 4846
rect 36430 4898 36482 4910
rect 36430 4834 36482 4846
rect 41246 4898 41298 4910
rect 41246 4834 41298 4846
rect 42926 4898 42978 4910
rect 42926 4834 42978 4846
rect 1344 4730 48608 4764
rect 1344 4678 19838 4730
rect 19890 4678 19942 4730
rect 19994 4678 20046 4730
rect 20098 4678 48608 4730
rect 1344 4644 48608 4678
rect 25342 4562 25394 4574
rect 25342 4498 25394 4510
rect 26574 4562 26626 4574
rect 26574 4498 26626 4510
rect 31054 4562 31106 4574
rect 39890 4510 39902 4562
rect 39954 4510 39966 4562
rect 31054 4498 31106 4510
rect 26686 4450 26738 4462
rect 31166 4450 31218 4462
rect 19058 4398 19070 4450
rect 19122 4398 19134 4450
rect 28130 4398 28142 4450
rect 28194 4398 28206 4450
rect 33842 4398 33854 4450
rect 33906 4398 33918 4450
rect 38434 4398 38446 4450
rect 38498 4398 38510 4450
rect 41682 4398 41694 4450
rect 41746 4398 41758 4450
rect 46274 4398 46286 4450
rect 46338 4398 46350 4450
rect 26686 4386 26738 4398
rect 31166 4386 31218 4398
rect 47630 4338 47682 4350
rect 18274 4286 18286 4338
rect 18338 4286 18350 4338
rect 21634 4286 21646 4338
rect 21698 4286 21710 4338
rect 27346 4286 27358 4338
rect 27410 4286 27422 4338
rect 33170 4286 33182 4338
rect 33234 4286 33246 4338
rect 39218 4286 39230 4338
rect 39282 4286 39294 4338
rect 40114 4286 40126 4338
rect 40178 4286 40190 4338
rect 40898 4286 40910 4338
rect 40962 4286 40974 4338
rect 47058 4286 47070 4338
rect 47122 4286 47134 4338
rect 47630 4274 47682 4286
rect 48190 4338 48242 4350
rect 48190 4274 48242 4286
rect 21186 4174 21198 4226
rect 21250 4174 21262 4226
rect 22306 4174 22318 4226
rect 22370 4174 22382 4226
rect 24434 4174 24446 4226
rect 24498 4174 24510 4226
rect 30258 4174 30270 4226
rect 30322 4174 30334 4226
rect 35970 4174 35982 4226
rect 36034 4174 36046 4226
rect 36306 4174 36318 4226
rect 36370 4174 36382 4226
rect 43810 4174 43822 4226
rect 43874 4174 43886 4226
rect 44146 4174 44158 4226
rect 44210 4174 44222 4226
rect 1344 3946 48608 3980
rect 1344 3894 4478 3946
rect 4530 3894 4582 3946
rect 4634 3894 4686 3946
rect 4738 3894 35198 3946
rect 35250 3894 35302 3946
rect 35354 3894 35406 3946
rect 35458 3894 48608 3946
rect 1344 3860 48608 3894
rect 22766 3778 22818 3790
rect 22766 3714 22818 3726
rect 21534 3666 21586 3678
rect 21534 3602 21586 3614
rect 22878 3666 22930 3678
rect 22878 3602 22930 3614
rect 36318 3666 36370 3678
rect 36318 3602 36370 3614
rect 40014 3666 40066 3678
rect 40014 3602 40066 3614
rect 43934 3666 43986 3678
rect 43934 3602 43986 3614
rect 48302 3666 48354 3678
rect 48302 3602 48354 3614
rect 1344 3162 48608 3196
rect 1344 3110 19838 3162
rect 19890 3110 19942 3162
rect 19994 3110 20046 3162
rect 20098 3110 48608 3162
rect 1344 3076 48608 3110
<< via1 >>
rect 13470 57038 13522 57090
rect 14590 57038 14642 57090
rect 27134 57038 27186 57090
rect 28366 57038 28418 57090
rect 19838 56422 19890 56474
rect 19942 56422 19994 56474
rect 20046 56422 20098 56474
rect 3838 56254 3890 56306
rect 5518 56254 5570 56306
rect 6974 56254 7026 56306
rect 8542 56254 8594 56306
rect 10110 56254 10162 56306
rect 11678 56254 11730 56306
rect 12574 56254 12626 56306
rect 13470 56254 13522 56306
rect 15374 56254 15426 56306
rect 22094 56254 22146 56306
rect 27470 56254 27522 56306
rect 28366 56254 28418 56306
rect 40798 56254 40850 56306
rect 44606 56254 44658 56306
rect 47406 56254 47458 56306
rect 25342 56142 25394 56194
rect 42814 56142 42866 56194
rect 16046 56030 16098 56082
rect 16942 56030 16994 56082
rect 21086 56030 21138 56082
rect 27134 56030 27186 56082
rect 31614 56030 31666 56082
rect 35086 56030 35138 56082
rect 38782 56030 38834 56082
rect 39790 56030 39842 56082
rect 43822 56030 43874 56082
rect 46846 56030 46898 56082
rect 47630 56030 47682 56082
rect 47854 56030 47906 56082
rect 48190 56030 48242 56082
rect 17726 55918 17778 55970
rect 19854 55918 19906 55970
rect 30158 55918 30210 55970
rect 32174 55918 32226 55970
rect 34302 55918 34354 55970
rect 35982 55918 36034 55970
rect 38110 55918 38162 55970
rect 42926 55918 42978 55970
rect 43038 55806 43090 55858
rect 46510 55806 46562 55858
rect 46846 55806 46898 55858
rect 47630 55806 47682 55858
rect 4478 55638 4530 55690
rect 4582 55638 4634 55690
rect 4686 55638 4738 55690
rect 35198 55638 35250 55690
rect 35302 55638 35354 55690
rect 35406 55638 35458 55690
rect 22206 55470 22258 55522
rect 17502 55358 17554 55410
rect 20750 55358 20802 55410
rect 27022 55358 27074 55410
rect 32846 55358 32898 55410
rect 34190 55358 34242 55410
rect 42030 55358 42082 55410
rect 43598 55358 43650 55410
rect 45278 55358 45330 55410
rect 47406 55358 47458 55410
rect 9662 55246 9714 55298
rect 9886 55246 9938 55298
rect 10782 55246 10834 55298
rect 13806 55246 13858 55298
rect 14590 55246 14642 55298
rect 17950 55246 18002 55298
rect 22878 55246 22930 55298
rect 23438 55246 23490 55298
rect 24110 55246 24162 55298
rect 30046 55246 30098 55298
rect 33182 55246 33234 55298
rect 36878 55246 36930 55298
rect 37214 55246 37266 55298
rect 37998 55246 38050 55298
rect 38446 55246 38498 55298
rect 39118 55246 39170 55298
rect 42702 55246 42754 55298
rect 43374 55246 43426 55298
rect 44046 55246 44098 55298
rect 48078 55246 48130 55298
rect 9326 55134 9378 55186
rect 10110 55134 10162 55186
rect 11678 55134 11730 55186
rect 13470 55134 13522 55186
rect 14030 55134 14082 55186
rect 15374 55134 15426 55186
rect 18622 55134 18674 55186
rect 21870 55134 21922 55186
rect 22318 55134 22370 55186
rect 23102 55134 23154 55186
rect 23774 55134 23826 55186
rect 24894 55134 24946 55186
rect 27582 55134 27634 55186
rect 28030 55134 28082 55186
rect 28366 55134 28418 55186
rect 28590 55134 28642 55186
rect 29150 55134 29202 55186
rect 30718 55134 30770 55186
rect 36206 55134 36258 55186
rect 36318 55134 36370 55186
rect 37550 55134 37602 55186
rect 39902 55134 39954 55186
rect 43038 55134 43090 55186
rect 44942 55134 44994 55186
rect 9438 55022 9490 55074
rect 10894 55022 10946 55074
rect 11454 55022 11506 55074
rect 11566 55022 11618 55074
rect 12238 55022 12290 55074
rect 13694 55022 13746 55074
rect 22206 55022 22258 55074
rect 22542 55022 22594 55074
rect 22654 55022 22706 55074
rect 23662 55022 23714 55074
rect 27246 55022 27298 55074
rect 27470 55022 27522 55074
rect 28254 55022 28306 55074
rect 36542 55022 36594 55074
rect 37102 55022 37154 55074
rect 42478 55022 42530 55074
rect 42590 55022 42642 55074
rect 43710 55022 43762 55074
rect 44270 55022 44322 55074
rect 44830 55022 44882 55074
rect 19838 54854 19890 54906
rect 19942 54854 19994 54906
rect 20046 54854 20098 54906
rect 11678 54686 11730 54738
rect 18622 54686 18674 54738
rect 39342 54686 39394 54738
rect 40238 54686 40290 54738
rect 41246 54686 41298 54738
rect 45726 54686 45778 54738
rect 48190 54686 48242 54738
rect 6862 54574 6914 54626
rect 9886 54574 9938 54626
rect 13918 54574 13970 54626
rect 30158 54574 30210 54626
rect 37102 54574 37154 54626
rect 41022 54574 41074 54626
rect 43598 54574 43650 54626
rect 6190 54462 6242 54514
rect 10334 54462 10386 54514
rect 11118 54462 11170 54514
rect 12798 54462 12850 54514
rect 13134 54462 13186 54514
rect 19070 54462 19122 54514
rect 22542 54462 22594 54514
rect 23886 54462 23938 54514
rect 25790 54462 25842 54514
rect 27134 54462 27186 54514
rect 30942 54462 30994 54514
rect 35870 54462 35922 54514
rect 38670 54462 38722 54514
rect 39230 54462 39282 54514
rect 39454 54462 39506 54514
rect 39678 54462 39730 54514
rect 40910 54462 40962 54514
rect 44270 54462 44322 54514
rect 44718 54462 44770 54514
rect 47854 54462 47906 54514
rect 8990 54350 9042 54402
rect 12574 54350 12626 54402
rect 16046 54350 16098 54402
rect 16494 54350 16546 54402
rect 17726 54350 17778 54402
rect 18286 54350 18338 54402
rect 18734 54350 18786 54402
rect 19854 54350 19906 54402
rect 21982 54350 22034 54402
rect 22654 54350 22706 54402
rect 25454 54350 25506 54402
rect 26238 54350 26290 54402
rect 26910 54350 26962 54402
rect 27694 54350 27746 54402
rect 28030 54350 28082 54402
rect 31390 54350 31442 54402
rect 31838 54350 31890 54402
rect 32510 54350 32562 54402
rect 33070 54350 33122 54402
rect 35198 54350 35250 54402
rect 40350 54350 40402 54402
rect 41470 54350 41522 54402
rect 12462 54238 12514 54290
rect 24110 54238 24162 54290
rect 4478 54070 4530 54122
rect 4582 54070 4634 54122
rect 4686 54070 4738 54122
rect 35198 54070 35250 54122
rect 35302 54070 35354 54122
rect 35406 54070 35458 54122
rect 10334 53902 10386 53954
rect 16046 53902 16098 53954
rect 22990 53902 23042 53954
rect 23326 53902 23378 53954
rect 9662 53790 9714 53842
rect 10222 53790 10274 53842
rect 14030 53790 14082 53842
rect 21870 53790 21922 53842
rect 24222 53790 24274 53842
rect 25118 53790 25170 53842
rect 27694 53790 27746 53842
rect 29262 53790 29314 53842
rect 41358 53790 41410 53842
rect 45278 53790 45330 53842
rect 9998 53678 10050 53730
rect 12238 53678 12290 53730
rect 14702 53678 14754 53730
rect 16046 53678 16098 53730
rect 17950 53678 18002 53730
rect 22206 53678 22258 53730
rect 24334 53678 24386 53730
rect 24782 53678 24834 53730
rect 25342 53678 25394 53730
rect 25566 53678 25618 53730
rect 26014 53678 26066 53730
rect 26126 53678 26178 53730
rect 27246 53678 27298 53730
rect 28030 53678 28082 53730
rect 29150 53678 29202 53730
rect 32958 53678 33010 53730
rect 33630 53678 33682 53730
rect 37214 53678 37266 53730
rect 37326 53678 37378 53730
rect 37662 53678 37714 53730
rect 38446 53678 38498 53730
rect 39230 53678 39282 53730
rect 41694 53678 41746 53730
rect 44942 53678 44994 53730
rect 47406 53678 47458 53730
rect 48078 53678 48130 53730
rect 9550 53566 9602 53618
rect 10894 53566 10946 53618
rect 12462 53566 12514 53618
rect 14142 53566 14194 53618
rect 14926 53566 14978 53618
rect 15038 53566 15090 53618
rect 16382 53566 16434 53618
rect 22094 53566 22146 53618
rect 22430 53566 22482 53618
rect 23774 53566 23826 53618
rect 25006 53566 25058 53618
rect 27582 53566 27634 53618
rect 28254 53566 28306 53618
rect 28366 53566 28418 53618
rect 30830 53566 30882 53618
rect 31054 53566 31106 53618
rect 31390 53566 31442 53618
rect 37438 53566 37490 53618
rect 9214 53454 9266 53506
rect 11006 53454 11058 53506
rect 13582 53454 13634 53506
rect 13918 53454 13970 53506
rect 14366 53454 14418 53506
rect 15598 53454 15650 53506
rect 18958 53454 19010 53506
rect 21646 53454 21698 53506
rect 22654 53454 22706 53506
rect 23102 53454 23154 53506
rect 24110 53454 24162 53506
rect 25902 53454 25954 53506
rect 26350 53454 26402 53506
rect 27022 53454 27074 53506
rect 27806 53454 27858 53506
rect 29374 53454 29426 53506
rect 29598 53454 29650 53506
rect 30270 53454 30322 53506
rect 31278 53454 31330 53506
rect 33294 53454 33346 53506
rect 34638 53454 34690 53506
rect 37102 53454 37154 53506
rect 38110 53454 38162 53506
rect 42702 53454 42754 53506
rect 19838 53286 19890 53338
rect 19942 53286 19994 53338
rect 20046 53286 20098 53338
rect 15822 53118 15874 53170
rect 16382 53118 16434 53170
rect 20526 53118 20578 53170
rect 22542 53118 22594 53170
rect 23214 53118 23266 53170
rect 23438 53118 23490 53170
rect 24222 53118 24274 53170
rect 25790 53118 25842 53170
rect 27470 53118 27522 53170
rect 37438 53118 37490 53170
rect 39006 53118 39058 53170
rect 39454 53118 39506 53170
rect 41918 53118 41970 53170
rect 45614 53118 45666 53170
rect 7422 53006 7474 53058
rect 12014 53006 12066 53058
rect 23102 53006 23154 53058
rect 29374 53006 29426 53058
rect 31726 53006 31778 53058
rect 34302 53006 34354 53058
rect 38222 53006 38274 53058
rect 4174 52894 4226 52946
rect 7198 52894 7250 52946
rect 7534 52894 7586 52946
rect 7982 52894 8034 52946
rect 11230 52894 11282 52946
rect 15374 52894 15426 52946
rect 15710 52894 15762 52946
rect 16046 52894 16098 52946
rect 16270 52894 16322 52946
rect 16494 52894 16546 52946
rect 16830 52894 16882 52946
rect 19630 52894 19682 52946
rect 22430 52894 22482 52946
rect 25342 52894 25394 52946
rect 29262 52894 29314 52946
rect 29598 52894 29650 52946
rect 31054 52894 31106 52946
rect 35198 52894 35250 52946
rect 36206 52894 36258 52946
rect 36766 52894 36818 52946
rect 36990 52894 37042 52946
rect 37662 52894 37714 52946
rect 37998 52894 38050 52946
rect 38894 52894 38946 52946
rect 40014 52894 40066 52946
rect 41358 52894 41410 52946
rect 44606 52894 44658 52946
rect 47966 52894 48018 52946
rect 4846 52782 4898 52834
rect 6974 52782 7026 52834
rect 14142 52782 14194 52834
rect 14590 52782 14642 52834
rect 17502 52782 17554 52834
rect 23774 52782 23826 52834
rect 30830 52782 30882 52834
rect 33854 52782 33906 52834
rect 35870 52782 35922 52834
rect 37550 52782 37602 52834
rect 43822 52782 43874 52834
rect 44158 52782 44210 52834
rect 47518 52782 47570 52834
rect 22542 52670 22594 52722
rect 23774 52670 23826 52722
rect 24110 52670 24162 52722
rect 4478 52502 4530 52554
rect 4582 52502 4634 52554
rect 4686 52502 4738 52554
rect 35198 52502 35250 52554
rect 35302 52502 35354 52554
rect 35406 52502 35458 52554
rect 6750 52334 6802 52386
rect 27358 52334 27410 52386
rect 38670 52334 38722 52386
rect 39678 52334 39730 52386
rect 46622 52334 46674 52386
rect 6078 52222 6130 52274
rect 7646 52222 7698 52274
rect 8206 52222 8258 52274
rect 8990 52222 9042 52274
rect 10334 52222 10386 52274
rect 11118 52222 11170 52274
rect 15486 52222 15538 52274
rect 25230 52222 25282 52274
rect 26798 52222 26850 52274
rect 31614 52222 31666 52274
rect 34750 52222 34802 52274
rect 35534 52222 35586 52274
rect 36430 52222 36482 52274
rect 38558 52222 38610 52274
rect 5966 52110 6018 52162
rect 6862 52110 6914 52162
rect 7198 52110 7250 52162
rect 9662 52110 9714 52162
rect 14030 52110 14082 52162
rect 17614 52110 17666 52162
rect 18286 52110 18338 52162
rect 20078 52110 20130 52162
rect 22318 52110 22370 52162
rect 22654 52110 22706 52162
rect 23326 52110 23378 52162
rect 23550 52110 23602 52162
rect 24222 52110 24274 52162
rect 26462 52110 26514 52162
rect 27246 52110 27298 52162
rect 29262 52110 29314 52162
rect 29486 52110 29538 52162
rect 30158 52110 30210 52162
rect 30830 52110 30882 52162
rect 31390 52110 31442 52162
rect 32286 52110 32338 52162
rect 32734 52110 32786 52162
rect 32958 52110 33010 52162
rect 35086 52110 35138 52162
rect 35646 52110 35698 52162
rect 37102 52110 37154 52162
rect 37438 52110 37490 52162
rect 38334 52110 38386 52162
rect 39118 52110 39170 52162
rect 40462 52110 40514 52162
rect 41246 52110 41298 52162
rect 41694 52110 41746 52162
rect 42478 52110 42530 52162
rect 44270 52110 44322 52162
rect 45614 52110 45666 52162
rect 5630 51998 5682 52050
rect 6190 51998 6242 52050
rect 9326 51998 9378 52050
rect 10446 51998 10498 52050
rect 10670 51998 10722 52050
rect 19630 51998 19682 52050
rect 19742 51998 19794 52050
rect 20414 51998 20466 52050
rect 25342 51998 25394 52050
rect 25566 51998 25618 52050
rect 33630 51998 33682 52050
rect 36990 51998 37042 52050
rect 39790 51998 39842 52050
rect 40238 51998 40290 52050
rect 42142 51998 42194 52050
rect 43486 51998 43538 52050
rect 43934 51998 43986 52050
rect 44830 51998 44882 52050
rect 6750 51886 6802 51938
rect 7534 51886 7586 51938
rect 7758 51886 7810 51938
rect 8094 51886 8146 51938
rect 9438 51886 9490 51938
rect 14142 51886 14194 51938
rect 14366 51886 14418 51938
rect 19406 51886 19458 51938
rect 20302 51886 20354 51938
rect 21310 51886 21362 51938
rect 21646 51886 21698 51938
rect 22766 51886 22818 51938
rect 22878 51886 22930 51938
rect 35422 51886 35474 51938
rect 40350 51886 40402 51938
rect 42926 51886 42978 51938
rect 44046 51886 44098 51938
rect 45166 51886 45218 51938
rect 19838 51718 19890 51770
rect 19942 51718 19994 51770
rect 20046 51718 20098 51770
rect 5630 51550 5682 51602
rect 5742 51550 5794 51602
rect 11454 51550 11506 51602
rect 14030 51550 14082 51602
rect 25566 51550 25618 51602
rect 28030 51550 28082 51602
rect 35534 51550 35586 51602
rect 35982 51550 36034 51602
rect 36094 51550 36146 51602
rect 37662 51550 37714 51602
rect 39230 51550 39282 51602
rect 39342 51550 39394 51602
rect 40126 51550 40178 51602
rect 44942 51550 44994 51602
rect 6862 51438 6914 51490
rect 9886 51438 9938 51490
rect 12126 51438 12178 51490
rect 20862 51438 20914 51490
rect 22206 51438 22258 51490
rect 27022 51438 27074 51490
rect 28142 51438 28194 51490
rect 29598 51438 29650 51490
rect 31054 51438 31106 51490
rect 34638 51438 34690 51490
rect 36990 51438 37042 51490
rect 37214 51438 37266 51490
rect 38110 51438 38162 51490
rect 41246 51438 41298 51490
rect 43038 51438 43090 51490
rect 47406 51438 47458 51490
rect 5070 51326 5122 51378
rect 5518 51326 5570 51378
rect 6078 51326 6130 51378
rect 10334 51326 10386 51378
rect 11118 51326 11170 51378
rect 12350 51326 12402 51378
rect 13694 51326 13746 51378
rect 15038 51326 15090 51378
rect 15374 51326 15426 51378
rect 16046 51326 16098 51378
rect 17502 51326 17554 51378
rect 21982 51326 22034 51378
rect 23774 51326 23826 51378
rect 26014 51326 26066 51378
rect 28926 51326 28978 51378
rect 30606 51326 30658 51378
rect 31166 51326 31218 51378
rect 31502 51326 31554 51378
rect 32510 51326 32562 51378
rect 33966 51326 34018 51378
rect 39454 51326 39506 51378
rect 39790 51326 39842 51378
rect 41470 51326 41522 51378
rect 42254 51326 42306 51378
rect 42478 51326 42530 51378
rect 43486 51326 43538 51378
rect 44158 51326 44210 51378
rect 48190 51326 48242 51378
rect 1822 51214 1874 51266
rect 4846 51214 4898 51266
rect 8990 51214 9042 51266
rect 13358 51214 13410 51266
rect 18174 51214 18226 51266
rect 20302 51214 20354 51266
rect 20638 51214 20690 51266
rect 23326 51214 23378 51266
rect 27358 51214 27410 51266
rect 27918 51214 27970 51266
rect 28702 51214 28754 51266
rect 33182 51214 33234 51266
rect 34302 51214 34354 51266
rect 37102 51214 37154 51266
rect 38782 51214 38834 51266
rect 40126 51214 40178 51266
rect 40462 51214 40514 51266
rect 42814 51214 42866 51266
rect 43934 51214 43986 51266
rect 45278 51214 45330 51266
rect 16494 51102 16546 51154
rect 23662 51102 23714 51154
rect 35870 51102 35922 51154
rect 38670 51102 38722 51154
rect 44494 51102 44546 51154
rect 4478 50934 4530 50986
rect 4582 50934 4634 50986
rect 4686 50934 4738 50986
rect 35198 50934 35250 50986
rect 35302 50934 35354 50986
rect 35406 50934 35458 50986
rect 16494 50766 16546 50818
rect 18398 50766 18450 50818
rect 18734 50766 18786 50818
rect 19294 50766 19346 50818
rect 22094 50766 22146 50818
rect 22430 50766 22482 50818
rect 27470 50766 27522 50818
rect 28590 50766 28642 50818
rect 29262 50766 29314 50818
rect 29598 50766 29650 50818
rect 31614 50766 31666 50818
rect 37102 50766 37154 50818
rect 43822 50766 43874 50818
rect 47518 50766 47570 50818
rect 48190 50766 48242 50818
rect 5966 50654 6018 50706
rect 6302 50654 6354 50706
rect 7086 50654 7138 50706
rect 9438 50654 9490 50706
rect 10782 50654 10834 50706
rect 12910 50654 12962 50706
rect 14926 50654 14978 50706
rect 16046 50654 16098 50706
rect 16606 50654 16658 50706
rect 19182 50654 19234 50706
rect 21870 50654 21922 50706
rect 24894 50654 24946 50706
rect 27022 50654 27074 50706
rect 28030 50654 28082 50706
rect 30158 50654 30210 50706
rect 36094 50654 36146 50706
rect 37550 50654 37602 50706
rect 38670 50654 38722 50706
rect 40798 50654 40850 50706
rect 42030 50654 42082 50706
rect 47070 50654 47122 50706
rect 47518 50654 47570 50706
rect 48078 50654 48130 50706
rect 2270 50542 2322 50594
rect 5630 50542 5682 50594
rect 6974 50542 7026 50594
rect 8318 50542 8370 50594
rect 8654 50542 8706 50594
rect 8990 50542 9042 50594
rect 9886 50542 9938 50594
rect 14142 50542 14194 50594
rect 14814 50542 14866 50594
rect 15374 50542 15426 50594
rect 16830 50542 16882 50594
rect 19630 50542 19682 50594
rect 20526 50542 20578 50594
rect 21310 50542 21362 50594
rect 23102 50542 23154 50594
rect 23662 50542 23714 50594
rect 23774 50542 23826 50594
rect 24110 50542 24162 50594
rect 27582 50542 27634 50594
rect 28254 50542 28306 50594
rect 30270 50542 30322 50594
rect 32622 50542 32674 50594
rect 33518 50542 33570 50594
rect 34078 50542 34130 50594
rect 34638 50542 34690 50594
rect 35086 50542 35138 50594
rect 35646 50542 35698 50594
rect 35982 50542 36034 50594
rect 37886 50542 37938 50594
rect 42366 50542 42418 50594
rect 43598 50542 43650 50594
rect 45502 50542 45554 50594
rect 1710 50430 1762 50482
rect 4846 50430 4898 50482
rect 8430 50430 8482 50482
rect 9998 50430 10050 50482
rect 11006 50430 11058 50482
rect 12686 50430 12738 50482
rect 13582 50430 13634 50482
rect 15486 50430 15538 50482
rect 17390 50430 17442 50482
rect 20078 50430 20130 50482
rect 21422 50430 21474 50482
rect 21646 50430 21698 50482
rect 27470 50430 27522 50482
rect 29486 50430 29538 50482
rect 29934 50430 29986 50482
rect 31054 50430 31106 50482
rect 32734 50430 32786 50482
rect 34414 50430 34466 50482
rect 35198 50430 35250 50482
rect 36318 50430 36370 50482
rect 36990 50430 37042 50482
rect 41470 50430 41522 50482
rect 45166 50430 45218 50482
rect 46846 50430 46898 50482
rect 5854 50318 5906 50370
rect 18510 50318 18562 50370
rect 20526 50318 20578 50370
rect 33518 50318 33570 50370
rect 34190 50318 34242 50370
rect 34974 50318 35026 50370
rect 41134 50318 41186 50370
rect 19838 50150 19890 50202
rect 19942 50150 19994 50202
rect 20046 50150 20098 50202
rect 10894 49982 10946 50034
rect 11566 49982 11618 50034
rect 11678 49982 11730 50034
rect 13022 49982 13074 50034
rect 13918 49982 13970 50034
rect 14590 49982 14642 50034
rect 14814 49982 14866 50034
rect 15038 49982 15090 50034
rect 32398 49982 32450 50034
rect 36654 49982 36706 50034
rect 37438 49982 37490 50034
rect 38110 49982 38162 50034
rect 39230 49982 39282 50034
rect 39790 49982 39842 50034
rect 41582 49982 41634 50034
rect 5630 49870 5682 49922
rect 12014 49870 12066 49922
rect 13358 49870 13410 49922
rect 15150 49870 15202 49922
rect 22654 49870 22706 49922
rect 22878 49870 22930 49922
rect 23438 49870 23490 49922
rect 23886 49870 23938 49922
rect 23998 49870 24050 49922
rect 26686 49870 26738 49922
rect 28478 49870 28530 49922
rect 29374 49870 29426 49922
rect 32174 49870 32226 49922
rect 33854 49870 33906 49922
rect 42142 49870 42194 49922
rect 46398 49870 46450 49922
rect 47854 49870 47906 49922
rect 1822 49758 1874 49810
rect 6526 49758 6578 49810
rect 11118 49758 11170 49810
rect 11790 49758 11842 49810
rect 14254 49758 14306 49810
rect 22542 49758 22594 49810
rect 23550 49758 23602 49810
rect 26798 49758 26850 49810
rect 27358 49758 27410 49810
rect 27582 49758 27634 49810
rect 28702 49758 28754 49810
rect 29710 49758 29762 49810
rect 33182 49758 33234 49810
rect 36318 49758 36370 49810
rect 36542 49758 36594 49810
rect 36766 49758 36818 49810
rect 36990 49758 37042 49810
rect 39118 49758 39170 49810
rect 39454 49758 39506 49810
rect 39790 49758 39842 49810
rect 40014 49758 40066 49810
rect 41358 49758 41410 49810
rect 41918 49758 41970 49810
rect 42590 49758 42642 49810
rect 45838 49758 45890 49810
rect 46734 49758 46786 49810
rect 47742 49758 47794 49810
rect 2494 49646 2546 49698
rect 4622 49646 4674 49698
rect 5070 49646 5122 49698
rect 7198 49646 7250 49698
rect 7870 49646 7922 49698
rect 10670 49646 10722 49698
rect 25454 49646 25506 49698
rect 25790 49646 25842 49698
rect 26574 49646 26626 49698
rect 28254 49646 28306 49698
rect 30158 49646 30210 49698
rect 32510 49646 32562 49698
rect 35982 49646 36034 49698
rect 38222 49646 38274 49698
rect 38670 49646 38722 49698
rect 40350 49646 40402 49698
rect 42030 49646 42082 49698
rect 42926 49646 42978 49698
rect 45054 49646 45106 49698
rect 46286 49646 46338 49698
rect 47406 49646 47458 49698
rect 13582 49534 13634 49586
rect 23438 49534 23490 49586
rect 23998 49534 24050 49586
rect 25902 49534 25954 49586
rect 4478 49366 4530 49418
rect 4582 49366 4634 49418
rect 4686 49366 4738 49418
rect 35198 49366 35250 49418
rect 35302 49366 35354 49418
rect 35406 49366 35458 49418
rect 6414 49198 6466 49250
rect 7310 49198 7362 49250
rect 8766 49198 8818 49250
rect 26462 49198 26514 49250
rect 29598 49198 29650 49250
rect 35982 49198 36034 49250
rect 45054 49198 45106 49250
rect 45390 49198 45442 49250
rect 6190 49086 6242 49138
rect 7422 49086 7474 49138
rect 18510 49086 18562 49138
rect 19630 49086 19682 49138
rect 25342 49086 25394 49138
rect 30046 49086 30098 49138
rect 32846 49086 32898 49138
rect 33742 49086 33794 49138
rect 34638 49086 34690 49138
rect 37102 49086 37154 49138
rect 39006 49086 39058 49138
rect 39454 49086 39506 49138
rect 40126 49086 40178 49138
rect 42142 49086 42194 49138
rect 44270 49086 44322 49138
rect 4734 48974 4786 49026
rect 5518 48974 5570 49026
rect 6302 48974 6354 49026
rect 9102 48974 9154 49026
rect 9326 48974 9378 49026
rect 9774 48974 9826 49026
rect 14030 48974 14082 49026
rect 14366 48974 14418 49026
rect 16382 48974 16434 49026
rect 18734 48974 18786 49026
rect 24558 48974 24610 49026
rect 26350 48974 26402 49026
rect 27358 48974 27410 49026
rect 27918 48974 27970 49026
rect 29262 48974 29314 49026
rect 31502 48974 31554 49026
rect 34190 48974 34242 49026
rect 35198 48974 35250 49026
rect 41358 48974 41410 49026
rect 44830 48974 44882 49026
rect 47630 48974 47682 49026
rect 4958 48862 5010 48914
rect 5070 48862 5122 48914
rect 11566 48862 11618 48914
rect 12238 48862 12290 48914
rect 14142 48862 14194 48914
rect 16046 48862 16098 48914
rect 17502 48862 17554 48914
rect 18062 48862 18114 48914
rect 18286 48862 18338 48914
rect 19966 48862 20018 48914
rect 20302 48862 20354 48914
rect 22542 48862 22594 48914
rect 26014 48862 26066 48914
rect 28590 48862 28642 48914
rect 30270 48862 30322 48914
rect 35422 48862 35474 48914
rect 35534 48862 35586 48914
rect 36094 48862 36146 48914
rect 41022 48862 41074 48914
rect 46734 48862 46786 48914
rect 3726 48750 3778 48802
rect 7534 48750 7586 48802
rect 8430 48750 8482 48802
rect 9998 48750 10050 48802
rect 10446 48750 10498 48802
rect 11678 48750 11730 48802
rect 11902 48750 11954 48802
rect 17390 48750 17442 48802
rect 19742 48750 19794 48802
rect 20414 48750 20466 48802
rect 20638 48750 20690 48802
rect 22878 48750 22930 48802
rect 23438 48750 23490 48802
rect 24110 48750 24162 48802
rect 24334 48750 24386 48802
rect 25678 48750 25730 48802
rect 26462 48750 26514 48802
rect 29486 48750 29538 48802
rect 35982 48750 36034 48802
rect 37774 48750 37826 48802
rect 40574 48750 40626 48802
rect 40910 48750 40962 48802
rect 45838 48750 45890 48802
rect 46510 48750 46562 48802
rect 46622 48750 46674 48802
rect 47406 48750 47458 48802
rect 48190 48750 48242 48802
rect 19838 48582 19890 48634
rect 19942 48582 19994 48634
rect 20046 48582 20098 48634
rect 3054 48414 3106 48466
rect 4398 48414 4450 48466
rect 9438 48414 9490 48466
rect 10670 48414 10722 48466
rect 12014 48414 12066 48466
rect 12574 48414 12626 48466
rect 15822 48414 15874 48466
rect 16718 48414 16770 48466
rect 16830 48414 16882 48466
rect 30382 48414 30434 48466
rect 42478 48414 42530 48466
rect 42590 48414 42642 48466
rect 43374 48414 43426 48466
rect 44046 48414 44098 48466
rect 44494 48414 44546 48466
rect 44942 48414 44994 48466
rect 3390 48302 3442 48354
rect 3950 48302 4002 48354
rect 4846 48302 4898 48354
rect 9662 48302 9714 48354
rect 10110 48302 10162 48354
rect 11678 48302 11730 48354
rect 11790 48302 11842 48354
rect 11902 48302 11954 48354
rect 12910 48302 12962 48354
rect 15710 48302 15762 48354
rect 20862 48302 20914 48354
rect 22206 48302 22258 48354
rect 24222 48302 24274 48354
rect 26238 48302 26290 48354
rect 27918 48302 27970 48354
rect 40014 48302 40066 48354
rect 41022 48302 41074 48354
rect 41694 48302 41746 48354
rect 42366 48302 42418 48354
rect 42926 48302 42978 48354
rect 47406 48302 47458 48354
rect 2158 48190 2210 48242
rect 2382 48190 2434 48242
rect 2718 48190 2770 48242
rect 2942 48190 2994 48242
rect 3166 48190 3218 48242
rect 4174 48190 4226 48242
rect 4958 48190 5010 48242
rect 5854 48190 5906 48242
rect 9774 48190 9826 48242
rect 10334 48190 10386 48242
rect 12126 48190 12178 48242
rect 12462 48190 12514 48242
rect 12686 48190 12738 48242
rect 16158 48190 16210 48242
rect 16606 48190 16658 48242
rect 17502 48190 17554 48242
rect 23774 48190 23826 48242
rect 25566 48190 25618 48242
rect 26574 48190 26626 48242
rect 26910 48190 26962 48242
rect 27134 48190 27186 48242
rect 27358 48190 27410 48242
rect 27582 48190 27634 48242
rect 28030 48190 28082 48242
rect 29934 48190 29986 48242
rect 30494 48190 30546 48242
rect 31278 48190 31330 48242
rect 35534 48190 35586 48242
rect 39230 48190 39282 48242
rect 40350 48190 40402 48242
rect 41470 48190 41522 48242
rect 42702 48190 42754 48242
rect 48078 48190 48130 48242
rect 2494 48078 2546 48130
rect 4286 48078 4338 48130
rect 6526 48078 6578 48130
rect 8654 48078 8706 48130
rect 15374 48078 15426 48130
rect 18174 48078 18226 48130
rect 20302 48078 20354 48130
rect 20638 48078 20690 48130
rect 22766 48078 22818 48130
rect 23326 48078 23378 48130
rect 24670 48078 24722 48130
rect 25342 48078 25394 48130
rect 27022 48078 27074 48130
rect 35870 48078 35922 48130
rect 36318 48078 36370 48130
rect 38446 48078 38498 48130
rect 39678 48078 39730 48130
rect 45278 48078 45330 48130
rect 4846 47966 4898 48018
rect 15822 47966 15874 48018
rect 39566 47966 39618 48018
rect 4478 47798 4530 47850
rect 4582 47798 4634 47850
rect 4686 47798 4738 47850
rect 35198 47798 35250 47850
rect 35302 47798 35354 47850
rect 35406 47798 35458 47850
rect 12798 47630 12850 47682
rect 18286 47630 18338 47682
rect 18622 47630 18674 47682
rect 37550 47630 37602 47682
rect 46734 47630 46786 47682
rect 2494 47518 2546 47570
rect 4622 47518 4674 47570
rect 5070 47518 5122 47570
rect 8542 47518 8594 47570
rect 9438 47518 9490 47570
rect 12126 47518 12178 47570
rect 16494 47518 16546 47570
rect 19630 47518 19682 47570
rect 23998 47518 24050 47570
rect 27470 47518 27522 47570
rect 29710 47518 29762 47570
rect 30718 47518 30770 47570
rect 35086 47518 35138 47570
rect 38894 47518 38946 47570
rect 41022 47518 41074 47570
rect 42142 47518 42194 47570
rect 46846 47518 46898 47570
rect 1822 47406 1874 47458
rect 7086 47406 7138 47458
rect 8318 47406 8370 47458
rect 8878 47406 8930 47458
rect 9326 47406 9378 47458
rect 9550 47406 9602 47458
rect 11230 47406 11282 47458
rect 11566 47406 11618 47458
rect 12462 47406 12514 47458
rect 13694 47406 13746 47458
rect 18286 47406 18338 47458
rect 20078 47406 20130 47458
rect 20526 47406 20578 47458
rect 21646 47406 21698 47458
rect 23550 47406 23602 47458
rect 24558 47406 24610 47458
rect 27694 47406 27746 47458
rect 28030 47406 28082 47458
rect 28366 47406 28418 47458
rect 29822 47406 29874 47458
rect 31278 47406 31330 47458
rect 31502 47406 31554 47458
rect 32174 47406 32226 47458
rect 33406 47406 33458 47458
rect 34974 47406 35026 47458
rect 35422 47406 35474 47458
rect 35646 47406 35698 47458
rect 37550 47406 37602 47458
rect 38222 47406 38274 47458
rect 41582 47406 41634 47458
rect 44830 47406 44882 47458
rect 45054 47406 45106 47458
rect 46622 47406 46674 47458
rect 47406 47406 47458 47458
rect 47966 47406 48018 47458
rect 7310 47294 7362 47346
rect 7646 47294 7698 47346
rect 10222 47294 10274 47346
rect 10558 47294 10610 47346
rect 14366 47294 14418 47346
rect 19406 47294 19458 47346
rect 21310 47294 21362 47346
rect 22094 47294 22146 47346
rect 22766 47294 22818 47346
rect 23438 47294 23490 47346
rect 25342 47294 25394 47346
rect 27918 47294 27970 47346
rect 34526 47294 34578 47346
rect 37214 47294 37266 47346
rect 42478 47294 42530 47346
rect 42702 47294 42754 47346
rect 43038 47294 43090 47346
rect 47630 47294 47682 47346
rect 6862 47182 6914 47234
rect 7198 47182 7250 47234
rect 11342 47182 11394 47234
rect 17054 47182 17106 47234
rect 17390 47182 17442 47234
rect 21422 47182 21474 47234
rect 22430 47182 22482 47234
rect 22878 47182 22930 47234
rect 23102 47182 23154 47234
rect 32734 47182 32786 47234
rect 32846 47182 32898 47234
rect 32958 47182 33010 47234
rect 33742 47182 33794 47234
rect 34414 47182 34466 47234
rect 35198 47182 35250 47234
rect 36206 47182 36258 47234
rect 41358 47182 41410 47234
rect 42926 47182 42978 47234
rect 43486 47182 43538 47234
rect 44270 47182 44322 47234
rect 45390 47182 45442 47234
rect 47742 47182 47794 47234
rect 19838 47014 19890 47066
rect 19942 47014 19994 47066
rect 20046 47014 20098 47066
rect 5070 46846 5122 46898
rect 7758 46846 7810 46898
rect 10446 46846 10498 46898
rect 11678 46846 11730 46898
rect 14926 46846 14978 46898
rect 15934 46846 15986 46898
rect 16718 46846 16770 46898
rect 24670 46846 24722 46898
rect 25342 46846 25394 46898
rect 26462 46846 26514 46898
rect 28702 46846 28754 46898
rect 34750 46846 34802 46898
rect 38782 46846 38834 46898
rect 39678 46846 39730 46898
rect 41022 46846 41074 46898
rect 44718 46846 44770 46898
rect 2830 46734 2882 46786
rect 7310 46734 7362 46786
rect 7534 46734 7586 46786
rect 7870 46734 7922 46786
rect 10222 46734 10274 46786
rect 10782 46734 10834 46786
rect 11006 46734 11058 46786
rect 11342 46734 11394 46786
rect 11454 46734 11506 46786
rect 12238 46734 12290 46786
rect 15822 46734 15874 46786
rect 16046 46734 16098 46786
rect 17726 46734 17778 46786
rect 18398 46734 18450 46786
rect 19182 46734 19234 46786
rect 27806 46734 27858 46786
rect 29934 46734 29986 46786
rect 31950 46734 32002 46786
rect 32510 46734 32562 46786
rect 35310 46734 35362 46786
rect 3278 46622 3330 46674
rect 3726 46622 3778 46674
rect 4510 46622 4562 46674
rect 10110 46622 10162 46674
rect 10670 46622 10722 46674
rect 14702 46622 14754 46674
rect 15150 46622 15202 46674
rect 15374 46622 15426 46674
rect 16494 46622 16546 46674
rect 16830 46622 16882 46674
rect 18510 46622 18562 46674
rect 18958 46622 19010 46674
rect 20414 46622 20466 46674
rect 23102 46622 23154 46674
rect 24334 46622 24386 46674
rect 27358 46622 27410 46674
rect 29150 46622 29202 46674
rect 29374 46622 29426 46674
rect 29486 46622 29538 46674
rect 29710 46622 29762 46674
rect 30270 46622 30322 46674
rect 32286 46622 32338 46674
rect 33294 46622 33346 46674
rect 33742 46622 33794 46674
rect 34190 46622 34242 46674
rect 36318 46622 36370 46674
rect 38894 46622 38946 46674
rect 39230 46622 39282 46674
rect 39342 46622 39394 46674
rect 39902 46622 39954 46674
rect 44270 46622 44322 46674
rect 48078 46622 48130 46674
rect 9774 46510 9826 46562
rect 17838 46510 17890 46562
rect 21086 46510 21138 46562
rect 23214 46510 23266 46562
rect 23886 46510 23938 46562
rect 25790 46510 25842 46562
rect 27022 46510 27074 46562
rect 28142 46510 28194 46562
rect 30382 46510 30434 46562
rect 32062 46510 32114 46562
rect 36990 46510 37042 46562
rect 39566 46510 39618 46562
rect 40350 46510 40402 46562
rect 41358 46510 41410 46562
rect 43486 46510 43538 46562
rect 45278 46510 45330 46562
rect 47406 46510 47458 46562
rect 4734 46398 4786 46450
rect 12350 46398 12402 46450
rect 17950 46398 18002 46450
rect 18622 46398 18674 46450
rect 19294 46398 19346 46450
rect 28366 46398 28418 46450
rect 35086 46398 35138 46450
rect 35422 46398 35474 46450
rect 4478 46230 4530 46282
rect 4582 46230 4634 46282
rect 4686 46230 4738 46282
rect 35198 46230 35250 46282
rect 35302 46230 35354 46282
rect 35406 46230 35458 46282
rect 25342 46062 25394 46114
rect 27358 46062 27410 46114
rect 43150 46062 43202 46114
rect 43486 46062 43538 46114
rect 45950 46062 46002 46114
rect 46286 46062 46338 46114
rect 47070 46062 47122 46114
rect 10334 45950 10386 46002
rect 12798 45950 12850 46002
rect 15038 45950 15090 46002
rect 17390 45950 17442 46002
rect 20078 45950 20130 46002
rect 22094 45950 22146 46002
rect 22542 45950 22594 46002
rect 27918 45950 27970 46002
rect 31614 45950 31666 46002
rect 33742 45950 33794 46002
rect 36430 45950 36482 46002
rect 39902 45950 39954 46002
rect 41918 45950 41970 46002
rect 44830 45950 44882 46002
rect 46958 45950 47010 46002
rect 4398 45838 4450 45890
rect 6526 45838 6578 45890
rect 6974 45838 7026 45890
rect 7646 45838 7698 45890
rect 10782 45838 10834 45890
rect 12350 45838 12402 45890
rect 12686 45838 12738 45890
rect 13582 45838 13634 45890
rect 13918 45838 13970 45890
rect 15598 45838 15650 45890
rect 16046 45838 16098 45890
rect 19294 45838 19346 45890
rect 19630 45838 19682 45890
rect 20190 45838 20242 45890
rect 21870 45838 21922 45890
rect 23214 45838 23266 45890
rect 25006 45838 25058 45890
rect 27694 45838 27746 45890
rect 29598 45838 29650 45890
rect 30942 45838 30994 45890
rect 34862 45838 34914 45890
rect 35870 45838 35922 45890
rect 37102 45838 37154 45890
rect 40350 45838 40402 45890
rect 43262 45838 43314 45890
rect 43598 45838 43650 45890
rect 45278 45838 45330 45890
rect 45838 45838 45890 45890
rect 46174 45838 46226 45890
rect 46734 45838 46786 45890
rect 47630 45838 47682 45890
rect 2270 45726 2322 45778
rect 2606 45726 2658 45778
rect 2830 45726 2882 45778
rect 3614 45726 3666 45778
rect 4062 45726 4114 45778
rect 4734 45726 4786 45778
rect 4846 45726 4898 45778
rect 5966 45726 6018 45778
rect 6302 45726 6354 45778
rect 7982 45726 8034 45778
rect 11230 45726 11282 45778
rect 12910 45726 12962 45778
rect 20302 45726 20354 45778
rect 23998 45726 24050 45778
rect 25454 45726 25506 45778
rect 25678 45726 25730 45778
rect 26014 45726 26066 45778
rect 29934 45726 29986 45778
rect 34526 45726 34578 45778
rect 37774 45726 37826 45778
rect 45166 45726 45218 45778
rect 2494 45614 2546 45666
rect 3278 45614 3330 45666
rect 3502 45614 3554 45666
rect 3726 45614 3778 45666
rect 4174 45614 4226 45666
rect 4510 45614 4562 45666
rect 6078 45614 6130 45666
rect 6862 45614 6914 45666
rect 7086 45614 7138 45666
rect 7310 45614 7362 45666
rect 7870 45614 7922 45666
rect 11566 45614 11618 45666
rect 16158 45614 16210 45666
rect 16270 45614 16322 45666
rect 22878 45614 22930 45666
rect 24334 45614 24386 45666
rect 24446 45614 24498 45666
rect 24558 45614 24610 45666
rect 25342 45614 25394 45666
rect 25902 45614 25954 45666
rect 44158 45614 44210 45666
rect 48190 45614 48242 45666
rect 19838 45446 19890 45498
rect 19942 45446 19994 45498
rect 20046 45446 20098 45498
rect 3838 45278 3890 45330
rect 8094 45278 8146 45330
rect 21198 45278 21250 45330
rect 33742 45278 33794 45330
rect 34302 45278 34354 45330
rect 34414 45278 34466 45330
rect 34526 45278 34578 45330
rect 38670 45278 38722 45330
rect 40014 45278 40066 45330
rect 40910 45278 40962 45330
rect 44830 45278 44882 45330
rect 45390 45278 45442 45330
rect 47070 45278 47122 45330
rect 2382 45166 2434 45218
rect 3726 45166 3778 45218
rect 5518 45166 5570 45218
rect 8430 45166 8482 45218
rect 11454 45166 11506 45218
rect 13694 45166 13746 45218
rect 18174 45166 18226 45218
rect 26574 45166 26626 45218
rect 27582 45166 27634 45218
rect 29374 45166 29426 45218
rect 33406 45166 33458 45218
rect 33518 45166 33570 45218
rect 38558 45166 38610 45218
rect 3054 45054 3106 45106
rect 3950 45054 4002 45106
rect 4398 45054 4450 45106
rect 4846 45054 4898 45106
rect 7982 45054 8034 45106
rect 8206 45054 8258 45106
rect 8990 45054 9042 45106
rect 10782 45054 10834 45106
rect 12910 45054 12962 45106
rect 16270 45054 16322 45106
rect 16830 45054 16882 45106
rect 17502 45054 17554 45106
rect 21758 45054 21810 45106
rect 25454 45054 25506 45106
rect 25902 45054 25954 45106
rect 26798 45054 26850 45106
rect 27246 45054 27298 45106
rect 29262 45054 29314 45106
rect 29598 45054 29650 45106
rect 30270 45054 30322 45106
rect 31950 45054 32002 45106
rect 34078 45054 34130 45106
rect 34750 45054 34802 45106
rect 35310 45054 35362 45106
rect 38782 45054 38834 45106
rect 39118 45054 39170 45106
rect 39454 45054 39506 45106
rect 39678 45054 39730 45106
rect 40350 45054 40402 45106
rect 41134 45054 41186 45106
rect 41582 45054 41634 45106
rect 42814 45054 42866 45106
rect 43038 45054 43090 45106
rect 43934 45054 43986 45106
rect 44494 45054 44546 45106
rect 44830 45054 44882 45106
rect 45166 45054 45218 45106
rect 45614 45054 45666 45106
rect 46286 45054 46338 45106
rect 46510 45054 46562 45106
rect 46622 45054 46674 45106
rect 47966 45054 48018 45106
rect 3166 44942 3218 44994
rect 7646 44942 7698 44994
rect 9550 44942 9602 44994
rect 11118 44942 11170 44994
rect 15822 44942 15874 44994
rect 20302 44942 20354 44994
rect 20750 44942 20802 44994
rect 22542 44942 22594 44994
rect 24670 44942 24722 44994
rect 25230 44942 25282 44994
rect 29822 44942 29874 44994
rect 35982 44942 36034 44994
rect 38110 44942 38162 44994
rect 39566 44942 39618 44994
rect 42030 44942 42082 44994
rect 43598 44942 43650 44994
rect 47518 44942 47570 44994
rect 9774 44830 9826 44882
rect 10110 44830 10162 44882
rect 16494 44830 16546 44882
rect 29934 44830 29986 44882
rect 42702 44830 42754 44882
rect 43486 44830 43538 44882
rect 47406 44830 47458 44882
rect 47742 44830 47794 44882
rect 4478 44662 4530 44714
rect 4582 44662 4634 44714
rect 4686 44662 4738 44714
rect 35198 44662 35250 44714
rect 35302 44662 35354 44714
rect 35406 44662 35458 44714
rect 7758 44494 7810 44546
rect 11342 44494 11394 44546
rect 19854 44494 19906 44546
rect 20750 44494 20802 44546
rect 24894 44494 24946 44546
rect 26238 44494 26290 44546
rect 34638 44494 34690 44546
rect 35758 44494 35810 44546
rect 38110 44494 38162 44546
rect 41134 44494 41186 44546
rect 42926 44494 42978 44546
rect 2494 44382 2546 44434
rect 4622 44382 4674 44434
rect 6302 44382 6354 44434
rect 6750 44382 6802 44434
rect 14478 44382 14530 44434
rect 14702 44382 14754 44434
rect 15150 44382 15202 44434
rect 19854 44382 19906 44434
rect 20750 44382 20802 44434
rect 23550 44382 23602 44434
rect 24670 44382 24722 44434
rect 26014 44382 26066 44434
rect 29374 44382 29426 44434
rect 31502 44382 31554 44434
rect 32398 44382 32450 44434
rect 34526 44382 34578 44434
rect 35870 44382 35922 44434
rect 37214 44382 37266 44434
rect 38222 44382 38274 44434
rect 38670 44382 38722 44434
rect 43038 44382 43090 44434
rect 44158 44382 44210 44434
rect 45278 44382 45330 44434
rect 47406 44382 47458 44434
rect 1822 44270 1874 44322
rect 6862 44270 6914 44322
rect 10558 44270 10610 44322
rect 10782 44270 10834 44322
rect 12462 44270 12514 44322
rect 15374 44270 15426 44322
rect 18622 44270 18674 44322
rect 23438 44270 23490 44322
rect 23662 44270 23714 44322
rect 23998 44270 24050 44322
rect 24894 44270 24946 44322
rect 25342 44270 25394 44322
rect 27246 44270 27298 44322
rect 27694 44270 27746 44322
rect 27918 44270 27970 44322
rect 29598 44270 29650 44322
rect 30158 44270 30210 44322
rect 30606 44270 30658 44322
rect 30830 44270 30882 44322
rect 33854 44270 33906 44322
rect 36094 44270 36146 44322
rect 40798 44270 40850 44322
rect 41134 44270 41186 44322
rect 41582 44270 41634 44322
rect 41918 44270 41970 44322
rect 42366 44270 42418 44322
rect 44270 44270 44322 44322
rect 48078 44270 48130 44322
rect 5070 44046 5122 44098
rect 5742 44046 5794 44098
rect 7646 44102 7698 44154
rect 7758 44158 7810 44210
rect 8766 44158 8818 44210
rect 10894 44158 10946 44210
rect 12126 44158 12178 44210
rect 16830 44158 16882 44210
rect 34190 44158 34242 44210
rect 42590 44158 42642 44210
rect 43822 44158 43874 44210
rect 43934 44158 43986 44210
rect 44942 44158 44994 44210
rect 9102 44046 9154 44098
rect 9550 44046 9602 44098
rect 9886 44046 9938 44098
rect 12238 44046 12290 44098
rect 19406 44046 19458 44098
rect 20302 44046 20354 44098
rect 22766 44046 22818 44098
rect 26574 44046 26626 44098
rect 31838 44046 31890 44098
rect 34078 44046 34130 44098
rect 40238 44046 40290 44098
rect 41694 44046 41746 44098
rect 44046 44046 44098 44098
rect 19838 43878 19890 43930
rect 19942 43878 19994 43930
rect 20046 43878 20098 43930
rect 10334 43710 10386 43762
rect 12126 43710 12178 43762
rect 25342 43710 25394 43762
rect 28142 43710 28194 43762
rect 36430 43710 36482 43762
rect 38782 43710 38834 43762
rect 41470 43710 41522 43762
rect 47070 43710 47122 43762
rect 3838 43598 3890 43650
rect 5406 43598 5458 43650
rect 8094 43598 8146 43650
rect 11230 43598 11282 43650
rect 11454 43598 11506 43650
rect 15374 43598 15426 43650
rect 15822 43598 15874 43650
rect 16382 43598 16434 43650
rect 16494 43598 16546 43650
rect 20302 43598 20354 43650
rect 21870 43598 21922 43650
rect 25230 43598 25282 43650
rect 26798 43598 26850 43650
rect 27246 43598 27298 43650
rect 29710 43598 29762 43650
rect 31054 43598 31106 43650
rect 36318 43598 36370 43650
rect 37326 43598 37378 43650
rect 37774 43598 37826 43650
rect 40910 43598 40962 43650
rect 41022 43598 41074 43650
rect 43262 43598 43314 43650
rect 44382 43598 44434 43650
rect 47182 43598 47234 43650
rect 48302 43598 48354 43650
rect 4286 43486 4338 43538
rect 4958 43486 5010 43538
rect 5182 43486 5234 43538
rect 5518 43486 5570 43538
rect 7870 43486 7922 43538
rect 8206 43486 8258 43538
rect 10222 43486 10274 43538
rect 10446 43486 10498 43538
rect 10894 43486 10946 43538
rect 11118 43486 11170 43538
rect 11678 43486 11730 43538
rect 12014 43486 12066 43538
rect 12238 43486 12290 43538
rect 12574 43486 12626 43538
rect 15710 43486 15762 43538
rect 16270 43486 16322 43538
rect 16830 43486 16882 43538
rect 17950 43486 18002 43538
rect 20750 43486 20802 43538
rect 26350 43486 26402 43538
rect 26686 43486 26738 43538
rect 27694 43486 27746 43538
rect 28030 43486 28082 43538
rect 29150 43486 29202 43538
rect 30382 43486 30434 43538
rect 35870 43486 35922 43538
rect 36542 43486 36594 43538
rect 36878 43486 36930 43538
rect 38558 43486 38610 43538
rect 39006 43486 39058 43538
rect 39230 43486 39282 43538
rect 43598 43486 43650 43538
rect 46734 43486 46786 43538
rect 47294 43486 47346 43538
rect 4398 43374 4450 43426
rect 14926 43374 14978 43426
rect 19630 43374 19682 43426
rect 22318 43374 22370 43426
rect 29374 43374 29426 43426
rect 30718 43374 30770 43426
rect 33070 43374 33122 43426
rect 35198 43374 35250 43426
rect 38782 43374 38834 43426
rect 39790 43374 39842 43426
rect 40126 43374 40178 43426
rect 46510 43374 46562 43426
rect 12798 43262 12850 43314
rect 13134 43262 13186 43314
rect 15822 43262 15874 43314
rect 4478 43094 4530 43146
rect 4582 43094 4634 43146
rect 4686 43094 4738 43146
rect 35198 43094 35250 43146
rect 35302 43094 35354 43146
rect 35406 43094 35458 43146
rect 4734 42926 4786 42978
rect 8318 42926 8370 42978
rect 12238 42926 12290 42978
rect 24558 42926 24610 42978
rect 24782 42926 24834 42978
rect 11118 42814 11170 42866
rect 17166 42814 17218 42866
rect 21758 42814 21810 42866
rect 22654 42814 22706 42866
rect 24558 42814 24610 42866
rect 25902 42814 25954 42866
rect 30046 42814 30098 42866
rect 34190 42814 34242 42866
rect 36318 42814 36370 42866
rect 38110 42814 38162 42866
rect 40014 42814 40066 42866
rect 40238 42814 40290 42866
rect 40686 42814 40738 42866
rect 42030 42814 42082 42866
rect 44158 42814 44210 42866
rect 45054 42814 45106 42866
rect 3390 42702 3442 42754
rect 3838 42702 3890 42754
rect 4846 42702 4898 42754
rect 5742 42702 5794 42754
rect 5966 42702 6018 42754
rect 6302 42702 6354 42754
rect 7198 42702 7250 42754
rect 7758 42702 7810 42754
rect 8094 42702 8146 42754
rect 8654 42702 8706 42754
rect 8990 42702 9042 42754
rect 9326 42702 9378 42754
rect 10446 42702 10498 42754
rect 10894 42702 10946 42754
rect 11790 42702 11842 42754
rect 12014 42702 12066 42754
rect 14702 42702 14754 42754
rect 15038 42702 15090 42754
rect 15598 42702 15650 42754
rect 16270 42702 16322 42754
rect 16494 42702 16546 42754
rect 19966 42702 20018 42754
rect 20862 42702 20914 42754
rect 21982 42702 22034 42754
rect 23102 42702 23154 42754
rect 25678 42702 25730 42754
rect 26238 42702 26290 42754
rect 27134 42702 27186 42754
rect 27358 42702 27410 42754
rect 31390 42702 31442 42754
rect 32062 42702 32114 42754
rect 32958 42702 33010 42754
rect 33070 42702 33122 42754
rect 33294 42702 33346 42754
rect 33630 42702 33682 42754
rect 34078 42702 34130 42754
rect 34638 42702 34690 42754
rect 36990 42702 37042 42754
rect 37662 42702 37714 42754
rect 38222 42702 38274 42754
rect 38446 42702 38498 42754
rect 39006 42702 39058 42754
rect 39230 42702 39282 42754
rect 39342 42702 39394 42754
rect 41246 42702 41298 42754
rect 2830 42590 2882 42642
rect 3166 42590 3218 42642
rect 6638 42590 6690 42642
rect 16606 42590 16658 42642
rect 19294 42590 19346 42642
rect 20526 42590 20578 42642
rect 21422 42590 21474 42642
rect 23438 42590 23490 42642
rect 23774 42590 23826 42642
rect 23998 42590 24050 42642
rect 30494 42590 30546 42642
rect 33406 42590 33458 42642
rect 38670 42590 38722 42642
rect 39678 42590 39730 42642
rect 2606 42478 2658 42530
rect 2942 42478 2994 42530
rect 3726 42478 3778 42530
rect 3950 42478 4002 42530
rect 4174 42478 4226 42530
rect 4734 42478 4786 42530
rect 6078 42478 6130 42530
rect 6526 42478 6578 42530
rect 6750 42478 6802 42530
rect 9214 42478 9266 42530
rect 12686 42478 12738 42530
rect 14814 42478 14866 42530
rect 20638 42478 20690 42530
rect 21646 42478 21698 42530
rect 23886 42478 23938 42530
rect 27694 42478 27746 42530
rect 34302 42478 34354 42530
rect 34750 42478 34802 42530
rect 34974 42478 35026 42530
rect 37102 42478 37154 42530
rect 37214 42478 37266 42530
rect 38110 42478 38162 42530
rect 40014 42478 40066 42530
rect 46734 42478 46786 42530
rect 47182 42478 47234 42530
rect 48302 42478 48354 42530
rect 19838 42310 19890 42362
rect 19942 42310 19994 42362
rect 20046 42310 20098 42362
rect 18510 42142 18562 42194
rect 29486 42142 29538 42194
rect 33182 42142 33234 42194
rect 34526 42142 34578 42194
rect 34974 42142 35026 42194
rect 41022 42142 41074 42194
rect 2494 42030 2546 42082
rect 6078 42030 6130 42082
rect 9550 42030 9602 42082
rect 12238 42030 12290 42082
rect 17838 42030 17890 42082
rect 19070 42030 19122 42082
rect 30158 42030 30210 42082
rect 33294 42030 33346 42082
rect 34302 42030 34354 42082
rect 34862 42030 34914 42082
rect 40014 42030 40066 42082
rect 47070 42030 47122 42082
rect 1822 41918 1874 41970
rect 5406 41918 5458 41970
rect 8654 41918 8706 41970
rect 9662 41918 9714 41970
rect 10446 41918 10498 41970
rect 11006 41918 11058 41970
rect 11902 41918 11954 41970
rect 12574 41918 12626 41970
rect 16382 41918 16434 41970
rect 18286 41918 18338 41970
rect 19182 41918 19234 41970
rect 19742 41918 19794 41970
rect 20526 41918 20578 41970
rect 24222 41918 24274 41970
rect 24670 41918 24722 41970
rect 25342 41918 25394 41970
rect 25566 41918 25618 41970
rect 26238 41918 26290 41970
rect 27358 41918 27410 41970
rect 29262 41918 29314 41970
rect 29822 41918 29874 41970
rect 33966 41918 34018 41970
rect 35198 41918 35250 41970
rect 35534 41918 35586 41970
rect 36318 41918 36370 41970
rect 46510 41918 46562 41970
rect 48078 41918 48130 41970
rect 4622 41806 4674 41858
rect 8206 41806 8258 41858
rect 10334 41806 10386 41858
rect 10894 41806 10946 41858
rect 11566 41806 11618 41858
rect 13358 41806 13410 41858
rect 15486 41806 15538 41858
rect 15822 41806 15874 41858
rect 16718 41806 16770 41858
rect 17726 41806 17778 41858
rect 22654 41806 22706 41858
rect 26462 41806 26514 41858
rect 27470 41806 27522 41858
rect 28590 41806 28642 41858
rect 34414 41806 34466 41858
rect 38446 41806 38498 41858
rect 38894 41806 38946 41858
rect 39342 41806 39394 41858
rect 46398 41806 46450 41858
rect 10110 41694 10162 41746
rect 17614 41694 17666 41746
rect 18622 41694 18674 41746
rect 19070 41694 19122 41746
rect 33070 41694 33122 41746
rect 38894 41694 38946 41746
rect 39566 41694 39618 41746
rect 40126 41694 40178 41746
rect 45726 41694 45778 41746
rect 47182 41694 47234 41746
rect 47406 41694 47458 41746
rect 47518 41694 47570 41746
rect 4478 41526 4530 41578
rect 4582 41526 4634 41578
rect 4686 41526 4738 41578
rect 35198 41526 35250 41578
rect 35302 41526 35354 41578
rect 35406 41526 35458 41578
rect 12798 41358 12850 41410
rect 25678 41358 25730 41410
rect 26014 41358 26066 41410
rect 30158 41358 30210 41410
rect 43486 41358 43538 41410
rect 3054 41246 3106 41298
rect 3390 41246 3442 41298
rect 4958 41246 5010 41298
rect 6974 41246 7026 41298
rect 7310 41246 7362 41298
rect 8542 41246 8594 41298
rect 10782 41246 10834 41298
rect 11566 41246 11618 41298
rect 14030 41246 14082 41298
rect 14478 41246 14530 41298
rect 15150 41246 15202 41298
rect 21422 41246 21474 41298
rect 24558 41246 24610 41298
rect 25454 41246 25506 41298
rect 27806 41246 27858 41298
rect 29710 41246 29762 41298
rect 32510 41246 32562 41298
rect 33182 41246 33234 41298
rect 35310 41246 35362 41298
rect 39342 41246 39394 41298
rect 41470 41246 41522 41298
rect 42814 41246 42866 41298
rect 46062 41246 46114 41298
rect 48190 41246 48242 41298
rect 3502 41134 3554 41186
rect 4510 41134 4562 41186
rect 7646 41134 7698 41186
rect 10222 41134 10274 41186
rect 11230 41134 11282 41186
rect 12126 41134 12178 41186
rect 13806 41134 13858 41186
rect 15038 41134 15090 41186
rect 15598 41134 15650 41186
rect 16046 41134 16098 41186
rect 16606 41134 16658 41186
rect 17614 41134 17666 41186
rect 18398 41134 18450 41186
rect 19854 41134 19906 41186
rect 24670 41134 24722 41186
rect 25118 41134 25170 41186
rect 27470 41134 27522 41186
rect 29038 41134 29090 41186
rect 29822 41134 29874 41186
rect 32846 41134 32898 41186
rect 33518 41134 33570 41186
rect 33854 41134 33906 41186
rect 36990 41134 37042 41186
rect 38110 41134 38162 41186
rect 38782 41134 38834 41186
rect 42254 41134 42306 41186
rect 43150 41134 43202 41186
rect 45390 41134 45442 41186
rect 9886 41022 9938 41074
rect 12910 41022 12962 41074
rect 15374 41022 15426 41074
rect 17390 41022 17442 41074
rect 20526 41022 20578 41074
rect 20638 41022 20690 41074
rect 21646 41022 21698 41074
rect 23326 41022 23378 41074
rect 27246 41022 27298 41074
rect 33070 41022 33122 41074
rect 37102 41022 37154 41074
rect 37662 41022 37714 41074
rect 38446 41022 38498 41074
rect 4398 40910 4450 40962
rect 8990 40910 9042 40962
rect 12350 40910 12402 40962
rect 12798 40910 12850 40962
rect 15934 40910 15986 40962
rect 16158 40910 16210 40962
rect 18734 40910 18786 40962
rect 19630 40910 19682 40962
rect 20862 40910 20914 40962
rect 23438 40910 23490 40962
rect 33294 40910 33346 40962
rect 37774 40910 37826 40962
rect 38334 40910 38386 40962
rect 38558 40910 38610 40962
rect 43374 40910 43426 40962
rect 19838 40742 19890 40794
rect 19942 40742 19994 40794
rect 20046 40742 20098 40794
rect 8318 40574 8370 40626
rect 11118 40574 11170 40626
rect 16382 40574 16434 40626
rect 20862 40574 20914 40626
rect 21646 40574 21698 40626
rect 32174 40574 32226 40626
rect 34190 40574 34242 40626
rect 47518 40574 47570 40626
rect 4510 40462 4562 40514
rect 8878 40462 8930 40514
rect 8990 40462 9042 40514
rect 10782 40462 10834 40514
rect 12238 40462 12290 40514
rect 12686 40462 12738 40514
rect 13358 40462 13410 40514
rect 14030 40462 14082 40514
rect 14142 40462 14194 40514
rect 16270 40462 16322 40514
rect 17614 40462 17666 40514
rect 23886 40462 23938 40514
rect 30270 40462 30322 40514
rect 33182 40462 33234 40514
rect 33294 40462 33346 40514
rect 35758 40462 35810 40514
rect 38222 40462 38274 40514
rect 41918 40462 41970 40514
rect 43374 40462 43426 40514
rect 45950 40462 46002 40514
rect 48190 40462 48242 40514
rect 4286 40350 4338 40402
rect 4622 40350 4674 40402
rect 7870 40350 7922 40402
rect 8206 40350 8258 40402
rect 9886 40350 9938 40402
rect 10446 40350 10498 40402
rect 11566 40350 11618 40402
rect 11790 40350 11842 40402
rect 12574 40350 12626 40402
rect 13582 40350 13634 40402
rect 14366 40350 14418 40402
rect 15934 40350 15986 40402
rect 16830 40350 16882 40402
rect 17726 40350 17778 40402
rect 17950 40350 18002 40402
rect 19070 40350 19122 40402
rect 19518 40350 19570 40402
rect 20414 40350 20466 40402
rect 21086 40350 21138 40402
rect 21310 40350 21362 40402
rect 21982 40350 22034 40402
rect 22430 40350 22482 40402
rect 24446 40350 24498 40402
rect 27134 40350 27186 40402
rect 28926 40350 28978 40402
rect 29822 40350 29874 40402
rect 30046 40350 30098 40402
rect 30382 40350 30434 40402
rect 31838 40350 31890 40402
rect 32062 40350 32114 40402
rect 32286 40350 32338 40402
rect 33518 40350 33570 40402
rect 34526 40350 34578 40402
rect 36542 40350 36594 40402
rect 37438 40350 37490 40402
rect 40910 40350 40962 40402
rect 41470 40350 41522 40402
rect 42702 40350 42754 40402
rect 46734 40350 46786 40402
rect 46958 40350 47010 40402
rect 47070 40350 47122 40402
rect 15374 40238 15426 40290
rect 19742 40238 19794 40290
rect 21198 40238 21250 40290
rect 27470 40238 27522 40290
rect 27918 40238 27970 40290
rect 29038 40238 29090 40290
rect 35982 40238 36034 40290
rect 37102 40238 37154 40290
rect 40350 40238 40402 40290
rect 45502 40238 45554 40290
rect 46174 40238 46226 40290
rect 47854 40238 47906 40290
rect 8318 40126 8370 40178
rect 8878 40126 8930 40178
rect 45838 40126 45890 40178
rect 4478 39958 4530 40010
rect 4582 39958 4634 40010
rect 4686 39958 4738 40010
rect 35198 39958 35250 40010
rect 35302 39958 35354 40010
rect 35406 39958 35458 40010
rect 2830 39790 2882 39842
rect 3950 39790 4002 39842
rect 35646 39790 35698 39842
rect 35982 39790 36034 39842
rect 36206 39790 36258 39842
rect 36542 39790 36594 39842
rect 45614 39790 45666 39842
rect 3166 39678 3218 39730
rect 8542 39678 8594 39730
rect 10894 39678 10946 39730
rect 12126 39678 12178 39730
rect 12910 39678 12962 39730
rect 13918 39678 13970 39730
rect 17950 39678 18002 39730
rect 20078 39678 20130 39730
rect 20750 39678 20802 39730
rect 22206 39678 22258 39730
rect 24110 39678 24162 39730
rect 29262 39678 29314 39730
rect 31726 39678 31778 39730
rect 33182 39678 33234 39730
rect 35310 39678 35362 39730
rect 36990 39678 37042 39730
rect 41134 39678 41186 39730
rect 42478 39678 42530 39730
rect 43374 39678 43426 39730
rect 47182 39678 47234 39730
rect 3614 39566 3666 39618
rect 3838 39566 3890 39618
rect 4510 39566 4562 39618
rect 5742 39566 5794 39618
rect 9550 39566 9602 39618
rect 12238 39566 12290 39618
rect 13470 39566 13522 39618
rect 13806 39566 13858 39618
rect 14030 39566 14082 39618
rect 14814 39566 14866 39618
rect 15374 39566 15426 39618
rect 16046 39566 16098 39618
rect 19518 39566 19570 39618
rect 21982 39566 22034 39618
rect 22318 39566 22370 39618
rect 23774 39566 23826 39618
rect 24670 39566 24722 39618
rect 25006 39566 25058 39618
rect 26014 39566 26066 39618
rect 26126 39566 26178 39618
rect 28030 39566 28082 39618
rect 28590 39566 28642 39618
rect 30718 39566 30770 39618
rect 32398 39566 32450 39618
rect 39118 39566 39170 39618
rect 42030 39566 42082 39618
rect 45838 39566 45890 39618
rect 47070 39566 47122 39618
rect 47406 39566 47458 39618
rect 47630 39566 47682 39618
rect 3054 39454 3106 39506
rect 6414 39454 6466 39506
rect 10446 39454 10498 39506
rect 15486 39454 15538 39506
rect 15822 39454 15874 39506
rect 18398 39454 18450 39506
rect 21422 39454 21474 39506
rect 21758 39454 21810 39506
rect 22654 39454 22706 39506
rect 23550 39454 23602 39506
rect 25566 39454 25618 39506
rect 26462 39454 26514 39506
rect 27918 39454 27970 39506
rect 29710 39454 29762 39506
rect 37550 39454 37602 39506
rect 37998 39454 38050 39506
rect 41694 39454 41746 39506
rect 42366 39454 42418 39506
rect 42702 39454 42754 39506
rect 42926 39454 42978 39506
rect 46398 39454 46450 39506
rect 46734 39454 46786 39506
rect 8990 39342 9042 39394
rect 17166 39342 17218 39394
rect 17614 39342 17666 39394
rect 24558 39342 24610 39394
rect 26350 39342 26402 39394
rect 28478 39342 28530 39394
rect 35870 39342 35922 39394
rect 36430 39342 36482 39394
rect 38334 39342 38386 39394
rect 41806 39342 41858 39394
rect 45278 39342 45330 39394
rect 46062 39342 46114 39394
rect 46286 39342 46338 39394
rect 48190 39342 48242 39394
rect 19838 39174 19890 39226
rect 19942 39174 19994 39226
rect 20046 39174 20098 39226
rect 6302 39006 6354 39058
rect 6414 39006 6466 39058
rect 6974 39006 7026 39058
rect 7422 39006 7474 39058
rect 7982 39006 8034 39058
rect 8318 39006 8370 39058
rect 8654 39006 8706 39058
rect 11790 39006 11842 39058
rect 12574 39006 12626 39058
rect 14030 39006 14082 39058
rect 17950 39006 18002 39058
rect 18286 39006 18338 39058
rect 22654 39006 22706 39058
rect 28926 39006 28978 39058
rect 30382 39006 30434 39058
rect 33070 39006 33122 39058
rect 33182 39006 33234 39058
rect 33294 39006 33346 39058
rect 45390 39006 45442 39058
rect 6526 38894 6578 38946
rect 7646 38894 7698 38946
rect 8990 38894 9042 38946
rect 10894 38894 10946 38946
rect 12910 38894 12962 38946
rect 16606 38894 16658 38946
rect 19070 38894 19122 38946
rect 24670 38894 24722 38946
rect 27358 38894 27410 38946
rect 28814 38894 28866 38946
rect 32286 38894 32338 38946
rect 33966 38894 34018 38946
rect 34078 38894 34130 38946
rect 36878 38894 36930 38946
rect 38446 38894 38498 38946
rect 39678 38894 39730 38946
rect 41806 38894 41858 38946
rect 45502 38894 45554 38946
rect 47518 38894 47570 38946
rect 4622 38782 4674 38834
rect 5294 38782 5346 38834
rect 9438 38782 9490 38834
rect 10222 38782 10274 38834
rect 11790 38782 11842 38834
rect 12798 38782 12850 38834
rect 13694 38782 13746 38834
rect 14814 38782 14866 38834
rect 15374 38782 15426 38834
rect 16382 38782 16434 38834
rect 17390 38782 17442 38834
rect 18510 38782 18562 38834
rect 18846 38782 18898 38834
rect 19182 38782 19234 38834
rect 20414 38782 20466 38834
rect 21758 38782 21810 38834
rect 22990 38782 23042 38834
rect 23214 38782 23266 38834
rect 23998 38782 24050 38834
rect 24558 38782 24610 38834
rect 28142 38782 28194 38834
rect 29150 38782 29202 38834
rect 30942 38782 30994 38834
rect 31726 38782 31778 38834
rect 33742 38782 33794 38834
rect 34302 38782 34354 38834
rect 37550 38782 37602 38834
rect 39006 38782 39058 38834
rect 41134 38782 41186 38834
rect 45950 38782 46002 38834
rect 48078 38782 48130 38834
rect 1710 38670 1762 38722
rect 3838 38670 3890 38722
rect 5070 38670 5122 38722
rect 5742 38670 5794 38722
rect 7534 38670 7586 38722
rect 10110 38670 10162 38722
rect 13918 38670 13970 38722
rect 19630 38670 19682 38722
rect 19742 38670 19794 38722
rect 21310 38670 21362 38722
rect 22094 38670 22146 38722
rect 25230 38670 25282 38722
rect 31502 38670 31554 38722
rect 34750 38670 34802 38722
rect 38110 38670 38162 38722
rect 40350 38670 40402 38722
rect 43934 38670 43986 38722
rect 4958 38558 5010 38610
rect 39566 38558 39618 38610
rect 39902 38558 39954 38610
rect 4478 38390 4530 38442
rect 4582 38390 4634 38442
rect 4686 38390 4738 38442
rect 35198 38390 35250 38442
rect 35302 38390 35354 38442
rect 35406 38390 35458 38442
rect 8094 38222 8146 38274
rect 12686 38222 12738 38274
rect 17838 38222 17890 38274
rect 22430 38222 22482 38274
rect 24558 38222 24610 38274
rect 24894 38222 24946 38274
rect 36094 38222 36146 38274
rect 42030 38222 42082 38274
rect 43822 38222 43874 38274
rect 43934 38222 43986 38274
rect 44158 38222 44210 38274
rect 3950 38110 4002 38162
rect 6414 38110 6466 38162
rect 8654 38110 8706 38162
rect 9998 38110 10050 38162
rect 11230 38110 11282 38162
rect 15262 38110 15314 38162
rect 16494 38110 16546 38162
rect 18398 38110 18450 38162
rect 24334 38110 24386 38162
rect 26014 38110 26066 38162
rect 28366 38110 28418 38162
rect 29262 38110 29314 38162
rect 31390 38110 31442 38162
rect 33070 38110 33122 38162
rect 34862 38110 34914 38162
rect 39454 38110 39506 38162
rect 41582 38110 41634 38162
rect 42366 38110 42418 38162
rect 2606 37998 2658 38050
rect 3502 37998 3554 38050
rect 4510 37998 4562 38050
rect 6190 37998 6242 38050
rect 6526 37998 6578 38050
rect 6862 37998 6914 38050
rect 7310 37998 7362 38050
rect 8430 37998 8482 38050
rect 9102 37998 9154 38050
rect 9886 37998 9938 38050
rect 10782 37998 10834 38050
rect 12014 37998 12066 38050
rect 12686 37998 12738 38050
rect 14254 37998 14306 38050
rect 14366 37998 14418 38050
rect 15150 37998 15202 38050
rect 16158 37998 16210 38050
rect 17166 37998 17218 38050
rect 18174 37998 18226 38050
rect 20078 37998 20130 38050
rect 20526 37998 20578 38050
rect 21646 37998 21698 38050
rect 23102 37998 23154 38050
rect 26126 37998 26178 38050
rect 29150 37998 29202 38050
rect 30158 37998 30210 38050
rect 32174 37998 32226 38050
rect 32398 37998 32450 38050
rect 33630 37998 33682 38050
rect 34750 37998 34802 38050
rect 35534 37998 35586 38050
rect 36206 37998 36258 38050
rect 36990 37998 37042 38050
rect 38782 37998 38834 38050
rect 42814 37998 42866 38050
rect 46062 37998 46114 38050
rect 46846 37998 46898 38050
rect 47630 37998 47682 38050
rect 2046 37886 2098 37938
rect 7422 37886 7474 37938
rect 9662 37886 9714 37938
rect 13694 37886 13746 37938
rect 15822 37886 15874 37938
rect 16270 37886 16322 37938
rect 19182 37886 19234 37938
rect 19294 37886 19346 37938
rect 20750 37886 20802 37938
rect 22094 37886 22146 37938
rect 23326 37886 23378 37938
rect 24110 37886 24162 37938
rect 29262 37886 29314 37938
rect 30606 37886 30658 37938
rect 30942 37886 30994 37938
rect 34302 37886 34354 37938
rect 36094 37886 36146 37938
rect 44270 37886 44322 37938
rect 45390 37886 45442 37938
rect 4174 37774 4226 37826
rect 4398 37774 4450 37826
rect 4958 37774 5010 37826
rect 7198 37774 7250 37826
rect 7646 37774 7698 37826
rect 13918 37774 13970 37826
rect 14142 37774 14194 37826
rect 18846 37774 18898 37826
rect 19518 37774 19570 37826
rect 19742 37774 19794 37826
rect 21422 37774 21474 37826
rect 21534 37774 21586 37826
rect 22318 37774 22370 37826
rect 25678 37774 25730 37826
rect 25902 37774 25954 37826
rect 26574 37774 26626 37826
rect 33406 37774 33458 37826
rect 33518 37774 33570 37826
rect 33854 37774 33906 37826
rect 37550 37774 37602 37826
rect 37886 37774 37938 37826
rect 38222 37774 38274 37826
rect 46062 37774 46114 37826
rect 19838 37606 19890 37658
rect 19942 37606 19994 37658
rect 20046 37606 20098 37658
rect 8766 37438 8818 37490
rect 8878 37438 8930 37490
rect 10222 37438 10274 37490
rect 19854 37438 19906 37490
rect 20190 37438 20242 37490
rect 21198 37438 21250 37490
rect 21646 37438 21698 37490
rect 22990 37438 23042 37490
rect 23550 37438 23602 37490
rect 24782 37438 24834 37490
rect 25454 37438 25506 37490
rect 26014 37438 26066 37490
rect 28030 37438 28082 37490
rect 36094 37438 36146 37490
rect 37886 37438 37938 37490
rect 38222 37438 38274 37490
rect 38558 37438 38610 37490
rect 39230 37438 39282 37490
rect 41918 37438 41970 37490
rect 2830 37326 2882 37378
rect 2942 37326 2994 37378
rect 3390 37326 3442 37378
rect 5854 37326 5906 37378
rect 10334 37326 10386 37378
rect 10782 37326 10834 37378
rect 11902 37326 11954 37378
rect 12574 37326 12626 37378
rect 14478 37326 14530 37378
rect 15150 37326 15202 37378
rect 20862 37326 20914 37378
rect 21086 37326 21138 37378
rect 25342 37326 25394 37378
rect 27806 37326 27858 37378
rect 28814 37326 28866 37378
rect 33630 37326 33682 37378
rect 34638 37326 34690 37378
rect 41470 37326 41522 37378
rect 42366 37326 42418 37378
rect 43598 37326 43650 37378
rect 44606 37326 44658 37378
rect 47182 37326 47234 37378
rect 3726 37214 3778 37266
rect 4398 37214 4450 37266
rect 5182 37214 5234 37266
rect 8206 37214 8258 37266
rect 8654 37214 8706 37266
rect 9662 37214 9714 37266
rect 11006 37214 11058 37266
rect 11566 37214 11618 37266
rect 12350 37214 12402 37266
rect 14702 37214 14754 37266
rect 15374 37214 15426 37266
rect 16270 37214 16322 37266
rect 17950 37214 18002 37266
rect 18286 37214 18338 37266
rect 18398 37214 18450 37266
rect 18734 37214 18786 37266
rect 19182 37214 19234 37266
rect 19294 37214 19346 37266
rect 19742 37214 19794 37266
rect 19966 37214 20018 37266
rect 20526 37214 20578 37266
rect 21870 37214 21922 37266
rect 22318 37214 22370 37266
rect 23438 37214 23490 37266
rect 23662 37214 23714 37266
rect 23998 37214 24050 37266
rect 25230 37214 25282 37266
rect 26462 37214 26514 37266
rect 27694 37214 27746 37266
rect 29374 37214 29426 37266
rect 30046 37214 30098 37266
rect 32510 37214 32562 37266
rect 32958 37214 33010 37266
rect 33294 37214 33346 37266
rect 34750 37214 34802 37266
rect 35646 37214 35698 37266
rect 38894 37214 38946 37266
rect 39790 37214 39842 37266
rect 41582 37214 41634 37266
rect 42142 37214 42194 37266
rect 42702 37214 42754 37266
rect 43822 37214 43874 37266
rect 47070 37214 47122 37266
rect 47966 37214 48018 37266
rect 3502 37102 3554 37154
rect 7982 37102 8034 37154
rect 16046 37102 16098 37154
rect 16718 37102 16770 37154
rect 18958 37102 19010 37154
rect 21758 37102 21810 37154
rect 27470 37102 27522 37154
rect 30718 37102 30770 37154
rect 33182 37102 33234 37154
rect 40238 37102 40290 37154
rect 42926 37102 42978 37154
rect 46734 37102 46786 37154
rect 47182 37102 47234 37154
rect 2830 36990 2882 37042
rect 10110 36990 10162 37042
rect 22654 36990 22706 37042
rect 22878 36990 22930 37042
rect 22990 36990 23042 37042
rect 25790 36990 25842 37042
rect 26574 36990 26626 37042
rect 41470 36990 41522 37042
rect 42254 36990 42306 37042
rect 43150 36990 43202 37042
rect 4478 36822 4530 36874
rect 4582 36822 4634 36874
rect 4686 36822 4738 36874
rect 35198 36822 35250 36874
rect 35302 36822 35354 36874
rect 35406 36822 35458 36874
rect 4958 36654 5010 36706
rect 20302 36654 20354 36706
rect 24670 36654 24722 36706
rect 25678 36654 25730 36706
rect 26798 36654 26850 36706
rect 30158 36654 30210 36706
rect 34526 36654 34578 36706
rect 34862 36654 34914 36706
rect 36094 36654 36146 36706
rect 4622 36542 4674 36594
rect 5070 36542 5122 36594
rect 5742 36542 5794 36594
rect 6190 36542 6242 36594
rect 7086 36542 7138 36594
rect 11006 36542 11058 36594
rect 12462 36542 12514 36594
rect 18398 36542 18450 36594
rect 18846 36542 18898 36594
rect 21982 36542 22034 36594
rect 23326 36542 23378 36594
rect 24222 36542 24274 36594
rect 25566 36542 25618 36594
rect 27582 36542 27634 36594
rect 28366 36542 28418 36594
rect 29486 36542 29538 36594
rect 34190 36542 34242 36594
rect 38558 36542 38610 36594
rect 41806 36542 41858 36594
rect 47742 36542 47794 36594
rect 1822 36430 1874 36482
rect 6638 36430 6690 36482
rect 8542 36430 8594 36482
rect 10670 36430 10722 36482
rect 13582 36430 13634 36482
rect 15262 36430 15314 36482
rect 17278 36430 17330 36482
rect 18286 36430 18338 36482
rect 18510 36430 18562 36482
rect 19406 36430 19458 36482
rect 20078 36430 20130 36482
rect 21422 36430 21474 36482
rect 22318 36430 22370 36482
rect 22878 36430 22930 36482
rect 23550 36430 23602 36482
rect 27022 36430 27074 36482
rect 27806 36430 27858 36482
rect 29598 36430 29650 36482
rect 31278 36430 31330 36482
rect 32062 36430 32114 36482
rect 35198 36430 35250 36482
rect 35534 36430 35586 36482
rect 38894 36430 38946 36482
rect 42254 36430 42306 36482
rect 42814 36430 42866 36482
rect 47294 36430 47346 36482
rect 47630 36430 47682 36482
rect 47854 36430 47906 36482
rect 2494 36318 2546 36370
rect 10446 36318 10498 36370
rect 11678 36318 11730 36370
rect 13470 36318 13522 36370
rect 17614 36318 17666 36370
rect 18062 36318 18114 36370
rect 21534 36318 21586 36370
rect 24670 36318 24722 36370
rect 24782 36318 24834 36370
rect 25230 36318 25282 36370
rect 34750 36318 34802 36370
rect 35310 36318 35362 36370
rect 36318 36318 36370 36370
rect 39678 36318 39730 36370
rect 42142 36318 42194 36370
rect 46622 36318 46674 36370
rect 8318 36206 8370 36258
rect 9886 36206 9938 36258
rect 11006 36206 11058 36258
rect 11230 36206 11282 36258
rect 13694 36206 13746 36258
rect 20638 36206 20690 36258
rect 30718 36206 30770 36258
rect 36206 36206 36258 36258
rect 37102 36206 37154 36258
rect 45726 36206 45778 36258
rect 46958 36206 47010 36258
rect 19838 36038 19890 36090
rect 19942 36038 19994 36090
rect 20046 36038 20098 36090
rect 3726 35870 3778 35922
rect 4734 35870 4786 35922
rect 8206 35870 8258 35922
rect 8990 35870 9042 35922
rect 12574 35870 12626 35922
rect 16494 35870 16546 35922
rect 19406 35870 19458 35922
rect 22430 35870 22482 35922
rect 47406 35870 47458 35922
rect 4286 35758 4338 35810
rect 7086 35758 7138 35810
rect 10110 35758 10162 35810
rect 13022 35758 13074 35810
rect 16718 35758 16770 35810
rect 17502 35758 17554 35810
rect 21534 35758 21586 35810
rect 22542 35758 22594 35810
rect 26014 35758 26066 35810
rect 27134 35758 27186 35810
rect 29598 35758 29650 35810
rect 37774 35758 37826 35810
rect 39902 35758 39954 35810
rect 40126 35758 40178 35810
rect 47630 35758 47682 35810
rect 2942 35646 2994 35698
rect 4062 35646 4114 35698
rect 6190 35646 6242 35698
rect 8766 35646 8818 35698
rect 9886 35646 9938 35698
rect 10334 35646 10386 35698
rect 11006 35646 11058 35698
rect 11678 35646 11730 35698
rect 12014 35646 12066 35698
rect 13358 35646 13410 35698
rect 14254 35646 14306 35698
rect 15822 35646 15874 35698
rect 16830 35646 16882 35698
rect 17390 35646 17442 35698
rect 18622 35646 18674 35698
rect 20414 35646 20466 35698
rect 20638 35646 20690 35698
rect 21086 35646 21138 35698
rect 21870 35646 21922 35698
rect 22206 35646 22258 35698
rect 22990 35646 23042 35698
rect 24110 35646 24162 35698
rect 25790 35646 25842 35698
rect 28590 35646 28642 35698
rect 28926 35646 28978 35698
rect 29486 35646 29538 35698
rect 31166 35646 31218 35698
rect 31502 35646 31554 35698
rect 31726 35646 31778 35698
rect 38558 35646 38610 35698
rect 38894 35646 38946 35698
rect 42702 35646 42754 35698
rect 46286 35646 46338 35698
rect 2270 35534 2322 35586
rect 3054 35534 3106 35586
rect 5518 35534 5570 35586
rect 7646 35534 7698 35586
rect 10894 35534 10946 35586
rect 17502 35534 17554 35586
rect 18174 35534 18226 35586
rect 20750 35534 20802 35586
rect 23662 35534 23714 35586
rect 28366 35534 28418 35586
rect 29710 35534 29762 35586
rect 30830 35534 30882 35586
rect 31614 35534 31666 35586
rect 34414 35534 34466 35586
rect 35646 35534 35698 35586
rect 39342 35534 39394 35586
rect 39790 35534 39842 35586
rect 43374 35534 43426 35586
rect 45502 35534 45554 35586
rect 46062 35534 46114 35586
rect 47294 35534 47346 35586
rect 9662 35422 9714 35474
rect 10446 35422 10498 35474
rect 24110 35422 24162 35474
rect 45950 35422 46002 35474
rect 4478 35254 4530 35306
rect 4582 35254 4634 35306
rect 4686 35254 4738 35306
rect 35198 35254 35250 35306
rect 35302 35254 35354 35306
rect 35406 35254 35458 35306
rect 2606 35086 2658 35138
rect 4398 35086 4450 35138
rect 6526 35086 6578 35138
rect 11006 35086 11058 35138
rect 11342 35086 11394 35138
rect 18846 35086 18898 35138
rect 29374 35086 29426 35138
rect 2830 34974 2882 35026
rect 14478 34974 14530 35026
rect 16382 34974 16434 35026
rect 18510 34974 18562 35026
rect 20526 34974 20578 35026
rect 21422 34974 21474 35026
rect 23550 34974 23602 35026
rect 25118 34974 25170 35026
rect 28030 34974 28082 35026
rect 29150 34974 29202 35026
rect 33182 34974 33234 35026
rect 33630 34974 33682 35026
rect 43822 34974 43874 35026
rect 46062 34974 46114 35026
rect 48190 34974 48242 35026
rect 2942 34862 2994 34914
rect 4958 34862 5010 34914
rect 5854 34862 5906 34914
rect 6414 34862 6466 34914
rect 7198 34862 7250 34914
rect 7758 34862 7810 34914
rect 8766 34862 8818 34914
rect 9998 34862 10050 34914
rect 11678 34862 11730 34914
rect 12126 34862 12178 34914
rect 12910 34862 12962 34914
rect 13806 34862 13858 34914
rect 14142 34862 14194 34914
rect 15710 34862 15762 34914
rect 19406 34862 19458 34914
rect 19630 34862 19682 34914
rect 22766 34862 22818 34914
rect 23214 34862 23266 34914
rect 25342 34862 25394 34914
rect 27582 34862 27634 34914
rect 27918 34862 27970 34914
rect 29710 34862 29762 34914
rect 30382 34862 30434 34914
rect 36990 34862 37042 34914
rect 37438 34862 37490 34914
rect 38446 34862 38498 34914
rect 44046 34862 44098 34914
rect 44270 34862 44322 34914
rect 45390 34862 45442 34914
rect 3614 34750 3666 34802
rect 4174 34750 4226 34802
rect 5070 34750 5122 34802
rect 7422 34750 7474 34802
rect 8654 34750 8706 34802
rect 12798 34750 12850 34802
rect 15038 34750 15090 34802
rect 15374 34750 15426 34802
rect 19294 34750 19346 34802
rect 21310 34750 21362 34802
rect 31054 34750 31106 34802
rect 38782 34750 38834 34802
rect 39118 34750 39170 34802
rect 43150 34750 43202 34802
rect 43710 34750 43762 34802
rect 2382 34638 2434 34690
rect 3278 34638 3330 34690
rect 3502 34638 3554 34690
rect 4286 34638 4338 34690
rect 4846 34638 4898 34690
rect 13806 34638 13858 34690
rect 15150 34638 15202 34690
rect 19966 34638 20018 34690
rect 21534 34638 21586 34690
rect 21758 34638 21810 34690
rect 28702 34638 28754 34690
rect 37886 34638 37938 34690
rect 39566 34638 39618 34690
rect 43262 34638 43314 34690
rect 43486 34638 43538 34690
rect 19838 34470 19890 34522
rect 19942 34470 19994 34522
rect 20046 34470 20098 34522
rect 7198 34302 7250 34354
rect 7422 34302 7474 34354
rect 8878 34302 8930 34354
rect 10782 34302 10834 34354
rect 13694 34302 13746 34354
rect 21870 34302 21922 34354
rect 24222 34302 24274 34354
rect 25454 34302 25506 34354
rect 25566 34302 25618 34354
rect 25678 34302 25730 34354
rect 25790 34302 25842 34354
rect 29374 34302 29426 34354
rect 31054 34302 31106 34354
rect 31950 34302 32002 34354
rect 36094 34302 36146 34354
rect 3390 34190 3442 34242
rect 4846 34190 4898 34242
rect 7534 34190 7586 34242
rect 8318 34190 8370 34242
rect 11342 34190 11394 34242
rect 14254 34190 14306 34242
rect 15598 34190 15650 34242
rect 15934 34190 15986 34242
rect 16718 34190 16770 34242
rect 17278 34190 17330 34242
rect 17838 34190 17890 34242
rect 18174 34190 18226 34242
rect 19966 34190 20018 34242
rect 20638 34190 20690 34242
rect 26014 34190 26066 34242
rect 30046 34190 30098 34242
rect 31278 34190 31330 34242
rect 31502 34190 31554 34242
rect 31838 34190 31890 34242
rect 33070 34190 33122 34242
rect 34862 34190 34914 34242
rect 37326 34190 37378 34242
rect 3614 34078 3666 34130
rect 4062 34078 4114 34130
rect 8206 34078 8258 34130
rect 8990 34078 9042 34130
rect 10558 34078 10610 34130
rect 12238 34078 12290 34130
rect 15262 34078 15314 34130
rect 15710 34078 15762 34130
rect 17502 34078 17554 34130
rect 19406 34078 19458 34130
rect 20526 34078 20578 34130
rect 22318 34078 22370 34130
rect 23102 34078 23154 34130
rect 24110 34078 24162 34130
rect 24334 34078 24386 34130
rect 24670 34078 24722 34130
rect 26574 34078 26626 34130
rect 28366 34078 28418 34130
rect 29262 34078 29314 34130
rect 29598 34078 29650 34130
rect 30830 34078 30882 34130
rect 33742 34078 33794 34130
rect 34526 34078 34578 34130
rect 34750 34078 34802 34130
rect 35086 34078 35138 34130
rect 37214 34078 37266 34130
rect 41022 34078 41074 34130
rect 44046 34078 44098 34130
rect 44382 34078 44434 34130
rect 44606 34078 44658 34130
rect 45390 34078 45442 34130
rect 6974 33966 7026 34018
rect 13470 33966 13522 34018
rect 19182 33966 19234 34018
rect 20862 33966 20914 34018
rect 21310 33966 21362 34018
rect 22542 33966 22594 34018
rect 23214 33966 23266 34018
rect 26350 33966 26402 34018
rect 28478 33966 28530 34018
rect 28814 33966 28866 34018
rect 33854 33966 33906 34018
rect 35534 33966 35586 34018
rect 41694 33966 41746 34018
rect 43822 33966 43874 34018
rect 44270 33966 44322 34018
rect 46062 33966 46114 34018
rect 48190 33966 48242 34018
rect 21534 33854 21586 33906
rect 26910 33854 26962 33906
rect 29822 33854 29874 33906
rect 30158 33854 30210 33906
rect 31950 33854 32002 33906
rect 37326 33854 37378 33906
rect 4478 33686 4530 33738
rect 4582 33686 4634 33738
rect 4686 33686 4738 33738
rect 35198 33686 35250 33738
rect 35302 33686 35354 33738
rect 35406 33686 35458 33738
rect 2718 33518 2770 33570
rect 3502 33518 3554 33570
rect 14030 33518 14082 33570
rect 26574 33518 26626 33570
rect 28702 33518 28754 33570
rect 30830 33518 30882 33570
rect 44942 33518 44994 33570
rect 2606 33406 2658 33458
rect 3614 33406 3666 33458
rect 5742 33406 5794 33458
rect 6638 33406 6690 33458
rect 9998 33406 10050 33458
rect 12350 33406 12402 33458
rect 18062 33406 18114 33458
rect 20302 33406 20354 33458
rect 26798 33406 26850 33458
rect 30606 33406 30658 33458
rect 33182 33406 33234 33458
rect 36430 33406 36482 33458
rect 36990 33406 37042 33458
rect 43150 33406 43202 33458
rect 3278 33294 3330 33346
rect 3726 33294 3778 33346
rect 5070 33294 5122 33346
rect 9102 33294 9154 33346
rect 10782 33294 10834 33346
rect 12462 33294 12514 33346
rect 13918 33294 13970 33346
rect 15262 33294 15314 33346
rect 17054 33294 17106 33346
rect 17390 33294 17442 33346
rect 19070 33294 19122 33346
rect 22094 33294 22146 33346
rect 22318 33294 22370 33346
rect 24782 33294 24834 33346
rect 25230 33294 25282 33346
rect 25678 33294 25730 33346
rect 26350 33294 26402 33346
rect 27470 33294 27522 33346
rect 27806 33294 27858 33346
rect 28254 33294 28306 33346
rect 29934 33294 29986 33346
rect 31054 33294 31106 33346
rect 32286 33294 32338 33346
rect 32734 33294 32786 33346
rect 33630 33294 33682 33346
rect 39902 33294 39954 33346
rect 40350 33294 40402 33346
rect 43934 33294 43986 33346
rect 45726 33294 45778 33346
rect 46174 33294 46226 33346
rect 46622 33294 46674 33346
rect 2494 33182 2546 33234
rect 4734 33182 4786 33234
rect 7422 33182 7474 33234
rect 8878 33182 8930 33234
rect 10670 33182 10722 33234
rect 12910 33182 12962 33234
rect 16046 33182 16098 33234
rect 17950 33182 18002 33234
rect 20302 33182 20354 33234
rect 20750 33182 20802 33234
rect 22878 33182 22930 33234
rect 27918 33182 27970 33234
rect 28142 33182 28194 33234
rect 29150 33182 29202 33234
rect 34302 33182 34354 33234
rect 39118 33182 39170 33234
rect 41022 33182 41074 33234
rect 43598 33182 43650 33234
rect 44830 33182 44882 33234
rect 44942 33182 44994 33234
rect 46398 33182 46450 33234
rect 46846 33182 46898 33234
rect 46958 33182 47010 33234
rect 4846 33070 4898 33122
rect 6302 33070 6354 33122
rect 7086 33070 7138 33122
rect 7758 33070 7810 33122
rect 8318 33070 8370 33122
rect 9662 33070 9714 33122
rect 13694 33070 13746 33122
rect 14030 33070 14082 33122
rect 15150 33070 15202 33122
rect 20526 33070 20578 33122
rect 23774 33070 23826 33122
rect 24446 33070 24498 33122
rect 29486 33070 29538 33122
rect 31838 33070 31890 33122
rect 43710 33070 43762 33122
rect 46062 33070 46114 33122
rect 47630 33070 47682 33122
rect 47854 33070 47906 33122
rect 48190 33070 48242 33122
rect 19838 32902 19890 32954
rect 19942 32902 19994 32954
rect 20046 32902 20098 32954
rect 5070 32734 5122 32786
rect 6974 32734 7026 32786
rect 8878 32734 8930 32786
rect 17726 32734 17778 32786
rect 20862 32734 20914 32786
rect 20974 32734 21026 32786
rect 33406 32734 33458 32786
rect 34638 32734 34690 32786
rect 35758 32734 35810 32786
rect 37550 32734 37602 32786
rect 40014 32734 40066 32786
rect 43822 32734 43874 32786
rect 45390 32734 45442 32786
rect 45614 32734 45666 32786
rect 46958 32734 47010 32786
rect 9774 32622 9826 32674
rect 10894 32622 10946 32674
rect 13134 32622 13186 32674
rect 19182 32622 19234 32674
rect 21198 32622 21250 32674
rect 21310 32622 21362 32674
rect 30158 32622 30210 32674
rect 33294 32622 33346 32674
rect 33854 32622 33906 32674
rect 34078 32622 34130 32674
rect 34750 32622 34802 32674
rect 35870 32622 35922 32674
rect 37438 32622 37490 32674
rect 41246 32622 41298 32674
rect 43486 32622 43538 32674
rect 43598 32622 43650 32674
rect 44046 32622 44098 32674
rect 44830 32622 44882 32674
rect 44942 32622 44994 32674
rect 45278 32622 45330 32674
rect 47406 32622 47458 32674
rect 47518 32622 47570 32674
rect 3838 32510 3890 32562
rect 4622 32510 4674 32562
rect 6078 32510 6130 32562
rect 6190 32510 6242 32562
rect 6526 32510 6578 32562
rect 8990 32510 9042 32562
rect 9998 32510 10050 32562
rect 11006 32510 11058 32562
rect 11342 32510 11394 32562
rect 12350 32510 12402 32562
rect 13582 32510 13634 32562
rect 14926 32510 14978 32562
rect 16606 32510 16658 32562
rect 18622 32510 18674 32562
rect 19630 32510 19682 32562
rect 20190 32510 20242 32562
rect 20414 32510 20466 32562
rect 22094 32510 22146 32562
rect 22654 32510 22706 32562
rect 22990 32510 23042 32562
rect 23214 32510 23266 32562
rect 24558 32510 24610 32562
rect 25566 32510 25618 32562
rect 26574 32510 26626 32562
rect 28366 32510 28418 32562
rect 29038 32510 29090 32562
rect 31054 32510 31106 32562
rect 32398 32510 32450 32562
rect 37774 32510 37826 32562
rect 39678 32510 39730 32562
rect 40238 32510 40290 32562
rect 44270 32510 44322 32562
rect 44606 32510 44658 32562
rect 46734 32510 46786 32562
rect 47070 32510 47122 32562
rect 1710 32398 1762 32450
rect 6414 32398 6466 32450
rect 7758 32398 7810 32450
rect 7982 32398 8034 32450
rect 8430 32398 8482 32450
rect 10894 32398 10946 32450
rect 11678 32398 11730 32450
rect 12014 32398 12066 32450
rect 16494 32398 16546 32450
rect 18286 32398 18338 32450
rect 21982 32398 22034 32450
rect 25902 32398 25954 32450
rect 29598 32398 29650 32450
rect 31726 32398 31778 32450
rect 32062 32398 32114 32450
rect 32286 32398 32338 32450
rect 34190 32398 34242 32450
rect 36654 32398 36706 32450
rect 7422 32286 7474 32338
rect 8878 32286 8930 32338
rect 15374 32286 15426 32338
rect 18062 32286 18114 32338
rect 23438 32286 23490 32338
rect 24222 32286 24274 32338
rect 24558 32286 24610 32338
rect 33406 32286 33458 32338
rect 34526 32286 34578 32338
rect 39902 32286 39954 32338
rect 41470 32286 41522 32338
rect 41806 32286 41858 32338
rect 47518 32286 47570 32338
rect 4478 32118 4530 32170
rect 4582 32118 4634 32170
rect 4686 32118 4738 32170
rect 35198 32118 35250 32170
rect 35302 32118 35354 32170
rect 35406 32118 35458 32170
rect 8878 31950 8930 32002
rect 19966 31950 20018 32002
rect 20190 31950 20242 32002
rect 23998 31950 24050 32002
rect 25454 31950 25506 32002
rect 28478 31950 28530 32002
rect 33406 31950 33458 32002
rect 34862 31950 34914 32002
rect 4958 31838 5010 31890
rect 7310 31838 7362 31890
rect 7870 31838 7922 31890
rect 11006 31838 11058 31890
rect 14366 31838 14418 31890
rect 16158 31838 16210 31890
rect 16942 31838 16994 31890
rect 20414 31838 20466 31890
rect 20750 31838 20802 31890
rect 21534 31838 21586 31890
rect 25230 31838 25282 31890
rect 29150 31838 29202 31890
rect 30158 31838 30210 31890
rect 32286 31838 32338 31890
rect 35758 31838 35810 31890
rect 38222 31838 38274 31890
rect 44158 31838 44210 31890
rect 48190 31838 48242 31890
rect 2606 31726 2658 31778
rect 4174 31726 4226 31778
rect 5742 31726 5794 31778
rect 6190 31726 6242 31778
rect 6414 31726 6466 31778
rect 6862 31726 6914 31778
rect 8318 31726 8370 31778
rect 9214 31726 9266 31778
rect 9774 31726 9826 31778
rect 9886 31726 9938 31778
rect 12462 31726 12514 31778
rect 14254 31726 14306 31778
rect 15038 31726 15090 31778
rect 16830 31726 16882 31778
rect 18286 31726 18338 31778
rect 20638 31726 20690 31778
rect 21982 31726 22034 31778
rect 22990 31726 23042 31778
rect 23438 31726 23490 31778
rect 23774 31726 23826 31778
rect 26798 31726 26850 31778
rect 28254 31726 28306 31778
rect 29598 31726 29650 31778
rect 33070 31726 33122 31778
rect 36094 31726 36146 31778
rect 38110 31726 38162 31778
rect 41358 31726 41410 31778
rect 45390 31726 45442 31778
rect 2046 31614 2098 31666
rect 3726 31614 3778 31666
rect 4510 31614 4562 31666
rect 9438 31614 9490 31666
rect 13582 31614 13634 31666
rect 16270 31614 16322 31666
rect 17502 31614 17554 31666
rect 21310 31614 21362 31666
rect 22430 31614 22482 31666
rect 22766 31614 22818 31666
rect 25678 31614 25730 31666
rect 28030 31614 28082 31666
rect 33742 31614 33794 31666
rect 34302 31614 34354 31666
rect 35198 31614 35250 31666
rect 37774 31614 37826 31666
rect 38334 31614 38386 31666
rect 38670 31614 38722 31666
rect 42030 31614 42082 31666
rect 46062 31614 46114 31666
rect 3614 31502 3666 31554
rect 4398 31502 4450 31554
rect 6302 31502 6354 31554
rect 15710 31502 15762 31554
rect 16046 31502 16098 31554
rect 33518 31502 33570 31554
rect 33966 31502 34018 31554
rect 34190 31502 34242 31554
rect 34974 31502 35026 31554
rect 37438 31502 37490 31554
rect 39006 31502 39058 31554
rect 19838 31334 19890 31386
rect 19942 31334 19994 31386
rect 20046 31334 20098 31386
rect 3390 31166 3442 31218
rect 7310 31166 7362 31218
rect 7534 31166 7586 31218
rect 7982 31166 8034 31218
rect 8990 31166 9042 31218
rect 9886 31166 9938 31218
rect 11230 31166 11282 31218
rect 15374 31166 15426 31218
rect 18510 31166 18562 31218
rect 30942 31166 30994 31218
rect 36990 31166 37042 31218
rect 37214 31166 37266 31218
rect 38110 31166 38162 31218
rect 39678 31166 39730 31218
rect 42478 31166 42530 31218
rect 43822 31166 43874 31218
rect 44494 31166 44546 31218
rect 44718 31166 44770 31218
rect 45278 31166 45330 31218
rect 46958 31166 47010 31218
rect 47854 31166 47906 31218
rect 2718 31054 2770 31106
rect 2942 31054 2994 31106
rect 4958 31054 5010 31106
rect 7646 31054 7698 31106
rect 10222 31054 10274 31106
rect 11790 31054 11842 31106
rect 14590 31054 14642 31106
rect 15038 31054 15090 31106
rect 15150 31054 15202 31106
rect 20974 31054 21026 31106
rect 24558 31054 24610 31106
rect 28590 31054 28642 31106
rect 31278 31054 31330 31106
rect 31614 31054 31666 31106
rect 32398 31054 32450 31106
rect 32510 31054 32562 31106
rect 39230 31054 39282 31106
rect 41358 31054 41410 31106
rect 42814 31054 42866 31106
rect 43710 31054 43762 31106
rect 44046 31054 44098 31106
rect 44830 31054 44882 31106
rect 46398 31054 46450 31106
rect 47182 31054 47234 31106
rect 2382 30942 2434 30994
rect 3278 30942 3330 30994
rect 3502 30942 3554 30994
rect 3950 30942 4002 30994
rect 4286 30942 4338 30994
rect 9550 30942 9602 30994
rect 10782 30942 10834 30994
rect 11118 30942 11170 30994
rect 12350 30942 12402 30994
rect 12798 30942 12850 30994
rect 13470 30942 13522 30994
rect 13582 30942 13634 30994
rect 16606 30942 16658 30994
rect 17390 30942 17442 30994
rect 17950 30942 18002 30994
rect 18846 30942 18898 30994
rect 20078 30942 20130 30994
rect 20526 30942 20578 30994
rect 20638 30942 20690 30994
rect 21534 30942 21586 30994
rect 23886 30942 23938 30994
rect 25230 30942 25282 30994
rect 31838 30942 31890 30994
rect 33182 30942 33234 30994
rect 33854 30942 33906 30994
rect 37438 30942 37490 30994
rect 37662 30942 37714 30994
rect 38222 30942 38274 30994
rect 38334 30942 38386 30994
rect 38670 30942 38722 30994
rect 39006 30942 39058 30994
rect 41694 30942 41746 30994
rect 44270 30942 44322 30994
rect 45502 30942 45554 30994
rect 46062 30942 46114 30994
rect 46734 30942 46786 30994
rect 47294 30942 47346 30994
rect 47742 30942 47794 30994
rect 2494 30830 2546 30882
rect 7086 30830 7138 30882
rect 8542 30830 8594 30882
rect 12462 30830 12514 30882
rect 18622 30830 18674 30882
rect 19630 30830 19682 30882
rect 20862 30830 20914 30882
rect 21870 30830 21922 30882
rect 24670 30830 24722 30882
rect 35982 30830 36034 30882
rect 36542 30830 36594 30882
rect 37102 30830 37154 30882
rect 39118 30830 39170 30882
rect 39566 30830 39618 30882
rect 41582 30830 41634 30882
rect 8318 30718 8370 30770
rect 13022 30718 13074 30770
rect 15822 30718 15874 30770
rect 22318 30718 22370 30770
rect 24334 30718 24386 30770
rect 32398 30718 32450 30770
rect 47854 30718 47906 30770
rect 4478 30550 4530 30602
rect 4582 30550 4634 30602
rect 4686 30550 4738 30602
rect 35198 30550 35250 30602
rect 35302 30550 35354 30602
rect 35406 30550 35458 30602
rect 9550 30382 9602 30434
rect 22206 30382 22258 30434
rect 2494 30270 2546 30322
rect 4622 30270 4674 30322
rect 7198 30270 7250 30322
rect 9214 30270 9266 30322
rect 10558 30270 10610 30322
rect 11118 30270 11170 30322
rect 12686 30270 12738 30322
rect 13918 30270 13970 30322
rect 18958 30270 19010 30322
rect 27022 30270 27074 30322
rect 29038 30270 29090 30322
rect 33630 30270 33682 30322
rect 34862 30270 34914 30322
rect 35758 30270 35810 30322
rect 37550 30270 37602 30322
rect 39678 30270 39730 30322
rect 40798 30270 40850 30322
rect 1822 30158 1874 30210
rect 5182 30158 5234 30210
rect 7646 30158 7698 30210
rect 11454 30158 11506 30210
rect 12014 30158 12066 30210
rect 12574 30158 12626 30210
rect 13694 30158 13746 30210
rect 14590 30158 14642 30210
rect 15486 30158 15538 30210
rect 16046 30158 16098 30210
rect 19630 30158 19682 30210
rect 20414 30158 20466 30210
rect 20750 30158 20802 30210
rect 21422 30158 21474 30210
rect 21870 30158 21922 30210
rect 22318 30158 22370 30210
rect 22990 30158 23042 30210
rect 23550 30158 23602 30210
rect 24782 30158 24834 30210
rect 26686 30158 26738 30210
rect 28590 30158 28642 30210
rect 30158 30158 30210 30210
rect 30494 30158 30546 30210
rect 31502 30158 31554 30210
rect 31950 30158 32002 30210
rect 32398 30158 32450 30210
rect 32846 30158 32898 30210
rect 35534 30158 35586 30210
rect 40462 30158 40514 30210
rect 41022 30158 41074 30210
rect 42254 30158 42306 30210
rect 42702 30158 42754 30210
rect 43822 30158 43874 30210
rect 47070 30158 47122 30210
rect 47406 30158 47458 30210
rect 7310 30046 7362 30098
rect 8430 30046 8482 30098
rect 8990 30046 9042 30098
rect 14254 30046 14306 30098
rect 14926 30046 14978 30098
rect 16830 30046 16882 30098
rect 20078 30046 20130 30098
rect 23662 30046 23714 30098
rect 25118 30046 25170 30098
rect 28478 30046 28530 30098
rect 29486 30046 29538 30098
rect 29934 30046 29986 30098
rect 34526 30046 34578 30098
rect 46734 30046 46786 30098
rect 7086 29934 7138 29986
rect 7758 29934 7810 29986
rect 7982 29934 8034 29986
rect 23102 29934 23154 29986
rect 30942 29934 30994 29986
rect 31054 29934 31106 29986
rect 31166 29934 31218 29986
rect 33518 29934 33570 29986
rect 33742 29934 33794 29986
rect 33966 29934 34018 29986
rect 36430 29934 36482 29986
rect 41358 29934 41410 29986
rect 42030 29934 42082 29986
rect 43038 29934 43090 29986
rect 43486 29934 43538 29986
rect 43710 29934 43762 29986
rect 47182 29934 47234 29986
rect 19838 29766 19890 29818
rect 19942 29766 19994 29818
rect 20046 29766 20098 29818
rect 1710 29598 1762 29650
rect 8766 29598 8818 29650
rect 14590 29598 14642 29650
rect 16830 29598 16882 29650
rect 17502 29598 17554 29650
rect 18734 29598 18786 29650
rect 20750 29598 20802 29650
rect 24558 29598 24610 29650
rect 26686 29598 26738 29650
rect 33182 29598 33234 29650
rect 36094 29598 36146 29650
rect 7758 29486 7810 29538
rect 9662 29486 9714 29538
rect 10110 29486 10162 29538
rect 11566 29486 11618 29538
rect 12798 29486 12850 29538
rect 13694 29486 13746 29538
rect 18846 29486 18898 29538
rect 19742 29486 19794 29538
rect 24110 29486 24162 29538
rect 25790 29486 25842 29538
rect 29710 29486 29762 29538
rect 30382 29486 30434 29538
rect 30606 29486 30658 29538
rect 31278 29486 31330 29538
rect 33630 29486 33682 29538
rect 35086 29486 35138 29538
rect 42814 29486 42866 29538
rect 43150 29486 43202 29538
rect 45614 29486 45666 29538
rect 5518 29374 5570 29426
rect 6302 29374 6354 29426
rect 6862 29374 6914 29426
rect 7982 29374 8034 29426
rect 9774 29374 9826 29426
rect 11118 29374 11170 29426
rect 12014 29374 12066 29426
rect 12574 29374 12626 29426
rect 14702 29374 14754 29426
rect 16046 29374 16098 29426
rect 17390 29374 17442 29426
rect 18398 29374 18450 29426
rect 18622 29374 18674 29426
rect 19182 29374 19234 29426
rect 20974 29374 21026 29426
rect 24670 29374 24722 29426
rect 26798 29374 26850 29426
rect 27022 29374 27074 29426
rect 28590 29374 28642 29426
rect 29150 29374 29202 29426
rect 29934 29374 29986 29426
rect 31614 29374 31666 29426
rect 32510 29374 32562 29426
rect 32958 29374 33010 29426
rect 33294 29374 33346 29426
rect 34078 29374 34130 29426
rect 34526 29374 34578 29426
rect 35422 29374 35474 29426
rect 35870 29374 35922 29426
rect 36766 29374 36818 29426
rect 37102 29374 37154 29426
rect 38110 29374 38162 29426
rect 43262 29374 43314 29426
rect 44830 29374 44882 29426
rect 2270 29262 2322 29314
rect 5966 29262 6018 29314
rect 8430 29262 8482 29314
rect 14926 29262 14978 29314
rect 22878 29262 22930 29314
rect 28814 29262 28866 29314
rect 29262 29262 29314 29314
rect 31502 29262 31554 29314
rect 41022 29262 41074 29314
rect 42926 29262 42978 29314
rect 44494 29262 44546 29314
rect 47742 29262 47794 29314
rect 9662 29150 9714 29202
rect 10334 29150 10386 29202
rect 40798 29150 40850 29202
rect 41022 29150 41074 29202
rect 4478 28982 4530 29034
rect 4582 28982 4634 29034
rect 4686 28982 4738 29034
rect 35198 28982 35250 29034
rect 35302 28982 35354 29034
rect 35406 28982 35458 29034
rect 6974 28814 7026 28866
rect 9550 28814 9602 28866
rect 23438 28814 23490 28866
rect 35646 28814 35698 28866
rect 35982 28814 36034 28866
rect 37550 28814 37602 28866
rect 47070 28814 47122 28866
rect 1822 28702 1874 28754
rect 4958 28702 5010 28754
rect 7198 28702 7250 28754
rect 12462 28702 12514 28754
rect 14142 28702 14194 28754
rect 16382 28702 16434 28754
rect 19854 28702 19906 28754
rect 20302 28702 20354 28754
rect 21422 28702 21474 28754
rect 22990 28702 23042 28754
rect 23998 28702 24050 28754
rect 26910 28702 26962 28754
rect 32062 28702 32114 28754
rect 34190 28702 34242 28754
rect 34974 28702 35026 28754
rect 35422 28702 35474 28754
rect 36430 28702 36482 28754
rect 42142 28702 42194 28754
rect 44270 28702 44322 28754
rect 44942 28702 44994 28754
rect 4622 28590 4674 28642
rect 4846 28590 4898 28642
rect 5182 28590 5234 28642
rect 5966 28590 6018 28642
rect 6750 28590 6802 28642
rect 8430 28590 8482 28642
rect 9438 28590 9490 28642
rect 9774 28590 9826 28642
rect 10446 28590 10498 28642
rect 11230 28590 11282 28642
rect 12910 28590 12962 28642
rect 17054 28590 17106 28642
rect 17726 28590 17778 28642
rect 17950 28590 18002 28642
rect 18174 28590 18226 28642
rect 18958 28590 19010 28642
rect 20750 28590 20802 28642
rect 21758 28590 21810 28642
rect 22430 28590 22482 28642
rect 23774 28590 23826 28642
rect 24446 28590 24498 28642
rect 26014 28590 26066 28642
rect 27022 28590 27074 28642
rect 27806 28590 27858 28642
rect 29486 28590 29538 28642
rect 30606 28590 30658 28642
rect 31390 28590 31442 28642
rect 34638 28590 34690 28642
rect 36990 28590 37042 28642
rect 37214 28590 37266 28642
rect 37886 28590 37938 28642
rect 39006 28590 39058 28642
rect 39230 28590 39282 28642
rect 41358 28590 41410 28642
rect 45726 28590 45778 28642
rect 46398 28590 46450 28642
rect 11342 28478 11394 28530
rect 17502 28478 17554 28530
rect 22878 28478 22930 28530
rect 23102 28478 23154 28530
rect 24334 28478 24386 28530
rect 29150 28478 29202 28530
rect 29822 28478 29874 28530
rect 30158 28478 30210 28530
rect 30942 28478 30994 28530
rect 39902 28478 39954 28530
rect 45950 28478 46002 28530
rect 47070 28478 47122 28530
rect 10446 28366 10498 28418
rect 11454 28366 11506 28418
rect 18398 28366 18450 28418
rect 19294 28366 19346 28418
rect 38222 28366 38274 28418
rect 46510 28366 46562 28418
rect 46734 28366 46786 28418
rect 47182 28422 47234 28474
rect 47630 28478 47682 28530
rect 47742 28478 47794 28530
rect 47406 28366 47458 28418
rect 19838 28198 19890 28250
rect 19942 28198 19994 28250
rect 20046 28198 20098 28250
rect 15038 28030 15090 28082
rect 17390 28030 17442 28082
rect 21982 28030 22034 28082
rect 22206 28030 22258 28082
rect 22430 28030 22482 28082
rect 22766 28030 22818 28082
rect 23662 28030 23714 28082
rect 32958 28030 33010 28082
rect 33070 28030 33122 28082
rect 34078 28030 34130 28082
rect 35646 28030 35698 28082
rect 40910 28030 40962 28082
rect 41918 28030 41970 28082
rect 44606 28030 44658 28082
rect 4510 27918 4562 27970
rect 10670 27918 10722 27970
rect 11230 27918 11282 27970
rect 12014 27918 12066 27970
rect 12238 27918 12290 27970
rect 12910 27918 12962 27970
rect 14030 27918 14082 27970
rect 16830 27918 16882 27970
rect 23326 27918 23378 27970
rect 23438 27918 23490 27970
rect 25566 27918 25618 27970
rect 31838 27918 31890 27970
rect 32174 27918 32226 27970
rect 42142 27918 42194 27970
rect 42814 27918 42866 27970
rect 42926 27918 42978 27970
rect 44942 27918 44994 27970
rect 4286 27806 4338 27858
rect 6414 27806 6466 27858
rect 7198 27806 7250 27858
rect 9774 27806 9826 27858
rect 10110 27806 10162 27858
rect 10894 27806 10946 27858
rect 11790 27806 11842 27858
rect 14926 27806 14978 27858
rect 15262 27806 15314 27858
rect 16494 27806 16546 27858
rect 18622 27806 18674 27858
rect 19406 27806 19458 27858
rect 21870 27806 21922 27858
rect 24334 27806 24386 27858
rect 26126 27806 26178 27858
rect 27358 27806 27410 27858
rect 27806 27806 27858 27858
rect 29710 27806 29762 27858
rect 32510 27806 32562 27858
rect 33294 27806 33346 27858
rect 33518 27806 33570 27858
rect 34750 27806 34802 27858
rect 39118 27806 39170 27858
rect 41134 27806 41186 27858
rect 41582 27806 41634 27858
rect 41694 27806 41746 27858
rect 42254 27806 42306 27858
rect 48078 27806 48130 27858
rect 6302 27694 6354 27746
rect 17838 27694 17890 27746
rect 21534 27694 21586 27746
rect 23886 27694 23938 27746
rect 26238 27694 26290 27746
rect 26910 27694 26962 27746
rect 27918 27694 27970 27746
rect 29374 27694 29426 27746
rect 30382 27694 30434 27746
rect 31278 27694 31330 27746
rect 34414 27694 34466 27746
rect 36206 27694 36258 27746
rect 38334 27694 38386 27746
rect 39566 27694 39618 27746
rect 41022 27694 41074 27746
rect 44270 27694 44322 27746
rect 45278 27694 45330 27746
rect 47406 27694 47458 27746
rect 34750 27582 34802 27634
rect 35086 27582 35138 27634
rect 42814 27582 42866 27634
rect 4478 27414 4530 27466
rect 4582 27414 4634 27466
rect 4686 27414 4738 27466
rect 35198 27414 35250 27466
rect 35302 27414 35354 27466
rect 35406 27414 35458 27466
rect 6414 27246 6466 27298
rect 8990 27246 9042 27298
rect 13806 27246 13858 27298
rect 29710 27246 29762 27298
rect 5070 27134 5122 27186
rect 19182 27190 19234 27242
rect 38222 27246 38274 27298
rect 8654 27134 8706 27186
rect 11118 27134 11170 27186
rect 13918 27134 13970 27186
rect 24334 27134 24386 27186
rect 31278 27134 31330 27186
rect 31726 27134 31778 27186
rect 33294 27134 33346 27186
rect 35422 27134 35474 27186
rect 35870 27134 35922 27186
rect 40238 27134 40290 27186
rect 42366 27134 42418 27186
rect 43598 27134 43650 27186
rect 47294 27134 47346 27186
rect 4622 27022 4674 27074
rect 6750 27022 6802 27074
rect 7086 27022 7138 27074
rect 9774 27022 9826 27074
rect 10558 27022 10610 27074
rect 12126 27022 12178 27074
rect 13694 27022 13746 27074
rect 14478 27022 14530 27074
rect 14702 27022 14754 27074
rect 16270 27022 16322 27074
rect 19518 27022 19570 27074
rect 20190 27022 20242 27074
rect 21422 27022 21474 27074
rect 26574 27022 26626 27074
rect 26798 27022 26850 27074
rect 28142 27022 28194 27074
rect 29150 27022 29202 27074
rect 30718 27022 30770 27074
rect 32622 27022 32674 27074
rect 36990 27022 37042 27074
rect 37102 27022 37154 27074
rect 37886 27022 37938 27074
rect 39566 27022 39618 27074
rect 44830 27022 44882 27074
rect 46286 27022 46338 27074
rect 47070 27022 47122 27074
rect 47518 27022 47570 27074
rect 9326 26910 9378 26962
rect 9550 26910 9602 26962
rect 12462 26910 12514 26962
rect 12910 26910 12962 26962
rect 15486 26910 15538 26962
rect 15598 26910 15650 26962
rect 15822 26910 15874 26962
rect 17054 26910 17106 26962
rect 19854 26910 19906 26962
rect 20526 26910 20578 26962
rect 22094 26910 22146 26962
rect 26014 26910 26066 26962
rect 27918 26910 27970 26962
rect 32174 26910 32226 26962
rect 38110 26910 38162 26962
rect 42926 26910 42978 26962
rect 46398 26910 46450 26962
rect 46846 26910 46898 26962
rect 47854 26910 47906 26962
rect 48190 26910 48242 26962
rect 25118 26798 25170 26850
rect 35758 26798 35810 26850
rect 35982 26798 36034 26850
rect 36206 26798 36258 26850
rect 37214 26798 37266 26850
rect 37438 26798 37490 26850
rect 43038 26798 43090 26850
rect 43262 26798 43314 26850
rect 45166 26798 45218 26850
rect 46622 26798 46674 26850
rect 19838 26630 19890 26682
rect 19942 26630 19994 26682
rect 20046 26630 20098 26682
rect 8094 26462 8146 26514
rect 9102 26462 9154 26514
rect 10110 26462 10162 26514
rect 10894 26462 10946 26514
rect 15598 26462 15650 26514
rect 15822 26462 15874 26514
rect 17950 26462 18002 26514
rect 18286 26462 18338 26514
rect 19070 26462 19122 26514
rect 19518 26462 19570 26514
rect 20302 26462 20354 26514
rect 23550 26462 23602 26514
rect 23886 26462 23938 26514
rect 26014 26462 26066 26514
rect 27470 26462 27522 26514
rect 28478 26462 28530 26514
rect 33070 26462 33122 26514
rect 34862 26462 34914 26514
rect 35198 26462 35250 26514
rect 37102 26462 37154 26514
rect 37998 26462 38050 26514
rect 39118 26462 39170 26514
rect 42366 26462 42418 26514
rect 45614 26462 45666 26514
rect 48302 26462 48354 26514
rect 7198 26350 7250 26402
rect 8990 26350 9042 26402
rect 18622 26350 18674 26402
rect 18958 26350 19010 26402
rect 20190 26350 20242 26402
rect 20862 26350 20914 26402
rect 25566 26350 25618 26402
rect 32510 26350 32562 26402
rect 39342 26350 39394 26402
rect 41022 26350 41074 26402
rect 41246 26350 41298 26402
rect 43374 26350 43426 26402
rect 43710 26350 43762 26402
rect 45278 26350 45330 26402
rect 8206 26238 8258 26290
rect 8430 26238 8482 26290
rect 8766 26238 8818 26290
rect 9550 26238 9602 26290
rect 14702 26238 14754 26290
rect 15150 26238 15202 26290
rect 15710 26238 15762 26290
rect 16606 26238 16658 26290
rect 17390 26238 17442 26290
rect 19630 26238 19682 26290
rect 20974 26238 21026 26290
rect 25342 26238 25394 26290
rect 27022 26238 27074 26290
rect 27358 26238 27410 26290
rect 28142 26238 28194 26290
rect 29262 26238 29314 26290
rect 35758 26238 35810 26290
rect 39454 26238 39506 26290
rect 41806 26238 41858 26290
rect 42590 26238 42642 26290
rect 46622 26238 46674 26290
rect 46958 26238 47010 26290
rect 47182 26238 47234 26290
rect 6414 26126 6466 26178
rect 11678 26126 11730 26178
rect 14030 26126 14082 26178
rect 16158 26126 16210 26178
rect 21758 26126 21810 26178
rect 22318 26126 22370 26178
rect 22654 26126 22706 26178
rect 23102 26126 23154 26178
rect 24670 26126 24722 26178
rect 27918 26126 27970 26178
rect 29934 26126 29986 26178
rect 32062 26126 32114 26178
rect 33518 26126 33570 26178
rect 34078 26126 34130 26178
rect 36206 26126 36258 26178
rect 36654 26126 36706 26178
rect 37550 26126 37602 26178
rect 41134 26126 41186 26178
rect 46846 26126 46898 26178
rect 19518 26014 19570 26066
rect 20302 26014 20354 26066
rect 20862 26014 20914 26066
rect 21758 26014 21810 26066
rect 23102 26014 23154 26066
rect 32398 26014 32450 26066
rect 35534 26014 35586 26066
rect 36430 26014 36482 26066
rect 37550 26014 37602 26066
rect 41582 26014 41634 26066
rect 4478 25846 4530 25898
rect 4582 25846 4634 25898
rect 4686 25846 4738 25898
rect 35198 25846 35250 25898
rect 35302 25846 35354 25898
rect 35406 25846 35458 25898
rect 18622 25678 18674 25730
rect 37438 25678 37490 25730
rect 41918 25678 41970 25730
rect 42254 25678 42306 25730
rect 10782 25566 10834 25618
rect 18286 25566 18338 25618
rect 19294 25566 19346 25618
rect 21870 25566 21922 25618
rect 23326 25566 23378 25618
rect 26126 25566 26178 25618
rect 27134 25566 27186 25618
rect 27470 25566 27522 25618
rect 28254 25566 28306 25618
rect 28590 25566 28642 25618
rect 29934 25566 29986 25618
rect 33630 25566 33682 25618
rect 34078 25566 34130 25618
rect 34526 25566 34578 25618
rect 38222 25566 38274 25618
rect 40350 25566 40402 25618
rect 46062 25566 46114 25618
rect 48190 25566 48242 25618
rect 4846 25454 4898 25506
rect 9662 25454 9714 25506
rect 10558 25454 10610 25506
rect 11790 25454 11842 25506
rect 12798 25454 12850 25506
rect 13694 25454 13746 25506
rect 14030 25454 14082 25506
rect 15374 25454 15426 25506
rect 25678 25454 25730 25506
rect 25790 25454 25842 25506
rect 26910 25454 26962 25506
rect 27694 25454 27746 25506
rect 30718 25454 30770 25506
rect 35534 25454 35586 25506
rect 36990 25454 37042 25506
rect 37214 25454 37266 25506
rect 41134 25454 41186 25506
rect 41918 25454 41970 25506
rect 43374 25454 43426 25506
rect 43486 25454 43538 25506
rect 43934 25454 43986 25506
rect 45390 25454 45442 25506
rect 4510 25342 4562 25394
rect 5070 25342 5122 25394
rect 8430 25342 8482 25394
rect 13806 25342 13858 25394
rect 14366 25342 14418 25394
rect 14926 25342 14978 25394
rect 16158 25342 16210 25394
rect 18734 25342 18786 25394
rect 19294 25342 19346 25394
rect 19406 25342 19458 25394
rect 19518 25342 19570 25394
rect 20302 25342 20354 25394
rect 20414 25342 20466 25394
rect 21646 25342 21698 25394
rect 21870 25342 21922 25394
rect 21982 25342 22034 25394
rect 22766 25342 22818 25394
rect 22878 25342 22930 25394
rect 22990 25342 23042 25394
rect 23550 25342 23602 25394
rect 23774 25342 23826 25394
rect 23886 25342 23938 25394
rect 24446 25342 24498 25394
rect 24558 25342 24610 25394
rect 29822 25342 29874 25394
rect 29934 25342 29986 25394
rect 30046 25342 30098 25394
rect 31502 25342 31554 25394
rect 34638 25342 34690 25394
rect 34862 25342 34914 25394
rect 35646 25342 35698 25394
rect 35870 25342 35922 25394
rect 35982 25342 36034 25394
rect 36430 25342 36482 25394
rect 37550 25342 37602 25394
rect 4734 25230 4786 25282
rect 6302 25230 6354 25282
rect 19070 25230 19122 25282
rect 20078 25230 20130 25282
rect 22206 25230 22258 25282
rect 22542 25230 22594 25282
rect 24782 25230 24834 25282
rect 25566 25230 25618 25282
rect 30270 25230 30322 25282
rect 36206 25230 36258 25282
rect 41582 25230 41634 25282
rect 43598 25230 43650 25282
rect 44942 25230 44994 25282
rect 19838 25062 19890 25114
rect 19942 25062 19994 25114
rect 20046 25062 20098 25114
rect 6526 24894 6578 24946
rect 9438 24894 9490 24946
rect 16046 24894 16098 24946
rect 19406 24894 19458 24946
rect 26014 24894 26066 24946
rect 26798 24894 26850 24946
rect 28590 24894 28642 24946
rect 29934 24894 29986 24946
rect 30718 24894 30770 24946
rect 31502 24894 31554 24946
rect 31614 24894 31666 24946
rect 44830 24894 44882 24946
rect 47294 24894 47346 24946
rect 47630 24894 47682 24946
rect 6974 24782 7026 24834
rect 9662 24782 9714 24834
rect 9774 24782 9826 24834
rect 11006 24782 11058 24834
rect 18174 24782 18226 24834
rect 18286 24782 18338 24834
rect 19518 24782 19570 24834
rect 19630 24782 19682 24834
rect 20526 24782 20578 24834
rect 23326 24782 23378 24834
rect 24446 24782 24498 24834
rect 24558 24782 24610 24834
rect 29710 24782 29762 24834
rect 31054 24782 31106 24834
rect 31838 24782 31890 24834
rect 33854 24782 33906 24834
rect 38446 24782 38498 24834
rect 43486 24782 43538 24834
rect 45054 24782 45106 24834
rect 45166 24782 45218 24834
rect 45614 24782 45666 24834
rect 47070 24782 47122 24834
rect 6078 24670 6130 24722
rect 7870 24670 7922 24722
rect 11454 24670 11506 24722
rect 12126 24670 12178 24722
rect 13134 24670 13186 24722
rect 17726 24670 17778 24722
rect 18510 24670 18562 24722
rect 18958 24670 19010 24722
rect 19294 24670 19346 24722
rect 20078 24670 20130 24722
rect 20302 24670 20354 24722
rect 20638 24670 20690 24722
rect 24110 24670 24162 24722
rect 25790 24670 25842 24722
rect 26126 24670 26178 24722
rect 28142 24670 28194 24722
rect 29598 24670 29650 24722
rect 30494 24670 30546 24722
rect 30830 24670 30882 24722
rect 31390 24670 31442 24722
rect 33182 24670 33234 24722
rect 39230 24670 39282 24722
rect 44270 24670 44322 24722
rect 45726 24670 45778 24722
rect 46958 24670 47010 24722
rect 47518 24670 47570 24722
rect 3166 24558 3218 24610
rect 5294 24558 5346 24610
rect 8206 24558 8258 24610
rect 10558 24558 10610 24610
rect 13806 24558 13858 24610
rect 16718 24558 16770 24610
rect 18174 24558 18226 24610
rect 21198 24558 21250 24610
rect 26238 24558 26290 24610
rect 27246 24558 27298 24610
rect 27694 24558 27746 24610
rect 29038 24558 29090 24610
rect 32398 24558 32450 24610
rect 35982 24558 36034 24610
rect 36318 24558 36370 24610
rect 39678 24558 39730 24610
rect 41358 24558 41410 24610
rect 46174 24558 46226 24610
rect 16830 24446 16882 24498
rect 24558 24446 24610 24498
rect 45614 24446 45666 24498
rect 47630 24446 47682 24498
rect 4478 24278 4530 24330
rect 4582 24278 4634 24330
rect 4686 24278 4738 24330
rect 35198 24278 35250 24330
rect 35302 24278 35354 24330
rect 35406 24278 35458 24330
rect 8654 24110 8706 24162
rect 12798 24110 12850 24162
rect 7198 23998 7250 24050
rect 8430 23998 8482 24050
rect 14142 23998 14194 24050
rect 14814 23998 14866 24050
rect 15934 23998 15986 24050
rect 22318 23998 22370 24050
rect 24558 23998 24610 24050
rect 27806 23998 27858 24050
rect 29710 23998 29762 24050
rect 7534 23886 7586 23938
rect 8654 23886 8706 23938
rect 10894 23886 10946 23938
rect 12350 23886 12402 23938
rect 12686 23886 12738 23938
rect 18846 23886 18898 23938
rect 19294 23886 19346 23938
rect 20190 23886 20242 23938
rect 21646 23886 21698 23938
rect 22654 23886 22706 23938
rect 24894 23886 24946 23938
rect 29262 23886 29314 23938
rect 31054 24110 31106 24162
rect 35086 23998 35138 24050
rect 35982 23998 36034 24050
rect 40686 23998 40738 24050
rect 44830 23998 44882 24050
rect 30382 23886 30434 23938
rect 30606 23886 30658 23938
rect 31614 23886 31666 23938
rect 34638 23886 34690 23938
rect 34974 23886 35026 23938
rect 35758 23886 35810 23938
rect 36094 23886 36146 23938
rect 36318 23886 36370 23938
rect 37886 23886 37938 23938
rect 47742 23886 47794 23938
rect 6526 23774 6578 23826
rect 11566 23774 11618 23826
rect 12126 23774 12178 23826
rect 12798 23774 12850 23826
rect 13694 23774 13746 23826
rect 13918 23774 13970 23826
rect 14254 23774 14306 23826
rect 14926 23774 14978 23826
rect 15150 23774 15202 23826
rect 18062 23774 18114 23826
rect 19518 23774 19570 23826
rect 21310 23774 21362 23826
rect 23102 23774 23154 23826
rect 23214 23774 23266 23826
rect 23998 23774 24050 23826
rect 24110 23774 24162 23826
rect 24222 23774 24274 23826
rect 25678 23774 25730 23826
rect 28478 23774 28530 23826
rect 31278 23774 31330 23826
rect 32062 23774 32114 23826
rect 35646 23774 35698 23826
rect 38558 23774 38610 23826
rect 46958 23774 47010 23826
rect 5070 23662 5122 23714
rect 5966 23662 6018 23714
rect 12014 23662 12066 23714
rect 14030 23662 14082 23714
rect 14590 23662 14642 23714
rect 14814 23662 14866 23714
rect 19966 23662 20018 23714
rect 20750 23662 20802 23714
rect 23326 23662 23378 23714
rect 23438 23662 23490 23714
rect 23774 23662 23826 23714
rect 28142 23662 28194 23714
rect 29150 23662 29202 23714
rect 30046 23662 30098 23714
rect 30830 23662 30882 23714
rect 37102 23662 37154 23714
rect 41134 23662 41186 23714
rect 44270 23662 44322 23714
rect 19838 23494 19890 23546
rect 19942 23494 19994 23546
rect 20046 23494 20098 23546
rect 10222 23326 10274 23378
rect 18286 23326 18338 23378
rect 18398 23326 18450 23378
rect 19070 23326 19122 23378
rect 21534 23326 21586 23378
rect 22206 23326 22258 23378
rect 22990 23326 23042 23378
rect 23214 23326 23266 23378
rect 27918 23326 27970 23378
rect 39566 23326 39618 23378
rect 44942 23326 44994 23378
rect 45614 23326 45666 23378
rect 11230 23214 11282 23266
rect 12686 23214 12738 23266
rect 18174 23214 18226 23266
rect 44606 23214 44658 23266
rect 44718 23214 44770 23266
rect 45166 23214 45218 23266
rect 45950 23214 46002 23266
rect 46174 23214 46226 23266
rect 46286 23214 46338 23266
rect 46622 23214 46674 23266
rect 48078 23214 48130 23266
rect 6302 23102 6354 23154
rect 7982 23102 8034 23154
rect 8430 23102 8482 23154
rect 12126 23102 12178 23154
rect 12574 23102 12626 23154
rect 13470 23102 13522 23154
rect 13918 23102 13970 23154
rect 16382 23102 16434 23154
rect 17614 23102 17666 23154
rect 17950 23102 18002 23154
rect 19406 23102 19458 23154
rect 19742 23102 19794 23154
rect 21310 23102 21362 23154
rect 21870 23102 21922 23154
rect 23326 23102 23378 23154
rect 28254 23102 28306 23154
rect 40910 23102 40962 23154
rect 45502 23102 45554 23154
rect 45838 23102 45890 23154
rect 46958 23102 47010 23154
rect 47294 23102 47346 23154
rect 47406 23102 47458 23154
rect 47742 23102 47794 23154
rect 3502 22990 3554 23042
rect 5630 22990 5682 23042
rect 8878 22990 8930 23042
rect 10446 22990 10498 23042
rect 15822 22990 15874 23042
rect 20302 22990 20354 23042
rect 20750 22990 20802 23042
rect 22654 22990 22706 23042
rect 23886 22990 23938 23042
rect 24334 22990 24386 23042
rect 25342 22990 25394 23042
rect 29038 22990 29090 23042
rect 31166 22990 31218 23042
rect 31614 22990 31666 23042
rect 36766 22990 36818 23042
rect 39118 22990 39170 23042
rect 40462 22990 40514 23042
rect 41694 22990 41746 23042
rect 43822 22990 43874 23042
rect 44270 22990 44322 23042
rect 47070 22990 47122 23042
rect 47630 22990 47682 23042
rect 7422 22878 7474 22930
rect 19854 22878 19906 22930
rect 4478 22710 4530 22762
rect 4582 22710 4634 22762
rect 4686 22710 4738 22762
rect 35198 22710 35250 22762
rect 35302 22710 35354 22762
rect 35406 22710 35458 22762
rect 35198 22542 35250 22594
rect 44718 22542 44770 22594
rect 45054 22542 45106 22594
rect 4734 22430 4786 22482
rect 6078 22430 6130 22482
rect 7086 22430 7138 22482
rect 7198 22430 7250 22482
rect 11118 22430 11170 22482
rect 16382 22430 16434 22482
rect 16942 22430 16994 22482
rect 21422 22430 21474 22482
rect 22430 22430 22482 22482
rect 23662 22430 23714 22482
rect 25790 22430 25842 22482
rect 28478 22430 28530 22482
rect 29486 22430 29538 22482
rect 34190 22430 34242 22482
rect 36318 22430 36370 22482
rect 40462 22430 40514 22482
rect 40910 22430 40962 22482
rect 43150 22430 43202 22482
rect 45278 22430 45330 22482
rect 47406 22430 47458 22482
rect 4958 22318 5010 22370
rect 5854 22318 5906 22370
rect 8990 22318 9042 22370
rect 9326 22318 9378 22370
rect 12686 22318 12738 22370
rect 13582 22318 13634 22370
rect 16718 22318 16770 22370
rect 17614 22318 17666 22370
rect 18174 22318 18226 22370
rect 18622 22318 18674 22370
rect 19630 22318 19682 22370
rect 19966 22318 20018 22370
rect 20190 22318 20242 22370
rect 22990 22318 23042 22370
rect 27022 22318 27074 22370
rect 27582 22318 27634 22370
rect 28030 22318 28082 22370
rect 30382 22318 30434 22370
rect 30606 22318 30658 22370
rect 31726 22318 31778 22370
rect 32286 22318 32338 22370
rect 32622 22318 32674 22370
rect 33854 22318 33906 22370
rect 34638 22318 34690 22370
rect 34862 22318 34914 22370
rect 35086 22318 35138 22370
rect 37550 22318 37602 22370
rect 42254 22318 42306 22370
rect 48190 22318 48242 22370
rect 7982 22206 8034 22258
rect 10334 22206 10386 22258
rect 12350 22206 12402 22258
rect 12798 22206 12850 22258
rect 14254 22206 14306 22258
rect 18510 22206 18562 22258
rect 19182 22206 19234 22258
rect 20526 22206 20578 22258
rect 27694 22206 27746 22258
rect 29374 22206 29426 22258
rect 29710 22206 29762 22258
rect 29934 22206 29986 22258
rect 35534 22206 35586 22258
rect 38334 22206 38386 22258
rect 42478 22206 42530 22258
rect 43598 22206 43650 22258
rect 9438 22094 9490 22146
rect 13022 22094 13074 22146
rect 19854 22094 19906 22146
rect 20414 22094 20466 22146
rect 21982 22094 22034 22146
rect 26238 22094 26290 22146
rect 27134 22094 27186 22146
rect 27358 22094 27410 22146
rect 30494 22094 30546 22146
rect 30830 22094 30882 22146
rect 31390 22094 31442 22146
rect 32958 22094 33010 22146
rect 33406 22094 33458 22146
rect 35870 22094 35922 22146
rect 37102 22094 37154 22146
rect 41582 22094 41634 22146
rect 41694 22094 41746 22146
rect 41806 22094 41858 22146
rect 42590 22094 42642 22146
rect 42814 22094 42866 22146
rect 43486 22094 43538 22146
rect 44158 22094 44210 22146
rect 44942 22094 44994 22146
rect 19838 21926 19890 21978
rect 19942 21926 19994 21978
rect 20046 21926 20098 21978
rect 8206 21758 8258 21810
rect 10894 21758 10946 21810
rect 12910 21758 12962 21810
rect 13918 21758 13970 21810
rect 14590 21758 14642 21810
rect 15150 21758 15202 21810
rect 15598 21758 15650 21810
rect 15934 21758 15986 21810
rect 18286 21758 18338 21810
rect 18734 21758 18786 21810
rect 20078 21758 20130 21810
rect 21310 21758 21362 21810
rect 21646 21758 21698 21810
rect 22206 21758 22258 21810
rect 22878 21758 22930 21810
rect 23438 21758 23490 21810
rect 24334 21758 24386 21810
rect 26350 21758 26402 21810
rect 29150 21758 29202 21810
rect 40350 21758 40402 21810
rect 41134 21758 41186 21810
rect 46622 21758 46674 21810
rect 46846 21758 46898 21810
rect 47182 21758 47234 21810
rect 9550 21646 9602 21698
rect 10670 21646 10722 21698
rect 10782 21646 10834 21698
rect 11678 21646 11730 21698
rect 12574 21646 12626 21698
rect 14142 21646 14194 21698
rect 21086 21646 21138 21698
rect 23102 21646 23154 21698
rect 23886 21646 23938 21698
rect 31054 21646 31106 21698
rect 31390 21646 31442 21698
rect 31614 21646 31666 21698
rect 39566 21646 39618 21698
rect 41470 21646 41522 21698
rect 46510 21646 46562 21698
rect 47070 21646 47122 21698
rect 47854 21646 47906 21698
rect 4846 21534 4898 21586
rect 9886 21534 9938 21586
rect 11118 21534 11170 21586
rect 11454 21534 11506 21586
rect 11902 21534 11954 21586
rect 12238 21534 12290 21586
rect 13358 21534 13410 21586
rect 13694 21534 13746 21586
rect 14702 21534 14754 21586
rect 14926 21534 14978 21586
rect 15262 21534 15314 21586
rect 16270 21534 16322 21586
rect 17726 21534 17778 21586
rect 17950 21534 18002 21586
rect 19966 21534 20018 21586
rect 20190 21534 20242 21586
rect 20974 21534 21026 21586
rect 21758 21534 21810 21586
rect 22766 21534 22818 21586
rect 23662 21534 23714 21586
rect 23998 21534 24050 21586
rect 24670 21534 24722 21586
rect 25342 21534 25394 21586
rect 26686 21534 26738 21586
rect 27358 21534 27410 21586
rect 27582 21534 27634 21586
rect 32062 21534 32114 21586
rect 35198 21534 35250 21586
rect 38558 21534 38610 21586
rect 39342 21534 39394 21586
rect 39790 21534 39842 21586
rect 40014 21534 40066 21586
rect 40798 21534 40850 21586
rect 41134 21534 41186 21586
rect 41918 21534 41970 21586
rect 48190 21534 48242 21586
rect 5518 21422 5570 21474
rect 9102 21422 9154 21474
rect 10334 21422 10386 21474
rect 11790 21422 11842 21474
rect 14030 21422 14082 21474
rect 16718 21422 16770 21474
rect 19294 21422 19346 21474
rect 20414 21422 20466 21474
rect 25678 21422 25730 21474
rect 28030 21422 28082 21474
rect 28702 21422 28754 21474
rect 29598 21422 29650 21474
rect 31278 21422 31330 21474
rect 32286 21422 32338 21474
rect 35982 21422 36034 21474
rect 38110 21422 38162 21474
rect 38894 21422 38946 21474
rect 42590 21422 42642 21474
rect 44718 21422 44770 21474
rect 46286 21422 46338 21474
rect 14590 21310 14642 21362
rect 20638 21310 20690 21362
rect 21646 21310 21698 21362
rect 28142 21310 28194 21362
rect 32398 21310 32450 21362
rect 47182 21310 47234 21362
rect 4478 21142 4530 21194
rect 4582 21142 4634 21194
rect 4686 21142 4738 21194
rect 35198 21142 35250 21194
rect 35302 21142 35354 21194
rect 35406 21142 35458 21194
rect 4958 20974 5010 21026
rect 6862 20974 6914 21026
rect 19966 20974 20018 21026
rect 21422 20974 21474 21026
rect 26462 20974 26514 21026
rect 27134 20974 27186 21026
rect 28030 20974 28082 21026
rect 28702 20974 28754 21026
rect 35758 20974 35810 21026
rect 4846 20862 4898 20914
rect 9662 20862 9714 20914
rect 10670 20862 10722 20914
rect 14142 20862 14194 20914
rect 17950 20862 18002 20914
rect 19406 20862 19458 20914
rect 20526 20862 20578 20914
rect 22542 20862 22594 20914
rect 22654 20862 22706 20914
rect 27358 20862 27410 20914
rect 28030 20862 28082 20914
rect 29822 20862 29874 20914
rect 32286 20862 32338 20914
rect 34414 20862 34466 20914
rect 36094 20862 36146 20914
rect 37662 20862 37714 20914
rect 39342 20862 39394 20914
rect 41918 20862 41970 20914
rect 42814 20862 42866 20914
rect 44942 20862 44994 20914
rect 45278 20862 45330 20914
rect 47406 20862 47458 20914
rect 4734 20750 4786 20802
rect 8766 20750 8818 20802
rect 11006 20750 11058 20802
rect 11902 20750 11954 20802
rect 17054 20750 17106 20802
rect 17726 20750 17778 20802
rect 19630 20750 19682 20802
rect 20190 20750 20242 20802
rect 20414 20750 20466 20802
rect 20638 20750 20690 20802
rect 21534 20750 21586 20802
rect 23998 20750 24050 20802
rect 25118 20750 25170 20802
rect 26126 20750 26178 20802
rect 26910 20750 26962 20802
rect 31502 20750 31554 20802
rect 35982 20750 36034 20802
rect 38222 20750 38274 20802
rect 40014 20750 40066 20802
rect 48078 20750 48130 20802
rect 11566 20638 11618 20690
rect 11678 20638 11730 20690
rect 12462 20638 12514 20690
rect 12574 20638 12626 20690
rect 13470 20638 13522 20690
rect 16270 20638 16322 20690
rect 21422 20638 21474 20690
rect 22094 20638 22146 20690
rect 22206 20638 22258 20690
rect 23438 20638 23490 20690
rect 23886 20638 23938 20690
rect 24334 20638 24386 20690
rect 24446 20638 24498 20690
rect 24894 20638 24946 20690
rect 26574 20638 26626 20690
rect 27470 20638 27522 20690
rect 34862 20638 34914 20690
rect 35310 20638 35362 20690
rect 35534 20638 35586 20690
rect 36206 20638 36258 20690
rect 36990 20638 37042 20690
rect 37102 20638 37154 20690
rect 38558 20638 38610 20690
rect 39006 20638 39058 20690
rect 42702 20638 42754 20690
rect 43038 20638 43090 20690
rect 43150 20638 43202 20690
rect 43934 20638 43986 20690
rect 6302 20526 6354 20578
rect 12686 20526 12738 20578
rect 12798 20526 12850 20578
rect 12910 20526 12962 20578
rect 13806 20526 13858 20578
rect 18286 20526 18338 20578
rect 18958 20526 19010 20578
rect 19070 20526 19122 20578
rect 19182 20526 19234 20578
rect 21870 20526 21922 20578
rect 23102 20526 23154 20578
rect 23662 20526 23714 20578
rect 25790 20526 25842 20578
rect 28366 20526 28418 20578
rect 39230 20526 39282 20578
rect 39454 20526 39506 20578
rect 42926 20526 42978 20578
rect 19838 20358 19890 20410
rect 19942 20358 19994 20410
rect 20046 20358 20098 20410
rect 14478 20190 14530 20242
rect 15822 20190 15874 20242
rect 16830 20190 16882 20242
rect 17614 20190 17666 20242
rect 20414 20190 20466 20242
rect 21310 20190 21362 20242
rect 23326 20190 23378 20242
rect 24782 20190 24834 20242
rect 39118 20190 39170 20242
rect 39566 20190 39618 20242
rect 5406 20078 5458 20130
rect 9662 20078 9714 20130
rect 9774 20078 9826 20130
rect 10446 20078 10498 20130
rect 11902 20078 11954 20130
rect 12014 20078 12066 20130
rect 12462 20078 12514 20130
rect 13246 20078 13298 20130
rect 15262 20078 15314 20130
rect 15374 20078 15426 20130
rect 16494 20078 16546 20130
rect 17390 20078 17442 20130
rect 20526 20078 20578 20130
rect 22094 20078 22146 20130
rect 22318 20078 22370 20130
rect 22654 20078 22706 20130
rect 22766 20078 22818 20130
rect 23886 20078 23938 20130
rect 25566 20078 25618 20130
rect 30718 20078 30770 20130
rect 31166 20078 31218 20130
rect 32174 20078 32226 20130
rect 32510 20078 32562 20130
rect 33742 20078 33794 20130
rect 33966 20078 34018 20130
rect 34750 20078 34802 20130
rect 35086 20078 35138 20130
rect 35646 20078 35698 20130
rect 38782 20078 38834 20130
rect 41806 20078 41858 20130
rect 42254 20078 42306 20130
rect 43262 20078 43314 20130
rect 47518 20078 47570 20130
rect 47854 20078 47906 20130
rect 5070 19966 5122 20018
rect 8654 19966 8706 20018
rect 10670 19966 10722 20018
rect 11454 19966 11506 20018
rect 11678 19966 11730 20018
rect 12126 19966 12178 20018
rect 13582 19966 13634 20018
rect 14702 19966 14754 20018
rect 17838 19966 17890 20018
rect 18062 19966 18114 20018
rect 19182 19966 19234 20018
rect 19966 19966 20018 20018
rect 20190 19966 20242 20018
rect 20638 19966 20690 20018
rect 21534 19966 21586 20018
rect 21982 19966 22034 20018
rect 23550 19966 23602 20018
rect 26910 19966 26962 20018
rect 30158 19966 30210 20018
rect 30382 19966 30434 20018
rect 31054 19966 31106 20018
rect 31278 19966 31330 20018
rect 31726 19966 31778 20018
rect 35870 19966 35922 20018
rect 40798 19966 40850 20018
rect 41134 19966 41186 20018
rect 41358 19966 41410 20018
rect 41918 19966 41970 20018
rect 42030 19966 42082 20018
rect 43710 19966 43762 20018
rect 45054 19966 45106 20018
rect 45726 19966 45778 20018
rect 46174 19966 46226 20018
rect 4958 19854 5010 19906
rect 5742 19854 5794 19906
rect 7870 19854 7922 19906
rect 14030 19854 14082 19906
rect 15710 19854 15762 19906
rect 17502 19854 17554 19906
rect 18622 19854 18674 19906
rect 19630 19854 19682 19906
rect 26574 19854 26626 19906
rect 27694 19854 27746 19906
rect 29822 19854 29874 19906
rect 30270 19854 30322 19906
rect 33854 19854 33906 19906
rect 34414 19854 34466 19906
rect 37102 19854 37154 19906
rect 40014 19854 40066 19906
rect 41022 19854 41074 19906
rect 42366 19854 42418 19906
rect 9774 19742 9826 19794
rect 15262 19742 15314 19794
rect 22654 19742 22706 19794
rect 42814 19854 42866 19906
rect 44270 19854 44322 19906
rect 44606 19854 44658 19906
rect 43262 19742 43314 19794
rect 4478 19574 4530 19626
rect 4582 19574 4634 19626
rect 4686 19574 4738 19626
rect 35198 19574 35250 19626
rect 35302 19574 35354 19626
rect 35406 19574 35458 19626
rect 6750 19406 6802 19458
rect 8318 19294 8370 19346
rect 12126 19294 12178 19346
rect 12910 19294 12962 19346
rect 16046 19294 16098 19346
rect 17838 19294 17890 19346
rect 18174 19294 18226 19346
rect 20302 19294 20354 19346
rect 23662 19294 23714 19346
rect 28142 19294 28194 19346
rect 29934 19294 29986 19346
rect 32062 19294 32114 19346
rect 33182 19294 33234 19346
rect 34526 19294 34578 19346
rect 35310 19294 35362 19346
rect 36206 19294 36258 19346
rect 39118 19294 39170 19346
rect 40238 19294 40290 19346
rect 42366 19294 42418 19346
rect 45166 19294 45218 19346
rect 46846 19294 46898 19346
rect 7310 19182 7362 19234
rect 11454 19182 11506 19234
rect 11678 19182 11730 19234
rect 12014 19182 12066 19234
rect 12462 19182 12514 19234
rect 14142 19182 14194 19234
rect 14254 19182 14306 19234
rect 14590 19182 14642 19234
rect 16382 19182 16434 19234
rect 16718 19182 16770 19234
rect 17278 19182 17330 19234
rect 17838 19182 17890 19234
rect 18734 19182 18786 19234
rect 21534 19182 21586 19234
rect 22094 19182 22146 19234
rect 25118 19182 25170 19234
rect 25454 19182 25506 19234
rect 26238 19182 26290 19234
rect 27918 19182 27970 19234
rect 28254 19182 28306 19234
rect 29262 19182 29314 19234
rect 32398 19182 32450 19234
rect 33294 19182 33346 19234
rect 34750 19182 34802 19234
rect 35198 19182 35250 19234
rect 35758 19182 35810 19234
rect 36878 19182 36930 19234
rect 37214 19182 37266 19234
rect 39566 19182 39618 19234
rect 43598 19182 43650 19234
rect 43822 19182 43874 19234
rect 44830 19182 44882 19234
rect 45950 19182 46002 19234
rect 10558 19070 10610 19122
rect 13694 19070 13746 19122
rect 14478 19070 14530 19122
rect 15150 19070 15202 19122
rect 16942 19070 16994 19122
rect 21758 19070 21810 19122
rect 25790 19070 25842 19122
rect 28590 19070 28642 19122
rect 34414 19070 34466 19122
rect 35422 19070 35474 19122
rect 36094 19070 36146 19122
rect 36318 19070 36370 19122
rect 37550 19070 37602 19122
rect 38222 19070 38274 19122
rect 43374 19070 43426 19122
rect 44942 19070 44994 19122
rect 46398 19070 46450 19122
rect 46510 19070 46562 19122
rect 46734 19070 46786 19122
rect 12238 18958 12290 19010
rect 13470 18958 13522 19010
rect 13582 18958 13634 19010
rect 15710 18958 15762 19010
rect 16494 18958 16546 19010
rect 17390 18958 17442 19010
rect 17502 18958 17554 19010
rect 25454 18958 25506 19010
rect 27806 18958 27858 19010
rect 34190 18958 34242 19010
rect 37102 18958 37154 19010
rect 37886 18958 37938 19010
rect 38670 18958 38722 19010
rect 42926 18958 42978 19010
rect 43486 18958 43538 19010
rect 46286 18958 46338 19010
rect 19838 18790 19890 18842
rect 19942 18790 19994 18842
rect 20046 18790 20098 18842
rect 8878 18622 8930 18674
rect 14590 18622 14642 18674
rect 17614 18622 17666 18674
rect 18734 18622 18786 18674
rect 24110 18622 24162 18674
rect 24670 18622 24722 18674
rect 28814 18622 28866 18674
rect 33182 18622 33234 18674
rect 35870 18622 35922 18674
rect 16270 18510 16322 18562
rect 16830 18510 16882 18562
rect 19070 18510 19122 18562
rect 21646 18510 21698 18562
rect 28926 18510 28978 18562
rect 40014 18510 40066 18562
rect 41246 18510 41298 18562
rect 42478 18510 42530 18562
rect 44270 18510 44322 18562
rect 46062 18510 46114 18562
rect 10222 18398 10274 18450
rect 10894 18398 10946 18450
rect 11678 18398 11730 18450
rect 12350 18398 12402 18450
rect 15150 18398 15202 18450
rect 15598 18398 15650 18450
rect 16606 18398 16658 18450
rect 17726 18398 17778 18450
rect 17838 18398 17890 18450
rect 18286 18398 18338 18450
rect 20078 18398 20130 18450
rect 22206 18398 22258 18450
rect 22654 18398 22706 18450
rect 22990 18398 23042 18450
rect 23214 18398 23266 18450
rect 23438 18398 23490 18450
rect 23886 18398 23938 18450
rect 23998 18398 24050 18450
rect 25230 18398 25282 18450
rect 26014 18398 26066 18450
rect 28702 18398 28754 18450
rect 29262 18398 29314 18450
rect 31950 18398 32002 18450
rect 32958 18398 33010 18450
rect 33294 18398 33346 18450
rect 33630 18398 33682 18450
rect 35086 18398 35138 18450
rect 35534 18398 35586 18450
rect 36094 18398 36146 18450
rect 36878 18398 36930 18450
rect 40350 18398 40402 18450
rect 40910 18398 40962 18450
rect 41470 18398 41522 18450
rect 42142 18398 42194 18450
rect 42702 18398 42754 18450
rect 42926 18398 42978 18450
rect 43262 18398 43314 18450
rect 43598 18398 43650 18450
rect 44606 18398 44658 18450
rect 44830 18398 44882 18450
rect 45390 18398 45442 18450
rect 16382 18286 16434 18338
rect 22766 18286 22818 18338
rect 28142 18286 28194 18338
rect 29374 18286 29426 18338
rect 29710 18286 29762 18338
rect 32510 18286 32562 18338
rect 34638 18286 34690 18338
rect 39006 18286 39058 18338
rect 39454 18286 39506 18338
rect 41022 18286 41074 18338
rect 42590 18286 42642 18338
rect 43150 18286 43202 18338
rect 43934 18286 43986 18338
rect 44942 18286 44994 18338
rect 48190 18286 48242 18338
rect 29710 18174 29762 18226
rect 32286 18174 32338 18226
rect 44046 18174 44098 18226
rect 4478 18006 4530 18058
rect 4582 18006 4634 18058
rect 4686 18006 4738 18058
rect 35198 18006 35250 18058
rect 35302 18006 35354 18058
rect 35406 18006 35458 18058
rect 19070 17838 19122 17890
rect 19294 17838 19346 17890
rect 20078 17838 20130 17890
rect 33182 17838 33234 17890
rect 33518 17838 33570 17890
rect 35086 17838 35138 17890
rect 35310 17838 35362 17890
rect 37214 17838 37266 17890
rect 9998 17726 10050 17778
rect 10670 17726 10722 17778
rect 11566 17726 11618 17778
rect 12462 17726 12514 17778
rect 13582 17726 13634 17778
rect 14814 17726 14866 17778
rect 16942 17726 16994 17778
rect 17390 17726 17442 17778
rect 17950 17726 18002 17778
rect 19742 17726 19794 17778
rect 20190 17726 20242 17778
rect 20526 17726 20578 17778
rect 21422 17726 21474 17778
rect 22542 17726 22594 17778
rect 24670 17726 24722 17778
rect 26126 17726 26178 17778
rect 31054 17726 31106 17778
rect 32958 17726 33010 17778
rect 36206 17726 36258 17778
rect 37774 17726 37826 17778
rect 40350 17726 40402 17778
rect 44270 17726 44322 17778
rect 44830 17726 44882 17778
rect 48190 17726 48242 17778
rect 9550 17614 9602 17666
rect 10894 17614 10946 17666
rect 11118 17614 11170 17666
rect 14030 17614 14082 17666
rect 21870 17614 21922 17666
rect 25006 17614 25058 17666
rect 26014 17614 26066 17666
rect 26238 17614 26290 17666
rect 27134 17614 27186 17666
rect 28590 17614 28642 17666
rect 29374 17614 29426 17666
rect 29710 17614 29762 17666
rect 29934 17614 29986 17666
rect 30382 17614 30434 17666
rect 30606 17614 30658 17666
rect 33966 17614 34018 17666
rect 34862 17614 34914 17666
rect 36094 17614 36146 17666
rect 36318 17614 36370 17666
rect 37998 17614 38050 17666
rect 38222 17614 38274 17666
rect 38446 17614 38498 17666
rect 39118 17614 39170 17666
rect 42926 17614 42978 17666
rect 43262 17614 43314 17666
rect 43374 17614 43426 17666
rect 43934 17614 43986 17666
rect 44158 17614 44210 17666
rect 45390 17614 45442 17666
rect 10558 17502 10610 17554
rect 18734 17502 18786 17554
rect 25342 17502 25394 17554
rect 28478 17502 28530 17554
rect 29150 17502 29202 17554
rect 31390 17502 31442 17554
rect 34302 17502 34354 17554
rect 34526 17502 34578 17554
rect 35422 17502 35474 17554
rect 35758 17502 35810 17554
rect 37102 17502 37154 17554
rect 38894 17502 38946 17554
rect 39230 17502 39282 17554
rect 41806 17502 41858 17554
rect 43710 17502 43762 17554
rect 44942 17502 44994 17554
rect 46062 17502 46114 17554
rect 13022 17390 13074 17442
rect 18174 17390 18226 17442
rect 19182 17390 19234 17442
rect 26462 17390 26514 17442
rect 26910 17390 26962 17442
rect 27694 17390 27746 17442
rect 28142 17390 28194 17442
rect 28366 17390 28418 17442
rect 29598 17390 29650 17442
rect 30158 17390 30210 17442
rect 30942 17390 30994 17442
rect 31166 17390 31218 17442
rect 34190 17390 34242 17442
rect 37214 17390 37266 17442
rect 19838 17222 19890 17274
rect 19942 17222 19994 17274
rect 20046 17222 20098 17274
rect 12014 17054 12066 17106
rect 12798 17054 12850 17106
rect 13582 17054 13634 17106
rect 17502 17054 17554 17106
rect 18062 17054 18114 17106
rect 21534 17054 21586 17106
rect 25342 17054 25394 17106
rect 30830 17054 30882 17106
rect 31726 17054 31778 17106
rect 34190 17054 34242 17106
rect 34414 17054 34466 17106
rect 35422 17054 35474 17106
rect 36318 17054 36370 17106
rect 43598 17054 43650 17106
rect 43822 17054 43874 17106
rect 45054 17054 45106 17106
rect 45614 17054 45666 17106
rect 47854 17054 47906 17106
rect 14702 16942 14754 16994
rect 18622 16942 18674 16994
rect 19630 16942 19682 16994
rect 21646 16942 21698 16994
rect 26910 16942 26962 16994
rect 29374 16942 29426 16994
rect 33294 16942 33346 16994
rect 36094 16942 36146 16994
rect 36430 16942 36482 16994
rect 37438 16942 37490 16994
rect 38334 16942 38386 16994
rect 38894 16942 38946 16994
rect 41134 16942 41186 16994
rect 42366 16942 42418 16994
rect 11566 16830 11618 16882
rect 14030 16830 14082 16882
rect 18734 16830 18786 16882
rect 19070 16830 19122 16882
rect 22766 16830 22818 16882
rect 26574 16830 26626 16882
rect 30158 16830 30210 16882
rect 31390 16830 31442 16882
rect 33518 16830 33570 16882
rect 34974 16830 35026 16882
rect 36654 16830 36706 16882
rect 37662 16830 37714 16882
rect 37886 16830 37938 16882
rect 38558 16830 38610 16882
rect 38782 16830 38834 16882
rect 39566 16830 39618 16882
rect 39790 16830 39842 16882
rect 40910 16830 40962 16882
rect 41582 16830 41634 16882
rect 41694 16830 41746 16882
rect 42030 16830 42082 16882
rect 42702 16830 42754 16882
rect 42926 16830 42978 16882
rect 44158 16830 44210 16882
rect 44494 16830 44546 16882
rect 45390 16830 45442 16882
rect 46062 16830 46114 16882
rect 46286 16830 46338 16882
rect 47182 16830 47234 16882
rect 47406 16830 47458 16882
rect 16830 16718 16882 16770
rect 27246 16718 27298 16770
rect 37998 16718 38050 16770
rect 40238 16718 40290 16770
rect 41022 16718 41074 16770
rect 41918 16718 41970 16770
rect 43710 16718 43762 16770
rect 44718 16718 44770 16770
rect 45502 16718 45554 16770
rect 46734 16718 46786 16770
rect 46958 16718 47010 16770
rect 30830 16606 30882 16658
rect 31614 16606 31666 16658
rect 36990 16606 37042 16658
rect 37102 16606 37154 16658
rect 39230 16606 39282 16658
rect 43262 16606 43314 16658
rect 4478 16438 4530 16490
rect 4582 16438 4634 16490
rect 4686 16438 4738 16490
rect 35198 16438 35250 16490
rect 35302 16438 35354 16490
rect 35406 16438 35458 16490
rect 19742 16270 19794 16322
rect 36094 16270 36146 16322
rect 36430 16270 36482 16322
rect 43822 16270 43874 16322
rect 45950 16270 46002 16322
rect 46286 16270 46338 16322
rect 14590 16158 14642 16210
rect 14926 16158 14978 16210
rect 16270 16158 16322 16210
rect 16830 16158 16882 16210
rect 23102 16158 23154 16210
rect 26462 16158 26514 16210
rect 30158 16158 30210 16210
rect 32286 16158 32338 16210
rect 35198 16158 35250 16210
rect 39230 16158 39282 16210
rect 41806 16158 41858 16210
rect 44270 16158 44322 16210
rect 46734 16158 46786 16210
rect 17502 16046 17554 16098
rect 21646 16046 21698 16098
rect 22206 16046 22258 16098
rect 23662 16046 23714 16098
rect 29374 16046 29426 16098
rect 33518 16046 33570 16098
rect 33966 16046 34018 16098
rect 35534 16046 35586 16098
rect 35870 16046 35922 16098
rect 37550 16046 37602 16098
rect 39902 16046 39954 16098
rect 42926 16046 42978 16098
rect 43150 16046 43202 16098
rect 43710 16046 43762 16098
rect 45054 16046 45106 16098
rect 45390 16046 45442 16098
rect 45726 16046 45778 16098
rect 17166 15934 17218 15986
rect 17726 15934 17778 15986
rect 18510 15934 18562 15986
rect 17278 15822 17330 15874
rect 18846 15822 18898 15874
rect 19182 15822 19234 15874
rect 19630 15878 19682 15930
rect 19742 15934 19794 15986
rect 20414 15934 20466 15986
rect 20750 15934 20802 15986
rect 21310 15934 21362 15986
rect 21870 15934 21922 15986
rect 22542 15934 22594 15986
rect 24334 15934 24386 15986
rect 34302 15934 34354 15986
rect 34638 15934 34690 15986
rect 36318 15934 36370 15986
rect 44942 15934 44994 15986
rect 47854 15934 47906 15986
rect 48190 15934 48242 15986
rect 21422 15822 21474 15874
rect 35646 15822 35698 15874
rect 43038 15822 43090 15874
rect 43374 15822 43426 15874
rect 44830 15822 44882 15874
rect 47630 15822 47682 15874
rect 19838 15654 19890 15706
rect 19942 15654 19994 15706
rect 20046 15654 20098 15706
rect 17614 15486 17666 15538
rect 18062 15486 18114 15538
rect 20526 15486 20578 15538
rect 25230 15486 25282 15538
rect 26574 15486 26626 15538
rect 27134 15486 27186 15538
rect 29598 15486 29650 15538
rect 31614 15486 31666 15538
rect 33294 15486 33346 15538
rect 33854 15486 33906 15538
rect 40238 15486 40290 15538
rect 41582 15486 41634 15538
rect 16606 15374 16658 15426
rect 19182 15374 19234 15426
rect 22206 15374 22258 15426
rect 30718 15374 30770 15426
rect 38446 15374 38498 15426
rect 38894 15374 38946 15426
rect 39454 15374 39506 15426
rect 41470 15374 41522 15426
rect 41694 15374 41746 15426
rect 42030 15374 42082 15426
rect 43598 15374 43650 15426
rect 16270 15262 16322 15314
rect 16830 15262 16882 15314
rect 17950 15262 18002 15314
rect 18174 15262 18226 15314
rect 18622 15262 18674 15314
rect 19070 15262 19122 15314
rect 22766 15262 22818 15314
rect 24110 15262 24162 15314
rect 25790 15262 25842 15314
rect 26014 15262 26066 15314
rect 26350 15262 26402 15314
rect 26798 15262 26850 15314
rect 27246 15262 27298 15314
rect 27470 15262 27522 15314
rect 30158 15262 30210 15314
rect 30942 15262 30994 15314
rect 31278 15262 31330 15314
rect 32174 15262 32226 15314
rect 35086 15262 35138 15314
rect 39006 15262 39058 15314
rect 39118 15262 39170 15314
rect 39678 15262 39730 15314
rect 39790 15262 39842 15314
rect 42254 15262 42306 15314
rect 42366 15262 42418 15314
rect 42702 15262 42754 15314
rect 43038 15262 43090 15314
rect 43262 15262 43314 15314
rect 43710 15262 43762 15314
rect 44158 15262 44210 15314
rect 44830 15262 44882 15314
rect 16382 15150 16434 15202
rect 23886 15150 23938 15202
rect 25566 15150 25618 15202
rect 26238 15150 26290 15202
rect 27918 15150 27970 15202
rect 30830 15150 30882 15202
rect 35870 15150 35922 15202
rect 37998 15150 38050 15202
rect 38334 15150 38386 15202
rect 46958 15150 47010 15202
rect 17278 15038 17330 15090
rect 17614 15038 17666 15090
rect 24558 15038 24610 15090
rect 31950 15038 32002 15090
rect 33070 15038 33122 15090
rect 33406 15038 33458 15090
rect 4478 14870 4530 14922
rect 4582 14870 4634 14922
rect 4686 14870 4738 14922
rect 35198 14870 35250 14922
rect 35302 14870 35354 14922
rect 35406 14870 35458 14922
rect 30270 14702 30322 14754
rect 31054 14702 31106 14754
rect 16046 14590 16098 14642
rect 18174 14590 18226 14642
rect 18846 14590 18898 14642
rect 20638 14590 20690 14642
rect 25678 14590 25730 14642
rect 27806 14590 27858 14642
rect 29598 14590 29650 14642
rect 30494 14590 30546 14642
rect 31390 14590 31442 14642
rect 33518 14590 33570 14642
rect 35534 14590 35586 14642
rect 36430 14590 36482 14642
rect 38110 14590 38162 14642
rect 41358 14590 41410 14642
rect 44942 14590 44994 14642
rect 15262 14478 15314 14530
rect 19182 14478 19234 14530
rect 19294 14478 19346 14530
rect 19742 14478 19794 14530
rect 23886 14478 23938 14530
rect 24782 14478 24834 14530
rect 25006 14478 25058 14530
rect 28590 14478 28642 14530
rect 34302 14478 34354 14530
rect 34526 14478 34578 14530
rect 37326 14478 37378 14530
rect 41022 14478 41074 14530
rect 44158 14478 44210 14530
rect 20526 14366 20578 14418
rect 22094 14366 22146 14418
rect 25342 14366 25394 14418
rect 35086 14366 35138 14418
rect 37662 14366 37714 14418
rect 40238 14366 40290 14418
rect 43486 14366 43538 14418
rect 19518 14254 19570 14306
rect 20302 14254 20354 14306
rect 20750 14254 20802 14306
rect 24334 14254 24386 14306
rect 25006 14254 25058 14306
rect 30046 14254 30098 14306
rect 31054 14254 31106 14306
rect 34862 14254 34914 14306
rect 35198 14254 35250 14306
rect 19838 14086 19890 14138
rect 19942 14086 19994 14138
rect 20046 14086 20098 14138
rect 17726 13918 17778 13970
rect 19518 13918 19570 13970
rect 23550 13918 23602 13970
rect 26798 13918 26850 13970
rect 27694 13918 27746 13970
rect 30830 13918 30882 13970
rect 33630 13918 33682 13970
rect 35422 13918 35474 13970
rect 36206 13918 36258 13970
rect 36990 13918 37042 13970
rect 39230 13918 39282 13970
rect 41470 13918 41522 13970
rect 41918 13918 41970 13970
rect 43038 13918 43090 13970
rect 43374 13918 43426 13970
rect 43822 13918 43874 13970
rect 46174 13918 46226 13970
rect 14702 13806 14754 13858
rect 17838 13806 17890 13858
rect 20750 13806 20802 13858
rect 23886 13806 23938 13858
rect 27246 13806 27298 13858
rect 32510 13806 32562 13858
rect 33406 13806 33458 13858
rect 33742 13806 33794 13858
rect 35534 13806 35586 13858
rect 35758 13806 35810 13858
rect 39118 13806 39170 13858
rect 42366 13806 42418 13858
rect 45614 13806 45666 13858
rect 45726 13806 45778 13858
rect 14030 13694 14082 13746
rect 17950 13694 18002 13746
rect 18398 13694 18450 13746
rect 18958 13694 19010 13746
rect 19406 13694 19458 13746
rect 19630 13694 19682 13746
rect 20078 13694 20130 13746
rect 23662 13694 23714 13746
rect 23998 13694 24050 13746
rect 24334 13694 24386 13746
rect 25230 13694 25282 13746
rect 25454 13694 25506 13746
rect 25902 13694 25954 13746
rect 26686 13694 26738 13746
rect 27022 13694 27074 13746
rect 29934 13694 29986 13746
rect 31838 13694 31890 13746
rect 33966 13694 34018 13746
rect 34414 13694 34466 13746
rect 35086 13694 35138 13746
rect 41134 13694 41186 13746
rect 44494 13694 44546 13746
rect 44942 13694 44994 13746
rect 45054 13694 45106 13746
rect 45390 13694 45442 13746
rect 16830 13582 16882 13634
rect 18734 13582 18786 13634
rect 22878 13582 22930 13634
rect 25342 13582 25394 13634
rect 26126 13582 26178 13634
rect 27694 13582 27746 13634
rect 30270 13582 30322 13634
rect 31950 13582 32002 13634
rect 44270 13582 44322 13634
rect 44718 13582 44770 13634
rect 26238 13470 26290 13522
rect 27806 13470 27858 13522
rect 28030 13470 28082 13522
rect 34526 13470 34578 13522
rect 34750 13470 34802 13522
rect 34862 13470 34914 13522
rect 42478 13470 42530 13522
rect 42702 13470 42754 13522
rect 43486 13470 43538 13522
rect 4478 13302 4530 13354
rect 4582 13302 4634 13354
rect 4686 13302 4738 13354
rect 35198 13302 35250 13354
rect 35302 13302 35354 13354
rect 35406 13302 35458 13354
rect 17054 13022 17106 13074
rect 24222 13022 24274 13074
rect 25678 13022 25730 13074
rect 27694 13022 27746 13074
rect 32174 13022 32226 13074
rect 34190 13022 34242 13074
rect 45614 13022 45666 13074
rect 47742 13022 47794 13074
rect 18734 12910 18786 12962
rect 21310 12910 21362 12962
rect 25118 12910 25170 12962
rect 29374 12910 29426 12962
rect 34414 12910 34466 12962
rect 34638 12910 34690 12962
rect 43934 12910 43986 12962
rect 44270 12910 44322 12962
rect 44830 12910 44882 12962
rect 18174 12798 18226 12850
rect 22094 12798 22146 12850
rect 30046 12798 30098 12850
rect 34078 12798 34130 12850
rect 35086 12798 35138 12850
rect 17838 12686 17890 12738
rect 18958 12686 19010 12738
rect 41918 12686 41970 12738
rect 42366 12686 42418 12738
rect 43710 12686 43762 12738
rect 44046 12686 44098 12738
rect 19838 12518 19890 12570
rect 19942 12518 19994 12570
rect 20046 12518 20098 12570
rect 17502 12350 17554 12402
rect 17838 12350 17890 12402
rect 18734 12350 18786 12402
rect 19070 12350 19122 12402
rect 20526 12350 20578 12402
rect 26574 12350 26626 12402
rect 29598 12350 29650 12402
rect 38110 12350 38162 12402
rect 39790 12350 39842 12402
rect 44494 12350 44546 12402
rect 16270 12238 16322 12290
rect 16606 12238 16658 12290
rect 16830 12238 16882 12290
rect 19742 12238 19794 12290
rect 27134 12238 27186 12290
rect 28142 12238 28194 12290
rect 28478 12238 28530 12290
rect 28814 12238 28866 12290
rect 30158 12238 30210 12290
rect 30382 12238 30434 12290
rect 17950 12126 18002 12178
rect 30494 12182 30546 12234
rect 31166 12238 31218 12290
rect 31614 12238 31666 12290
rect 31726 12238 31778 12290
rect 32174 12238 32226 12290
rect 35310 12238 35362 12290
rect 38782 12238 38834 12290
rect 39118 12238 39170 12290
rect 40126 12238 40178 12290
rect 18062 12126 18114 12178
rect 18398 12126 18450 12178
rect 20302 12126 20354 12178
rect 24558 12126 24610 12178
rect 25790 12126 25842 12178
rect 26126 12126 26178 12178
rect 26798 12126 26850 12178
rect 27918 12126 27970 12178
rect 30718 12126 30770 12178
rect 30942 12126 30994 12178
rect 31278 12126 31330 12178
rect 33854 12126 33906 12178
rect 34526 12126 34578 12178
rect 37774 12126 37826 12178
rect 38558 12126 38610 12178
rect 39342 12126 39394 12178
rect 40910 12126 40962 12178
rect 16382 12014 16434 12066
rect 21758 12014 21810 12066
rect 23886 12014 23938 12066
rect 25342 12014 25394 12066
rect 30382 12014 30434 12066
rect 34078 12014 34130 12066
rect 37438 12014 37490 12066
rect 41694 12014 41746 12066
rect 43822 12014 43874 12066
rect 26798 11902 26850 11954
rect 34190 11902 34242 11954
rect 4478 11734 4530 11786
rect 4582 11734 4634 11786
rect 4686 11734 4738 11786
rect 35198 11734 35250 11786
rect 35302 11734 35354 11786
rect 35406 11734 35458 11786
rect 23438 11566 23490 11618
rect 23774 11566 23826 11618
rect 24446 11566 24498 11618
rect 27022 11566 27074 11618
rect 27806 11566 27858 11618
rect 32734 11566 32786 11618
rect 34190 11566 34242 11618
rect 15598 11454 15650 11506
rect 17726 11454 17778 11506
rect 23214 11454 23266 11506
rect 34302 11454 34354 11506
rect 41246 11454 41298 11506
rect 43038 11454 43090 11506
rect 14926 11342 14978 11394
rect 18286 11342 18338 11394
rect 18846 11342 18898 11394
rect 19966 11342 20018 11394
rect 20414 11342 20466 11394
rect 21870 11342 21922 11394
rect 22990 11342 23042 11394
rect 24334 11342 24386 11394
rect 25230 11342 25282 11394
rect 25678 11342 25730 11394
rect 25790 11342 25842 11394
rect 26014 11342 26066 11394
rect 26238 11342 26290 11394
rect 26686 11342 26738 11394
rect 27806 11342 27858 11394
rect 28366 11342 28418 11394
rect 31166 11342 31218 11394
rect 32510 11342 32562 11394
rect 33070 11342 33122 11394
rect 33406 11342 33458 11394
rect 34638 11342 34690 11394
rect 34974 11342 35026 11394
rect 35646 11342 35698 11394
rect 38110 11342 38162 11394
rect 38894 11342 38946 11394
rect 39118 11342 39170 11394
rect 39902 11342 39954 11394
rect 40014 11342 40066 11394
rect 41134 11342 41186 11394
rect 41358 11342 41410 11394
rect 42254 11342 42306 11394
rect 43374 11342 43426 11394
rect 20638 11230 20690 11282
rect 21422 11230 21474 11282
rect 24222 11230 24274 11282
rect 28030 11230 28082 11282
rect 28590 11230 28642 11282
rect 36094 11230 36146 11282
rect 37102 11230 37154 11282
rect 38558 11230 38610 11282
rect 41694 11230 41746 11282
rect 42590 11230 42642 11282
rect 42702 11230 42754 11282
rect 43486 11230 43538 11282
rect 44942 11230 44994 11282
rect 18062 11118 18114 11170
rect 19070 11118 19122 11170
rect 19406 11118 19458 11170
rect 19742 11118 19794 11170
rect 20190 11118 20242 11170
rect 21310 11118 21362 11170
rect 21534 11118 21586 11170
rect 24894 11118 24946 11170
rect 25678 11118 25730 11170
rect 27134 11118 27186 11170
rect 28142 11118 28194 11170
rect 29150 11118 29202 11170
rect 29262 11118 29314 11170
rect 29374 11118 29426 11170
rect 29598 11118 29650 11170
rect 30718 11118 30770 11170
rect 30942 11118 30994 11170
rect 31054 11118 31106 11170
rect 33742 11118 33794 11170
rect 35758 11118 35810 11170
rect 35870 11118 35922 11170
rect 36990 11118 37042 11170
rect 37662 11118 37714 11170
rect 38670 11118 38722 11170
rect 39566 11118 39618 11170
rect 39790 11118 39842 11170
rect 40574 11118 40626 11170
rect 42478 11118 42530 11170
rect 43598 11118 43650 11170
rect 43822 11118 43874 11170
rect 44830 11118 44882 11170
rect 19838 10950 19890 11002
rect 19942 10950 19994 11002
rect 20046 10950 20098 11002
rect 16046 10782 16098 10834
rect 17614 10782 17666 10834
rect 17950 10782 18002 10834
rect 23662 10782 23714 10834
rect 25342 10782 25394 10834
rect 30158 10782 30210 10834
rect 37998 10782 38050 10834
rect 38446 10782 38498 10834
rect 38894 10782 38946 10834
rect 39454 10782 39506 10834
rect 41470 10782 41522 10834
rect 42254 10782 42306 10834
rect 47518 10782 47570 10834
rect 16270 10670 16322 10722
rect 16606 10670 16658 10722
rect 16830 10670 16882 10722
rect 19966 10670 20018 10722
rect 24334 10670 24386 10722
rect 26686 10670 26738 10722
rect 29486 10670 29538 10722
rect 33182 10670 33234 10722
rect 33518 10670 33570 10722
rect 37662 10670 37714 10722
rect 39678 10670 39730 10722
rect 41918 10670 41970 10722
rect 42030 10670 42082 10722
rect 43262 10670 43314 10722
rect 18062 10558 18114 10610
rect 18174 10558 18226 10610
rect 18510 10558 18562 10610
rect 19182 10558 19234 10610
rect 23550 10558 23602 10610
rect 23886 10558 23938 10610
rect 25454 10558 25506 10610
rect 25902 10558 25954 10610
rect 29150 10558 29202 10610
rect 29710 10558 29762 10610
rect 30046 10558 30098 10610
rect 30270 10558 30322 10610
rect 30718 10558 30770 10610
rect 30830 10558 30882 10610
rect 31278 10558 31330 10610
rect 31390 10558 31442 10610
rect 31950 10558 32002 10610
rect 34414 10558 34466 10610
rect 40014 10558 40066 10610
rect 40238 10558 40290 10610
rect 40798 10558 40850 10610
rect 41246 10558 41298 10610
rect 41358 10558 41410 10610
rect 42478 10558 42530 10610
rect 16382 10446 16434 10498
rect 22094 10446 22146 10498
rect 22654 10446 22706 10498
rect 23102 10446 23154 10498
rect 28814 10446 28866 10498
rect 29262 10446 29314 10498
rect 31054 10446 31106 10498
rect 35198 10446 35250 10498
rect 37326 10446 37378 10498
rect 39790 10446 39842 10498
rect 45390 10446 45442 10498
rect 47630 10446 47682 10498
rect 22542 10334 22594 10386
rect 24110 10334 24162 10386
rect 24446 10334 24498 10386
rect 25342 10334 25394 10386
rect 4478 10166 4530 10218
rect 4582 10166 4634 10218
rect 4686 10166 4738 10218
rect 35198 10166 35250 10218
rect 35302 10166 35354 10218
rect 35406 10166 35458 10218
rect 25454 9998 25506 10050
rect 25566 9998 25618 10050
rect 15710 9886 15762 9938
rect 17838 9886 17890 9938
rect 18286 9886 18338 9938
rect 22094 9886 22146 9938
rect 24222 9886 24274 9938
rect 24670 9886 24722 9938
rect 26126 9886 26178 9938
rect 27358 9886 27410 9938
rect 28702 9886 28754 9938
rect 32398 9886 32450 9938
rect 35310 9886 35362 9938
rect 36094 9886 36146 9938
rect 36542 9886 36594 9938
rect 37998 9886 38050 9938
rect 40126 9886 40178 9938
rect 41246 9886 41298 9938
rect 41806 9886 41858 9938
rect 45838 9886 45890 9938
rect 15038 9774 15090 9826
rect 21310 9774 21362 9826
rect 26910 9774 26962 9826
rect 29598 9774 29650 9826
rect 34638 9774 34690 9826
rect 34862 9774 34914 9826
rect 35086 9774 35138 9826
rect 35534 9774 35586 9826
rect 37214 9774 37266 9826
rect 42702 9774 42754 9826
rect 43374 9774 43426 9826
rect 43934 9774 43986 9826
rect 44830 9774 44882 9826
rect 45166 9774 45218 9826
rect 24670 9662 24722 9714
rect 24894 9662 24946 9714
rect 25230 9662 25282 9714
rect 26574 9662 26626 9714
rect 30270 9662 30322 9714
rect 40910 9662 40962 9714
rect 44270 9662 44322 9714
rect 45390 9662 45442 9714
rect 47854 9662 47906 9714
rect 48190 9662 48242 9714
rect 34974 9550 35026 9602
rect 42142 9550 42194 9602
rect 42254 9550 42306 9602
rect 42366 9550 42418 9602
rect 43262 9550 43314 9602
rect 45278 9550 45330 9602
rect 47630 9550 47682 9602
rect 19838 9382 19890 9434
rect 19942 9382 19994 9434
rect 20046 9382 20098 9434
rect 18286 9214 18338 9266
rect 19070 9214 19122 9266
rect 19854 9214 19906 9266
rect 21198 9214 21250 9266
rect 23214 9214 23266 9266
rect 23662 9214 23714 9266
rect 24558 9214 24610 9266
rect 35086 9214 35138 9266
rect 35646 9214 35698 9266
rect 37326 9214 37378 9266
rect 39566 9214 39618 9266
rect 18398 9102 18450 9154
rect 20078 9102 20130 9154
rect 20414 9102 20466 9154
rect 20638 9102 20690 9154
rect 21310 9102 21362 9154
rect 27470 9102 27522 9154
rect 34078 9102 34130 9154
rect 34190 9102 34242 9154
rect 38670 9102 38722 9154
rect 41694 9102 41746 9154
rect 46622 9102 46674 9154
rect 17950 8990 18002 9042
rect 18622 8990 18674 9042
rect 21086 8990 21138 9042
rect 21646 8990 21698 9042
rect 22990 8990 23042 9042
rect 23438 8990 23490 9042
rect 23774 8990 23826 9042
rect 24110 8990 24162 9042
rect 26686 8990 26738 9042
rect 33182 8990 33234 9042
rect 33406 8990 33458 9042
rect 33742 8990 33794 9042
rect 33854 8990 33906 9042
rect 34750 8990 34802 9042
rect 35870 8990 35922 9042
rect 39006 8990 39058 9042
rect 41022 8990 41074 9042
rect 47294 8990 47346 9042
rect 20190 8878 20242 8930
rect 25790 8878 25842 8930
rect 29598 8878 29650 8930
rect 33518 8878 33570 8930
rect 37774 8878 37826 8930
rect 43822 8878 43874 8930
rect 44494 8878 44546 8930
rect 24222 8766 24274 8818
rect 24782 8766 24834 8818
rect 4478 8598 4530 8650
rect 4582 8598 4634 8650
rect 4686 8598 4738 8650
rect 35198 8598 35250 8650
rect 35302 8598 35354 8650
rect 35406 8598 35458 8650
rect 25006 8430 25058 8482
rect 43598 8430 43650 8482
rect 44942 8430 44994 8482
rect 45502 8430 45554 8482
rect 18174 8318 18226 8370
rect 18846 8318 18898 8370
rect 19742 8318 19794 8370
rect 31502 8318 31554 8370
rect 33630 8318 33682 8370
rect 46062 8318 46114 8370
rect 15374 8206 15426 8258
rect 18734 8206 18786 8258
rect 18958 8206 19010 8258
rect 23774 8206 23826 8258
rect 23998 8206 24050 8258
rect 24334 8206 24386 8258
rect 24782 8206 24834 8258
rect 25230 8206 25282 8258
rect 25454 8206 25506 8258
rect 30270 8206 30322 8258
rect 31166 8206 31218 8258
rect 34414 8206 34466 8258
rect 34638 8206 34690 8258
rect 37550 8206 37602 8258
rect 39678 8206 39730 8258
rect 42478 8206 42530 8258
rect 43150 8206 43202 8258
rect 43822 8206 43874 8258
rect 44046 8206 44098 8258
rect 44830 8206 44882 8258
rect 45614 8206 45666 8258
rect 16046 8094 16098 8146
rect 19182 8094 19234 8146
rect 26686 8094 26738 8146
rect 30494 8094 30546 8146
rect 35086 8094 35138 8146
rect 35310 8094 35362 8146
rect 35646 8094 35698 8146
rect 37662 8094 37714 8146
rect 40238 8094 40290 8146
rect 42142 8094 42194 8146
rect 42702 8094 42754 8146
rect 44270 8094 44322 8146
rect 44942 8094 44994 8146
rect 23886 7982 23938 8034
rect 25902 7982 25954 8034
rect 27022 7982 27074 8034
rect 31054 7982 31106 8034
rect 34862 7982 34914 8034
rect 35982 7982 36034 8034
rect 36430 7982 36482 8034
rect 41246 7982 41298 8034
rect 42254 7982 42306 8034
rect 45502 7982 45554 8034
rect 19838 7814 19890 7866
rect 19942 7814 19994 7866
rect 20046 7814 20098 7866
rect 16382 7646 16434 7698
rect 17950 7646 18002 7698
rect 18062 7646 18114 7698
rect 27022 7646 27074 7698
rect 33406 7646 33458 7698
rect 35646 7646 35698 7698
rect 37550 7646 37602 7698
rect 38558 7646 38610 7698
rect 38894 7646 38946 7698
rect 39902 7646 39954 7698
rect 45390 7646 45442 7698
rect 16830 7534 16882 7586
rect 19966 7534 20018 7586
rect 23662 7534 23714 7586
rect 27470 7534 27522 7586
rect 28926 7534 28978 7586
rect 33182 7534 33234 7586
rect 33742 7534 33794 7586
rect 34078 7534 34130 7586
rect 34190 7534 34242 7586
rect 34750 7534 34802 7586
rect 34862 7534 34914 7586
rect 35422 7534 35474 7586
rect 36430 7534 36482 7586
rect 37886 7534 37938 7586
rect 40014 7534 40066 7586
rect 42590 7534 42642 7586
rect 42814 7534 42866 7586
rect 43486 7534 43538 7586
rect 16270 7422 16322 7474
rect 16606 7422 16658 7474
rect 18174 7422 18226 7474
rect 18510 7422 18562 7474
rect 19294 7422 19346 7474
rect 23886 7422 23938 7474
rect 24222 7422 24274 7474
rect 25454 7422 25506 7474
rect 27918 7422 27970 7474
rect 30046 7422 30098 7474
rect 31054 7422 31106 7474
rect 31502 7422 31554 7474
rect 31614 7422 31666 7474
rect 31950 7422 32002 7474
rect 32174 7422 32226 7474
rect 33070 7422 33122 7474
rect 34414 7422 34466 7474
rect 34526 7422 34578 7474
rect 35758 7422 35810 7474
rect 35982 7422 36034 7474
rect 36654 7422 36706 7474
rect 38110 7422 38162 7474
rect 39566 7422 39618 7474
rect 40238 7422 40290 7474
rect 41582 7422 41634 7474
rect 41806 7422 41858 7474
rect 42926 7422 42978 7474
rect 43150 7422 43202 7474
rect 43710 7422 43762 7474
rect 44046 7422 44098 7474
rect 17502 7310 17554 7362
rect 22094 7310 22146 7362
rect 22542 7310 22594 7362
rect 23774 7310 23826 7362
rect 30382 7310 30434 7362
rect 31838 7310 31890 7362
rect 43598 7310 43650 7362
rect 44494 7310 44546 7362
rect 44942 7310 44994 7362
rect 30606 7198 30658 7250
rect 30830 7198 30882 7250
rect 36878 7198 36930 7250
rect 37102 7198 37154 7250
rect 41246 7198 41298 7250
rect 42142 7198 42194 7250
rect 42254 7198 42306 7250
rect 4478 7030 4530 7082
rect 4582 7030 4634 7082
rect 4686 7030 4738 7082
rect 35198 7030 35250 7082
rect 35302 7030 35354 7082
rect 35406 7030 35458 7082
rect 22766 6862 22818 6914
rect 25790 6862 25842 6914
rect 31390 6862 31442 6914
rect 34638 6862 34690 6914
rect 42366 6862 42418 6914
rect 42478 6862 42530 6914
rect 19294 6750 19346 6802
rect 24334 6750 24386 6802
rect 25118 6750 25170 6802
rect 34414 6750 34466 6802
rect 35646 6750 35698 6802
rect 40686 6750 40738 6802
rect 41918 6750 41970 6802
rect 43374 6750 43426 6802
rect 44830 6750 44882 6802
rect 16494 6638 16546 6690
rect 17166 6638 17218 6690
rect 19742 6638 19794 6690
rect 20302 6638 20354 6690
rect 21982 6638 22034 6690
rect 22990 6638 23042 6690
rect 23886 6638 23938 6690
rect 24222 6638 24274 6690
rect 24894 6638 24946 6690
rect 25230 6638 25282 6690
rect 25566 6638 25618 6690
rect 26126 6638 26178 6690
rect 27022 6638 27074 6690
rect 27470 6638 27522 6690
rect 27694 6638 27746 6690
rect 28366 6638 28418 6690
rect 28590 6638 28642 6690
rect 29038 6638 29090 6690
rect 29262 6638 29314 6690
rect 29486 6638 29538 6690
rect 30046 6638 30098 6690
rect 31614 6638 31666 6690
rect 31950 6638 32002 6690
rect 32174 6638 32226 6690
rect 33182 6638 33234 6690
rect 35310 6638 35362 6690
rect 35870 6638 35922 6690
rect 37326 6638 37378 6690
rect 37998 6638 38050 6690
rect 40126 6638 40178 6690
rect 40462 6638 40514 6690
rect 41470 6638 41522 6690
rect 41806 6638 41858 6690
rect 42030 6638 42082 6690
rect 43038 6638 43090 6690
rect 43262 6638 43314 6690
rect 43822 6638 43874 6690
rect 47630 6638 47682 6690
rect 24670 6526 24722 6578
rect 29710 6526 29762 6578
rect 30270 6526 30322 6578
rect 31054 6526 31106 6578
rect 34862 6526 34914 6578
rect 37550 6526 37602 6578
rect 37774 6526 37826 6578
rect 38782 6526 38834 6578
rect 44158 6526 44210 6578
rect 44270 6526 44322 6578
rect 46958 6526 47010 6578
rect 21534 6414 21586 6466
rect 22094 6414 22146 6466
rect 22430 6414 22482 6466
rect 23438 6414 23490 6466
rect 23662 6414 23714 6466
rect 23774 6414 23826 6466
rect 27358 6414 27410 6466
rect 28030 6414 28082 6466
rect 30158 6414 30210 6466
rect 30494 6414 30546 6466
rect 32062 6414 32114 6466
rect 32398 6414 32450 6466
rect 32846 6414 32898 6466
rect 34750 6414 34802 6466
rect 36542 6414 36594 6466
rect 38334 6414 38386 6466
rect 38558 6414 38610 6466
rect 38670 6414 38722 6466
rect 39678 6414 39730 6466
rect 39902 6414 39954 6466
rect 40014 6414 40066 6466
rect 41022 6414 41074 6466
rect 42814 6414 42866 6466
rect 19838 6246 19890 6298
rect 19942 6246 19994 6298
rect 20046 6246 20098 6298
rect 18398 6078 18450 6130
rect 20638 6078 20690 6130
rect 24670 6078 24722 6130
rect 27918 6078 27970 6130
rect 32622 6078 32674 6130
rect 33070 6078 33122 6130
rect 42254 6078 42306 6130
rect 19518 5966 19570 6018
rect 19854 5966 19906 6018
rect 22094 5966 22146 6018
rect 26686 5966 26738 6018
rect 27022 5966 27074 6018
rect 27246 5966 27298 6018
rect 29262 5966 29314 6018
rect 29598 5966 29650 6018
rect 31278 5966 31330 6018
rect 31502 5966 31554 6018
rect 33742 5966 33794 6018
rect 34078 5966 34130 6018
rect 34974 5966 35026 6018
rect 35534 5966 35586 6018
rect 36318 5966 36370 6018
rect 37438 5966 37490 6018
rect 37774 5966 37826 6018
rect 38222 5966 38274 6018
rect 38670 5966 38722 6018
rect 41246 5966 41298 6018
rect 41582 5966 41634 6018
rect 18622 5854 18674 5906
rect 18846 5854 18898 5906
rect 19294 5854 19346 5906
rect 19966 5854 20018 5906
rect 20414 5854 20466 5906
rect 20526 5854 20578 5906
rect 20974 5854 21026 5906
rect 21310 5854 21362 5906
rect 26014 5854 26066 5906
rect 27134 5854 27186 5906
rect 27694 5854 27746 5906
rect 28366 5854 28418 5906
rect 29038 5854 29090 5906
rect 29150 5854 29202 5906
rect 29822 5854 29874 5906
rect 29934 5854 29986 5906
rect 31054 5854 31106 5906
rect 31166 5854 31218 5906
rect 31838 5854 31890 5906
rect 31950 5854 32002 5906
rect 33406 5854 33458 5906
rect 34638 5854 34690 5906
rect 34750 5854 34802 5906
rect 35310 5854 35362 5906
rect 35422 5854 35474 5906
rect 36094 5854 36146 5906
rect 36654 5854 36706 5906
rect 36766 5854 36818 5906
rect 36990 5854 37042 5906
rect 38446 5854 38498 5906
rect 39006 5854 39058 5906
rect 39118 5854 39170 5906
rect 39454 5854 39506 5906
rect 39790 5854 39842 5906
rect 40014 5854 40066 5906
rect 40910 5854 40962 5906
rect 41022 5854 41074 5906
rect 41806 5854 41858 5906
rect 42590 5854 42642 5906
rect 42814 5854 42866 5906
rect 19070 5742 19122 5794
rect 19630 5742 19682 5794
rect 24222 5742 24274 5794
rect 25454 5742 25506 5794
rect 26350 5742 26402 5794
rect 27806 5742 27858 5794
rect 38110 5742 38162 5794
rect 41918 5742 41970 5794
rect 25790 5630 25842 5682
rect 26462 5630 26514 5682
rect 35982 5630 36034 5682
rect 4478 5462 4530 5514
rect 4582 5462 4634 5514
rect 4686 5462 4738 5514
rect 35198 5462 35250 5514
rect 35302 5462 35354 5514
rect 35406 5462 35458 5514
rect 24222 5294 24274 5346
rect 41470 5294 41522 5346
rect 41806 5294 41858 5346
rect 18622 5182 18674 5234
rect 20750 5182 20802 5234
rect 21422 5182 21474 5234
rect 22318 5182 22370 5234
rect 25006 5182 25058 5234
rect 28366 5182 28418 5234
rect 29262 5182 29314 5234
rect 32734 5182 32786 5234
rect 33518 5182 33570 5234
rect 36318 5182 36370 5234
rect 37214 5182 37266 5234
rect 37438 5182 37490 5234
rect 37886 5182 37938 5234
rect 41134 5182 41186 5234
rect 41694 5182 41746 5234
rect 42814 5182 42866 5234
rect 44046 5182 44098 5234
rect 17950 5070 18002 5122
rect 21870 5070 21922 5122
rect 23326 5070 23378 5122
rect 23438 5070 23490 5122
rect 23774 5070 23826 5122
rect 24110 5070 24162 5122
rect 25118 5070 25170 5122
rect 25566 5070 25618 5122
rect 29934 5070 29986 5122
rect 33182 5070 33234 5122
rect 35422 5070 35474 5122
rect 35534 5070 35586 5122
rect 37550 5070 37602 5122
rect 40014 5070 40066 5122
rect 40798 5070 40850 5122
rect 21310 4958 21362 5010
rect 21534 4958 21586 5010
rect 23214 4958 23266 5010
rect 24558 4958 24610 5010
rect 24782 4958 24834 5010
rect 26238 4958 26290 5010
rect 29150 4958 29202 5010
rect 30606 4958 30658 5010
rect 35646 4958 35698 5010
rect 33630 4846 33682 4898
rect 35870 4846 35922 4898
rect 36430 4846 36482 4898
rect 41246 4846 41298 4898
rect 42926 4846 42978 4898
rect 19838 4678 19890 4730
rect 19942 4678 19994 4730
rect 20046 4678 20098 4730
rect 25342 4510 25394 4562
rect 26574 4510 26626 4562
rect 31054 4510 31106 4562
rect 39902 4510 39954 4562
rect 19070 4398 19122 4450
rect 26686 4398 26738 4450
rect 28142 4398 28194 4450
rect 31166 4398 31218 4450
rect 33854 4398 33906 4450
rect 38446 4398 38498 4450
rect 41694 4398 41746 4450
rect 46286 4398 46338 4450
rect 18286 4286 18338 4338
rect 21646 4286 21698 4338
rect 27358 4286 27410 4338
rect 33182 4286 33234 4338
rect 39230 4286 39282 4338
rect 40126 4286 40178 4338
rect 40910 4286 40962 4338
rect 47070 4286 47122 4338
rect 47630 4286 47682 4338
rect 48190 4286 48242 4338
rect 21198 4174 21250 4226
rect 22318 4174 22370 4226
rect 24446 4174 24498 4226
rect 30270 4174 30322 4226
rect 35982 4174 36034 4226
rect 36318 4174 36370 4226
rect 43822 4174 43874 4226
rect 44158 4174 44210 4226
rect 4478 3894 4530 3946
rect 4582 3894 4634 3946
rect 4686 3894 4738 3946
rect 35198 3894 35250 3946
rect 35302 3894 35354 3946
rect 35406 3894 35458 3946
rect 22766 3726 22818 3778
rect 21534 3614 21586 3666
rect 22878 3614 22930 3666
rect 36318 3614 36370 3666
rect 40014 3614 40066 3666
rect 43934 3614 43986 3666
rect 48302 3614 48354 3666
rect 19838 3110 19890 3162
rect 19942 3110 19994 3162
rect 20046 3110 20098 3162
<< metal2 >>
rect 3584 59200 3696 60000
rect 5152 59200 5264 60000
rect 6720 59200 6832 60000
rect 8288 59200 8400 60000
rect 9856 59200 9968 60000
rect 11424 59200 11536 60000
rect 12992 59200 13104 60000
rect 14560 59200 14672 60000
rect 16128 59200 16240 60000
rect 17696 59200 17808 60000
rect 19264 59200 19376 60000
rect 20832 59200 20944 60000
rect 22400 59200 22512 60000
rect 23968 59200 24080 60000
rect 25536 59200 25648 60000
rect 27104 59200 27216 60000
rect 28672 59200 28784 60000
rect 30240 59200 30352 60000
rect 31808 59200 31920 60000
rect 33376 59200 33488 60000
rect 34944 59200 35056 60000
rect 36512 59200 36624 60000
rect 38080 59200 38192 60000
rect 39648 59200 39760 60000
rect 41216 59200 41328 60000
rect 42784 59200 42896 60000
rect 44352 59200 44464 60000
rect 44716 59276 45220 59332
rect 3612 56308 3668 59200
rect 5180 57764 5236 59200
rect 5180 57708 5572 57764
rect 3836 56308 3892 56318
rect 3612 56306 3892 56308
rect 3612 56254 3838 56306
rect 3890 56254 3892 56306
rect 3612 56252 3892 56254
rect 3836 56242 3892 56252
rect 5516 56306 5572 57708
rect 5516 56254 5518 56306
rect 5570 56254 5572 56306
rect 5516 56242 5572 56254
rect 6748 56308 6804 59200
rect 6972 56308 7028 56318
rect 6748 56306 7028 56308
rect 6748 56254 6974 56306
rect 7026 56254 7028 56306
rect 6748 56252 7028 56254
rect 8316 56308 8372 59200
rect 8540 56308 8596 56318
rect 8316 56306 8596 56308
rect 8316 56254 8542 56306
rect 8594 56254 8596 56306
rect 8316 56252 8596 56254
rect 9884 56308 9940 59200
rect 10108 56308 10164 56318
rect 9884 56306 10164 56308
rect 9884 56254 10110 56306
rect 10162 56254 10164 56306
rect 9884 56252 10164 56254
rect 11452 56308 11508 59200
rect 13020 57764 13076 59200
rect 12572 57708 13076 57764
rect 11676 56308 11732 56318
rect 11452 56306 11732 56308
rect 11452 56254 11678 56306
rect 11730 56254 11732 56306
rect 11452 56252 11732 56254
rect 6972 56242 7028 56252
rect 8540 56242 8596 56252
rect 10108 56242 10164 56252
rect 11676 56242 11732 56252
rect 12572 56306 12628 57708
rect 12572 56254 12574 56306
rect 12626 56254 12628 56306
rect 12572 56242 12628 56254
rect 13468 57090 13524 57102
rect 13468 57038 13470 57090
rect 13522 57038 13524 57090
rect 13468 56306 13524 57038
rect 14588 57090 14644 59200
rect 14588 57038 14590 57090
rect 14642 57038 14644 57090
rect 14588 57026 14644 57038
rect 13468 56254 13470 56306
rect 13522 56254 13524 56306
rect 13468 56242 13524 56254
rect 15372 56308 15428 56318
rect 15372 56214 15428 56252
rect 16156 56308 16212 59200
rect 17724 56308 17780 59200
rect 17724 56252 18228 56308
rect 16156 56242 16212 56252
rect 16044 56082 16100 56094
rect 16044 56030 16046 56082
rect 16098 56030 16100 56082
rect 4476 55692 4740 55702
rect 4532 55636 4580 55692
rect 4636 55636 4684 55692
rect 4476 55626 4740 55636
rect 13804 55356 14532 55412
rect 9660 55300 9716 55310
rect 9884 55300 9940 55310
rect 10780 55300 10836 55310
rect 9660 55298 9940 55300
rect 9660 55246 9662 55298
rect 9714 55246 9886 55298
rect 9938 55246 9940 55298
rect 9660 55244 9940 55246
rect 9660 55234 9716 55244
rect 9884 55234 9940 55244
rect 10220 55298 10836 55300
rect 10220 55246 10782 55298
rect 10834 55246 10836 55298
rect 10220 55244 10836 55246
rect 9324 55186 9380 55198
rect 9324 55134 9326 55186
rect 9378 55134 9380 55186
rect 6860 55076 6916 55086
rect 6860 54626 6916 55020
rect 9324 54852 9380 55134
rect 10108 55186 10164 55198
rect 10108 55134 10110 55186
rect 10162 55134 10164 55186
rect 9436 55076 9492 55086
rect 9436 55074 10052 55076
rect 9436 55022 9438 55074
rect 9490 55022 10052 55074
rect 9436 55020 10052 55022
rect 9436 55010 9492 55020
rect 9324 54786 9380 54796
rect 6860 54574 6862 54626
rect 6914 54574 6916 54626
rect 6860 54562 6916 54574
rect 9884 54626 9940 54638
rect 9884 54574 9886 54626
rect 9938 54574 9940 54626
rect 6188 54514 6244 54526
rect 6188 54462 6190 54514
rect 6242 54462 6244 54514
rect 4476 54124 4740 54134
rect 4532 54068 4580 54124
rect 4636 54068 4684 54124
rect 4476 54058 4740 54068
rect 4172 52948 4228 52958
rect 1596 52388 1652 52398
rect 1484 48804 1540 48814
rect 1484 21812 1540 48748
rect 1484 21746 1540 21756
rect 1596 19460 1652 52332
rect 1820 51268 1876 51278
rect 1708 51266 1876 51268
rect 1708 51214 1822 51266
rect 1874 51214 1876 51266
rect 1708 51212 1876 51214
rect 1708 50482 1764 51212
rect 1820 51202 1876 51212
rect 3724 51268 3780 51278
rect 2268 50594 2324 50606
rect 2268 50542 2270 50594
rect 2322 50542 2324 50594
rect 1708 50430 1710 50482
rect 1762 50430 1764 50482
rect 1708 49812 1764 50430
rect 1708 49746 1764 49756
rect 1820 50484 1876 50494
rect 1820 49810 1876 50428
rect 2156 50036 2212 50046
rect 1820 49758 1822 49810
rect 1874 49758 1876 49810
rect 1820 47572 1876 49758
rect 1820 47458 1876 47516
rect 1820 47406 1822 47458
rect 1874 47406 1876 47458
rect 1820 47394 1876 47406
rect 2044 49980 2156 50036
rect 1820 44322 1876 44334
rect 1820 44270 1822 44322
rect 1874 44270 1876 44322
rect 1820 41972 1876 44270
rect 2044 43708 2100 49980
rect 2156 49970 2212 49980
rect 2268 48804 2324 50542
rect 2492 49698 2548 49710
rect 2492 49646 2494 49698
rect 2546 49646 2548 49698
rect 2492 49252 2548 49646
rect 2492 49186 2548 49196
rect 2268 48738 2324 48748
rect 3724 48802 3780 51212
rect 4172 50484 4228 52892
rect 6188 52948 6244 54462
rect 8988 54402 9044 54414
rect 8988 54350 8990 54402
rect 9042 54350 9044 54402
rect 8988 53844 9044 54350
rect 9660 53844 9716 53854
rect 9884 53844 9940 54574
rect 8988 53842 9940 53844
rect 8988 53790 9662 53842
rect 9714 53790 9940 53842
rect 8988 53788 9940 53790
rect 9660 53778 9716 53788
rect 9996 53732 10052 55020
rect 9772 53730 10052 53732
rect 9772 53678 9998 53730
rect 10050 53678 10052 53730
rect 9772 53676 10052 53678
rect 9548 53620 9604 53630
rect 9772 53620 9828 53676
rect 9996 53666 10052 53676
rect 9548 53618 9828 53620
rect 9548 53566 9550 53618
rect 9602 53566 9828 53618
rect 9548 53564 9828 53566
rect 10108 53620 10164 55134
rect 10220 53842 10276 55244
rect 10780 55234 10836 55244
rect 13804 55298 13860 55356
rect 13804 55246 13806 55298
rect 13858 55246 13860 55298
rect 13804 55234 13860 55246
rect 10892 55188 10948 55198
rect 10892 55074 10948 55132
rect 11676 55186 11732 55198
rect 11676 55134 11678 55186
rect 11730 55134 11732 55186
rect 10892 55022 10894 55074
rect 10946 55022 10948 55074
rect 10332 54852 10388 54862
rect 10332 54514 10388 54796
rect 10332 54462 10334 54514
rect 10386 54462 10388 54514
rect 10332 53956 10388 54462
rect 10332 53954 10612 53956
rect 10332 53902 10334 53954
rect 10386 53902 10612 53954
rect 10332 53900 10612 53902
rect 10332 53890 10388 53900
rect 10220 53790 10222 53842
rect 10274 53790 10276 53842
rect 10220 53778 10276 53790
rect 9548 53554 9604 53564
rect 9212 53506 9268 53518
rect 9212 53454 9214 53506
rect 9266 53454 9268 53506
rect 7420 53058 7476 53070
rect 7420 53006 7422 53058
rect 7474 53006 7476 53058
rect 6188 52882 6244 52892
rect 7196 52948 7252 52958
rect 7196 52946 7364 52948
rect 7196 52894 7198 52946
rect 7250 52894 7364 52946
rect 7196 52892 7364 52894
rect 7196 52882 7252 52892
rect 4844 52834 4900 52846
rect 4844 52782 4846 52834
rect 4898 52782 4900 52834
rect 4476 52556 4740 52566
rect 4532 52500 4580 52556
rect 4636 52500 4684 52556
rect 4476 52490 4740 52500
rect 4844 52276 4900 52782
rect 6972 52834 7028 52846
rect 6972 52782 6974 52834
rect 7026 52782 7028 52834
rect 6972 52724 7028 52782
rect 6972 52658 7028 52668
rect 6748 52388 6804 52398
rect 6748 52386 7252 52388
rect 6748 52334 6750 52386
rect 6802 52334 7252 52386
rect 6748 52332 7252 52334
rect 6748 52322 6804 52332
rect 4844 52210 4900 52220
rect 6076 52276 6132 52286
rect 6076 52182 6132 52220
rect 5964 52162 6020 52174
rect 5964 52110 5966 52162
rect 6018 52110 6020 52162
rect 5628 52050 5684 52062
rect 5628 51998 5630 52050
rect 5682 51998 5684 52050
rect 5628 51602 5684 51998
rect 5628 51550 5630 51602
rect 5682 51550 5684 51602
rect 5628 51538 5684 51550
rect 5740 51604 5796 51614
rect 5740 51510 5796 51548
rect 5068 51378 5124 51390
rect 5068 51326 5070 51378
rect 5122 51326 5124 51378
rect 4844 51268 4900 51278
rect 5068 51268 5124 51326
rect 5516 51380 5572 51390
rect 5516 51286 5572 51324
rect 5964 51380 6020 52110
rect 6860 52164 6916 52174
rect 6860 52162 7028 52164
rect 6860 52110 6862 52162
rect 6914 52110 7028 52162
rect 6860 52108 7028 52110
rect 6860 52098 6916 52108
rect 6188 52050 6244 52062
rect 6188 51998 6190 52050
rect 6242 51998 6244 52050
rect 6188 51604 6244 51998
rect 6748 51938 6804 51950
rect 6748 51886 6750 51938
rect 6802 51886 6804 51938
rect 6244 51548 6356 51604
rect 6188 51538 6244 51548
rect 5964 51314 6020 51324
rect 6076 51378 6132 51390
rect 6076 51326 6078 51378
rect 6130 51326 6132 51378
rect 4900 51212 5124 51268
rect 4844 51174 4900 51212
rect 4476 50988 4740 50998
rect 4532 50932 4580 50988
rect 4636 50932 4684 50988
rect 4476 50922 4740 50932
rect 5964 50708 6020 50718
rect 5740 50706 6020 50708
rect 5740 50654 5966 50706
rect 6018 50654 6020 50706
rect 5740 50652 6020 50654
rect 5628 50594 5684 50606
rect 5628 50542 5630 50594
rect 5682 50542 5684 50594
rect 4172 50418 4228 50428
rect 4844 50484 4900 50522
rect 4844 50418 4900 50428
rect 5628 49922 5684 50542
rect 5628 49870 5630 49922
rect 5682 49870 5684 49922
rect 4620 49700 4676 49710
rect 4620 49606 4676 49644
rect 4956 49700 5012 49710
rect 4476 49420 4740 49430
rect 4532 49364 4580 49420
rect 4636 49364 4684 49420
rect 4476 49354 4740 49364
rect 4732 49028 4788 49038
rect 4732 48934 4788 48972
rect 4956 48914 5012 49644
rect 4956 48862 4958 48914
rect 5010 48862 5012 48914
rect 4956 48850 5012 48862
rect 5068 49698 5124 49710
rect 5068 49646 5070 49698
rect 5122 49646 5124 49698
rect 5068 48916 5124 49646
rect 5628 49700 5684 49870
rect 5628 49634 5684 49644
rect 5516 49028 5572 49038
rect 5516 48934 5572 48972
rect 5068 48850 5124 48860
rect 5740 48916 5796 50652
rect 5964 50642 6020 50652
rect 6076 50484 6132 51326
rect 6300 50706 6356 51548
rect 6300 50654 6302 50706
rect 6354 50654 6356 50706
rect 6300 50642 6356 50654
rect 6412 51380 6468 51390
rect 6748 51380 6804 51886
rect 6860 51940 6916 51950
rect 6972 51940 7028 52108
rect 7196 52162 7252 52332
rect 7196 52110 7198 52162
rect 7250 52110 7252 52162
rect 7196 52098 7252 52110
rect 7308 51940 7364 52892
rect 6972 51884 7364 51940
rect 6860 51490 6916 51884
rect 7420 51828 7476 53006
rect 7532 52948 7588 52958
rect 7980 52948 8036 52958
rect 7532 52946 7812 52948
rect 7532 52894 7534 52946
rect 7586 52894 7812 52946
rect 7532 52892 7812 52894
rect 7532 52882 7588 52892
rect 7644 52388 7700 52398
rect 7644 52274 7700 52332
rect 7644 52222 7646 52274
rect 7698 52222 7700 52274
rect 7644 52210 7700 52222
rect 7532 51940 7588 51950
rect 7532 51828 7588 51884
rect 6860 51438 6862 51490
rect 6914 51438 6916 51490
rect 6860 51426 6916 51438
rect 6972 51772 7588 51828
rect 7756 51938 7812 52892
rect 7980 52854 8036 52892
rect 8988 52948 9044 52958
rect 9212 52948 9268 53454
rect 10108 53396 10164 53564
rect 9044 52892 9268 52948
rect 9996 53340 10164 53396
rect 8092 52724 8148 52734
rect 8148 52668 8260 52724
rect 8092 52658 8148 52668
rect 8204 52274 8260 52668
rect 8204 52222 8206 52274
rect 8258 52222 8260 52274
rect 8204 52210 8260 52222
rect 8988 52274 9044 52892
rect 8988 52222 8990 52274
rect 9042 52222 9044 52274
rect 8988 52210 9044 52222
rect 9660 52164 9716 52174
rect 9660 52162 9828 52164
rect 9660 52110 9662 52162
rect 9714 52110 9828 52162
rect 9660 52108 9828 52110
rect 9660 52098 9716 52108
rect 9324 52050 9380 52062
rect 9324 51998 9326 52050
rect 9378 51998 9380 52050
rect 7756 51886 7758 51938
rect 7810 51886 7812 51938
rect 6468 51324 6804 51380
rect 6076 50418 6132 50428
rect 5852 50370 5908 50382
rect 5852 50318 5854 50370
rect 5906 50318 5908 50370
rect 5852 49140 5908 50318
rect 6412 49250 6468 51324
rect 6972 50594 7028 51772
rect 6972 50542 6974 50594
rect 7026 50542 7028 50594
rect 6972 50530 7028 50542
rect 7084 50706 7140 50718
rect 7084 50654 7086 50706
rect 7138 50654 7140 50706
rect 7084 50428 7140 50654
rect 6748 50372 7140 50428
rect 7756 50428 7812 51886
rect 8092 51940 8148 51950
rect 8092 51846 8148 51884
rect 8316 51380 8372 51390
rect 8316 50594 8372 51324
rect 9324 51380 9380 51998
rect 9324 51314 9380 51324
rect 9436 51938 9492 51950
rect 9436 51886 9438 51938
rect 9490 51886 9492 51938
rect 8988 51268 9044 51278
rect 8988 51156 9044 51212
rect 8316 50542 8318 50594
rect 8370 50542 8372 50594
rect 8316 50530 8372 50542
rect 8540 51100 9044 51156
rect 8428 50484 8484 50494
rect 8540 50484 8596 51100
rect 8652 50764 9044 50820
rect 8652 50594 8708 50764
rect 8652 50542 8654 50594
rect 8706 50542 8708 50594
rect 8652 50530 8708 50542
rect 8876 50596 8932 50606
rect 8428 50482 8596 50484
rect 8428 50430 8430 50482
rect 8482 50430 8596 50482
rect 8428 50428 8596 50430
rect 7756 50372 8036 50428
rect 8428 50418 8484 50428
rect 6748 50306 6804 50316
rect 7980 50306 8036 50316
rect 6412 49198 6414 49250
rect 6466 49198 6468 49250
rect 6412 49186 6468 49198
rect 6524 49810 6580 49822
rect 6524 49758 6526 49810
rect 6578 49758 6580 49810
rect 6188 49140 6244 49150
rect 5852 49138 6244 49140
rect 5852 49086 6190 49138
rect 6242 49086 6244 49138
rect 5852 49084 6244 49086
rect 6188 49074 6244 49084
rect 5740 48850 5796 48860
rect 6300 49028 6356 49038
rect 6524 49028 6580 49758
rect 7196 49700 7252 49710
rect 7196 49698 7364 49700
rect 7196 49646 7198 49698
rect 7250 49646 7364 49698
rect 7196 49644 7364 49646
rect 7196 49634 7252 49644
rect 7308 49250 7364 49644
rect 7308 49198 7310 49250
rect 7362 49198 7364 49250
rect 7308 49186 7364 49198
rect 7868 49698 7924 49710
rect 7868 49646 7870 49698
rect 7922 49646 7924 49698
rect 7420 49140 7476 49150
rect 7420 49046 7476 49084
rect 6300 49026 6580 49028
rect 6300 48974 6302 49026
rect 6354 48974 6580 49026
rect 6300 48972 6580 48974
rect 3724 48750 3726 48802
rect 3778 48750 3780 48802
rect 3052 48468 3108 48478
rect 2156 48466 3108 48468
rect 2156 48414 3054 48466
rect 3106 48414 3108 48466
rect 2156 48412 3108 48414
rect 2156 48242 2212 48412
rect 3052 48402 3108 48412
rect 3388 48356 3444 48366
rect 3724 48356 3780 48750
rect 5068 48692 5124 48702
rect 4396 48524 5012 48580
rect 4396 48466 4452 48524
rect 4396 48414 4398 48466
rect 4450 48414 4452 48466
rect 4396 48402 4452 48414
rect 3388 48354 3780 48356
rect 3388 48302 3390 48354
rect 3442 48302 3780 48354
rect 3388 48300 3780 48302
rect 3948 48354 4004 48366
rect 3948 48302 3950 48354
rect 4002 48302 4004 48354
rect 2156 48190 2158 48242
rect 2210 48190 2212 48242
rect 2156 48178 2212 48190
rect 2380 48244 2436 48254
rect 2380 48150 2436 48188
rect 2716 48244 2772 48254
rect 2940 48244 2996 48254
rect 2716 48242 2996 48244
rect 2716 48190 2718 48242
rect 2770 48190 2942 48242
rect 2994 48190 2996 48242
rect 2716 48188 2996 48190
rect 2716 48178 2772 48188
rect 2492 48130 2548 48142
rect 2492 48078 2494 48130
rect 2546 48078 2548 48130
rect 2492 47570 2548 48078
rect 2492 47518 2494 47570
rect 2546 47518 2548 47570
rect 2492 47506 2548 47518
rect 2828 46786 2884 48188
rect 2940 48178 2996 48188
rect 3164 48244 3220 48254
rect 3164 48150 3220 48188
rect 2828 46734 2830 46786
rect 2882 46734 2884 46786
rect 2828 46722 2884 46734
rect 3276 47460 3332 47470
rect 3276 46674 3332 47404
rect 3276 46622 3278 46674
rect 3330 46622 3332 46674
rect 3276 46610 3332 46622
rect 2268 45778 2324 45790
rect 2268 45726 2270 45778
rect 2322 45726 2324 45778
rect 2268 45220 2324 45726
rect 2604 45778 2660 45790
rect 2604 45726 2606 45778
rect 2658 45726 2660 45778
rect 2492 45666 2548 45678
rect 2492 45614 2494 45666
rect 2546 45614 2548 45666
rect 2380 45220 2436 45230
rect 2268 45164 2380 45220
rect 2380 45126 2436 45164
rect 2492 44434 2548 45614
rect 2604 45108 2660 45726
rect 2828 45778 2884 45790
rect 2828 45726 2830 45778
rect 2882 45726 2884 45778
rect 2828 45332 2884 45726
rect 2828 45266 2884 45276
rect 3276 45666 3332 45678
rect 3276 45614 3278 45666
rect 3330 45614 3332 45666
rect 2604 45042 2660 45052
rect 3052 45106 3108 45118
rect 3052 45054 3054 45106
rect 3106 45054 3108 45106
rect 3052 44996 3108 45054
rect 3276 45108 3332 45614
rect 3276 45042 3332 45052
rect 3052 44930 3108 44940
rect 3164 44994 3220 45006
rect 3164 44942 3166 44994
rect 3218 44942 3220 44994
rect 3164 44884 3220 44942
rect 3276 44884 3332 44894
rect 3164 44828 3276 44884
rect 3276 44818 3332 44828
rect 3388 44772 3444 48300
rect 3948 48244 4004 48302
rect 4844 48354 4900 48366
rect 4844 48302 4846 48354
rect 4898 48302 4900 48354
rect 3948 47236 4004 48188
rect 4172 48244 4228 48254
rect 4172 47460 4228 48188
rect 4844 48244 4900 48302
rect 4844 48178 4900 48188
rect 4956 48242 5012 48524
rect 4956 48190 4958 48242
rect 5010 48190 5012 48242
rect 4172 47394 4228 47404
rect 4284 48130 4340 48142
rect 4284 48078 4286 48130
rect 4338 48078 4340 48130
rect 3948 47180 4228 47236
rect 3724 46676 3780 46686
rect 3724 46582 3780 46620
rect 4172 45892 4228 47180
rect 4284 46452 4340 48078
rect 4844 48018 4900 48030
rect 4844 47966 4846 48018
rect 4898 47966 4900 48018
rect 4476 47852 4740 47862
rect 4532 47796 4580 47852
rect 4636 47796 4684 47852
rect 4476 47786 4740 47796
rect 4620 47570 4676 47582
rect 4620 47518 4622 47570
rect 4674 47518 4676 47570
rect 4620 47460 4676 47518
rect 4620 47394 4676 47404
rect 4844 47236 4900 47966
rect 4508 47180 4900 47236
rect 4508 46674 4564 47180
rect 4508 46622 4510 46674
rect 4562 46622 4564 46674
rect 4508 46610 4564 46622
rect 4844 46676 4900 46686
rect 4956 46676 5012 48190
rect 5068 47572 5124 48636
rect 5852 48692 5908 48702
rect 5852 48242 5908 48636
rect 5852 48190 5854 48242
rect 5906 48190 5908 48242
rect 5852 48178 5908 48190
rect 5068 47478 5124 47516
rect 5068 46900 5124 46910
rect 6300 46900 6356 48972
rect 7532 48804 7588 48814
rect 7868 48804 7924 49646
rect 8764 49252 8820 49262
rect 8876 49252 8932 50540
rect 8988 50594 9044 50764
rect 9436 50706 9492 51886
rect 9772 51268 9828 52108
rect 9884 51490 9940 51502
rect 9884 51438 9886 51490
rect 9938 51438 9940 51490
rect 9884 51268 9940 51438
rect 9828 51212 9940 51268
rect 9772 51202 9828 51212
rect 9436 50654 9438 50706
rect 9490 50654 9492 50706
rect 9436 50642 9492 50654
rect 8988 50542 8990 50594
rect 9042 50542 9044 50594
rect 8988 50530 9044 50542
rect 9884 50596 9940 50606
rect 9884 50502 9940 50540
rect 9996 50482 10052 53340
rect 10332 52274 10388 52286
rect 10332 52222 10334 52274
rect 10386 52222 10388 52274
rect 10332 52164 10388 52222
rect 10332 52098 10388 52108
rect 10444 52276 10500 52286
rect 10444 52050 10500 52220
rect 10444 51998 10446 52050
rect 10498 51998 10500 52050
rect 10444 51986 10500 51998
rect 10556 51604 10612 53900
rect 10892 53618 10948 55022
rect 11452 55074 11508 55086
rect 11452 55022 11454 55074
rect 11506 55022 11508 55074
rect 11452 54964 11508 55022
rect 11564 55076 11620 55086
rect 11564 54982 11620 55020
rect 11452 54898 11508 54908
rect 11676 54738 11732 55134
rect 13468 55188 13524 55198
rect 13468 55094 13524 55132
rect 14028 55186 14084 55198
rect 14028 55134 14030 55186
rect 14082 55134 14084 55186
rect 11676 54686 11678 54738
rect 11730 54686 11732 54738
rect 11676 54674 11732 54686
rect 12236 55074 12292 55086
rect 12236 55022 12238 55074
rect 12290 55022 12292 55074
rect 12236 54964 12292 55022
rect 12236 54628 12292 54908
rect 13692 55074 13748 55086
rect 13692 55022 13694 55074
rect 13746 55022 13748 55074
rect 13692 54740 13748 55022
rect 13692 54684 13972 54740
rect 12236 54572 12740 54628
rect 11116 54514 11172 54526
rect 11116 54462 11118 54514
rect 11170 54462 11172 54514
rect 10892 53566 10894 53618
rect 10946 53566 10948 53618
rect 10892 53554 10948 53566
rect 11004 54292 11060 54302
rect 11004 53506 11060 54236
rect 11116 53620 11172 54462
rect 12684 54516 12740 54572
rect 13916 54626 13972 54684
rect 13916 54574 13918 54626
rect 13970 54574 13972 54626
rect 13916 54562 13972 54574
rect 12796 54516 12852 54526
rect 12684 54514 12852 54516
rect 12684 54462 12798 54514
rect 12850 54462 12852 54514
rect 12684 54460 12852 54462
rect 12572 54402 12628 54414
rect 12572 54350 12574 54402
rect 12626 54350 12628 54402
rect 12460 54292 12516 54302
rect 12460 54198 12516 54236
rect 11116 53554 11172 53564
rect 11228 53732 11284 53742
rect 11004 53454 11006 53506
rect 11058 53454 11060 53506
rect 11004 53442 11060 53454
rect 11228 52948 11284 53676
rect 12236 53730 12292 53742
rect 12236 53678 12238 53730
rect 12290 53678 12292 53730
rect 12236 53396 12292 53678
rect 12460 53620 12516 53630
rect 12460 53526 12516 53564
rect 12236 53330 12292 53340
rect 12572 53172 12628 54350
rect 12796 53508 12852 54460
rect 13132 54514 13188 54526
rect 13132 54462 13134 54514
rect 13186 54462 13188 54514
rect 13132 53844 13188 54462
rect 13804 54404 13860 54414
rect 13132 53778 13188 53788
rect 13692 53844 13748 53854
rect 13804 53844 13860 54348
rect 13748 53788 13860 53844
rect 13692 53778 13748 53788
rect 12796 53442 12852 53452
rect 13580 53508 13636 53518
rect 12012 53116 12628 53172
rect 12012 53058 12068 53116
rect 12012 53006 12014 53058
rect 12066 53006 12068 53058
rect 12012 52994 12068 53006
rect 11228 52854 11284 52892
rect 11116 52276 11172 52286
rect 11116 52182 11172 52220
rect 13580 52276 13636 53452
rect 10668 52052 10724 52062
rect 10668 52050 11060 52052
rect 10668 51998 10670 52050
rect 10722 51998 11060 52050
rect 10668 51996 11060 51998
rect 10668 51986 10724 51996
rect 11004 51716 11060 51996
rect 11004 51660 11508 51716
rect 10556 51548 11060 51604
rect 11004 51492 11060 51548
rect 11452 51602 11508 51660
rect 11452 51550 11454 51602
rect 11506 51550 11508 51602
rect 11452 51538 11508 51550
rect 13580 51604 13636 52220
rect 13580 51538 13636 51548
rect 13804 52836 13860 53788
rect 14028 53842 14084 55134
rect 14476 54180 14532 55356
rect 14588 55298 14644 55310
rect 14588 55246 14590 55298
rect 14642 55246 14644 55298
rect 14588 54404 14644 55246
rect 15372 55188 15428 55198
rect 15372 55186 15988 55188
rect 15372 55134 15374 55186
rect 15426 55134 15988 55186
rect 15372 55132 15988 55134
rect 15372 55122 15428 55132
rect 14588 54338 14644 54348
rect 14476 54124 14756 54180
rect 14028 53790 14030 53842
rect 14082 53790 14084 53842
rect 14028 53778 14084 53790
rect 14700 53730 14756 54124
rect 15932 53956 15988 55132
rect 16044 54402 16100 56030
rect 16940 56082 16996 56094
rect 16940 56030 16942 56082
rect 16994 56030 16996 56082
rect 16044 54350 16046 54402
rect 16098 54350 16100 54402
rect 16044 54338 16100 54350
rect 16492 54404 16548 54414
rect 16492 54310 16548 54348
rect 16940 54404 16996 56030
rect 17724 55972 17780 55982
rect 17724 55878 17780 55916
rect 16940 54338 16996 54348
rect 17500 55410 17556 55422
rect 17500 55358 17502 55410
rect 17554 55358 17556 55410
rect 16044 53956 16100 53966
rect 15932 53954 16100 53956
rect 15932 53902 16046 53954
rect 16098 53902 16100 53954
rect 15932 53900 16100 53902
rect 16044 53890 16100 53900
rect 16044 53732 16100 53742
rect 14700 53678 14702 53730
rect 14754 53678 14756 53730
rect 14700 53666 14756 53678
rect 15820 53730 16100 53732
rect 15820 53678 16046 53730
rect 16098 53678 16100 53730
rect 15820 53676 16100 53678
rect 17500 53732 17556 55358
rect 17948 55300 18004 55310
rect 17948 55298 18116 55300
rect 17948 55246 17950 55298
rect 18002 55246 18116 55298
rect 17948 55244 18116 55246
rect 17948 55234 18004 55244
rect 18060 54516 18116 55244
rect 17724 54404 17780 54414
rect 17724 54310 17780 54348
rect 17948 53732 18004 53742
rect 17500 53730 18004 53732
rect 17500 53678 17950 53730
rect 18002 53678 18004 53730
rect 17500 53676 18004 53678
rect 14140 53620 14196 53630
rect 9996 50430 9998 50482
rect 10050 50430 10052 50482
rect 9996 50418 10052 50430
rect 10332 51380 10388 51390
rect 8764 49250 8932 49252
rect 8764 49198 8766 49250
rect 8818 49198 8932 49250
rect 8764 49196 8932 49198
rect 8764 49186 8820 49196
rect 9100 49028 9156 49038
rect 9100 49026 9268 49028
rect 9100 48974 9102 49026
rect 9154 48974 9268 49026
rect 9100 48972 9268 48974
rect 9100 48962 9156 48972
rect 7420 48802 7924 48804
rect 7420 48750 7534 48802
rect 7586 48750 7924 48802
rect 7420 48748 7924 48750
rect 8428 48802 8484 48814
rect 8428 48750 8430 48802
rect 8482 48750 8484 48802
rect 6524 48130 6580 48142
rect 6524 48078 6526 48130
rect 6578 48078 6580 48130
rect 6524 47012 6580 48078
rect 7084 47460 7140 47470
rect 7084 47366 7140 47404
rect 7308 47348 7364 47358
rect 7308 47254 7364 47292
rect 6524 46946 6580 46956
rect 6860 47234 6916 47246
rect 6860 47182 6862 47234
rect 6914 47182 6916 47234
rect 5068 46898 6356 46900
rect 5068 46846 5070 46898
rect 5122 46846 6356 46898
rect 5068 46844 6356 46846
rect 5068 46834 5124 46844
rect 4900 46620 5012 46676
rect 4844 46610 4900 46620
rect 4732 46452 4788 46462
rect 4284 46450 4788 46452
rect 4284 46398 4734 46450
rect 4786 46398 4788 46450
rect 4284 46396 4788 46398
rect 4732 46386 4788 46396
rect 4476 46284 4740 46294
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4476 46218 4740 46228
rect 6860 46116 6916 47182
rect 7196 47234 7252 47246
rect 7196 47182 7198 47234
rect 7250 47182 7252 47234
rect 7196 46788 7252 47182
rect 7308 46788 7364 46798
rect 7196 46786 7364 46788
rect 7196 46734 7310 46786
rect 7362 46734 7364 46786
rect 7196 46732 7364 46734
rect 7308 46722 7364 46732
rect 6860 46060 7252 46116
rect 4396 45892 4452 45902
rect 6524 45892 6580 45902
rect 6972 45892 7028 45902
rect 4172 45836 4340 45892
rect 3612 45780 3668 45790
rect 3612 45686 3668 45724
rect 4060 45778 4116 45790
rect 4060 45726 4062 45778
rect 4114 45726 4116 45778
rect 3500 45666 3556 45678
rect 3500 45614 3502 45666
rect 3554 45614 3556 45666
rect 3500 44996 3556 45614
rect 3724 45668 3780 45678
rect 4060 45668 4116 45726
rect 3724 45666 4116 45668
rect 3724 45614 3726 45666
rect 3778 45614 4116 45666
rect 3724 45612 4116 45614
rect 3724 45602 3780 45612
rect 3836 45332 3892 45342
rect 3836 45238 3892 45276
rect 3724 45220 3780 45230
rect 3724 45126 3780 45164
rect 3500 44930 3556 44940
rect 3836 45108 3892 45118
rect 3948 45108 4004 45118
rect 3892 45106 4004 45108
rect 3892 45054 3950 45106
rect 4002 45054 4004 45106
rect 3892 45052 4004 45054
rect 3388 44706 3444 44716
rect 2492 44382 2494 44434
rect 2546 44382 2548 44434
rect 2492 44370 2548 44382
rect 2044 43652 2212 43708
rect 1820 41878 1876 41916
rect 1708 40516 1764 40526
rect 1708 38724 1764 40460
rect 1708 38722 2100 38724
rect 1708 38670 1710 38722
rect 1762 38670 2100 38722
rect 1708 38668 2100 38670
rect 1708 38658 1764 38668
rect 2044 37938 2100 38668
rect 2044 37886 2046 37938
rect 2098 37886 2100 37938
rect 2044 37874 2100 37886
rect 1820 36708 1876 36718
rect 1820 36482 1876 36652
rect 1820 36430 1822 36482
rect 1874 36430 1876 36482
rect 1820 36418 1876 36430
rect 1708 33684 1764 33694
rect 1708 32450 1764 33628
rect 1708 32398 1710 32450
rect 1762 32398 1764 32450
rect 1708 31948 1764 32398
rect 1708 31892 2100 31948
rect 2044 31666 2100 31892
rect 2044 31614 2046 31666
rect 2098 31614 2100 31666
rect 2044 31602 2100 31614
rect 1820 30996 1876 31006
rect 1820 30210 1876 30940
rect 1820 30158 1822 30210
rect 1874 30158 1876 30210
rect 1820 30146 1876 30158
rect 1708 29876 1764 29886
rect 1708 29652 1764 29820
rect 1708 29650 1876 29652
rect 1708 29598 1710 29650
rect 1762 29598 1876 29650
rect 1708 29596 1876 29598
rect 1708 29586 1764 29596
rect 1820 28754 1876 29596
rect 1820 28702 1822 28754
rect 1874 28702 1876 28754
rect 1820 28690 1876 28702
rect 2156 22148 2212 43652
rect 3836 43650 3892 45052
rect 3948 45042 4004 45052
rect 4060 44884 4116 45612
rect 4060 44818 4116 44828
rect 4172 45666 4228 45678
rect 4172 45614 4174 45666
rect 4226 45614 4228 45666
rect 4172 44996 4228 45614
rect 4284 45668 4340 45836
rect 4396 45890 4788 45892
rect 4396 45838 4398 45890
rect 4450 45838 4788 45890
rect 4396 45836 4788 45838
rect 4396 45826 4452 45836
rect 4732 45778 4788 45836
rect 6524 45890 7028 45892
rect 6524 45838 6526 45890
rect 6578 45838 6974 45890
rect 7026 45838 7028 45890
rect 6524 45836 7028 45838
rect 6524 45826 6580 45836
rect 6972 45826 7028 45836
rect 4732 45726 4734 45778
rect 4786 45726 4788 45778
rect 4732 45714 4788 45726
rect 4844 45780 4900 45790
rect 4844 45686 4900 45724
rect 5964 45778 6020 45790
rect 5964 45726 5966 45778
rect 6018 45726 6020 45778
rect 4508 45668 4564 45678
rect 4284 45666 4564 45668
rect 4284 45614 4510 45666
rect 4562 45614 4564 45666
rect 4284 45612 4564 45614
rect 4508 45602 4564 45612
rect 5964 45668 6020 45726
rect 6300 45780 6356 45790
rect 6300 45686 6356 45724
rect 7084 45780 7140 45790
rect 5964 45602 6020 45612
rect 6076 45666 6132 45678
rect 6076 45614 6078 45666
rect 6130 45614 6132 45666
rect 6076 45332 6132 45614
rect 5516 45276 6132 45332
rect 6412 45668 6468 45678
rect 5516 45218 5572 45276
rect 6412 45220 6468 45612
rect 6860 45668 6916 45678
rect 6860 45574 6916 45612
rect 7084 45666 7140 45724
rect 7084 45614 7086 45666
rect 7138 45614 7140 45666
rect 5516 45166 5518 45218
rect 5570 45166 5572 45218
rect 5516 45154 5572 45166
rect 6300 45164 6468 45220
rect 7084 45220 7140 45614
rect 7196 45668 7252 46060
rect 7308 45668 7364 45678
rect 7196 45666 7364 45668
rect 7196 45614 7310 45666
rect 7362 45614 7364 45666
rect 7196 45612 7364 45614
rect 4396 45106 4452 45118
rect 4396 45054 4398 45106
rect 4450 45054 4452 45106
rect 4396 44996 4452 45054
rect 4844 45108 4900 45118
rect 4844 45014 4900 45052
rect 4172 44436 4228 44940
rect 4284 44940 4396 44996
rect 4284 44772 4340 44940
rect 4396 44930 4452 44940
rect 5740 44996 5796 45006
rect 4284 44706 4340 44716
rect 4476 44716 4740 44726
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4476 44650 4740 44660
rect 4620 44436 4676 44446
rect 4172 44434 4676 44436
rect 4172 44382 4622 44434
rect 4674 44382 4676 44434
rect 4172 44380 4676 44382
rect 4620 44370 4676 44380
rect 5068 44098 5124 44110
rect 5068 44046 5070 44098
rect 5122 44046 5124 44098
rect 3836 43598 3838 43650
rect 3890 43598 3892 43650
rect 3836 43586 3892 43598
rect 4284 43652 4340 43662
rect 4284 43538 4340 43596
rect 4284 43486 4286 43538
rect 4338 43486 4340 43538
rect 3500 43428 3556 43438
rect 3500 42980 3556 43372
rect 3276 42924 3556 42980
rect 2828 42642 2884 42654
rect 2828 42590 2830 42642
rect 2882 42590 2884 42642
rect 2604 42530 2660 42542
rect 2604 42478 2606 42530
rect 2658 42478 2660 42530
rect 2604 42420 2660 42478
rect 2828 42532 2884 42590
rect 3164 42644 3220 42654
rect 3164 42550 3220 42588
rect 2828 42466 2884 42476
rect 2940 42530 2996 42542
rect 2940 42478 2942 42530
rect 2994 42478 2996 42530
rect 2604 42354 2660 42364
rect 2940 42196 2996 42478
rect 2492 42140 2996 42196
rect 3052 42532 3108 42542
rect 2492 42082 2548 42140
rect 2492 42030 2494 42082
rect 2546 42030 2548 42082
rect 2492 42018 2548 42030
rect 3052 41298 3108 42476
rect 3276 42420 3332 42924
rect 4172 42868 4228 42878
rect 3388 42756 3444 42766
rect 3836 42756 3892 42766
rect 3388 42754 3892 42756
rect 3388 42702 3390 42754
rect 3442 42702 3838 42754
rect 3890 42702 3892 42754
rect 3388 42700 3892 42702
rect 3388 42690 3444 42700
rect 3836 42690 3892 42700
rect 3724 42532 3780 42542
rect 3724 42438 3780 42476
rect 3948 42532 4004 42542
rect 4172 42532 4228 42812
rect 3276 42364 3444 42420
rect 3052 41246 3054 41298
rect 3106 41246 3108 41298
rect 3052 41234 3108 41246
rect 3388 41298 3444 42364
rect 3388 41246 3390 41298
rect 3442 41246 3444 41298
rect 3388 41234 3444 41246
rect 3500 42084 3556 42094
rect 3500 41186 3556 42028
rect 3500 41134 3502 41186
rect 3554 41134 3556 41186
rect 3500 41122 3556 41134
rect 3164 40516 3220 40526
rect 3052 40460 3164 40516
rect 2828 40404 2884 40414
rect 2828 39844 2884 40348
rect 2604 39842 2884 39844
rect 2604 39790 2830 39842
rect 2882 39790 2884 39842
rect 2604 39788 2884 39790
rect 2604 38050 2660 39788
rect 2828 39778 2884 39788
rect 3052 39506 3108 40460
rect 3164 40450 3220 40460
rect 3948 39842 4004 42476
rect 3948 39790 3950 39842
rect 4002 39790 4004 39842
rect 3948 39778 4004 39790
rect 4060 42530 4228 42532
rect 4060 42478 4174 42530
rect 4226 42478 4228 42530
rect 4060 42476 4228 42478
rect 4060 42420 4116 42476
rect 4172 42466 4228 42476
rect 3164 39732 3220 39742
rect 3164 39730 3668 39732
rect 3164 39678 3166 39730
rect 3218 39678 3668 39730
rect 3164 39676 3668 39678
rect 3164 39666 3220 39676
rect 3612 39618 3668 39676
rect 3836 39620 3892 39630
rect 3612 39566 3614 39618
rect 3666 39566 3668 39618
rect 3612 39554 3668 39566
rect 3724 39618 3892 39620
rect 3724 39566 3838 39618
rect 3890 39566 3892 39618
rect 3724 39564 3892 39566
rect 3052 39454 3054 39506
rect 3106 39454 3108 39506
rect 3052 39442 3108 39454
rect 3724 38668 3780 39564
rect 3836 39554 3892 39564
rect 2604 37998 2606 38050
rect 2658 37998 2660 38050
rect 2604 37986 2660 37998
rect 3500 38612 3780 38668
rect 3836 38724 3892 38762
rect 3836 38658 3892 38668
rect 3500 38050 3556 38612
rect 4060 38388 4116 42364
rect 4284 42084 4340 43486
rect 4956 43538 5012 43550
rect 4956 43486 4958 43538
rect 5010 43486 5012 43538
rect 4396 43428 4452 43438
rect 4396 43334 4452 43372
rect 4476 43148 4740 43158
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4476 43082 4740 43092
rect 4732 42980 4788 42990
rect 4956 42980 5012 43486
rect 4732 42978 5012 42980
rect 4732 42926 4734 42978
rect 4786 42926 5012 42978
rect 4732 42924 5012 42926
rect 4732 42914 4788 42924
rect 4844 42756 4900 42766
rect 4844 42662 4900 42700
rect 4732 42532 4788 42542
rect 4732 42438 4788 42476
rect 4284 41972 4340 42028
rect 5068 41972 5124 44046
rect 5740 44100 5796 44940
rect 6300 44434 6356 45164
rect 7084 45154 7140 45164
rect 6300 44382 6302 44434
rect 6354 44382 6356 44434
rect 6300 44370 6356 44382
rect 6748 44434 6804 44446
rect 6748 44382 6750 44434
rect 6802 44382 6804 44434
rect 6748 44100 6804 44382
rect 6860 44324 6916 44334
rect 6860 44230 6916 44268
rect 5740 44098 5908 44100
rect 5740 44046 5742 44098
rect 5794 44046 5908 44098
rect 5740 44044 5908 44046
rect 5740 44034 5796 44044
rect 5404 43652 5460 43662
rect 5404 43558 5460 43596
rect 5180 43538 5236 43550
rect 5180 43486 5182 43538
rect 5234 43486 5236 43538
rect 5180 42756 5236 43486
rect 5516 43538 5572 43550
rect 5516 43486 5518 43538
rect 5570 43486 5572 43538
rect 5516 43428 5572 43486
rect 5516 42980 5572 43372
rect 5516 42914 5572 42924
rect 5180 42690 5236 42700
rect 5740 42754 5796 42766
rect 5740 42702 5742 42754
rect 5794 42702 5796 42754
rect 5740 42644 5796 42702
rect 5740 42578 5796 42588
rect 5404 41972 5460 41982
rect 4172 41916 4340 41972
rect 4956 41916 5404 41972
rect 4172 40964 4228 41916
rect 4620 41860 4676 41870
rect 4284 41858 4676 41860
rect 4284 41806 4622 41858
rect 4674 41806 4676 41858
rect 4284 41804 4676 41806
rect 4284 41188 4340 41804
rect 4620 41794 4676 41804
rect 4476 41580 4740 41590
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4476 41514 4740 41524
rect 4956 41298 5012 41916
rect 4956 41246 4958 41298
rect 5010 41246 5012 41298
rect 4956 41234 5012 41246
rect 4508 41188 4564 41198
rect 4284 41186 4564 41188
rect 4284 41134 4510 41186
rect 4562 41134 4564 41186
rect 4284 41132 4564 41134
rect 4508 41122 4564 41132
rect 4396 40964 4452 40974
rect 4172 40962 4452 40964
rect 4172 40910 4398 40962
rect 4450 40910 4452 40962
rect 4172 40908 4452 40910
rect 4396 40898 4452 40908
rect 4172 40628 4228 40638
rect 4172 39732 4228 40572
rect 4508 40516 4564 40526
rect 4732 40516 4788 40526
rect 4508 40422 4564 40460
rect 4620 40460 4732 40516
rect 4284 40402 4340 40414
rect 4284 40350 4286 40402
rect 4338 40350 4340 40402
rect 4284 39844 4340 40350
rect 4620 40402 4676 40460
rect 4732 40450 4788 40460
rect 4620 40350 4622 40402
rect 4674 40350 4676 40402
rect 4620 40338 4676 40350
rect 4476 40012 4740 40022
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4476 39946 4740 39956
rect 4284 39788 4564 39844
rect 4172 39676 4340 39732
rect 3500 37998 3502 38050
rect 3554 37998 3556 38050
rect 2828 37378 2884 37390
rect 2828 37326 2830 37378
rect 2882 37326 2884 37378
rect 2828 37268 2884 37326
rect 2940 37380 2996 37390
rect 2940 37286 2996 37324
rect 3388 37378 3444 37390
rect 3388 37326 3390 37378
rect 3442 37326 3444 37378
rect 2828 37202 2884 37212
rect 2828 37044 2884 37054
rect 2828 37042 3108 37044
rect 2828 36990 2830 37042
rect 2882 36990 3108 37042
rect 2828 36988 3108 36990
rect 2828 36978 2884 36988
rect 2492 36372 2548 36382
rect 2492 36370 2884 36372
rect 2492 36318 2494 36370
rect 2546 36318 2884 36370
rect 2492 36316 2884 36318
rect 2492 36306 2548 36316
rect 2268 35588 2324 35598
rect 2268 35586 2660 35588
rect 2268 35534 2270 35586
rect 2322 35534 2660 35586
rect 2268 35532 2660 35534
rect 2268 35522 2324 35532
rect 2604 35138 2660 35532
rect 2604 35086 2606 35138
rect 2658 35086 2660 35138
rect 2604 35074 2660 35086
rect 2828 35026 2884 36316
rect 2940 35698 2996 35710
rect 2940 35646 2942 35698
rect 2994 35646 2996 35698
rect 2940 35364 2996 35646
rect 3052 35586 3108 36988
rect 3052 35534 3054 35586
rect 3106 35534 3108 35586
rect 3052 35522 3108 35534
rect 3388 35364 3444 37326
rect 3500 37154 3556 37998
rect 3836 38332 4116 38388
rect 4172 38612 4228 38622
rect 3500 37102 3502 37154
rect 3554 37102 3556 37154
rect 3500 37090 3556 37102
rect 3724 37268 3780 37278
rect 3724 35922 3780 37212
rect 3724 35870 3726 35922
rect 3778 35870 3780 35922
rect 3724 35858 3780 35870
rect 2940 35308 3444 35364
rect 2828 34974 2830 35026
rect 2882 34974 2884 35026
rect 2828 34962 2884 34974
rect 2940 34914 2996 34926
rect 2940 34862 2942 34914
rect 2994 34862 2996 34914
rect 2380 34690 2436 34702
rect 2380 34638 2382 34690
rect 2434 34638 2436 34690
rect 2380 34580 2436 34638
rect 2380 34514 2436 34524
rect 2492 34692 2548 34702
rect 2492 33684 2548 34636
rect 2940 34580 2996 34862
rect 2940 34514 2996 34524
rect 3276 34690 3332 34702
rect 3276 34638 3278 34690
rect 3330 34638 3332 34690
rect 2492 33234 2548 33628
rect 2716 34132 2772 34142
rect 2716 33570 2772 34076
rect 2716 33518 2718 33570
rect 2770 33518 2772 33570
rect 2716 33506 2772 33518
rect 2604 33460 2660 33470
rect 2604 33366 2660 33404
rect 3276 33346 3332 34638
rect 3388 34468 3444 35308
rect 3612 34804 3668 34814
rect 3500 34692 3556 34702
rect 3500 34598 3556 34636
rect 3388 34412 3556 34468
rect 3276 33294 3278 33346
rect 3330 33294 3332 33346
rect 3276 33282 3332 33294
rect 3388 34242 3444 34254
rect 3388 34190 3390 34242
rect 3442 34190 3444 34242
rect 2492 33182 2494 33234
rect 2546 33182 2548 33234
rect 2492 33170 2548 33182
rect 2604 33124 2660 33134
rect 2604 31778 2660 33068
rect 3388 33124 3444 34190
rect 3500 33570 3556 34412
rect 3612 34132 3668 34748
rect 3612 34038 3668 34076
rect 3500 33518 3502 33570
rect 3554 33518 3556 33570
rect 3500 33506 3556 33518
rect 3612 33460 3668 33470
rect 3612 33366 3668 33404
rect 3724 33346 3780 33358
rect 3724 33294 3726 33346
rect 3778 33294 3780 33346
rect 3388 33058 3444 33068
rect 3612 33236 3668 33246
rect 2604 31726 2606 31778
rect 2658 31726 2660 31778
rect 2604 31714 2660 31726
rect 3612 31554 3668 33180
rect 3724 31780 3780 33294
rect 3836 32788 3892 38332
rect 3948 38164 4004 38174
rect 4172 38164 4228 38556
rect 3948 38162 4228 38164
rect 3948 38110 3950 38162
rect 4002 38110 4228 38162
rect 3948 38108 4228 38110
rect 3948 38098 4004 38108
rect 4284 38052 4340 39676
rect 4508 39618 4564 39788
rect 4508 39566 4510 39618
rect 4562 39566 4564 39618
rect 4508 39554 4564 39566
rect 4844 39620 4900 39630
rect 4620 38836 4676 38846
rect 4844 38836 4900 39564
rect 4620 38834 4900 38836
rect 4620 38782 4622 38834
rect 4674 38782 4900 38834
rect 4620 38780 4900 38782
rect 4620 38770 4676 38780
rect 4476 38444 4740 38454
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4476 38378 4740 38388
rect 4508 38052 4564 38062
rect 4060 38050 4564 38052
rect 4060 37998 4510 38050
rect 4562 37998 4564 38050
rect 4060 37996 4564 37998
rect 3948 36708 4004 36718
rect 3948 34132 4004 36652
rect 4060 35698 4116 37996
rect 4508 37986 4564 37996
rect 4172 37826 4228 37838
rect 4396 37828 4452 37838
rect 4172 37774 4174 37826
rect 4226 37774 4228 37826
rect 4172 37380 4228 37774
rect 4172 37044 4228 37324
rect 4172 36978 4228 36988
rect 4284 37826 4452 37828
rect 4284 37774 4398 37826
rect 4450 37774 4452 37826
rect 4284 37772 4452 37774
rect 4844 37828 4900 38780
rect 5180 39172 5236 39182
rect 5068 38724 5124 38762
rect 5068 38658 5124 38668
rect 4956 38612 5012 38622
rect 4956 38518 5012 38556
rect 4956 37828 5012 37838
rect 4844 37826 5012 37828
rect 4844 37774 4958 37826
rect 5010 37774 5012 37826
rect 4844 37772 5012 37774
rect 4284 36596 4340 37772
rect 4396 37762 4452 37772
rect 4396 37268 4452 37278
rect 4956 37268 5012 37772
rect 5180 37492 5236 39116
rect 5292 38834 5348 38846
rect 5292 38782 5294 38834
rect 5346 38782 5348 38834
rect 5292 38612 5348 38782
rect 5404 38668 5460 41916
rect 5740 40292 5796 40302
rect 5740 39620 5796 40236
rect 5740 39526 5796 39564
rect 5740 38722 5796 38734
rect 5740 38670 5742 38722
rect 5794 38670 5796 38722
rect 5404 38612 5572 38668
rect 5292 38546 5348 38556
rect 5516 38388 5572 38612
rect 5404 38332 5572 38388
rect 5740 38612 5796 38670
rect 5180 37436 5348 37492
rect 5180 37268 5236 37278
rect 4396 37266 4900 37268
rect 4396 37214 4398 37266
rect 4450 37214 4900 37266
rect 4396 37212 4900 37214
rect 4956 37212 5180 37268
rect 4396 37202 4452 37212
rect 4476 36876 4740 36886
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4476 36810 4740 36820
rect 4844 36708 4900 37212
rect 5180 37174 5236 37212
rect 5068 37044 5124 37054
rect 4956 36708 5012 36718
rect 4844 36706 5012 36708
rect 4844 36654 4958 36706
rect 5010 36654 5012 36706
rect 4844 36652 5012 36654
rect 4956 36642 5012 36652
rect 4620 36596 4676 36606
rect 4284 36594 4676 36596
rect 4284 36542 4622 36594
rect 4674 36542 4676 36594
rect 4284 36540 4676 36542
rect 4060 35646 4062 35698
rect 4114 35646 4116 35698
rect 4060 35634 4116 35646
rect 4172 35924 4228 35934
rect 4172 34802 4228 35868
rect 4284 35810 4340 36540
rect 4620 36530 4676 36540
rect 5068 36594 5124 36988
rect 5068 36542 5070 36594
rect 5122 36542 5124 36594
rect 5068 36530 5124 36542
rect 5292 36260 5348 37436
rect 5404 36708 5460 38332
rect 5740 37716 5796 38556
rect 5404 36642 5460 36652
rect 5516 37660 5796 37716
rect 5516 36596 5572 37660
rect 5852 37604 5908 44044
rect 6748 44034 6804 44044
rect 5964 42754 6020 42766
rect 5964 42702 5966 42754
rect 6018 42702 6020 42754
rect 5964 42084 6020 42702
rect 6300 42754 6356 42766
rect 6300 42702 6302 42754
rect 6354 42702 6356 42754
rect 5964 42018 6020 42028
rect 6076 42530 6132 42542
rect 6076 42478 6078 42530
rect 6130 42478 6132 42530
rect 6076 42082 6132 42478
rect 6300 42532 6356 42702
rect 7196 42756 7252 42766
rect 7308 42756 7364 45612
rect 7196 42754 7364 42756
rect 7196 42702 7198 42754
rect 7250 42702 7364 42754
rect 7196 42700 7364 42702
rect 6636 42644 6692 42654
rect 6636 42550 6692 42588
rect 6524 42532 6580 42542
rect 6300 42530 6580 42532
rect 6300 42478 6526 42530
rect 6578 42478 6580 42530
rect 6300 42476 6580 42478
rect 6076 42030 6078 42082
rect 6130 42030 6132 42082
rect 6076 42018 6132 42030
rect 6524 41300 6580 42476
rect 6748 42530 6804 42542
rect 6748 42478 6750 42530
rect 6802 42478 6804 42530
rect 6748 42084 6804 42478
rect 6748 42018 6804 42028
rect 6972 41300 7028 41310
rect 6524 41298 7028 41300
rect 6524 41246 6974 41298
rect 7026 41246 7028 41298
rect 6524 41244 7028 41246
rect 6972 41234 7028 41244
rect 6412 39506 6468 39518
rect 6412 39454 6414 39506
rect 6466 39454 6468 39506
rect 6300 39172 6356 39182
rect 6300 39058 6356 39116
rect 6300 39006 6302 39058
rect 6354 39006 6356 39058
rect 6300 38994 6356 39006
rect 6412 39058 6468 39454
rect 6412 39006 6414 39058
rect 6466 39006 6468 39058
rect 6412 38994 6468 39006
rect 6524 39396 6580 39406
rect 6524 38946 6580 39340
rect 6972 39172 7028 39182
rect 6972 39058 7028 39116
rect 6972 39006 6974 39058
rect 7026 39006 7028 39058
rect 6972 38994 7028 39006
rect 6524 38894 6526 38946
rect 6578 38894 6580 38946
rect 6524 38882 6580 38894
rect 7196 38500 7252 42700
rect 7308 41300 7364 41310
rect 7308 41206 7364 41244
rect 7420 41076 7476 48748
rect 7532 48738 7588 48748
rect 8428 48692 8484 48750
rect 8428 48626 8484 48636
rect 8652 48356 8708 48366
rect 8652 48132 8708 48300
rect 8316 48130 8708 48132
rect 8316 48078 8654 48130
rect 8706 48078 8708 48130
rect 8316 48076 8708 48078
rect 7532 47460 7588 47470
rect 7532 46786 7588 47404
rect 8316 47458 8372 48076
rect 8652 48066 8708 48076
rect 9100 48356 9156 48366
rect 8540 47572 8596 47582
rect 8540 47478 8596 47516
rect 8316 47406 8318 47458
rect 8370 47406 8372 47458
rect 8316 47394 8372 47406
rect 8876 47460 8932 47470
rect 9100 47460 9156 48300
rect 9212 48132 9268 48972
rect 9324 49026 9380 49038
rect 9324 48974 9326 49026
rect 9378 48974 9380 49026
rect 9324 48468 9380 48974
rect 9772 49028 9828 49038
rect 9772 49026 9940 49028
rect 9772 48974 9774 49026
rect 9826 48974 9940 49026
rect 9772 48972 9940 48974
rect 9772 48962 9828 48972
rect 9884 48804 9940 48972
rect 9436 48468 9492 48478
rect 9324 48466 9492 48468
rect 9324 48414 9438 48466
rect 9490 48414 9492 48466
rect 9324 48412 9492 48414
rect 9436 48402 9492 48412
rect 9660 48356 9716 48366
rect 9660 48262 9716 48300
rect 9772 48242 9828 48254
rect 9772 48190 9774 48242
rect 9826 48190 9828 48242
rect 9212 48076 9492 48132
rect 9436 47570 9492 48076
rect 9436 47518 9438 47570
rect 9490 47518 9492 47570
rect 9436 47506 9492 47518
rect 9548 47572 9604 47582
rect 9772 47572 9828 48190
rect 9604 47516 9828 47572
rect 9324 47460 9380 47470
rect 9100 47458 9380 47460
rect 9100 47406 9326 47458
rect 9378 47406 9380 47458
rect 9100 47404 9380 47406
rect 8876 47366 8932 47404
rect 9324 47394 9380 47404
rect 9548 47458 9604 47516
rect 9548 47406 9550 47458
rect 9602 47406 9604 47458
rect 9548 47394 9604 47406
rect 7644 47348 7700 47358
rect 7700 47292 7924 47348
rect 7644 47254 7700 47292
rect 7756 47012 7812 47022
rect 7756 46898 7812 46956
rect 7756 46846 7758 46898
rect 7810 46846 7812 46898
rect 7756 46834 7812 46846
rect 7532 46734 7534 46786
rect 7586 46734 7588 46786
rect 7532 45892 7588 46734
rect 7868 46786 7924 47292
rect 9772 47124 9828 47516
rect 9772 47058 9828 47068
rect 7868 46734 7870 46786
rect 7922 46734 7924 46786
rect 7868 46722 7924 46734
rect 9772 46564 9828 46574
rect 9884 46564 9940 48748
rect 9996 48916 10052 48926
rect 9996 48804 10052 48860
rect 9996 48802 10164 48804
rect 9996 48750 9998 48802
rect 10050 48750 10164 48802
rect 9996 48748 10164 48750
rect 9996 48738 10052 48748
rect 10108 48354 10164 48748
rect 10108 48302 10110 48354
rect 10162 48302 10164 48354
rect 10108 48290 10164 48302
rect 10332 48244 10388 51324
rect 10780 50706 10836 50718
rect 10780 50654 10782 50706
rect 10834 50654 10836 50706
rect 10668 49700 10724 49710
rect 10780 49700 10836 50654
rect 11004 50482 11060 51436
rect 12124 51492 12180 51502
rect 12124 51398 12180 51436
rect 11116 51378 11172 51390
rect 11116 51326 11118 51378
rect 11170 51326 11172 51378
rect 11116 50596 11172 51326
rect 11116 50530 11172 50540
rect 12348 51378 12404 51390
rect 12348 51326 12350 51378
rect 12402 51326 12404 51378
rect 11004 50430 11006 50482
rect 11058 50430 11060 50482
rect 11004 50418 11060 50430
rect 12348 50428 12404 51326
rect 12908 51380 12964 51390
rect 12908 50706 12964 51324
rect 13692 51378 13748 51390
rect 13692 51326 13694 51378
rect 13746 51326 13748 51378
rect 12908 50654 12910 50706
rect 12962 50654 12964 50706
rect 12908 50642 12964 50654
rect 13356 51268 13412 51278
rect 13692 51268 13748 51326
rect 13356 51266 13748 51268
rect 13356 51214 13358 51266
rect 13410 51214 13748 51266
rect 13356 51212 13748 51214
rect 10892 50372 10948 50382
rect 10892 50034 10948 50316
rect 10892 49982 10894 50034
rect 10946 49982 10948 50034
rect 10892 49970 10948 49982
rect 11564 50372 11620 50382
rect 11564 50034 11620 50316
rect 11900 50372 12404 50428
rect 12684 50482 12740 50494
rect 12684 50430 12686 50482
rect 12738 50430 12740 50482
rect 11788 50148 11844 50158
rect 11564 49982 11566 50034
rect 11618 49982 11620 50034
rect 11564 49970 11620 49982
rect 11676 50036 11732 50046
rect 11788 50036 11844 50092
rect 11676 50034 11844 50036
rect 11676 49982 11678 50034
rect 11730 49982 11844 50034
rect 11676 49980 11844 49982
rect 11676 49970 11732 49980
rect 11116 49810 11172 49822
rect 11788 49812 11844 49822
rect 11900 49812 11956 50372
rect 11116 49758 11118 49810
rect 11170 49758 11172 49810
rect 11116 49700 11172 49758
rect 10668 49698 11172 49700
rect 10668 49646 10670 49698
rect 10722 49646 11172 49698
rect 10668 49644 11172 49646
rect 10668 49634 10724 49644
rect 11116 48916 11172 49644
rect 11676 49810 11956 49812
rect 11676 49758 11790 49810
rect 11842 49758 11956 49810
rect 11676 49756 11956 49758
rect 12012 49922 12068 49934
rect 12012 49870 12014 49922
rect 12066 49870 12068 49922
rect 11116 48850 11172 48860
rect 11564 48916 11620 48926
rect 11564 48822 11620 48860
rect 10444 48804 10500 48814
rect 10444 48710 10500 48748
rect 11676 48804 11732 49756
rect 11788 49746 11844 49756
rect 11900 48804 11956 48814
rect 11676 48710 11732 48748
rect 11788 48802 11956 48804
rect 11788 48750 11902 48802
rect 11954 48750 11956 48802
rect 11788 48748 11956 48750
rect 11788 48580 11844 48748
rect 11900 48738 11956 48748
rect 11676 48524 11844 48580
rect 10668 48466 10724 48478
rect 10668 48414 10670 48466
rect 10722 48414 10724 48466
rect 10668 48356 10724 48414
rect 10668 48290 10724 48300
rect 11228 48356 11284 48366
rect 10332 48242 10612 48244
rect 10332 48190 10334 48242
rect 10386 48190 10612 48242
rect 10332 48188 10612 48190
rect 10332 48178 10388 48188
rect 10220 47348 10276 47358
rect 9772 46562 9884 46564
rect 9772 46510 9774 46562
rect 9826 46510 9884 46562
rect 9772 46508 9884 46510
rect 9772 46498 9828 46508
rect 7644 45892 7700 45902
rect 7532 45890 7700 45892
rect 7532 45838 7646 45890
rect 7698 45838 7700 45890
rect 7532 45836 7700 45838
rect 7644 45826 7700 45836
rect 7980 45780 8036 45790
rect 7980 45778 8148 45780
rect 7980 45726 7982 45778
rect 8034 45726 8148 45778
rect 7980 45724 8148 45726
rect 7980 45714 8036 45724
rect 7868 45666 7924 45678
rect 7868 45614 7870 45666
rect 7922 45614 7924 45666
rect 7644 44994 7700 45006
rect 7644 44942 7646 44994
rect 7698 44942 7700 44994
rect 7644 44324 7700 44942
rect 7756 44548 7812 44558
rect 7868 44548 7924 45614
rect 8092 45330 8148 45724
rect 8092 45278 8094 45330
rect 8146 45278 8148 45330
rect 8092 45266 8148 45278
rect 8316 45220 8372 45230
rect 8428 45220 8484 45230
rect 8372 45218 8484 45220
rect 8372 45166 8430 45218
rect 8482 45166 8484 45218
rect 8372 45164 8484 45166
rect 7756 44546 7924 44548
rect 7756 44494 7758 44546
rect 7810 44494 7924 44546
rect 7756 44492 7924 44494
rect 7980 45106 8036 45118
rect 8204 45108 8260 45118
rect 7980 45054 7982 45106
rect 8034 45054 8036 45106
rect 7756 44482 7812 44492
rect 7700 44268 7812 44324
rect 7644 44258 7700 44268
rect 7756 44210 7812 44268
rect 7644 44154 7700 44166
rect 7644 44102 7646 44154
rect 7698 44102 7700 44154
rect 7644 44100 7700 44102
rect 7644 44034 7700 44044
rect 7756 44158 7758 44210
rect 7810 44158 7812 44210
rect 7756 43876 7812 44158
rect 7980 44100 8036 45054
rect 7980 44034 8036 44044
rect 8092 45106 8260 45108
rect 8092 45054 8206 45106
rect 8258 45054 8260 45106
rect 8092 45052 8260 45054
rect 8092 43876 8148 45052
rect 8204 45042 8260 45052
rect 7756 43820 8148 43876
rect 8092 43650 8148 43662
rect 8092 43598 8094 43650
rect 8146 43598 8148 43650
rect 7868 43540 7924 43550
rect 7756 43538 7924 43540
rect 7756 43486 7870 43538
rect 7922 43486 7924 43538
rect 7756 43484 7924 43486
rect 7756 42754 7812 43484
rect 7868 43474 7924 43484
rect 8092 42980 8148 43598
rect 8204 43540 8260 43550
rect 8204 43446 8260 43484
rect 8092 42924 8260 42980
rect 7756 42702 7758 42754
rect 7810 42702 7812 42754
rect 7756 42690 7812 42702
rect 8092 42754 8148 42766
rect 8092 42702 8094 42754
rect 8146 42702 8148 42754
rect 8092 41748 8148 42702
rect 8204 42084 8260 42924
rect 8316 42978 8372 45164
rect 8428 45154 8484 45164
rect 8988 45108 9044 45118
rect 8988 45014 9044 45052
rect 9548 44994 9604 45006
rect 9548 44942 9550 44994
rect 9602 44942 9604 44994
rect 8764 44884 8820 44894
rect 8764 44210 8820 44828
rect 8764 44158 8766 44210
rect 8818 44158 8820 44210
rect 8764 44146 8820 44158
rect 9100 44098 9156 44110
rect 9100 44046 9102 44098
rect 9154 44046 9156 44098
rect 8988 43540 9044 43550
rect 8316 42926 8318 42978
rect 8370 42926 8372 42978
rect 8316 42914 8372 42926
rect 8540 42980 8596 42990
rect 8204 42018 8260 42028
rect 8204 41860 8260 41870
rect 8204 41766 8260 41804
rect 7644 41188 7700 41198
rect 8092 41188 8148 41692
rect 7644 41186 8148 41188
rect 7644 41134 7646 41186
rect 7698 41134 8148 41186
rect 7644 41132 8148 41134
rect 8204 41412 8260 41422
rect 7644 41122 7700 41132
rect 7308 41020 7476 41076
rect 7308 39172 7364 41020
rect 8204 40628 8260 41356
rect 8540 41298 8596 42924
rect 8652 42756 8708 42766
rect 8652 42662 8708 42700
rect 8988 42754 9044 43484
rect 8988 42702 8990 42754
rect 9042 42702 9044 42754
rect 8988 42690 9044 42702
rect 9100 42532 9156 44046
rect 9548 44100 9604 44942
rect 9772 44884 9828 44894
rect 9772 44790 9828 44828
rect 9884 44660 9940 46508
rect 10108 47346 10276 47348
rect 10108 47294 10222 47346
rect 10274 47294 10276 47346
rect 10108 47292 10276 47294
rect 10108 46674 10164 47292
rect 10220 47282 10276 47292
rect 10556 47346 10612 48188
rect 11228 47458 11284 48300
rect 11676 48354 11732 48524
rect 12012 48466 12068 49870
rect 12236 48916 12292 48926
rect 12236 48822 12292 48860
rect 12012 48414 12014 48466
rect 12066 48414 12068 48466
rect 12012 48402 12068 48414
rect 12572 48468 12628 48478
rect 12684 48468 12740 50430
rect 13020 50036 13076 50046
rect 13356 50036 13412 51212
rect 13804 51156 13860 52780
rect 13916 53506 13972 53518
rect 13916 53454 13918 53506
rect 13970 53454 13972 53506
rect 13916 53396 13972 53454
rect 13916 52164 13972 53340
rect 14140 52834 14196 53564
rect 14924 53620 14980 53630
rect 14924 53526 14980 53564
rect 15036 53618 15092 53630
rect 15036 53566 15038 53618
rect 15090 53566 15092 53618
rect 14364 53508 14420 53518
rect 14364 53414 14420 53452
rect 15036 53396 15092 53566
rect 15596 53508 15652 53518
rect 15596 53414 15652 53452
rect 15036 53330 15092 53340
rect 15820 53170 15876 53676
rect 16044 53666 16100 53676
rect 17948 53666 18004 53676
rect 15820 53118 15822 53170
rect 15874 53118 15876 53170
rect 15820 53106 15876 53118
rect 16380 53618 16436 53630
rect 16380 53566 16382 53618
rect 16434 53566 16436 53618
rect 16380 53170 16436 53566
rect 16380 53118 16382 53170
rect 16434 53118 16436 53170
rect 16380 53106 16436 53118
rect 15372 52946 15428 52958
rect 15708 52948 15764 52958
rect 15372 52894 15374 52946
rect 15426 52894 15428 52946
rect 14140 52782 14142 52834
rect 14194 52782 14196 52834
rect 14140 52770 14196 52782
rect 14588 52836 14644 52846
rect 14588 52742 14644 52780
rect 15372 52500 15428 52894
rect 15372 52434 15428 52444
rect 15484 52892 15708 52948
rect 15484 52276 15540 52892
rect 15708 52854 15764 52892
rect 16044 52948 16100 52958
rect 16268 52948 16324 52958
rect 16044 52946 16324 52948
rect 16044 52894 16046 52946
rect 16098 52894 16270 52946
rect 16322 52894 16324 52946
rect 16044 52892 16324 52894
rect 16044 52882 16100 52892
rect 15148 52274 15540 52276
rect 15148 52222 15486 52274
rect 15538 52222 15540 52274
rect 15148 52220 15540 52222
rect 14028 52164 14084 52174
rect 15148 52164 15204 52220
rect 15484 52210 15540 52220
rect 16044 52500 16100 52510
rect 13916 52162 14532 52164
rect 13916 52110 14030 52162
rect 14082 52110 14532 52162
rect 13916 52108 14532 52110
rect 14028 52098 14084 52108
rect 14140 51938 14196 51950
rect 14140 51886 14142 51938
rect 14194 51886 14196 51938
rect 14140 51828 14196 51886
rect 14364 51940 14420 51950
rect 14364 51846 14420 51884
rect 14028 51772 14140 51828
rect 14028 51602 14084 51772
rect 14140 51762 14196 51772
rect 14028 51550 14030 51602
rect 14082 51550 14084 51602
rect 14028 51538 14084 51550
rect 13692 51100 13860 51156
rect 13580 50482 13636 50494
rect 13580 50430 13582 50482
rect 13634 50430 13636 50482
rect 13580 50428 13636 50430
rect 13076 49980 13412 50036
rect 13020 49942 13076 49980
rect 13356 49922 13412 49980
rect 13356 49870 13358 49922
rect 13410 49870 13412 49922
rect 13356 49858 13412 49870
rect 13468 50372 13636 50428
rect 13468 49700 13524 50372
rect 13356 49644 13524 49700
rect 13244 48916 13300 48926
rect 13356 48916 13412 49644
rect 13580 49588 13636 49598
rect 13300 48860 13412 48916
rect 13468 49532 13580 49588
rect 13020 48804 13076 48814
rect 12572 48466 12740 48468
rect 12572 48414 12574 48466
rect 12626 48414 12740 48466
rect 12572 48412 12740 48414
rect 12796 48692 12852 48702
rect 12572 48402 12628 48412
rect 11676 48302 11678 48354
rect 11730 48302 11732 48354
rect 11676 48290 11732 48302
rect 11788 48356 11844 48366
rect 11788 48262 11844 48300
rect 11900 48354 11956 48366
rect 11900 48302 11902 48354
rect 11954 48302 11956 48354
rect 11900 48244 11956 48302
rect 11676 47796 11732 47806
rect 11228 47406 11230 47458
rect 11282 47406 11284 47458
rect 11228 47394 11284 47406
rect 11564 47460 11620 47470
rect 11564 47366 11620 47404
rect 10556 47294 10558 47346
rect 10610 47294 10612 47346
rect 10556 47282 10612 47294
rect 11340 47234 11396 47246
rect 11340 47182 11342 47234
rect 11394 47182 11396 47234
rect 10332 47124 10388 47134
rect 10108 46622 10110 46674
rect 10162 46622 10164 46674
rect 10108 45220 10164 46622
rect 10220 46786 10276 46798
rect 10220 46734 10222 46786
rect 10274 46734 10276 46786
rect 10220 46564 10276 46734
rect 10220 46498 10276 46508
rect 10332 46002 10388 47068
rect 11340 47012 11396 47182
rect 10668 46956 11396 47012
rect 10444 46900 10500 46910
rect 10668 46900 10724 46956
rect 10444 46898 10724 46900
rect 10444 46846 10446 46898
rect 10498 46846 10724 46898
rect 10444 46844 10724 46846
rect 10444 46834 10500 46844
rect 10780 46788 10836 46798
rect 10780 46694 10836 46732
rect 11004 46788 11060 46798
rect 11004 46694 11060 46732
rect 11340 46786 11396 46956
rect 11676 46898 11732 47740
rect 11676 46846 11678 46898
rect 11730 46846 11732 46898
rect 11676 46834 11732 46846
rect 11340 46734 11342 46786
rect 11394 46734 11396 46786
rect 11340 46722 11396 46734
rect 11452 46788 11508 46798
rect 11452 46694 11508 46732
rect 10668 46676 10724 46686
rect 11900 46676 11956 48188
rect 12124 48244 12180 48254
rect 12460 48244 12516 48254
rect 12124 48242 12516 48244
rect 12124 48190 12126 48242
rect 12178 48190 12462 48242
rect 12514 48190 12516 48242
rect 12124 48188 12516 48190
rect 12124 47796 12180 48188
rect 12460 48178 12516 48188
rect 12684 48244 12740 48254
rect 12684 48150 12740 48188
rect 12124 47730 12180 47740
rect 12796 47682 12852 48636
rect 12908 48356 12964 48366
rect 12908 48262 12964 48300
rect 12796 47630 12798 47682
rect 12850 47630 12852 47682
rect 12796 47618 12852 47630
rect 12124 47570 12180 47582
rect 12124 47518 12126 47570
rect 12178 47518 12180 47570
rect 12124 47460 12180 47518
rect 12124 47394 12180 47404
rect 12460 47460 12516 47470
rect 12460 47458 12852 47460
rect 12460 47406 12462 47458
rect 12514 47406 12852 47458
rect 12460 47404 12852 47406
rect 12460 47394 12516 47404
rect 12236 46788 12292 46798
rect 12236 46694 12292 46732
rect 10668 46564 10724 46620
rect 11676 46620 11956 46676
rect 10668 46508 10948 46564
rect 10332 45950 10334 46002
rect 10386 45950 10388 46002
rect 10332 45938 10388 45950
rect 10108 45154 10164 45164
rect 10668 45892 10724 45902
rect 10108 44884 10164 44894
rect 10108 44882 10500 44884
rect 10108 44830 10110 44882
rect 10162 44830 10500 44882
rect 10108 44828 10500 44830
rect 10108 44818 10164 44828
rect 9548 44006 9604 44044
rect 9772 44604 9940 44660
rect 9324 43540 9380 43550
rect 9324 42756 9380 43484
rect 9324 42662 9380 42700
rect 8988 42476 9156 42532
rect 9212 42530 9268 42542
rect 9212 42478 9214 42530
rect 9266 42478 9268 42530
rect 8988 42196 9044 42476
rect 8988 42130 9044 42140
rect 9100 42308 9156 42318
rect 8652 41972 8708 41982
rect 8652 41878 8708 41916
rect 9100 41524 9156 42252
rect 9212 42084 9268 42478
rect 9548 42084 9604 42094
rect 9212 42082 9604 42084
rect 9212 42030 9550 42082
rect 9602 42030 9604 42082
rect 9212 42028 9604 42030
rect 9212 41748 9268 42028
rect 9548 42018 9604 42028
rect 9660 41970 9716 41982
rect 9660 41918 9662 41970
rect 9714 41918 9716 41970
rect 9660 41860 9716 41918
rect 9660 41794 9716 41804
rect 9212 41682 9268 41692
rect 9100 41468 9380 41524
rect 8540 41246 8542 41298
rect 8594 41246 8596 41298
rect 8540 41234 8596 41246
rect 8988 40964 9044 41002
rect 8988 40898 9044 40908
rect 7980 40572 8260 40628
rect 8316 40628 8372 40638
rect 8316 40626 8484 40628
rect 8316 40574 8318 40626
rect 8370 40574 8484 40626
rect 8316 40572 8484 40574
rect 7980 40516 8036 40572
rect 8316 40562 8372 40572
rect 7868 40404 7924 40414
rect 7868 40310 7924 40348
rect 7308 39106 7364 39116
rect 7420 39508 7476 39518
rect 7420 39058 7476 39452
rect 7420 39006 7422 39058
rect 7474 39006 7476 39058
rect 7420 38994 7476 39006
rect 7644 39284 7700 39294
rect 7644 38946 7700 39228
rect 7980 39058 8036 40460
rect 8204 40402 8260 40414
rect 8204 40350 8206 40402
rect 8258 40350 8260 40402
rect 8204 39284 8260 40350
rect 8428 40292 8484 40572
rect 8876 40516 8932 40526
rect 8428 40226 8484 40236
rect 8540 40514 8932 40516
rect 8540 40462 8878 40514
rect 8930 40462 8932 40514
rect 8540 40460 8932 40462
rect 8316 40180 8372 40190
rect 8316 40086 8372 40124
rect 8540 39956 8596 40460
rect 8876 40450 8932 40460
rect 8988 40516 9044 40526
rect 8204 39218 8260 39228
rect 8428 39900 8596 39956
rect 8652 40292 8708 40302
rect 7980 39006 7982 39058
rect 8034 39006 8036 39058
rect 7980 38994 8036 39006
rect 8316 39060 8372 39070
rect 8316 38966 8372 39004
rect 7644 38894 7646 38946
rect 7698 38894 7700 38946
rect 7644 38882 7700 38894
rect 8092 38836 8148 38846
rect 7532 38724 7588 38762
rect 7532 38658 7588 38668
rect 7196 38444 7700 38500
rect 5516 36530 5572 36540
rect 5628 37548 5908 37604
rect 5964 38220 6356 38276
rect 4732 36204 5348 36260
rect 4732 35924 4788 36204
rect 4732 35830 4788 35868
rect 4284 35758 4286 35810
rect 4338 35758 4340 35810
rect 4284 35746 4340 35758
rect 4396 35588 4452 35598
rect 4284 35532 4396 35588
rect 4284 35140 4340 35532
rect 4396 35522 4452 35532
rect 5516 35588 5572 35598
rect 5516 35494 5572 35532
rect 4476 35308 4740 35318
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4476 35242 4740 35252
rect 4396 35140 4452 35150
rect 4284 35138 4452 35140
rect 4284 35086 4398 35138
rect 4450 35086 4452 35138
rect 4284 35084 4452 35086
rect 4396 35074 4452 35084
rect 4956 34916 5012 34926
rect 4956 34822 5012 34860
rect 4172 34750 4174 34802
rect 4226 34750 4228 34802
rect 4172 34738 4228 34750
rect 5068 34802 5124 34814
rect 5068 34750 5070 34802
rect 5122 34750 5124 34802
rect 4284 34690 4340 34702
rect 4284 34638 4286 34690
rect 4338 34638 4340 34690
rect 4284 34356 4340 34638
rect 4844 34692 4900 34702
rect 4844 34598 4900 34636
rect 5068 34580 5124 34750
rect 5068 34514 5124 34524
rect 4284 34300 4900 34356
rect 4844 34242 4900 34300
rect 4844 34190 4846 34242
rect 4898 34190 4900 34242
rect 4844 34178 4900 34190
rect 4060 34132 4116 34142
rect 3948 34130 4116 34132
rect 3948 34078 4062 34130
rect 4114 34078 4116 34130
rect 3948 34076 4116 34078
rect 4060 32788 4116 34076
rect 4476 33740 4740 33750
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4476 33674 4740 33684
rect 5068 33684 5124 33694
rect 5068 33346 5124 33628
rect 5068 33294 5070 33346
rect 5122 33294 5124 33346
rect 5068 33282 5124 33294
rect 5628 33460 5684 37548
rect 5852 37380 5908 37390
rect 5964 37380 6020 38220
rect 6300 38164 6356 38220
rect 6412 38164 6468 38174
rect 6300 38162 6468 38164
rect 6300 38110 6414 38162
rect 6466 38110 6468 38162
rect 6300 38108 6468 38110
rect 6412 38098 6468 38108
rect 5852 37378 6020 37380
rect 5852 37326 5854 37378
rect 5906 37326 6020 37378
rect 5852 37324 6020 37326
rect 6188 38050 6244 38062
rect 6188 37998 6190 38050
rect 6242 37998 6244 38050
rect 6188 37828 6244 37998
rect 5852 37314 5908 37324
rect 5740 36708 5796 36718
rect 5740 36594 5796 36652
rect 5740 36542 5742 36594
rect 5794 36542 5796 36594
rect 5740 36530 5796 36542
rect 5852 36596 5908 36606
rect 5852 35812 5908 36540
rect 6188 36594 6244 37772
rect 6188 36542 6190 36594
rect 6242 36542 6244 36594
rect 6188 36530 6244 36542
rect 6524 38050 6580 38062
rect 6524 37998 6526 38050
rect 6578 37998 6580 38050
rect 6524 37940 6580 37998
rect 6860 38052 6916 38062
rect 7308 38052 7364 38062
rect 6860 38050 7364 38052
rect 6860 37998 6862 38050
rect 6914 37998 7310 38050
rect 7362 37998 7364 38050
rect 6860 37996 7364 37998
rect 6860 37986 6916 37996
rect 7308 37986 7364 37996
rect 4732 33236 4788 33246
rect 4732 33142 4788 33180
rect 4844 33122 4900 33134
rect 4844 33070 4846 33122
rect 4898 33070 4900 33122
rect 3836 32732 4004 32788
rect 3836 32564 3892 32574
rect 3836 32470 3892 32508
rect 3948 32004 4004 32732
rect 4060 32722 4116 32732
rect 4620 32788 4676 32798
rect 4620 32562 4676 32732
rect 4620 32510 4622 32562
rect 4674 32510 4676 32562
rect 4620 32498 4676 32510
rect 4732 32564 4788 32574
rect 4844 32564 4900 33070
rect 5068 32788 5124 32798
rect 5068 32694 5124 32732
rect 4788 32508 4900 32564
rect 4732 32498 4788 32508
rect 4956 32452 5012 32462
rect 4844 32396 4956 32452
rect 4476 32172 4740 32182
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4476 32106 4740 32116
rect 3948 31948 4340 32004
rect 4284 31892 4340 31948
rect 4172 31780 4228 31790
rect 3724 31778 4228 31780
rect 3724 31726 4174 31778
rect 4226 31726 4228 31778
rect 3724 31724 4228 31726
rect 3724 31666 3780 31724
rect 4172 31714 4228 31724
rect 3724 31614 3726 31666
rect 3778 31614 3780 31666
rect 3724 31602 3780 31614
rect 4284 31556 4340 31836
rect 4508 31666 4564 31678
rect 4508 31614 4510 31666
rect 4562 31614 4564 31666
rect 3612 31502 3614 31554
rect 3666 31502 3668 31554
rect 3612 31490 3668 31502
rect 3948 31500 4340 31556
rect 4396 31554 4452 31566
rect 4396 31502 4398 31554
rect 4450 31502 4452 31554
rect 3388 31220 3444 31230
rect 2940 31218 3444 31220
rect 2940 31166 3390 31218
rect 3442 31166 3444 31218
rect 2940 31164 3444 31166
rect 2716 31108 2772 31118
rect 2716 31014 2772 31052
rect 2940 31106 2996 31164
rect 3388 31154 3444 31164
rect 2940 31054 2942 31106
rect 2994 31054 2996 31106
rect 2940 31042 2996 31054
rect 3500 31108 3556 31118
rect 2380 30994 2436 31006
rect 2380 30942 2382 30994
rect 2434 30942 2436 30994
rect 2380 30884 2436 30942
rect 3276 30994 3332 31006
rect 3276 30942 3278 30994
rect 3330 30942 3332 30994
rect 2380 30818 2436 30828
rect 2492 30882 2548 30894
rect 2492 30830 2494 30882
rect 2546 30830 2548 30882
rect 2492 30322 2548 30830
rect 3276 30884 3332 30942
rect 3276 30818 3332 30828
rect 3500 30994 3556 31052
rect 3500 30942 3502 30994
rect 3554 30942 3556 30994
rect 3500 30884 3556 30942
rect 3948 30994 4004 31500
rect 3948 30942 3950 30994
rect 4002 30942 4004 30994
rect 3948 30930 4004 30942
rect 4284 31220 4340 31230
rect 4284 30994 4340 31164
rect 4284 30942 4286 30994
rect 4338 30942 4340 30994
rect 4284 30930 4340 30942
rect 3500 30818 3556 30828
rect 4396 30884 4452 31502
rect 4396 30772 4452 30828
rect 2492 30270 2494 30322
rect 2546 30270 2548 30322
rect 2492 30258 2548 30270
rect 4284 30716 4452 30772
rect 4508 31332 4564 31614
rect 4508 30772 4564 31276
rect 4844 31108 4900 32396
rect 4956 32386 5012 32396
rect 4956 31892 5012 31902
rect 4956 31798 5012 31836
rect 5628 31780 5684 33404
rect 5740 35756 5908 35812
rect 5740 34468 5796 35756
rect 6188 35698 6244 35710
rect 6188 35646 6190 35698
rect 6242 35646 6244 35698
rect 5852 34916 5908 34926
rect 6188 34916 6244 35646
rect 6524 35138 6580 37884
rect 7420 37940 7476 37950
rect 7420 37846 7476 37884
rect 7196 37828 7252 37838
rect 7196 37734 7252 37772
rect 7644 37826 7700 38444
rect 8092 38274 8148 38780
rect 8428 38668 8484 39900
rect 8540 39732 8596 39742
rect 8652 39732 8708 40236
rect 8876 40180 8932 40190
rect 8540 39730 8708 39732
rect 8540 39678 8542 39730
rect 8594 39678 8708 39730
rect 8540 39676 8708 39678
rect 8764 40178 8932 40180
rect 8764 40126 8878 40178
rect 8930 40126 8932 40178
rect 8764 40124 8932 40126
rect 8540 39508 8596 39676
rect 8540 39442 8596 39452
rect 8652 39284 8708 39294
rect 8652 39058 8708 39228
rect 8652 39006 8654 39058
rect 8706 39006 8708 39058
rect 8652 38994 8708 39006
rect 8764 38668 8820 40124
rect 8876 40114 8932 40124
rect 8988 39956 9044 40460
rect 8092 38222 8094 38274
rect 8146 38222 8148 38274
rect 8092 38210 8148 38222
rect 8316 38612 8484 38668
rect 8652 38612 8820 38668
rect 8876 39900 9044 39956
rect 7644 37774 7646 37826
rect 7698 37774 7700 37826
rect 7084 37716 7140 37726
rect 6636 37044 6692 37054
rect 6636 36482 6692 36988
rect 7084 36594 7140 37660
rect 7644 36596 7700 37774
rect 8204 37940 8260 37950
rect 8204 37266 8260 37884
rect 8204 37214 8206 37266
rect 8258 37214 8260 37266
rect 8204 37202 8260 37214
rect 8316 37268 8372 38612
rect 8652 38162 8708 38612
rect 8876 38388 8932 39900
rect 8988 39396 9044 39406
rect 8988 39302 9044 39340
rect 9212 39060 9268 39070
rect 8988 38948 9044 38958
rect 8988 38854 9044 38892
rect 8652 38110 8654 38162
rect 8706 38110 8708 38162
rect 8652 38098 8708 38110
rect 8764 38332 8932 38388
rect 8428 38052 8484 38062
rect 8428 38050 8596 38052
rect 8428 37998 8430 38050
rect 8482 37998 8596 38050
rect 8428 37996 8596 37998
rect 8428 37986 8484 37996
rect 8540 37492 8596 37996
rect 8652 37716 8708 37726
rect 8764 37716 8820 38332
rect 9100 38050 9156 38062
rect 9100 37998 9102 38050
rect 9154 37998 9156 38050
rect 8708 37660 8820 37716
rect 8988 37716 9044 37726
rect 8652 37650 8708 37660
rect 8764 37492 8820 37502
rect 8540 37490 8820 37492
rect 8540 37438 8766 37490
rect 8818 37438 8820 37490
rect 8540 37436 8820 37438
rect 8764 37426 8820 37436
rect 8876 37492 8932 37502
rect 8988 37492 9044 37660
rect 8876 37490 9044 37492
rect 8876 37438 8878 37490
rect 8930 37438 9044 37490
rect 8876 37436 9044 37438
rect 8876 37426 8932 37436
rect 8652 37268 8708 37278
rect 8316 37266 8708 37268
rect 8316 37214 8654 37266
rect 8706 37214 8708 37266
rect 8316 37212 8708 37214
rect 7980 37154 8036 37166
rect 7980 37102 7982 37154
rect 8034 37102 8036 37154
rect 7980 37044 8036 37102
rect 7980 36978 8036 36988
rect 8652 37044 8708 37212
rect 8652 36978 8708 36988
rect 8988 36820 9044 36830
rect 7084 36542 7086 36594
rect 7138 36542 7140 36594
rect 7084 36530 7140 36542
rect 7308 36540 7700 36596
rect 8204 36708 8260 36718
rect 6636 36430 6638 36482
rect 6690 36430 6692 36482
rect 6636 36418 6692 36430
rect 6524 35086 6526 35138
rect 6578 35086 6580 35138
rect 6524 35074 6580 35086
rect 7084 35810 7140 35822
rect 7084 35758 7086 35810
rect 7138 35758 7140 35810
rect 6412 34916 6468 34926
rect 6188 34914 6468 34916
rect 6188 34862 6414 34914
rect 6466 34862 6468 34914
rect 6188 34860 6468 34862
rect 5852 34822 5908 34860
rect 5740 33684 5796 34412
rect 5740 33458 5796 33628
rect 6412 33572 6468 34860
rect 6972 34692 7028 34702
rect 7084 34692 7140 35758
rect 7028 34636 7140 34692
rect 7196 34914 7252 34926
rect 7196 34862 7198 34914
rect 7250 34862 7252 34914
rect 6972 34356 7028 34636
rect 6972 34018 7028 34300
rect 7196 34354 7252 34862
rect 7196 34302 7198 34354
rect 7250 34302 7252 34354
rect 7196 34290 7252 34302
rect 6972 33966 6974 34018
rect 7026 33966 7028 34018
rect 6972 33954 7028 33966
rect 6412 33506 6468 33516
rect 7196 33572 7252 33582
rect 5740 33406 5742 33458
rect 5794 33406 5796 33458
rect 5740 33394 5796 33406
rect 6636 33460 6692 33470
rect 6692 33404 7028 33460
rect 6636 33366 6692 33404
rect 6300 33124 6356 33134
rect 6300 33030 6356 33068
rect 6972 32786 7028 33404
rect 6972 32734 6974 32786
rect 7026 32734 7028 32786
rect 6972 32722 7028 32734
rect 7084 33124 7140 33134
rect 6076 32562 6132 32574
rect 6076 32510 6078 32562
rect 6130 32510 6132 32562
rect 5740 31780 5796 31790
rect 5628 31778 5796 31780
rect 5628 31726 5742 31778
rect 5794 31726 5796 31778
rect 5628 31724 5796 31726
rect 5740 31714 5796 31724
rect 6076 31556 6132 32510
rect 6188 32562 6244 32574
rect 6188 32510 6190 32562
rect 6242 32510 6244 32562
rect 6188 31780 6244 32510
rect 6524 32562 6580 32574
rect 7084 32564 7140 33068
rect 6524 32510 6526 32562
rect 6578 32510 6580 32562
rect 6412 32452 6468 32462
rect 6412 32358 6468 32396
rect 6188 31686 6244 31724
rect 6412 32004 6468 32014
rect 6524 32004 6580 32510
rect 6468 31948 6580 32004
rect 6860 32508 7140 32564
rect 6412 31778 6468 31948
rect 6412 31726 6414 31778
rect 6466 31726 6468 31778
rect 6412 31714 6468 31726
rect 6860 31778 6916 32508
rect 6860 31726 6862 31778
rect 6914 31726 6916 31778
rect 6860 31714 6916 31726
rect 7084 31780 7140 31790
rect 6300 31556 6356 31566
rect 6076 31554 6356 31556
rect 6076 31502 6302 31554
rect 6354 31502 6356 31554
rect 6076 31500 6356 31502
rect 6300 31490 6356 31500
rect 5180 31220 5236 31230
rect 4956 31108 5012 31118
rect 4844 31106 5012 31108
rect 4844 31054 4958 31106
rect 5010 31054 5012 31106
rect 4844 31052 5012 31054
rect 4956 31042 5012 31052
rect 4284 30324 4340 30716
rect 4508 30706 4564 30716
rect 4476 30604 4740 30614
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4476 30538 4740 30548
rect 4620 30324 4676 30334
rect 4284 30322 4676 30324
rect 4284 30270 4622 30322
rect 4674 30270 4676 30322
rect 4284 30268 4676 30270
rect 4620 30258 4676 30268
rect 4956 30324 5012 30334
rect 4844 29988 4900 29998
rect 2268 29314 2324 29326
rect 2268 29262 2270 29314
rect 2322 29262 2324 29314
rect 2268 27636 2324 29262
rect 4476 29036 4740 29046
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4476 28970 4740 28980
rect 4508 28868 4564 28878
rect 4284 27972 4340 27982
rect 4284 27858 4340 27916
rect 4508 27970 4564 28812
rect 4620 28644 4676 28654
rect 4620 28550 4676 28588
rect 4844 28642 4900 29932
rect 4956 28754 5012 30268
rect 5180 30210 5236 31164
rect 5180 30158 5182 30210
rect 5234 30158 5236 30210
rect 5180 30146 5236 30158
rect 5740 31108 5796 31118
rect 5516 29426 5572 29438
rect 5516 29374 5518 29426
rect 5570 29374 5572 29426
rect 4956 28702 4958 28754
rect 5010 28702 5012 28754
rect 4956 28690 5012 28702
rect 5180 29204 5236 29214
rect 4844 28590 4846 28642
rect 4898 28590 4900 28642
rect 4508 27918 4510 27970
rect 4562 27918 4564 27970
rect 4508 27906 4564 27918
rect 4284 27806 4286 27858
rect 4338 27806 4340 27858
rect 4284 27794 4340 27806
rect 2268 27570 2324 27580
rect 4476 27468 4740 27478
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4476 27402 4740 27412
rect 4844 27188 4900 28590
rect 5180 28642 5236 29148
rect 5180 28590 5182 28642
rect 5234 28590 5236 28642
rect 5180 28578 5236 28590
rect 5180 27860 5236 27870
rect 5068 27188 5124 27198
rect 4844 27186 5124 27188
rect 4844 27134 5070 27186
rect 5122 27134 5124 27186
rect 4844 27132 5124 27134
rect 5068 27122 5124 27132
rect 4620 27076 4676 27086
rect 4620 27074 5012 27076
rect 4620 27022 4622 27074
rect 4674 27022 5012 27074
rect 4620 27020 5012 27022
rect 4620 27010 4676 27020
rect 4844 26180 4900 26190
rect 4476 25900 4740 25910
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4476 25834 4740 25844
rect 4732 25620 4788 25630
rect 4508 25394 4564 25406
rect 4508 25342 4510 25394
rect 4562 25342 4564 25394
rect 3164 24612 3220 24622
rect 3164 24518 3220 24556
rect 4508 24500 4564 25342
rect 4732 25282 4788 25564
rect 4844 25506 4900 26124
rect 4956 25620 5012 27020
rect 4956 25554 5012 25564
rect 4844 25454 4846 25506
rect 4898 25454 4900 25506
rect 4844 25442 4900 25454
rect 5068 25396 5124 25406
rect 5068 25302 5124 25340
rect 4732 25230 4734 25282
rect 4786 25230 4788 25282
rect 4732 25218 4788 25230
rect 4508 24434 4564 24444
rect 4476 24332 4740 24342
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4476 24266 4740 24276
rect 4284 23940 4340 23950
rect 5180 23940 5236 27804
rect 5516 26852 5572 29374
rect 5516 26786 5572 26796
rect 5404 25284 5460 25294
rect 3500 23044 3556 23054
rect 3500 22950 3556 22988
rect 4284 22484 4340 23884
rect 4844 23884 5236 23940
rect 5292 24610 5348 24622
rect 5292 24558 5294 24610
rect 5346 24558 5348 24610
rect 4476 22764 4740 22774
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4476 22698 4740 22708
rect 4732 22484 4788 22494
rect 4284 22482 4788 22484
rect 4284 22430 4734 22482
rect 4786 22430 4788 22482
rect 4284 22428 4788 22430
rect 4732 22418 4788 22428
rect 2156 22082 2212 22092
rect 4844 21924 4900 23884
rect 5068 23716 5124 23726
rect 5068 23714 5236 23716
rect 5068 23662 5070 23714
rect 5122 23662 5236 23714
rect 5068 23660 5236 23662
rect 5068 23650 5124 23660
rect 4956 23044 5012 23054
rect 4956 22370 5012 22988
rect 4956 22318 4958 22370
rect 5010 22318 5012 22370
rect 4956 22306 5012 22318
rect 4844 21868 5012 21924
rect 4844 21588 4900 21598
rect 4844 21494 4900 21532
rect 4476 21196 4740 21206
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4476 21130 4740 21140
rect 4732 21028 4788 21038
rect 4732 20802 4788 20972
rect 4956 21026 5012 21868
rect 5180 21588 5236 23660
rect 5292 23604 5348 24558
rect 5292 23538 5348 23548
rect 5180 21522 5236 21532
rect 4956 20974 4958 21026
rect 5010 20974 5012 21026
rect 4956 20962 5012 20974
rect 4844 20916 4900 20926
rect 4844 20822 4900 20860
rect 4732 20750 4734 20802
rect 4786 20750 4788 20802
rect 4732 20738 4788 20750
rect 5404 20130 5460 25228
rect 5628 23042 5684 23054
rect 5628 22990 5630 23042
rect 5682 22990 5684 23042
rect 5628 22036 5684 22990
rect 5628 21970 5684 21980
rect 5516 21474 5572 21486
rect 5516 21422 5518 21474
rect 5570 21422 5572 21474
rect 5516 20244 5572 21422
rect 5740 21028 5796 31052
rect 7084 30882 7140 31724
rect 7196 31668 7252 33516
rect 7308 33236 7364 36540
rect 8204 35922 8260 36652
rect 8540 36482 8596 36494
rect 8540 36430 8542 36482
rect 8594 36430 8596 36482
rect 8204 35870 8206 35922
rect 8258 35870 8260 35922
rect 8204 35858 8260 35870
rect 8316 36258 8372 36270
rect 8316 36206 8318 36258
rect 8370 36206 8372 36258
rect 7644 35588 7700 35598
rect 8316 35588 8372 36206
rect 7644 35586 8372 35588
rect 7644 35534 7646 35586
rect 7698 35534 8372 35586
rect 7644 35532 8372 35534
rect 7644 35522 7700 35532
rect 7756 34916 7812 34926
rect 7756 34822 7812 34860
rect 7420 34804 7476 34814
rect 7420 34710 7476 34748
rect 8316 34804 8372 34814
rect 8204 34692 8260 34702
rect 7532 34580 7588 34590
rect 7420 34356 7476 34366
rect 7420 34262 7476 34300
rect 7532 34242 7588 34524
rect 7532 34190 7534 34242
rect 7586 34190 7588 34242
rect 7532 34178 7588 34190
rect 7644 34244 7700 34254
rect 7420 33236 7476 33246
rect 7308 33234 7476 33236
rect 7308 33182 7422 33234
rect 7474 33182 7476 33234
rect 7308 33180 7476 33182
rect 7420 33170 7476 33180
rect 7644 32900 7700 34188
rect 8204 34130 8260 34636
rect 8316 34244 8372 34748
rect 8540 34580 8596 36430
rect 8988 35922 9044 36764
rect 8988 35870 8990 35922
rect 9042 35870 9044 35922
rect 8988 35858 9044 35870
rect 8764 35700 8820 35710
rect 8764 35606 8820 35644
rect 8764 34916 8820 34926
rect 8764 34822 8820 34860
rect 8316 34242 8484 34244
rect 8316 34190 8318 34242
rect 8370 34190 8484 34242
rect 8316 34188 8484 34190
rect 8316 34178 8372 34188
rect 8204 34078 8206 34130
rect 8258 34078 8260 34130
rect 8204 34066 8260 34078
rect 7756 33124 7812 33134
rect 8316 33124 8372 33134
rect 7812 33122 8372 33124
rect 7812 33070 8318 33122
rect 8370 33070 8372 33122
rect 7812 33068 8372 33070
rect 7756 33030 7812 33068
rect 7644 32844 7924 32900
rect 7756 32452 7812 32462
rect 7756 32358 7812 32396
rect 7420 32340 7476 32350
rect 7420 32338 7700 32340
rect 7420 32286 7422 32338
rect 7474 32286 7700 32338
rect 7420 32284 7700 32286
rect 7420 32274 7476 32284
rect 7644 32004 7700 32284
rect 7308 31892 7364 31902
rect 7308 31798 7364 31836
rect 7532 31780 7588 31790
rect 7196 31612 7364 31668
rect 7308 31218 7364 31612
rect 7308 31166 7310 31218
rect 7362 31166 7364 31218
rect 7308 31154 7364 31166
rect 7532 31218 7588 31724
rect 7532 31166 7534 31218
rect 7586 31166 7588 31218
rect 7532 31154 7588 31166
rect 7644 31106 7700 31948
rect 7868 31890 7924 32844
rect 7868 31838 7870 31890
rect 7922 31838 7924 31890
rect 7868 31826 7924 31838
rect 7980 32450 8036 32462
rect 7980 32398 7982 32450
rect 8034 32398 8036 32450
rect 7980 31892 8036 32398
rect 8316 32452 8372 33068
rect 8428 32788 8484 34188
rect 8540 33460 8596 34524
rect 8652 34802 8708 34814
rect 8652 34750 8654 34802
rect 8706 34750 8708 34802
rect 8652 33572 8708 34750
rect 8876 34692 8932 34702
rect 8764 34636 8876 34692
rect 8764 34132 8820 34636
rect 8876 34626 8932 34636
rect 8876 34356 8932 34366
rect 9100 34356 9156 37998
rect 8876 34354 9156 34356
rect 8876 34302 8878 34354
rect 8930 34302 9156 34354
rect 8876 34300 9156 34302
rect 8876 34290 8932 34300
rect 8764 34076 8932 34132
rect 8652 33506 8708 33516
rect 8876 33460 8932 34076
rect 8988 34130 9044 34142
rect 8988 34078 8990 34130
rect 9042 34078 9044 34130
rect 8988 33684 9044 34078
rect 8988 33618 9044 33628
rect 9100 33572 9156 33582
rect 9212 33572 9268 39004
rect 9324 38668 9380 41468
rect 9660 40964 9716 40974
rect 9436 40180 9492 40190
rect 9436 38834 9492 40124
rect 9436 38782 9438 38834
rect 9490 38782 9492 38834
rect 9436 38770 9492 38782
rect 9548 39618 9604 39630
rect 9548 39566 9550 39618
rect 9602 39566 9604 39618
rect 9548 38836 9604 39566
rect 9548 38770 9604 38780
rect 9660 38668 9716 40908
rect 9324 38612 9492 38668
rect 9324 37940 9380 37950
rect 9324 35700 9380 37884
rect 9324 34580 9380 35644
rect 9436 35252 9492 38612
rect 9548 38612 9716 38668
rect 9548 35252 9604 38612
rect 9660 37940 9716 37950
rect 9660 37846 9716 37884
rect 9660 37268 9716 37278
rect 9660 37174 9716 37212
rect 9660 35476 9716 35486
rect 9660 35382 9716 35420
rect 9772 35364 9828 44604
rect 10444 44324 10500 44828
rect 10556 44324 10612 44334
rect 10444 44322 10612 44324
rect 10444 44270 10558 44322
rect 10610 44270 10612 44322
rect 10444 44268 10612 44270
rect 10668 44324 10724 45836
rect 10780 45890 10836 45902
rect 10780 45838 10782 45890
rect 10834 45838 10836 45890
rect 10780 45108 10836 45838
rect 10892 45780 10948 46508
rect 11452 45892 11508 45902
rect 11228 45780 11284 45790
rect 10892 45778 11284 45780
rect 10892 45726 11230 45778
rect 11282 45726 11284 45778
rect 10892 45724 11284 45726
rect 11228 45714 11284 45724
rect 11452 45218 11508 45836
rect 11452 45166 11454 45218
rect 11506 45166 11508 45218
rect 11452 45154 11508 45166
rect 11564 45666 11620 45678
rect 11564 45614 11566 45666
rect 11618 45614 11620 45666
rect 10780 45106 11060 45108
rect 10780 45054 10782 45106
rect 10834 45054 11060 45106
rect 10780 45052 11060 45054
rect 10780 45042 10836 45052
rect 10780 44324 10836 44334
rect 10668 44322 10836 44324
rect 10668 44270 10782 44322
rect 10834 44270 10836 44322
rect 10668 44268 10836 44270
rect 10556 44258 10612 44268
rect 10780 44258 10836 44268
rect 10892 44210 10948 44222
rect 10892 44158 10894 44210
rect 10946 44158 10948 44210
rect 9884 44100 9940 44110
rect 10892 44100 10948 44158
rect 9884 44098 10052 44100
rect 9884 44046 9886 44098
rect 9938 44046 10052 44098
rect 9884 44044 10052 44046
rect 9884 44034 9940 44044
rect 9996 43652 10052 44044
rect 10332 44044 10948 44100
rect 10332 43762 10388 44044
rect 11004 43988 11060 45052
rect 11116 44996 11172 45006
rect 11564 44996 11620 45614
rect 11116 44994 11620 44996
rect 11116 44942 11118 44994
rect 11170 44942 11620 44994
rect 11116 44940 11620 44942
rect 11116 44324 11172 44940
rect 11340 44548 11396 44558
rect 11676 44548 11732 46620
rect 12348 46450 12404 46462
rect 12348 46398 12350 46450
rect 12402 46398 12404 46450
rect 12348 45890 12404 46398
rect 12796 46002 12852 47404
rect 12796 45950 12798 46002
rect 12850 45950 12852 46002
rect 12796 45938 12852 45950
rect 12348 45838 12350 45890
rect 12402 45838 12404 45890
rect 12348 45826 12404 45838
rect 12684 45892 12740 45902
rect 12684 45798 12740 45836
rect 12908 45780 12964 45790
rect 11340 44546 11732 44548
rect 11340 44494 11342 44546
rect 11394 44494 11732 44546
rect 11340 44492 11732 44494
rect 12796 45724 12908 45780
rect 11340 44482 11396 44492
rect 12460 44324 12516 44334
rect 12796 44324 12852 45724
rect 12908 45686 12964 45724
rect 12908 45108 12964 45118
rect 12908 45014 12964 45052
rect 11116 44268 11620 44324
rect 10892 43932 11060 43988
rect 11452 44100 11508 44110
rect 10892 43764 10948 43932
rect 11452 43876 11508 44044
rect 10332 43710 10334 43762
rect 10386 43710 10388 43762
rect 10332 43698 10388 43710
rect 10780 43708 10948 43764
rect 11004 43820 11508 43876
rect 9884 42756 9940 42766
rect 9884 41300 9940 42700
rect 9996 42308 10052 43596
rect 10220 43540 10276 43550
rect 10444 43540 10500 43550
rect 10220 43538 10388 43540
rect 10220 43486 10222 43538
rect 10274 43486 10388 43538
rect 10220 43484 10388 43486
rect 10220 43474 10276 43484
rect 10332 42980 10388 43484
rect 10444 43446 10500 43484
rect 10332 42914 10388 42924
rect 10444 42754 10500 42766
rect 10444 42702 10446 42754
rect 10498 42702 10500 42754
rect 9996 42242 10052 42252
rect 10332 42644 10388 42654
rect 10332 41858 10388 42588
rect 10444 42308 10500 42702
rect 10444 42242 10500 42252
rect 10332 41806 10334 41858
rect 10386 41806 10388 41858
rect 10332 41794 10388 41806
rect 10444 41970 10500 41982
rect 10444 41918 10446 41970
rect 10498 41918 10500 41970
rect 10108 41748 10164 41758
rect 9884 41074 9940 41244
rect 9884 41022 9886 41074
rect 9938 41022 9940 41074
rect 9884 41010 9940 41022
rect 9996 41746 10164 41748
rect 9996 41694 10110 41746
rect 10162 41694 10164 41746
rect 9996 41692 10164 41694
rect 9996 40964 10052 41692
rect 10108 41682 10164 41692
rect 10220 41188 10276 41198
rect 10444 41188 10500 41918
rect 10780 41524 10836 43708
rect 10892 43540 10948 43550
rect 11004 43540 11060 43820
rect 11228 43652 11284 43662
rect 11228 43558 11284 43596
rect 11452 43650 11508 43820
rect 11452 43598 11454 43650
rect 11506 43598 11508 43650
rect 11452 43586 11508 43598
rect 10892 43538 11060 43540
rect 10892 43486 10894 43538
rect 10946 43486 11060 43538
rect 10892 43484 11060 43486
rect 11116 43538 11172 43550
rect 11116 43486 11118 43538
rect 11170 43486 11172 43538
rect 10892 43474 10948 43484
rect 11116 43092 11172 43486
rect 11564 43428 11620 44268
rect 12460 44322 12852 44324
rect 12460 44270 12462 44322
rect 12514 44270 12852 44322
rect 12460 44268 12852 44270
rect 12460 44258 12516 44268
rect 12124 44210 12180 44222
rect 12124 44158 12126 44210
rect 12178 44158 12180 44210
rect 12124 43764 12180 44158
rect 12236 44100 12292 44110
rect 12236 44006 12292 44044
rect 12124 43762 12628 43764
rect 12124 43710 12126 43762
rect 12178 43710 12628 43762
rect 12124 43708 12628 43710
rect 12124 43698 12180 43708
rect 11004 43036 11172 43092
rect 11452 43372 11620 43428
rect 11676 43538 11732 43550
rect 11676 43486 11678 43538
rect 11730 43486 11732 43538
rect 10892 42756 10948 42766
rect 11004 42756 11060 43036
rect 11116 42868 11172 42878
rect 11116 42774 11172 42812
rect 10892 42754 11060 42756
rect 10892 42702 10894 42754
rect 10946 42702 11060 42754
rect 10892 42700 11060 42702
rect 10892 42196 10948 42700
rect 10892 42130 10948 42140
rect 11116 42084 11172 42094
rect 11004 41970 11060 41982
rect 11004 41918 11006 41970
rect 11058 41918 11060 41970
rect 10780 41458 10836 41468
rect 10892 41858 10948 41870
rect 10892 41806 10894 41858
rect 10946 41806 10948 41858
rect 10220 41186 10444 41188
rect 10220 41134 10222 41186
rect 10274 41134 10444 41186
rect 10220 41132 10444 41134
rect 10220 41122 10276 41132
rect 10444 41122 10500 41132
rect 10780 41298 10836 41310
rect 10780 41246 10782 41298
rect 10834 41246 10836 41298
rect 9996 40898 10052 40908
rect 10780 40964 10836 41246
rect 10780 40898 10836 40908
rect 9884 40628 9940 40638
rect 9884 40402 9940 40572
rect 10780 40516 10836 40554
rect 10780 40450 10836 40460
rect 9884 40350 9886 40402
rect 9938 40350 9940 40402
rect 9884 40338 9940 40350
rect 10444 40404 10500 40414
rect 10444 40402 10724 40404
rect 10444 40350 10446 40402
rect 10498 40350 10724 40402
rect 10444 40348 10724 40350
rect 10444 40338 10500 40348
rect 10444 39508 10500 39518
rect 10444 39414 10500 39452
rect 10220 38836 10276 38846
rect 10108 38724 10164 38762
rect 10220 38742 10276 38780
rect 10108 38658 10164 38668
rect 9996 38162 10052 38174
rect 9996 38110 9998 38162
rect 10050 38110 10052 38162
rect 9884 38050 9940 38062
rect 9884 37998 9886 38050
rect 9938 37998 9940 38050
rect 9884 37044 9940 37998
rect 9996 38052 10052 38110
rect 9996 37986 10052 37996
rect 10220 37828 10276 37838
rect 10220 37490 10276 37772
rect 10220 37438 10222 37490
rect 10274 37438 10276 37490
rect 10220 37426 10276 37438
rect 10332 37380 10388 37390
rect 10332 37378 10612 37380
rect 10332 37326 10334 37378
rect 10386 37326 10612 37378
rect 10332 37324 10612 37326
rect 10332 37314 10388 37324
rect 9884 36978 9940 36988
rect 10108 37042 10164 37054
rect 10108 36990 10110 37042
rect 10162 36990 10164 37042
rect 10108 36932 10164 36990
rect 9996 36876 10164 36932
rect 9996 36820 10052 36876
rect 9884 36764 10052 36820
rect 9884 36258 9940 36764
rect 10556 36708 10612 37324
rect 10668 37044 10724 40348
rect 10892 39730 10948 41806
rect 11004 41412 11060 41918
rect 11004 41346 11060 41356
rect 11116 41188 11172 42028
rect 11452 41636 11508 43372
rect 11676 42980 11732 43486
rect 12012 43538 12068 43550
rect 12236 43540 12292 43550
rect 12012 43486 12014 43538
rect 12066 43486 12068 43538
rect 12012 43204 12068 43486
rect 11676 42914 11732 42924
rect 11788 43148 12068 43204
rect 12124 43538 12292 43540
rect 12124 43486 12238 43538
rect 12290 43486 12292 43538
rect 12124 43484 12292 43486
rect 11788 42754 11844 43148
rect 11788 42702 11790 42754
rect 11842 42702 11844 42754
rect 11788 42644 11844 42702
rect 11788 42578 11844 42588
rect 12012 42756 12068 42766
rect 12124 42756 12180 43484
rect 12236 43474 12292 43484
rect 12572 43538 12628 43708
rect 12572 43486 12574 43538
rect 12626 43486 12628 43538
rect 12572 43474 12628 43486
rect 12684 43652 12740 43662
rect 12236 42980 12292 42990
rect 12236 42886 12292 42924
rect 12684 42756 12740 43596
rect 12012 42754 12180 42756
rect 12012 42702 12014 42754
rect 12066 42702 12180 42754
rect 12012 42700 12180 42702
rect 12572 42700 12740 42756
rect 12796 43314 12852 43326
rect 12796 43262 12798 43314
rect 12850 43262 12852 43314
rect 11900 41970 11956 41982
rect 11900 41918 11902 41970
rect 11954 41918 11956 41970
rect 11564 41860 11620 41870
rect 11564 41858 11844 41860
rect 11564 41806 11566 41858
rect 11618 41806 11844 41858
rect 11564 41804 11844 41806
rect 11564 41794 11620 41804
rect 11452 41580 11732 41636
rect 11564 41298 11620 41310
rect 11564 41246 11566 41298
rect 11618 41246 11620 41298
rect 10892 39678 10894 39730
rect 10946 39678 10948 39730
rect 10892 39284 10948 39678
rect 10892 39218 10948 39228
rect 11004 41132 11172 41188
rect 11228 41188 11284 41198
rect 10892 38948 10948 38958
rect 11004 38948 11060 41132
rect 11116 40628 11172 40638
rect 11116 40534 11172 40572
rect 10892 38946 11060 38948
rect 10892 38894 10894 38946
rect 10946 38894 11060 38946
rect 10892 38892 11060 38894
rect 10892 38882 10948 38892
rect 11228 38836 11284 41132
rect 11564 41188 11620 41246
rect 11564 40402 11620 41132
rect 11564 40350 11566 40402
rect 11618 40350 11620 40402
rect 11564 40338 11620 40350
rect 11116 38780 11284 38836
rect 11116 38668 11172 38780
rect 10892 38612 11172 38668
rect 10780 38052 10836 38062
rect 10780 37958 10836 37996
rect 10668 36978 10724 36988
rect 10780 37378 10836 37390
rect 10780 37326 10782 37378
rect 10834 37326 10836 37378
rect 10556 36642 10612 36652
rect 9884 36206 9886 36258
rect 9938 36206 9940 36258
rect 9884 36148 9940 36206
rect 9884 35698 9940 36092
rect 9884 35646 9886 35698
rect 9938 35646 9940 35698
rect 9884 35634 9940 35646
rect 9996 36484 10052 36494
rect 9772 35308 9940 35364
rect 9548 35196 9828 35252
rect 9436 35186 9492 35196
rect 9772 35028 9828 35196
rect 9772 34962 9828 34972
rect 9324 34524 9492 34580
rect 9212 33516 9380 33572
rect 8876 33404 9044 33460
rect 8540 33394 8596 33404
rect 8764 33348 8820 33358
rect 8764 33236 8820 33292
rect 8876 33236 8932 33246
rect 8764 33234 8932 33236
rect 8764 33182 8878 33234
rect 8930 33182 8932 33234
rect 8764 33180 8932 33182
rect 8876 33170 8932 33180
rect 8876 32788 8932 32798
rect 8988 32788 9044 33404
rect 8428 32732 8596 32788
rect 8540 32564 8596 32732
rect 8876 32786 9044 32788
rect 8876 32734 8878 32786
rect 8930 32734 9044 32786
rect 8876 32732 9044 32734
rect 9100 33346 9156 33516
rect 9100 33294 9102 33346
rect 9154 33294 9156 33346
rect 8876 32722 8932 32732
rect 8988 32564 9044 32574
rect 8540 32562 9044 32564
rect 8540 32510 8990 32562
rect 9042 32510 9044 32562
rect 8540 32508 9044 32510
rect 8988 32498 9044 32508
rect 8428 32452 8484 32462
rect 8316 32450 8484 32452
rect 8316 32398 8430 32450
rect 8482 32398 8484 32450
rect 8316 32396 8484 32398
rect 8428 32340 8484 32396
rect 8428 32274 8484 32284
rect 8876 32340 8932 32350
rect 9100 32340 9156 33294
rect 8876 32338 9156 32340
rect 8876 32286 8878 32338
rect 8930 32286 9156 32338
rect 8876 32284 9156 32286
rect 8876 32274 8932 32284
rect 8876 32004 8932 32014
rect 8876 31910 8932 31948
rect 7980 31826 8036 31836
rect 8316 31780 8372 31790
rect 8316 31686 8372 31724
rect 9212 31778 9268 31790
rect 9212 31726 9214 31778
rect 9266 31726 9268 31778
rect 8988 31668 9044 31678
rect 7980 31332 8036 31342
rect 7980 31218 8036 31276
rect 7980 31166 7982 31218
rect 8034 31166 8036 31218
rect 7980 31154 8036 31166
rect 8988 31220 9044 31612
rect 8988 31126 9044 31164
rect 7644 31054 7646 31106
rect 7698 31054 7700 31106
rect 7644 31042 7700 31054
rect 7084 30830 7086 30882
rect 7138 30830 7140 30882
rect 7084 30818 7140 30830
rect 8540 30882 8596 30894
rect 8540 30830 8542 30882
rect 8594 30830 8596 30882
rect 6972 30772 7028 30782
rect 6860 29540 6916 29550
rect 6300 29426 6356 29438
rect 6300 29374 6302 29426
rect 6354 29374 6356 29426
rect 5964 29316 6020 29326
rect 5964 29222 6020 29260
rect 5964 28644 6020 28654
rect 6300 28644 6356 29374
rect 6860 29426 6916 29484
rect 6860 29374 6862 29426
rect 6914 29374 6916 29426
rect 6860 29362 6916 29374
rect 6972 28866 7028 30716
rect 8316 30772 8372 30782
rect 8316 30678 8372 30716
rect 7196 30324 7252 30334
rect 7196 30322 7700 30324
rect 7196 30270 7198 30322
rect 7250 30270 7700 30322
rect 7196 30268 7700 30270
rect 7196 30258 7252 30268
rect 7644 30210 7700 30268
rect 7644 30158 7646 30210
rect 7698 30158 7700 30210
rect 7644 30146 7700 30158
rect 8540 30212 8596 30830
rect 9212 30772 9268 31726
rect 9212 30706 9268 30716
rect 9212 30324 9268 30334
rect 9212 30230 9268 30268
rect 7308 30098 7364 30110
rect 7308 30046 7310 30098
rect 7362 30046 7364 30098
rect 7084 29986 7140 29998
rect 7084 29934 7086 29986
rect 7138 29934 7140 29986
rect 7084 29540 7140 29934
rect 7084 29474 7140 29484
rect 6972 28814 6974 28866
rect 7026 28814 7028 28866
rect 6972 28802 7028 28814
rect 7196 28754 7252 28766
rect 7196 28702 7198 28754
rect 7250 28702 7252 28754
rect 5964 28642 6356 28644
rect 5964 28590 5966 28642
rect 6018 28590 6356 28642
rect 5964 28588 6356 28590
rect 6748 28644 6804 28654
rect 5964 26292 6020 28588
rect 6748 28550 6804 28588
rect 6972 28644 7028 28654
rect 6412 27858 6468 27870
rect 6412 27806 6414 27858
rect 6466 27806 6468 27858
rect 6300 27746 6356 27758
rect 6300 27694 6302 27746
rect 6354 27694 6356 27746
rect 6300 26908 6356 27694
rect 6412 27298 6468 27806
rect 6412 27246 6414 27298
rect 6466 27246 6468 27298
rect 6412 27234 6468 27246
rect 6748 27074 6804 27086
rect 6748 27022 6750 27074
rect 6802 27022 6804 27074
rect 6300 26852 6580 26908
rect 6300 26786 6356 26796
rect 5964 25284 6020 26236
rect 6412 26180 6468 26190
rect 6412 26086 6468 26124
rect 5964 25218 6020 25228
rect 6300 25282 6356 25294
rect 6300 25230 6302 25282
rect 6354 25230 6356 25282
rect 6076 24724 6132 24734
rect 6300 24724 6356 25230
rect 6524 24946 6580 26852
rect 6748 25732 6804 27022
rect 6524 24894 6526 24946
rect 6578 24894 6580 24946
rect 6524 24882 6580 24894
rect 6636 25676 6804 25732
rect 6860 26852 6916 26862
rect 6076 24722 6356 24724
rect 6076 24670 6078 24722
rect 6130 24670 6356 24722
rect 6076 24668 6356 24670
rect 5852 24500 5908 24510
rect 5852 23716 5908 24444
rect 5964 23716 6020 23726
rect 5852 23714 6020 23716
rect 5852 23662 5966 23714
rect 6018 23662 6020 23714
rect 5852 23660 6020 23662
rect 5852 22370 5908 23660
rect 5964 23650 6020 23660
rect 5964 23380 6020 23390
rect 5964 23044 6020 23324
rect 6076 23156 6132 24668
rect 6524 23828 6580 23838
rect 6636 23828 6692 25676
rect 6580 23772 6692 23828
rect 6748 25508 6804 25518
rect 6524 23734 6580 23772
rect 6300 23156 6356 23166
rect 6076 23154 6356 23156
rect 6076 23102 6302 23154
rect 6354 23102 6356 23154
rect 6076 23100 6356 23102
rect 5964 22988 6132 23044
rect 6076 22482 6132 22988
rect 6076 22430 6078 22482
rect 6130 22430 6132 22482
rect 6076 22418 6132 22430
rect 5852 22318 5854 22370
rect 5906 22318 5908 22370
rect 5852 22306 5908 22318
rect 6300 21588 6356 23100
rect 5740 20972 5908 21028
rect 5516 20178 5572 20188
rect 5404 20078 5406 20130
rect 5458 20078 5460 20130
rect 5404 20066 5460 20078
rect 5068 20018 5124 20030
rect 5068 19966 5070 20018
rect 5122 19966 5124 20018
rect 4956 19906 5012 19918
rect 4956 19854 4958 19906
rect 5010 19854 5012 19906
rect 4956 19796 5012 19854
rect 5068 19908 5124 19966
rect 5068 19842 5124 19852
rect 5740 19908 5796 19918
rect 4956 19730 5012 19740
rect 4476 19628 4740 19638
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4476 19562 4740 19572
rect 1596 19394 1652 19404
rect 5740 19124 5796 19852
rect 5740 19058 5796 19068
rect 4476 18060 4740 18070
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4476 17994 4740 18004
rect 4476 16492 4740 16502
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4476 16426 4740 16436
rect 5852 15148 5908 20972
rect 6300 20578 6356 21532
rect 6748 21028 6804 25452
rect 6860 25396 6916 26796
rect 6860 24836 6916 25340
rect 6972 25060 7028 28588
rect 7196 27858 7252 28702
rect 7308 28644 7364 30046
rect 8428 30098 8484 30110
rect 8428 30046 8430 30098
rect 8482 30046 8484 30098
rect 7756 29988 7812 29998
rect 7812 29932 7924 29988
rect 7756 29894 7812 29932
rect 7756 29538 7812 29550
rect 7756 29486 7758 29538
rect 7810 29486 7812 29538
rect 7756 29092 7812 29486
rect 7756 29026 7812 29036
rect 7308 28578 7364 28588
rect 7868 28532 7924 29932
rect 7980 29986 8036 29998
rect 7980 29934 7982 29986
rect 8034 29934 8036 29986
rect 7980 29426 8036 29934
rect 7980 29374 7982 29426
rect 8034 29374 8036 29426
rect 7980 29362 8036 29374
rect 8428 29316 8484 30046
rect 8428 29222 8484 29260
rect 8428 28868 8484 28878
rect 8540 28868 8596 30156
rect 8988 30100 9044 30110
rect 8988 30006 9044 30044
rect 8764 29652 8820 29662
rect 8764 29558 8820 29596
rect 8484 28812 8596 28868
rect 8428 28642 8484 28812
rect 8428 28590 8430 28642
rect 8482 28590 8484 28642
rect 8428 28578 8484 28590
rect 7868 28466 7924 28476
rect 9324 28420 9380 33516
rect 9436 32004 9492 34524
rect 9660 33124 9716 33134
rect 9660 33030 9716 33068
rect 9884 32900 9940 35308
rect 9996 34914 10052 36428
rect 10668 36482 10724 36494
rect 10668 36430 10670 36482
rect 10722 36430 10724 36482
rect 10444 36372 10500 36382
rect 10444 36278 10500 36316
rect 10108 35812 10164 35822
rect 10108 35718 10164 35756
rect 9996 34862 9998 34914
rect 10050 34862 10052 34914
rect 9996 34850 10052 34862
rect 10332 35698 10388 35710
rect 10332 35646 10334 35698
rect 10386 35646 10388 35698
rect 10332 33572 10388 35646
rect 10444 35476 10500 35486
rect 10444 35382 10500 35420
rect 10332 33506 10388 33516
rect 10444 34916 10500 34926
rect 9996 33460 10052 33470
rect 9996 33366 10052 33404
rect 9436 31938 9492 31948
rect 9660 32844 9940 32900
rect 9436 31668 9492 31678
rect 9436 30212 9492 31612
rect 9548 30994 9604 31006
rect 9548 30942 9550 30994
rect 9602 30942 9604 30994
rect 9548 30772 9604 30942
rect 9548 30706 9604 30716
rect 9548 30436 9604 30446
rect 9660 30436 9716 32844
rect 9772 32676 9828 32686
rect 9772 32674 9940 32676
rect 9772 32622 9774 32674
rect 9826 32622 9940 32674
rect 9772 32620 9940 32622
rect 9772 32610 9828 32620
rect 9772 32452 9828 32462
rect 9772 31778 9828 32396
rect 9884 32116 9940 32620
rect 9884 32050 9940 32060
rect 9996 32562 10052 32574
rect 9996 32510 9998 32562
rect 10050 32510 10052 32562
rect 9772 31726 9774 31778
rect 9826 31726 9828 31778
rect 9772 31714 9828 31726
rect 9884 31892 9940 31902
rect 9884 31778 9940 31836
rect 9884 31726 9886 31778
rect 9938 31726 9940 31778
rect 9884 31714 9940 31726
rect 9884 31220 9940 31230
rect 9996 31220 10052 32510
rect 9884 31218 10052 31220
rect 9884 31166 9886 31218
rect 9938 31166 10052 31218
rect 9884 31164 10052 31166
rect 9884 31154 9940 31164
rect 9548 30434 9716 30436
rect 9548 30382 9550 30434
rect 9602 30382 9716 30434
rect 9548 30380 9716 30382
rect 10220 31106 10276 31118
rect 10220 31054 10222 31106
rect 10274 31054 10276 31106
rect 9548 30370 9604 30380
rect 10220 30324 10276 31054
rect 9436 30146 9492 30156
rect 9996 30268 10276 30324
rect 9996 29988 10052 30268
rect 9660 29540 9716 29550
rect 9660 29446 9716 29484
rect 9772 29428 9828 29438
rect 9772 29426 9940 29428
rect 9772 29374 9774 29426
rect 9826 29374 9940 29426
rect 9772 29372 9940 29374
rect 9772 29362 9828 29372
rect 9660 29202 9716 29214
rect 9660 29150 9662 29202
rect 9714 29150 9716 29202
rect 9548 28868 9604 28878
rect 9548 28774 9604 28812
rect 7196 27806 7198 27858
rect 7250 27806 7252 27858
rect 7084 27074 7140 27086
rect 7084 27022 7086 27074
rect 7138 27022 7140 27074
rect 7084 26852 7140 27022
rect 7084 26786 7140 26796
rect 7196 26628 7252 27806
rect 8988 28364 9380 28420
rect 9436 28642 9492 28654
rect 9436 28590 9438 28642
rect 9490 28590 9492 28642
rect 8988 27298 9044 28364
rect 9436 27972 9492 28590
rect 9660 28420 9716 29150
rect 9772 28644 9828 28654
rect 9772 28550 9828 28588
rect 9660 28354 9716 28364
rect 9492 27916 9716 27972
rect 9436 27906 9492 27916
rect 8988 27246 8990 27298
rect 9042 27246 9044 27298
rect 8988 27234 9044 27246
rect 8652 27188 8708 27198
rect 8652 27094 8708 27132
rect 9100 27132 9604 27188
rect 7196 26562 7252 26572
rect 8652 26628 8708 26638
rect 8092 26514 8148 26526
rect 8092 26462 8094 26514
rect 8146 26462 8148 26514
rect 7196 26402 7252 26414
rect 7196 26350 7198 26402
rect 7250 26350 7252 26402
rect 6972 25004 7140 25060
rect 6972 24836 7028 24846
rect 6860 24834 7028 24836
rect 6860 24782 6974 24834
rect 7026 24782 7028 24834
rect 6860 24780 7028 24782
rect 6748 20962 6804 20972
rect 6860 24276 6916 24286
rect 6860 22260 6916 24220
rect 6972 22260 7028 24780
rect 7084 22482 7140 25004
rect 7196 24276 7252 26350
rect 7196 24210 7252 24220
rect 7420 26180 7476 26190
rect 7420 24500 7476 26124
rect 8092 25508 8148 26462
rect 8204 26292 8260 26302
rect 8204 26290 8372 26292
rect 8204 26238 8206 26290
rect 8258 26238 8372 26290
rect 8204 26236 8372 26238
rect 8204 26226 8260 26236
rect 8092 25442 8148 25452
rect 7868 24722 7924 24734
rect 7868 24670 7870 24722
rect 7922 24670 7924 24722
rect 7868 24500 7924 24670
rect 7420 24444 7924 24500
rect 8204 24610 8260 24622
rect 8204 24558 8206 24610
rect 8258 24558 8260 24610
rect 7084 22430 7086 22482
rect 7138 22430 7140 22482
rect 7084 22418 7140 22430
rect 7196 24052 7252 24062
rect 7420 24052 7476 24444
rect 7196 24050 7476 24052
rect 7196 23998 7198 24050
rect 7250 23998 7476 24050
rect 7196 23996 7476 23998
rect 7196 22482 7252 23996
rect 7532 23938 7588 23950
rect 7532 23886 7534 23938
rect 7586 23886 7588 23938
rect 7532 23044 7588 23886
rect 7980 23156 8036 23166
rect 7980 23154 8148 23156
rect 7980 23102 7982 23154
rect 8034 23102 8148 23154
rect 7980 23100 8148 23102
rect 7980 23090 8036 23100
rect 7532 22978 7588 22988
rect 7196 22430 7198 22482
rect 7250 22430 7252 22482
rect 7196 22418 7252 22430
rect 7420 22930 7476 22942
rect 7420 22878 7422 22930
rect 7474 22878 7476 22930
rect 7420 22260 7476 22878
rect 7980 22260 8036 22270
rect 6972 22258 8036 22260
rect 6972 22206 7982 22258
rect 8034 22206 8036 22258
rect 6972 22204 8036 22206
rect 6860 21026 6916 22204
rect 7980 22194 8036 22204
rect 6860 20974 6862 21026
rect 6914 20974 6916 21026
rect 6860 20962 6916 20974
rect 6300 20526 6302 20578
rect 6354 20526 6356 20578
rect 6300 20020 6356 20526
rect 6300 19954 6356 19964
rect 6748 20804 6804 20814
rect 6748 19796 6804 20748
rect 7980 20804 8036 20814
rect 8092 20804 8148 23100
rect 8204 21810 8260 24558
rect 8316 23380 8372 26236
rect 8428 26290 8484 26302
rect 8428 26238 8430 26290
rect 8482 26238 8484 26290
rect 8428 25620 8484 26238
rect 8428 25554 8484 25564
rect 8428 25394 8484 25406
rect 8428 25342 8430 25394
rect 8482 25342 8484 25394
rect 8428 24050 8484 25342
rect 8652 24162 8708 26572
rect 9100 26514 9156 27132
rect 9100 26462 9102 26514
rect 9154 26462 9156 26514
rect 9100 26450 9156 26462
rect 9324 26962 9380 26974
rect 9324 26910 9326 26962
rect 9378 26910 9380 26962
rect 8988 26402 9044 26414
rect 8988 26350 8990 26402
rect 9042 26350 9044 26402
rect 8764 26292 8820 26302
rect 8764 26198 8820 26236
rect 8652 24110 8654 24162
rect 8706 24110 8708 24162
rect 8652 24098 8708 24110
rect 8428 23998 8430 24050
rect 8482 23998 8484 24050
rect 8428 23940 8484 23998
rect 8428 23874 8484 23884
rect 8652 23940 8708 23950
rect 8652 23846 8708 23884
rect 8988 23828 9044 26350
rect 9324 24948 9380 26910
rect 9436 26964 9492 26974
rect 9436 26292 9492 26908
rect 9548 26962 9604 27132
rect 9548 26910 9550 26962
rect 9602 26910 9604 26962
rect 9548 26898 9604 26910
rect 9548 26292 9604 26302
rect 9436 26290 9604 26292
rect 9436 26238 9550 26290
rect 9602 26238 9604 26290
rect 9436 26236 9604 26238
rect 9548 26226 9604 26236
rect 9660 25506 9716 27916
rect 9772 27860 9828 27870
rect 9772 27766 9828 27804
rect 9884 27748 9940 29372
rect 9772 27076 9828 27086
rect 9884 27076 9940 27692
rect 9772 27074 9940 27076
rect 9772 27022 9774 27074
rect 9826 27022 9940 27074
rect 9772 27020 9940 27022
rect 9772 27010 9828 27020
rect 9996 26964 10052 29932
rect 10108 30100 10164 30110
rect 10444 30100 10500 34860
rect 10556 34468 10612 34478
rect 10556 34130 10612 34412
rect 10556 34078 10558 34130
rect 10610 34078 10612 34130
rect 10556 34066 10612 34078
rect 10556 33684 10612 33694
rect 10668 33684 10724 36430
rect 10780 36484 10836 37326
rect 10780 36418 10836 36428
rect 10892 35586 10948 38612
rect 11228 38164 11284 38174
rect 11228 38070 11284 38108
rect 11004 37940 11060 37950
rect 11004 37266 11060 37884
rect 11564 37268 11620 37278
rect 11004 37214 11006 37266
rect 11058 37214 11060 37266
rect 11004 37202 11060 37214
rect 11452 37266 11620 37268
rect 11452 37214 11566 37266
rect 11618 37214 11620 37266
rect 11452 37212 11620 37214
rect 11004 36932 11060 36942
rect 11004 36594 11060 36876
rect 11004 36542 11006 36594
rect 11058 36542 11060 36594
rect 11004 36530 11060 36542
rect 11004 36260 11060 36270
rect 11228 36260 11284 36270
rect 11004 36258 11172 36260
rect 11004 36206 11006 36258
rect 11058 36206 11172 36258
rect 11004 36204 11172 36206
rect 11004 36194 11060 36204
rect 10892 35534 10894 35586
rect 10946 35534 10948 35586
rect 10892 35522 10948 35534
rect 11004 35698 11060 35710
rect 11004 35646 11006 35698
rect 11058 35646 11060 35698
rect 10780 35364 10836 35374
rect 11004 35364 11060 35646
rect 10780 34354 10836 35308
rect 10780 34302 10782 34354
rect 10834 34302 10836 34354
rect 10780 34290 10836 34302
rect 10892 35308 11060 35364
rect 10612 33628 10724 33684
rect 10556 31220 10612 33628
rect 10780 33348 10836 33358
rect 10780 33254 10836 33292
rect 10668 33234 10724 33246
rect 10668 33182 10670 33234
rect 10722 33182 10724 33234
rect 10668 31444 10724 33182
rect 10780 33124 10836 33134
rect 10780 32452 10836 33068
rect 10892 32676 10948 35308
rect 11004 35140 11060 35150
rect 11004 35046 11060 35084
rect 11116 34692 11172 36204
rect 11228 36258 11396 36260
rect 11228 36206 11230 36258
rect 11282 36206 11396 36258
rect 11228 36204 11396 36206
rect 11228 36194 11284 36204
rect 11340 35138 11396 36204
rect 11452 35252 11508 37212
rect 11564 37202 11620 37212
rect 11676 36596 11732 41580
rect 11788 40516 11844 41804
rect 11788 40402 11844 40460
rect 11788 40350 11790 40402
rect 11842 40350 11844 40402
rect 11788 40338 11844 40350
rect 11788 39620 11844 39630
rect 11788 39060 11844 39564
rect 11788 38994 11844 39004
rect 11788 38836 11844 38846
rect 11788 38742 11844 38780
rect 11452 35186 11508 35196
rect 11564 36540 11732 36596
rect 11788 38276 11844 38286
rect 11340 35086 11342 35138
rect 11394 35086 11396 35138
rect 11340 34804 11396 35086
rect 11564 35028 11620 36540
rect 11676 36372 11732 36382
rect 11676 36278 11732 36316
rect 11676 36148 11732 36158
rect 11676 35698 11732 36092
rect 11676 35646 11678 35698
rect 11730 35646 11732 35698
rect 11676 35634 11732 35646
rect 11340 34738 11396 34748
rect 11452 34972 11620 35028
rect 11116 34626 11172 34636
rect 11340 34242 11396 34254
rect 11340 34190 11342 34242
rect 11394 34190 11396 34242
rect 11340 33908 11396 34190
rect 11452 34132 11508 34972
rect 11676 34914 11732 34926
rect 11676 34862 11678 34914
rect 11730 34862 11732 34914
rect 11676 34804 11732 34862
rect 11676 34738 11732 34748
rect 11788 34356 11844 38220
rect 11900 38052 11956 41918
rect 12012 40516 12068 42700
rect 12236 42082 12292 42094
rect 12236 42030 12238 42082
rect 12290 42030 12292 42082
rect 12124 41188 12180 41198
rect 12236 41188 12292 42030
rect 12572 41972 12628 42700
rect 12684 42532 12740 42542
rect 12796 42532 12852 43262
rect 12684 42530 12852 42532
rect 12684 42478 12686 42530
rect 12738 42478 12852 42530
rect 12684 42476 12852 42478
rect 12684 42466 12740 42476
rect 12572 41878 12628 41916
rect 12796 41412 12852 41422
rect 13020 41412 13076 48748
rect 13132 43316 13188 43326
rect 13132 43222 13188 43260
rect 12796 41410 13076 41412
rect 12796 41358 12798 41410
rect 12850 41358 13076 41410
rect 12796 41356 13076 41358
rect 12796 41346 12852 41356
rect 12124 41186 12292 41188
rect 12124 41134 12126 41186
rect 12178 41134 12292 41186
rect 12124 41132 12292 41134
rect 12124 41122 12180 41132
rect 12908 41076 12964 41086
rect 12908 41074 13076 41076
rect 12908 41022 12910 41074
rect 12962 41022 13076 41074
rect 12908 41020 13076 41022
rect 12908 41010 12964 41020
rect 12348 40962 12404 40974
rect 12348 40910 12350 40962
rect 12402 40910 12404 40962
rect 12348 40740 12404 40910
rect 12796 40962 12852 40974
rect 12796 40910 12798 40962
rect 12850 40910 12852 40962
rect 12348 40684 12740 40740
rect 12236 40516 12292 40526
rect 12012 40514 12292 40516
rect 12012 40462 12238 40514
rect 12290 40462 12292 40514
rect 12012 40460 12292 40462
rect 12236 40450 12292 40460
rect 12684 40514 12740 40684
rect 12684 40462 12686 40514
rect 12738 40462 12740 40514
rect 12684 40450 12740 40462
rect 12572 40402 12628 40414
rect 12572 40350 12574 40402
rect 12626 40350 12628 40402
rect 12572 40068 12628 40350
rect 12572 40002 12628 40012
rect 12796 39844 12852 40910
rect 12460 39788 12852 39844
rect 13020 39844 13076 41020
rect 12124 39730 12180 39742
rect 12124 39678 12126 39730
rect 12178 39678 12180 39730
rect 12124 38836 12180 39678
rect 12236 39620 12292 39630
rect 12460 39620 12516 39788
rect 13020 39778 13076 39788
rect 13132 40852 13188 40862
rect 12908 39732 12964 39742
rect 12908 39638 12964 39676
rect 12236 39526 12292 39564
rect 12348 39564 12516 39620
rect 12572 39620 12628 39630
rect 13132 39620 13188 40796
rect 11900 37986 11956 37996
rect 12012 38050 12068 38062
rect 12012 37998 12014 38050
rect 12066 37998 12068 38050
rect 11900 37378 11956 37390
rect 11900 37326 11902 37378
rect 11954 37326 11956 37378
rect 11900 36484 11956 37326
rect 12012 37044 12068 37998
rect 12012 36978 12068 36988
rect 12124 36932 12180 38780
rect 12348 37940 12404 39564
rect 12572 39058 12628 39564
rect 13020 39564 13188 39620
rect 12572 39006 12574 39058
rect 12626 39006 12628 39058
rect 12572 38994 12628 39006
rect 12796 39508 12852 39518
rect 12684 38948 12740 38958
rect 12348 37874 12404 37884
rect 12460 38836 12516 38846
rect 12348 37380 12404 37390
rect 12348 37266 12404 37324
rect 12348 37214 12350 37266
rect 12402 37214 12404 37266
rect 12348 37202 12404 37214
rect 12124 36876 12404 36932
rect 12012 36820 12068 36830
rect 12012 36596 12068 36764
rect 12012 36530 12068 36540
rect 11900 36418 11956 36428
rect 12348 35924 12404 36876
rect 12460 36594 12516 38780
rect 12684 38274 12740 38892
rect 12796 38834 12852 39452
rect 13020 39396 13076 39564
rect 12908 39340 13076 39396
rect 13132 39396 13188 39406
rect 12908 38946 12964 39340
rect 12908 38894 12910 38946
rect 12962 38894 12964 38946
rect 12908 38882 12964 38894
rect 12796 38782 12798 38834
rect 12850 38782 12852 38834
rect 12796 38770 12852 38782
rect 12684 38222 12686 38274
rect 12738 38222 12740 38274
rect 12684 38210 12740 38222
rect 12684 38052 12740 38062
rect 12684 37958 12740 37996
rect 13132 37828 13188 39340
rect 13132 37762 13188 37772
rect 12460 36542 12462 36594
rect 12514 36542 12516 36594
rect 12460 36530 12516 36542
rect 12572 37378 12628 37390
rect 12572 37326 12574 37378
rect 12626 37326 12628 37378
rect 12572 36596 12628 37326
rect 12572 36530 12628 36540
rect 12684 37380 12740 37390
rect 12572 35924 12628 35934
rect 12348 35922 12628 35924
rect 12348 35870 12574 35922
rect 12626 35870 12628 35922
rect 12348 35868 12628 35870
rect 12572 35858 12628 35868
rect 11676 34300 11844 34356
rect 11900 35700 11956 35710
rect 11452 34076 11620 34132
rect 11452 33908 11508 33918
rect 11340 33852 11452 33908
rect 11452 33842 11508 33852
rect 10892 32582 10948 32620
rect 11004 32562 11060 32574
rect 11004 32510 11006 32562
rect 11058 32510 11060 32562
rect 10892 32452 10948 32462
rect 10780 32450 10948 32452
rect 10780 32398 10894 32450
rect 10946 32398 10948 32450
rect 10780 32396 10948 32398
rect 10892 32386 10948 32396
rect 11004 32452 11060 32510
rect 11004 32386 11060 32396
rect 11340 32562 11396 32574
rect 11340 32510 11342 32562
rect 11394 32510 11396 32562
rect 10668 31378 10724 31388
rect 11004 31890 11060 31902
rect 11004 31838 11006 31890
rect 11058 31838 11060 31890
rect 10556 31164 10724 31220
rect 10556 30996 10612 31006
rect 10556 30322 10612 30940
rect 10556 30270 10558 30322
rect 10610 30270 10612 30322
rect 10556 30258 10612 30270
rect 10668 30212 10724 31164
rect 10780 30994 10836 31006
rect 10780 30942 10782 30994
rect 10834 30942 10836 30994
rect 10780 30436 10836 30942
rect 10780 30370 10836 30380
rect 11004 30324 11060 31838
rect 11116 31780 11172 31790
rect 11340 31780 11396 32510
rect 11172 31724 11396 31780
rect 11116 31220 11172 31724
rect 11116 30994 11172 31164
rect 11228 31556 11284 31566
rect 11228 31218 11284 31500
rect 11228 31166 11230 31218
rect 11282 31166 11284 31218
rect 11228 31154 11284 31166
rect 11116 30942 11118 30994
rect 11170 30942 11172 30994
rect 11116 30930 11172 30942
rect 11116 30324 11172 30334
rect 11004 30268 11116 30324
rect 11116 30230 11172 30268
rect 11452 30212 11508 30222
rect 10668 30156 10836 30212
rect 10444 30044 10724 30100
rect 10108 29538 10164 30044
rect 10108 29486 10110 29538
rect 10162 29486 10164 29538
rect 10108 28980 10164 29486
rect 10332 29204 10388 29214
rect 10332 29110 10388 29148
rect 10108 28914 10164 28924
rect 9996 26898 10052 26908
rect 10108 28756 10164 28766
rect 10108 27858 10164 28700
rect 10444 28644 10500 28654
rect 10108 27806 10110 27858
rect 10162 27806 10164 27858
rect 10108 26908 10164 27806
rect 10332 28642 10500 28644
rect 10332 28590 10446 28642
rect 10498 28590 10500 28642
rect 10332 28588 10500 28590
rect 10332 26908 10388 28588
rect 10444 28578 10500 28588
rect 10556 28644 10612 28654
rect 10444 28420 10500 28430
rect 10444 28326 10500 28364
rect 10556 27074 10612 28588
rect 10668 27970 10724 30044
rect 10668 27918 10670 27970
rect 10722 27918 10724 27970
rect 10668 27906 10724 27918
rect 10556 27022 10558 27074
rect 10610 27022 10612 27074
rect 10556 27010 10612 27022
rect 10108 26852 10276 26908
rect 10332 26852 10500 26908
rect 10108 26516 10164 26526
rect 10108 26422 10164 26460
rect 9660 25454 9662 25506
rect 9714 25454 9716 25506
rect 9436 24948 9492 24958
rect 9324 24946 9492 24948
rect 9324 24894 9438 24946
rect 9490 24894 9492 24946
rect 9324 24892 9492 24894
rect 9436 24882 9492 24892
rect 9660 24834 9716 25454
rect 9660 24782 9662 24834
rect 9714 24782 9716 24834
rect 8988 23772 9380 23828
rect 9324 23716 9380 23772
rect 8316 23314 8372 23324
rect 8988 23604 9044 23614
rect 8428 23154 8484 23166
rect 8428 23102 8430 23154
rect 8482 23102 8484 23154
rect 8316 23044 8372 23054
rect 8428 23044 8484 23102
rect 8372 22988 8484 23044
rect 8876 23042 8932 23054
rect 8876 22990 8878 23042
rect 8930 22990 8932 23042
rect 8316 22978 8372 22988
rect 8876 22932 8932 22990
rect 8876 22866 8932 22876
rect 8988 22370 9044 23548
rect 8988 22318 8990 22370
rect 9042 22318 9044 22370
rect 8988 22306 9044 22318
rect 9324 22370 9380 23660
rect 9324 22318 9326 22370
rect 9378 22318 9380 22370
rect 9324 22306 9380 22318
rect 9436 22148 9492 22158
rect 9436 22054 9492 22092
rect 8204 21758 8206 21810
rect 8258 21758 8260 21810
rect 8204 21700 8260 21758
rect 8204 21634 8260 21644
rect 9548 21698 9604 21710
rect 9548 21646 9550 21698
rect 9602 21646 9604 21698
rect 9100 21474 9156 21486
rect 9100 21422 9102 21474
rect 9154 21422 9156 21474
rect 9100 21364 9156 21422
rect 9100 21298 9156 21308
rect 8036 20748 8148 20804
rect 8764 20804 8820 20814
rect 7980 20738 8036 20748
rect 8764 20710 8820 20748
rect 9548 20692 9604 21646
rect 9660 20914 9716 24782
rect 9772 25284 9828 25294
rect 10220 25284 10276 26852
rect 10444 25284 10500 26852
rect 10780 25618 10836 30156
rect 11452 30118 11508 30156
rect 10892 29540 10948 29550
rect 10892 28868 10948 29484
rect 11564 29538 11620 34076
rect 11676 33124 11732 34300
rect 11676 33058 11732 33068
rect 11676 32452 11732 32462
rect 11676 32358 11732 32396
rect 11900 31556 11956 35644
rect 12012 35700 12068 35710
rect 12684 35700 12740 37324
rect 12012 35698 12740 35700
rect 12012 35646 12014 35698
rect 12066 35646 12740 35698
rect 12012 35644 12740 35646
rect 12796 36372 12852 36382
rect 12012 35634 12068 35644
rect 12236 35252 12292 35262
rect 12124 34914 12180 34926
rect 12124 34862 12126 34914
rect 12178 34862 12180 34914
rect 12124 34132 12180 34862
rect 12012 33572 12068 33582
rect 12012 32564 12068 33516
rect 12124 33460 12180 34076
rect 12236 34916 12292 35196
rect 12236 34130 12292 34860
rect 12796 34802 12852 36316
rect 13020 35812 13076 35822
rect 13020 35810 13188 35812
rect 13020 35758 13022 35810
rect 13074 35758 13188 35810
rect 13020 35756 13188 35758
rect 13020 35746 13076 35756
rect 12908 34916 12964 34926
rect 12908 34914 13076 34916
rect 12908 34862 12910 34914
rect 12962 34862 13076 34914
rect 12908 34860 13076 34862
rect 12908 34850 12964 34860
rect 12796 34750 12798 34802
rect 12850 34750 12852 34802
rect 12460 34468 12516 34478
rect 12236 34078 12238 34130
rect 12290 34078 12292 34130
rect 12236 34066 12292 34078
rect 12348 34412 12460 34468
rect 12124 33394 12180 33404
rect 12348 33458 12404 34412
rect 12460 34402 12516 34412
rect 12348 33406 12350 33458
rect 12402 33406 12404 33458
rect 12348 33394 12404 33406
rect 12460 33460 12516 33470
rect 12460 33346 12516 33404
rect 12460 33294 12462 33346
rect 12514 33294 12516 33346
rect 12460 33282 12516 33294
rect 12012 32450 12068 32508
rect 12012 32398 12014 32450
rect 12066 32398 12068 32450
rect 12012 32386 12068 32398
rect 12348 32562 12404 32574
rect 12348 32510 12350 32562
rect 12402 32510 12404 32562
rect 12348 31892 12404 32510
rect 12348 31826 12404 31836
rect 11900 31490 11956 31500
rect 12460 31778 12516 31790
rect 12460 31726 12462 31778
rect 12514 31726 12516 31778
rect 11788 31220 11844 31230
rect 11788 31106 11844 31164
rect 11788 31054 11790 31106
rect 11842 31054 11844 31106
rect 11788 31042 11844 31054
rect 12348 30994 12404 31006
rect 12348 30942 12350 30994
rect 12402 30942 12404 30994
rect 12348 30884 12404 30942
rect 12012 30436 12068 30446
rect 12012 30210 12068 30380
rect 12012 30158 12014 30210
rect 12066 30158 12068 30210
rect 12012 30146 12068 30158
rect 12348 30212 12404 30828
rect 12348 30146 12404 30156
rect 12460 30882 12516 31726
rect 12796 30996 12852 34750
rect 12908 33236 12964 33246
rect 12908 33142 12964 33180
rect 13020 32452 13076 34860
rect 13132 34020 13188 35756
rect 13132 33954 13188 33964
rect 13132 32676 13188 32686
rect 13132 32582 13188 32620
rect 13020 32386 13076 32396
rect 12796 30902 12852 30940
rect 13020 31780 13076 31790
rect 12460 30830 12462 30882
rect 12514 30830 12516 30882
rect 11564 29486 11566 29538
rect 11618 29486 11620 29538
rect 11564 29474 11620 29486
rect 12460 30100 12516 30830
rect 13020 30770 13076 31724
rect 13020 30718 13022 30770
rect 13074 30718 13076 30770
rect 13020 30706 13076 30718
rect 12684 30324 12740 30334
rect 12684 30230 12740 30268
rect 11116 29426 11172 29438
rect 11116 29374 11118 29426
rect 11170 29374 11172 29426
rect 11116 29316 11172 29374
rect 12012 29428 12068 29438
rect 12012 29426 12180 29428
rect 12012 29374 12014 29426
rect 12066 29374 12180 29426
rect 12012 29372 12180 29374
rect 12012 29362 12068 29372
rect 11116 29250 11172 29260
rect 11228 29204 11284 29214
rect 10892 27858 10948 28812
rect 10892 27806 10894 27858
rect 10946 27806 10948 27858
rect 10892 27794 10948 27806
rect 11004 29092 11060 29102
rect 10892 27636 10948 27646
rect 10892 26514 10948 27580
rect 10892 26462 10894 26514
rect 10946 26462 10948 26514
rect 10892 26450 10948 26462
rect 10780 25566 10782 25618
rect 10834 25566 10836 25618
rect 10780 25554 10836 25566
rect 10220 25228 10388 25284
rect 9772 24834 9828 25228
rect 9772 24782 9774 24834
rect 9826 24782 9828 24834
rect 9772 24770 9828 24782
rect 10220 23940 10276 23950
rect 10108 23884 10220 23940
rect 9996 23044 10052 23054
rect 9884 21586 9940 21598
rect 9884 21534 9886 21586
rect 9938 21534 9940 21586
rect 9884 21476 9940 21534
rect 9884 21410 9940 21420
rect 9660 20862 9662 20914
rect 9714 20862 9716 20914
rect 9660 20850 9716 20862
rect 9996 20916 10052 22988
rect 10108 21252 10164 23884
rect 10220 23874 10276 23884
rect 10220 23380 10276 23390
rect 10332 23380 10388 25228
rect 10444 25218 10500 25228
rect 10556 25506 10612 25518
rect 10556 25454 10558 25506
rect 10610 25454 10612 25506
rect 10556 25396 10612 25454
rect 11004 25396 11060 29036
rect 11228 28644 11284 29148
rect 11116 28642 11284 28644
rect 11116 28590 11230 28642
rect 11282 28590 11284 28642
rect 11116 28588 11284 28590
rect 11116 27186 11172 28588
rect 11228 28578 11284 28588
rect 11340 28532 11396 28542
rect 11340 28438 11396 28476
rect 12012 28532 12068 28542
rect 11452 28420 11508 28430
rect 11452 28326 11508 28364
rect 11116 27134 11118 27186
rect 11170 27134 11172 27186
rect 11116 27122 11172 27134
rect 11228 27970 11284 27982
rect 11228 27918 11230 27970
rect 11282 27918 11284 27970
rect 11228 26908 11284 27918
rect 12012 27970 12068 28476
rect 12012 27918 12014 27970
rect 12066 27918 12068 27970
rect 12012 27906 12068 27918
rect 11788 27858 11844 27870
rect 11788 27806 11790 27858
rect 11842 27806 11844 27858
rect 11788 27748 11844 27806
rect 11788 26908 11844 27692
rect 12124 27300 12180 29372
rect 12236 28980 12292 28990
rect 12236 28420 12292 28924
rect 12460 28754 12516 30044
rect 12572 30210 12628 30222
rect 12572 30158 12574 30210
rect 12626 30158 12628 30210
rect 12572 29652 12628 30158
rect 12572 29586 12628 29596
rect 12796 29538 12852 29550
rect 12796 29486 12798 29538
rect 12850 29486 12852 29538
rect 12460 28702 12462 28754
rect 12514 28702 12516 28754
rect 12460 28690 12516 28702
rect 12572 29426 12628 29438
rect 12572 29374 12574 29426
rect 12626 29374 12628 29426
rect 12572 28756 12628 29374
rect 12572 28690 12628 28700
rect 12796 28532 12852 29486
rect 12908 28756 12964 28766
rect 12908 28642 12964 28700
rect 12908 28590 12910 28642
rect 12962 28590 12964 28642
rect 12908 28578 12964 28590
rect 12796 28466 12852 28476
rect 12236 27970 12292 28364
rect 12236 27918 12238 27970
rect 12290 27918 12292 27970
rect 12236 27906 12292 27918
rect 12908 27972 12964 27982
rect 13244 27972 13300 48860
rect 13468 44884 13524 49532
rect 13580 49494 13636 49532
rect 13692 47458 13748 51100
rect 14140 50594 14196 50606
rect 14140 50542 14142 50594
rect 14194 50542 14196 50594
rect 14140 50428 14196 50542
rect 13804 50372 14196 50428
rect 14364 50596 14420 50606
rect 13804 50148 13860 50372
rect 13804 49028 13860 50092
rect 13916 50036 13972 50046
rect 13972 49980 14196 50036
rect 13916 49942 13972 49980
rect 14028 49028 14084 49038
rect 13804 49026 14084 49028
rect 13804 48974 14030 49026
rect 14082 48974 14084 49026
rect 13804 48972 14084 48974
rect 14028 48962 14084 48972
rect 14140 48914 14196 49980
rect 14252 49810 14308 49822
rect 14252 49758 14254 49810
rect 14306 49758 14308 49810
rect 14252 49588 14308 49758
rect 14252 49522 14308 49532
rect 14364 49026 14420 50540
rect 14476 50036 14532 52108
rect 15036 52108 15204 52164
rect 15036 51378 15092 52108
rect 15148 51940 15204 51950
rect 15204 51884 15316 51940
rect 15148 51874 15204 51884
rect 15036 51326 15038 51378
rect 15090 51326 15092 51378
rect 15036 51314 15092 51326
rect 14924 50708 14980 50718
rect 14924 50614 14980 50652
rect 14812 50594 14868 50606
rect 14812 50542 14814 50594
rect 14866 50542 14868 50594
rect 14588 50036 14644 50046
rect 14476 50034 14644 50036
rect 14476 49982 14590 50034
rect 14642 49982 14644 50034
rect 14476 49980 14644 49982
rect 14588 49970 14644 49980
rect 14812 50034 14868 50542
rect 15260 50428 15316 51884
rect 15372 51828 15428 51838
rect 15372 51378 15428 51772
rect 15372 51326 15374 51378
rect 15426 51326 15428 51378
rect 15372 51314 15428 51326
rect 16044 51378 16100 52444
rect 16156 51828 16212 52892
rect 16268 52882 16324 52892
rect 16492 52948 16548 52958
rect 16492 52854 16548 52892
rect 16828 52946 16884 52958
rect 16828 52894 16830 52946
rect 16882 52894 16884 52946
rect 16828 52612 16884 52894
rect 16828 52546 16884 52556
rect 17500 52834 17556 52846
rect 17500 52782 17502 52834
rect 17554 52782 17556 52834
rect 17500 52612 17556 52782
rect 17500 52546 17556 52556
rect 16156 51762 16212 51772
rect 16604 52164 16660 52174
rect 16044 51326 16046 51378
rect 16098 51326 16100 51378
rect 16044 51314 16100 51326
rect 16492 51154 16548 51166
rect 16492 51102 16494 51154
rect 16546 51102 16548 51154
rect 16492 50818 16548 51102
rect 16492 50766 16494 50818
rect 16546 50766 16548 50818
rect 16492 50754 16548 50766
rect 16044 50708 16100 50718
rect 16044 50614 16100 50652
rect 16604 50706 16660 52108
rect 17612 52164 17668 52174
rect 17612 52070 17668 52108
rect 18060 52164 18116 54460
rect 18172 53732 18228 56252
rect 18508 55972 18564 55982
rect 18284 54404 18340 54414
rect 18284 54310 18340 54348
rect 18284 53732 18340 53742
rect 18172 53676 18284 53732
rect 18284 53666 18340 53676
rect 18508 53172 18564 55916
rect 18620 55186 18676 55198
rect 18620 55134 18622 55186
rect 18674 55134 18676 55186
rect 18620 54738 18676 55134
rect 18620 54686 18622 54738
rect 18674 54686 18676 54738
rect 18620 54674 18676 54686
rect 19068 54516 19124 54526
rect 19068 54422 19124 54460
rect 18732 54404 18788 54414
rect 18732 54310 18788 54348
rect 18956 53732 19012 53742
rect 18956 53506 19012 53676
rect 18956 53454 18958 53506
rect 19010 53454 19012 53506
rect 18956 53442 19012 53454
rect 19292 53172 19348 59200
rect 19836 56476 20100 56486
rect 19892 56420 19940 56476
rect 19996 56420 20044 56476
rect 19836 56410 20100 56420
rect 20860 56308 20916 59200
rect 20860 56242 20916 56252
rect 22092 56308 22148 56318
rect 22092 56214 22148 56252
rect 22428 56196 22484 59200
rect 22428 56130 22484 56140
rect 21084 56084 21140 56094
rect 20748 56082 21140 56084
rect 20748 56030 21086 56082
rect 21138 56030 21140 56082
rect 20748 56028 21140 56030
rect 19852 55970 19908 55982
rect 19852 55918 19854 55970
rect 19906 55918 19908 55970
rect 19852 55076 19908 55918
rect 20748 55410 20804 56028
rect 21084 56018 21140 56028
rect 20748 55358 20750 55410
rect 20802 55358 20804 55410
rect 20748 55346 20804 55358
rect 22204 55522 22260 55534
rect 22204 55470 22206 55522
rect 22258 55470 22260 55522
rect 22204 55412 22260 55470
rect 23996 55412 24052 59200
rect 25564 56308 25620 59200
rect 27132 57090 27188 59200
rect 28700 57316 28756 59200
rect 28700 57260 29204 57316
rect 27132 57038 27134 57090
rect 27186 57038 27188 57090
rect 27132 57026 27188 57038
rect 28364 57090 28420 57102
rect 28364 57038 28366 57090
rect 28418 57038 28420 57090
rect 25564 56242 25620 56252
rect 27468 56308 27524 56318
rect 27468 56214 27524 56252
rect 28364 56306 28420 57038
rect 28364 56254 28366 56306
rect 28418 56254 28420 56306
rect 28364 56242 28420 56254
rect 25340 56196 25396 56206
rect 25340 56102 25396 56140
rect 27132 56082 27188 56094
rect 27132 56030 27134 56082
rect 27186 56030 27188 56082
rect 22204 55356 22484 55412
rect 22428 55300 22484 55356
rect 22988 55356 23268 55412
rect 22876 55300 22932 55310
rect 22428 55298 22932 55300
rect 22428 55246 22878 55298
rect 22930 55246 22932 55298
rect 22428 55244 22932 55246
rect 22876 55234 22932 55244
rect 21868 55188 21924 55198
rect 21868 55094 21924 55132
rect 22316 55186 22372 55198
rect 22316 55134 22318 55186
rect 22370 55134 22372 55186
rect 18508 53116 18676 53172
rect 18284 52164 18340 52174
rect 18060 52162 18340 52164
rect 18060 52110 18286 52162
rect 18338 52110 18340 52162
rect 18060 52108 18340 52110
rect 16604 50654 16606 50706
rect 16658 50654 16660 50706
rect 16604 50642 16660 50654
rect 17500 51380 17556 51390
rect 18060 51380 18116 52108
rect 18284 52098 18340 52108
rect 17500 51378 18116 51380
rect 17500 51326 17502 51378
rect 17554 51326 18116 51378
rect 17500 51324 18116 51326
rect 15372 50596 15428 50606
rect 15372 50502 15428 50540
rect 16828 50594 16884 50606
rect 16828 50542 16830 50594
rect 16882 50542 16884 50594
rect 15484 50482 15540 50494
rect 15484 50430 15486 50482
rect 15538 50430 15540 50482
rect 15484 50428 15540 50430
rect 15148 50372 15540 50428
rect 16828 50428 16884 50542
rect 17388 50482 17444 50494
rect 17388 50430 17390 50482
rect 17442 50430 17444 50482
rect 17388 50428 17444 50430
rect 16828 50372 17444 50428
rect 17500 50428 17556 51324
rect 18172 51268 18228 51278
rect 18172 51266 18452 51268
rect 18172 51214 18174 51266
rect 18226 51214 18452 51266
rect 18172 51212 18452 51214
rect 18172 51202 18228 51212
rect 18396 50818 18452 51212
rect 18396 50766 18398 50818
rect 18450 50766 18452 50818
rect 18396 50754 18452 50766
rect 17500 50372 17668 50428
rect 18508 50372 18564 50382
rect 14812 49982 14814 50034
rect 14866 49982 14868 50034
rect 14812 49970 14868 49982
rect 15036 50036 15092 50046
rect 15036 49942 15092 49980
rect 15148 49922 15204 50372
rect 15148 49870 15150 49922
rect 15202 49870 15204 49922
rect 15148 49858 15204 49870
rect 14364 48974 14366 49026
rect 14418 48974 14420 49026
rect 14364 48962 14420 48974
rect 16380 49026 16436 49038
rect 16380 48974 16382 49026
rect 16434 48974 16436 49026
rect 14140 48862 14142 48914
rect 14194 48862 14196 48914
rect 14140 48850 14196 48862
rect 16044 48914 16100 48926
rect 16044 48862 16046 48914
rect 16098 48862 16100 48914
rect 15708 48804 15764 48814
rect 15596 48748 15708 48804
rect 15372 48130 15428 48142
rect 15372 48078 15374 48130
rect 15426 48078 15428 48130
rect 15372 47796 15428 48078
rect 15596 48020 15652 48748
rect 15708 48738 15764 48748
rect 15708 48468 15764 48478
rect 15708 48354 15764 48412
rect 15820 48468 15876 48478
rect 16044 48468 16100 48862
rect 16380 48468 16436 48974
rect 15820 48466 16324 48468
rect 15820 48414 15822 48466
rect 15874 48414 16324 48466
rect 15820 48412 16324 48414
rect 15820 48402 15876 48412
rect 15708 48302 15710 48354
rect 15762 48302 15764 48354
rect 15708 48290 15764 48302
rect 16156 48242 16212 48254
rect 16156 48190 16158 48242
rect 16210 48190 16212 48242
rect 15820 48020 15876 48030
rect 15596 48018 15876 48020
rect 15596 47966 15822 48018
rect 15874 47966 15876 48018
rect 15596 47964 15876 47966
rect 15820 47954 15876 47964
rect 16156 47796 16212 48190
rect 16268 48244 16324 48412
rect 16380 48402 16436 48412
rect 16716 48916 16772 48926
rect 16716 48466 16772 48860
rect 16716 48414 16718 48466
rect 16770 48414 16772 48466
rect 16716 48402 16772 48414
rect 16828 48468 16884 48478
rect 16828 48374 16884 48412
rect 16604 48244 16660 48254
rect 16268 48242 16660 48244
rect 16268 48190 16606 48242
rect 16658 48190 16660 48242
rect 16268 48188 16660 48190
rect 13692 47406 13694 47458
rect 13746 47406 13748 47458
rect 13692 47124 13748 47406
rect 15260 47740 16212 47796
rect 13580 45892 13636 45902
rect 13580 45798 13636 45836
rect 13692 45668 13748 47068
rect 14364 47346 14420 47358
rect 14364 47294 14366 47346
rect 14418 47294 14420 47346
rect 14364 46900 14420 47294
rect 14924 46900 14980 46910
rect 15260 46900 15316 47740
rect 16044 47572 16100 47582
rect 14364 46834 14420 46844
rect 14476 46898 14980 46900
rect 14476 46846 14926 46898
rect 14978 46846 14980 46898
rect 14476 46844 14980 46846
rect 13916 45890 13972 45902
rect 13916 45838 13918 45890
rect 13970 45838 13972 45890
rect 13916 45780 13972 45838
rect 13916 45714 13972 45724
rect 13580 45612 13748 45668
rect 13580 45108 13636 45612
rect 14476 45556 14532 46844
rect 14924 46834 14980 46844
rect 15036 46844 15316 46900
rect 15932 46900 15988 46910
rect 13692 45500 14532 45556
rect 14700 46674 14756 46686
rect 14700 46622 14702 46674
rect 14754 46622 14756 46674
rect 13692 45218 13748 45500
rect 13692 45166 13694 45218
rect 13746 45166 13748 45218
rect 13692 45154 13748 45166
rect 13580 45042 13636 45052
rect 14476 45108 14532 45118
rect 13468 44828 13748 44884
rect 13356 41860 13412 41870
rect 13356 41766 13412 41804
rect 13580 40628 13636 40638
rect 13356 40514 13412 40526
rect 13356 40462 13358 40514
rect 13410 40462 13412 40514
rect 13356 39508 13412 40462
rect 13468 40516 13524 40526
rect 13468 39618 13524 40460
rect 13468 39566 13470 39618
rect 13522 39566 13524 39618
rect 13468 39554 13524 39566
rect 13580 40402 13636 40572
rect 13580 40350 13582 40402
rect 13634 40350 13636 40402
rect 13356 39442 13412 39452
rect 13356 39060 13412 39070
rect 13356 35698 13412 39004
rect 13580 38052 13636 40350
rect 13692 39396 13748 44828
rect 14476 44434 14532 45052
rect 14476 44382 14478 44434
rect 14530 44382 14532 44434
rect 14476 44370 14532 44382
rect 14700 44434 14756 46622
rect 15036 46452 15092 46844
rect 15932 46806 15988 46844
rect 15820 46786 15876 46798
rect 15820 46734 15822 46786
rect 15874 46734 15876 46786
rect 15148 46676 15204 46686
rect 15148 46582 15204 46620
rect 15372 46674 15428 46686
rect 15372 46622 15374 46674
rect 15426 46622 15428 46674
rect 15036 46396 15316 46452
rect 15036 46004 15092 46014
rect 15036 45910 15092 45948
rect 14700 44382 14702 44434
rect 14754 44382 14756 44434
rect 14700 43428 14756 44382
rect 15148 45332 15204 45342
rect 15148 44434 15204 45276
rect 15148 44382 15150 44434
rect 15202 44382 15204 44434
rect 15148 44370 15204 44382
rect 15260 43708 15316 46396
rect 15372 45108 15428 46622
rect 15596 46676 15652 46686
rect 15596 45892 15652 46620
rect 15820 46676 15876 46734
rect 16044 46786 16100 47516
rect 16492 47570 16548 48188
rect 16604 48178 16660 48188
rect 16492 47518 16494 47570
rect 16546 47518 16548 47570
rect 16492 47506 16548 47518
rect 17052 47236 17108 47246
rect 16940 47234 17108 47236
rect 16940 47182 17054 47234
rect 17106 47182 17108 47234
rect 16940 47180 17108 47182
rect 16716 46900 16772 46910
rect 16044 46734 16046 46786
rect 16098 46734 16100 46786
rect 16044 46722 16100 46734
rect 16156 46898 16772 46900
rect 16156 46846 16718 46898
rect 16770 46846 16772 46898
rect 16156 46844 16772 46846
rect 15820 46610 15876 46620
rect 16044 45892 16100 45902
rect 16156 45892 16212 46844
rect 16716 46834 16772 46844
rect 16492 46676 16548 46686
rect 16828 46676 16884 46686
rect 15596 45798 15652 45836
rect 15708 45890 16212 45892
rect 15708 45838 16046 45890
rect 16098 45838 16212 45890
rect 15708 45836 16212 45838
rect 16380 46674 16548 46676
rect 16380 46622 16494 46674
rect 16546 46622 16548 46674
rect 16380 46620 16548 46622
rect 15372 45042 15428 45052
rect 15708 44996 15764 45836
rect 16044 45826 16100 45836
rect 16156 45666 16212 45678
rect 16156 45614 16158 45666
rect 16210 45614 16212 45666
rect 15932 45108 15988 45118
rect 15988 45052 16100 45108
rect 15932 45042 15988 45052
rect 15820 44996 15876 45006
rect 15708 44994 15876 44996
rect 15708 44942 15822 44994
rect 15874 44942 15876 44994
rect 15708 44940 15876 44942
rect 15820 44772 15876 44940
rect 15372 44716 15876 44772
rect 15372 44322 15428 44716
rect 15372 44270 15374 44322
rect 15426 44270 15428 44322
rect 15372 44258 15428 44270
rect 14700 43362 14756 43372
rect 14924 43652 15316 43708
rect 16044 43708 16100 45052
rect 16156 44884 16212 45614
rect 16268 45666 16324 45678
rect 16268 45614 16270 45666
rect 16322 45614 16324 45666
rect 16268 45332 16324 45614
rect 16268 45266 16324 45276
rect 16268 45108 16324 45118
rect 16380 45108 16436 46620
rect 16492 46610 16548 46620
rect 16716 46674 16884 46676
rect 16716 46622 16830 46674
rect 16882 46622 16884 46674
rect 16716 46620 16884 46622
rect 16492 45892 16548 45902
rect 16548 45836 16660 45892
rect 16492 45826 16548 45836
rect 16268 45106 16436 45108
rect 16268 45054 16270 45106
rect 16322 45054 16436 45106
rect 16268 45052 16436 45054
rect 16268 45042 16324 45052
rect 16492 44884 16548 44894
rect 16156 44882 16548 44884
rect 16156 44830 16494 44882
rect 16546 44830 16548 44882
rect 16156 44828 16548 44830
rect 16492 44818 16548 44828
rect 15372 43652 15428 43662
rect 14924 43426 14980 43652
rect 15372 43558 15428 43596
rect 15820 43652 15876 43662
rect 16044 43652 16436 43708
rect 15820 43650 15988 43652
rect 15820 43598 15822 43650
rect 15874 43598 15988 43650
rect 15820 43596 15988 43598
rect 15820 43586 15876 43596
rect 14924 43374 14926 43426
rect 14978 43374 14980 43426
rect 14924 43204 14980 43374
rect 14924 43138 14980 43148
rect 15036 43540 15092 43550
rect 14700 42756 14756 42766
rect 14700 42662 14756 42700
rect 15036 42754 15092 43484
rect 15708 43540 15764 43550
rect 15708 43446 15764 43484
rect 15820 43316 15876 43326
rect 15036 42702 15038 42754
rect 15090 42702 15092 42754
rect 15036 42690 15092 42702
rect 15596 43314 15876 43316
rect 15596 43262 15822 43314
rect 15874 43262 15876 43314
rect 15596 43260 15876 43262
rect 15596 42754 15652 43260
rect 15820 43250 15876 43260
rect 15596 42702 15598 42754
rect 15650 42702 15652 42754
rect 15596 42690 15652 42702
rect 14812 42532 14868 42542
rect 14812 42438 14868 42476
rect 15932 42084 15988 43596
rect 16380 43650 16436 43652
rect 16380 43598 16382 43650
rect 16434 43598 16436 43650
rect 16380 43586 16436 43598
rect 16492 43652 16548 43662
rect 16604 43652 16660 45836
rect 16716 45332 16772 46620
rect 16828 46610 16884 46620
rect 16940 46676 16996 47180
rect 17052 47170 17108 47180
rect 16716 45266 16772 45276
rect 16828 45108 16884 45118
rect 16828 45014 16884 45052
rect 16828 44210 16884 44222
rect 16828 44158 16830 44210
rect 16882 44158 16884 44210
rect 16828 43708 16884 44158
rect 16492 43650 16660 43652
rect 16492 43598 16494 43650
rect 16546 43598 16660 43650
rect 16492 43596 16660 43598
rect 16492 43586 16548 43596
rect 16268 43540 16324 43550
rect 16268 43446 16324 43484
rect 15372 42028 15988 42084
rect 16268 42754 16324 42766
rect 16268 42702 16270 42754
rect 16322 42702 16324 42754
rect 16268 42532 16324 42702
rect 15148 41860 15204 41870
rect 14476 41412 14532 41422
rect 14028 41300 14084 41310
rect 13916 41298 14084 41300
rect 13916 41246 14030 41298
rect 14082 41246 14084 41298
rect 13916 41244 14084 41246
rect 13804 41188 13860 41198
rect 13804 41094 13860 41132
rect 13916 39730 13972 41244
rect 14028 41234 14084 41244
rect 14476 41298 14532 41356
rect 14476 41246 14478 41298
rect 14530 41246 14532 41298
rect 14476 41234 14532 41246
rect 15036 41300 15092 41310
rect 15036 41186 15092 41244
rect 15148 41298 15204 41804
rect 15148 41246 15150 41298
rect 15202 41246 15204 41298
rect 15148 41234 15204 41246
rect 15260 41636 15316 41646
rect 15260 41300 15316 41580
rect 15036 41134 15038 41186
rect 15090 41134 15092 41186
rect 15036 41122 15092 41134
rect 15260 40964 15316 41244
rect 15260 40898 15316 40908
rect 15372 41074 15428 42028
rect 16268 41972 16324 42476
rect 16492 42756 16548 42766
rect 16380 41972 16436 41982
rect 16268 41970 16436 41972
rect 16268 41918 16382 41970
rect 16434 41918 16436 41970
rect 16268 41916 16436 41918
rect 15484 41860 15540 41870
rect 15484 41858 15764 41860
rect 15484 41806 15486 41858
rect 15538 41806 15764 41858
rect 15484 41804 15764 41806
rect 15484 41794 15540 41804
rect 15708 41412 15764 41804
rect 15820 41858 15876 41870
rect 15820 41806 15822 41858
rect 15874 41806 15876 41858
rect 15820 41636 15876 41806
rect 15820 41570 15876 41580
rect 15708 41356 16324 41412
rect 15596 41188 15652 41198
rect 16044 41188 16100 41198
rect 15596 41186 16100 41188
rect 15596 41134 15598 41186
rect 15650 41134 16046 41186
rect 16098 41134 16100 41186
rect 15596 41132 16100 41134
rect 15596 41122 15652 41132
rect 16044 41122 16100 41132
rect 15372 41022 15374 41074
rect 15426 41022 15428 41074
rect 14140 40852 14196 40862
rect 14028 40740 14084 40750
rect 14028 40514 14084 40684
rect 14028 40462 14030 40514
rect 14082 40462 14084 40514
rect 14028 40450 14084 40462
rect 14140 40514 14196 40796
rect 14140 40462 14142 40514
rect 14194 40462 14196 40514
rect 14140 40450 14196 40462
rect 15372 40516 15428 41022
rect 15932 40964 15988 40974
rect 15932 40870 15988 40908
rect 16156 40962 16212 40974
rect 16156 40910 16158 40962
rect 16210 40910 16212 40962
rect 15372 40450 15428 40460
rect 16156 40516 16212 40910
rect 16156 40450 16212 40460
rect 16268 40514 16324 41356
rect 16380 40626 16436 41916
rect 16492 41860 16548 42700
rect 16604 42642 16660 43596
rect 16716 43652 16884 43708
rect 16716 43586 16772 43596
rect 16828 43538 16884 43550
rect 16828 43486 16830 43538
rect 16882 43486 16884 43538
rect 16828 43204 16884 43486
rect 16828 43138 16884 43148
rect 16604 42590 16606 42642
rect 16658 42590 16660 42642
rect 16604 42578 16660 42590
rect 16716 41860 16772 41870
rect 16492 41804 16716 41860
rect 16716 41766 16772 41804
rect 16380 40574 16382 40626
rect 16434 40574 16436 40626
rect 16380 40562 16436 40574
rect 16492 41524 16548 41534
rect 16268 40462 16270 40514
rect 16322 40462 16324 40514
rect 16268 40450 16324 40462
rect 14364 40402 14420 40414
rect 14364 40350 14366 40402
rect 14418 40350 14420 40402
rect 14028 39844 14084 39854
rect 14084 39788 14196 39844
rect 14028 39778 14084 39788
rect 13916 39678 13918 39730
rect 13970 39678 13972 39730
rect 13916 39666 13972 39678
rect 13692 39330 13748 39340
rect 13804 39618 13860 39630
rect 13804 39566 13806 39618
rect 13858 39566 13860 39618
rect 13692 38836 13748 38874
rect 13692 38770 13748 38780
rect 13804 38668 13860 39566
rect 14028 39620 14084 39630
rect 14028 39526 14084 39564
rect 14028 39060 14084 39070
rect 14140 39060 14196 39788
rect 14084 39004 14196 39060
rect 14028 38966 14084 39004
rect 13692 38612 13860 38668
rect 13692 38164 13748 38612
rect 13804 38546 13860 38556
rect 13916 38722 13972 38734
rect 13916 38670 13918 38722
rect 13970 38670 13972 38722
rect 13692 38098 13748 38108
rect 13916 38052 13972 38670
rect 13580 37716 13636 37996
rect 13804 37996 13972 38052
rect 14252 38052 14308 38062
rect 13692 37940 13748 37950
rect 13692 37846 13748 37884
rect 13580 37660 13748 37716
rect 13580 36484 13636 36494
rect 13580 36390 13636 36428
rect 13356 35646 13358 35698
rect 13410 35646 13412 35698
rect 13356 35634 13412 35646
rect 13468 36370 13524 36382
rect 13468 36318 13470 36370
rect 13522 36318 13524 36370
rect 13468 34468 13524 36318
rect 13692 36258 13748 37660
rect 13692 36206 13694 36258
rect 13746 36206 13748 36258
rect 13692 36194 13748 36206
rect 13804 36036 13860 37996
rect 14252 37958 14308 37996
rect 14364 38050 14420 40350
rect 15596 40404 15652 40414
rect 15372 40292 15428 40302
rect 15260 40290 15428 40292
rect 15260 40238 15374 40290
rect 15426 40238 15428 40290
rect 15260 40236 15428 40238
rect 14812 39618 14868 39630
rect 14812 39566 14814 39618
rect 14866 39566 14868 39618
rect 14812 38834 14868 39566
rect 14812 38782 14814 38834
rect 14866 38782 14868 38834
rect 14812 38612 14868 38782
rect 14812 38546 14868 38556
rect 15148 38612 15204 38622
rect 14364 37998 14366 38050
rect 14418 37998 14420 38050
rect 14364 37986 14420 37998
rect 15148 38050 15204 38556
rect 15260 38162 15316 40236
rect 15372 40226 15428 40236
rect 15372 39620 15428 39630
rect 15372 39526 15428 39564
rect 15484 39508 15540 39518
rect 15484 39414 15540 39452
rect 15372 39396 15428 39406
rect 15372 38948 15428 39340
rect 15372 38834 15428 38892
rect 15372 38782 15374 38834
rect 15426 38782 15428 38834
rect 15372 38770 15428 38782
rect 15596 38668 15652 40348
rect 15932 40404 15988 40414
rect 15932 40402 16100 40404
rect 15932 40350 15934 40402
rect 15986 40350 16100 40402
rect 15932 40348 16100 40350
rect 15932 40338 15988 40348
rect 15820 39620 15876 39630
rect 15820 39506 15876 39564
rect 15820 39454 15822 39506
rect 15874 39454 15876 39506
rect 15820 39442 15876 39454
rect 16044 39618 16100 40348
rect 16044 39566 16046 39618
rect 16098 39566 16100 39618
rect 16044 39396 16100 39566
rect 16044 39330 16100 39340
rect 15820 39172 15876 39182
rect 15596 38612 15764 38668
rect 15260 38110 15262 38162
rect 15314 38110 15316 38162
rect 15260 38098 15316 38110
rect 15148 37998 15150 38050
rect 15202 37998 15204 38050
rect 15148 37986 15204 37998
rect 13580 35980 13860 36036
rect 13916 37826 13972 37838
rect 14140 37828 14196 37838
rect 13916 37774 13918 37826
rect 13970 37774 13972 37826
rect 13580 34916 13636 35980
rect 13804 35588 13860 35598
rect 13580 34850 13636 34860
rect 13692 35532 13804 35588
rect 13468 34402 13524 34412
rect 13692 34354 13748 35532
rect 13804 35522 13860 35532
rect 13804 34916 13860 34954
rect 13804 34850 13860 34860
rect 13916 34804 13972 37774
rect 13916 34738 13972 34748
rect 14028 37826 14196 37828
rect 14028 37774 14142 37826
rect 14194 37774 14196 37826
rect 14028 37772 14196 37774
rect 13692 34302 13694 34354
rect 13746 34302 13748 34354
rect 13692 34290 13748 34302
rect 13804 34690 13860 34702
rect 13804 34638 13806 34690
rect 13858 34638 13860 34690
rect 13468 34020 13524 34030
rect 13468 33926 13524 33964
rect 13804 33348 13860 34638
rect 14028 34132 14084 37772
rect 14140 37762 14196 37772
rect 14476 37378 14532 37390
rect 14476 37326 14478 37378
rect 14530 37326 14532 37378
rect 14252 35700 14308 35710
rect 14252 35606 14308 35644
rect 14476 35026 14532 37326
rect 15148 37380 15204 37390
rect 15148 37286 15204 37324
rect 14476 34974 14478 35026
rect 14530 34974 14532 35026
rect 14476 34962 14532 34974
rect 14700 37268 14756 37278
rect 14140 34914 14196 34926
rect 14140 34862 14142 34914
rect 14194 34862 14196 34914
rect 14140 34244 14196 34862
rect 14700 34692 14756 37212
rect 15372 37268 15428 37278
rect 15372 37174 15428 37212
rect 15260 36482 15316 36494
rect 15260 36430 15262 36482
rect 15314 36430 15316 36482
rect 15260 35364 15316 36430
rect 15708 35924 15764 38612
rect 15820 37938 15876 39116
rect 16380 38834 16436 38846
rect 16380 38782 16382 38834
rect 16434 38782 16436 38834
rect 16380 38724 16436 38782
rect 16380 38658 16436 38668
rect 16492 38162 16548 41468
rect 16604 41186 16660 41198
rect 16604 41134 16606 41186
rect 16658 41134 16660 41186
rect 16604 40404 16660 41134
rect 16828 40404 16884 40414
rect 16604 40402 16884 40404
rect 16604 40350 16830 40402
rect 16882 40350 16884 40402
rect 16604 40348 16884 40350
rect 16604 39956 16660 39966
rect 16604 38946 16660 39900
rect 16604 38894 16606 38946
rect 16658 38894 16660 38946
rect 16604 38882 16660 38894
rect 16716 38948 16772 40348
rect 16828 40338 16884 40348
rect 16716 38892 16884 38948
rect 16492 38110 16494 38162
rect 16546 38110 16548 38162
rect 16492 38098 16548 38110
rect 16156 38052 16212 38062
rect 16156 37958 16212 37996
rect 16604 38052 16660 38062
rect 15820 37886 15822 37938
rect 15874 37886 15876 37938
rect 15820 37874 15876 37886
rect 16268 37938 16324 37950
rect 16268 37886 16270 37938
rect 16322 37886 16324 37938
rect 16268 37492 16324 37886
rect 16156 37436 16324 37492
rect 16044 37154 16100 37166
rect 16044 37102 16046 37154
rect 16098 37102 16100 37154
rect 16044 37044 16100 37102
rect 16044 36978 16100 36988
rect 15372 35476 15428 35486
rect 15428 35420 15540 35476
rect 15372 35410 15428 35420
rect 15260 35298 15316 35308
rect 15260 35028 15316 35038
rect 14476 34636 14756 34692
rect 15036 34802 15092 34814
rect 15036 34750 15038 34802
rect 15090 34750 15092 34802
rect 14140 34178 14196 34188
rect 14252 34244 14308 34254
rect 14252 34242 14420 34244
rect 14252 34190 14254 34242
rect 14306 34190 14420 34242
rect 14252 34188 14420 34190
rect 14252 34178 14308 34188
rect 14028 34066 14084 34076
rect 14140 34020 14196 34030
rect 14028 33796 14084 33806
rect 13804 33282 13860 33292
rect 13916 33572 13972 33582
rect 13916 33346 13972 33516
rect 14028 33570 14084 33740
rect 14028 33518 14030 33570
rect 14082 33518 14084 33570
rect 14028 33506 14084 33518
rect 13916 33294 13918 33346
rect 13970 33294 13972 33346
rect 13916 33282 13972 33294
rect 13692 33122 13748 33134
rect 13692 33070 13694 33122
rect 13746 33070 13748 33122
rect 13580 32564 13636 32574
rect 13468 32562 13636 32564
rect 13468 32510 13582 32562
rect 13634 32510 13636 32562
rect 13468 32508 13636 32510
rect 13356 31780 13412 31790
rect 13468 31780 13524 32508
rect 13580 32498 13636 32508
rect 13692 32340 13748 33070
rect 14028 33124 14084 33134
rect 14028 33030 14084 33068
rect 13412 31724 13524 31780
rect 13580 31892 13636 31902
rect 13356 31714 13412 31724
rect 13580 31666 13636 31836
rect 13580 31614 13582 31666
rect 13634 31614 13636 31666
rect 13580 31602 13636 31614
rect 13468 31444 13524 31454
rect 13468 30994 13524 31388
rect 13468 30942 13470 30994
rect 13522 30942 13524 30994
rect 13468 30930 13524 30942
rect 13580 30994 13636 31006
rect 13580 30942 13582 30994
rect 13634 30942 13636 30994
rect 13580 30436 13636 30942
rect 13692 30996 13748 32284
rect 13692 30930 13748 30940
rect 13916 32452 13972 32462
rect 13580 30370 13636 30380
rect 13804 30324 13860 30334
rect 13692 30212 13748 30222
rect 13692 30118 13748 30156
rect 13692 29540 13748 29550
rect 13804 29540 13860 30268
rect 13916 30322 13972 32396
rect 14140 31444 14196 33964
rect 14364 33236 14420 34188
rect 14364 33170 14420 33180
rect 14476 33908 14532 34636
rect 14364 31892 14420 31902
rect 14364 31798 14420 31836
rect 14252 31778 14308 31790
rect 14252 31726 14254 31778
rect 14306 31726 14308 31778
rect 14252 31668 14308 31726
rect 14252 31602 14308 31612
rect 14140 31388 14308 31444
rect 13916 30270 13918 30322
rect 13970 30270 13972 30322
rect 13916 30258 13972 30270
rect 14252 30098 14308 31388
rect 14252 30046 14254 30098
rect 14306 30046 14308 30098
rect 13692 29538 14084 29540
rect 13692 29486 13694 29538
rect 13746 29486 14084 29538
rect 13692 29484 14084 29486
rect 13692 29474 13748 29484
rect 12908 27970 13300 27972
rect 12908 27918 12910 27970
rect 12962 27918 13300 27970
rect 12908 27916 13300 27918
rect 13916 29316 13972 29326
rect 12908 27906 12964 27916
rect 12124 27234 12180 27244
rect 13804 27300 13860 27310
rect 13804 27206 13860 27244
rect 13916 27186 13972 29260
rect 14028 27970 14084 29484
rect 14140 29428 14196 29438
rect 14140 28756 14196 29372
rect 14140 28662 14196 28700
rect 14028 27918 14030 27970
rect 14082 27918 14084 27970
rect 14028 27906 14084 27918
rect 13916 27134 13918 27186
rect 13970 27134 13972 27186
rect 13916 27122 13972 27134
rect 12124 27074 12180 27086
rect 12124 27022 12126 27074
rect 12178 27022 12180 27074
rect 11228 26852 11620 26908
rect 11788 26852 12068 26908
rect 10556 25340 11060 25396
rect 10556 24610 10612 25340
rect 10556 24558 10558 24610
rect 10610 24558 10612 24610
rect 10556 24546 10612 24558
rect 11004 24834 11060 24846
rect 11004 24782 11006 24834
rect 11058 24782 11060 24834
rect 11004 24052 11060 24782
rect 11452 24722 11508 24734
rect 11452 24670 11454 24722
rect 11506 24670 11508 24722
rect 10892 23996 11004 24052
rect 10892 23938 10948 23996
rect 11004 23986 11060 23996
rect 11340 24052 11396 24062
rect 10892 23886 10894 23938
rect 10946 23886 10948 23938
rect 10892 23874 10948 23886
rect 10220 23378 10388 23380
rect 10220 23326 10222 23378
rect 10274 23326 10388 23378
rect 10220 23324 10388 23326
rect 10220 23314 10276 23324
rect 11228 23266 11284 23278
rect 11228 23214 11230 23266
rect 11282 23214 11284 23266
rect 11228 23156 11284 23214
rect 10444 23042 10500 23054
rect 10444 22990 10446 23042
rect 10498 22990 10500 23042
rect 10332 22260 10388 22270
rect 10332 22166 10388 22204
rect 10332 22036 10388 22046
rect 10332 21474 10388 21980
rect 10444 21700 10500 22990
rect 11116 22596 11172 22606
rect 11116 22482 11172 22540
rect 11116 22430 11118 22482
rect 11170 22430 11172 22482
rect 11004 22148 11060 22158
rect 10892 21812 10948 21822
rect 11004 21812 11060 22092
rect 11116 22036 11172 22430
rect 11228 22260 11284 23100
rect 11228 22194 11284 22204
rect 11116 21970 11172 21980
rect 10892 21810 11060 21812
rect 10892 21758 10894 21810
rect 10946 21758 11060 21810
rect 10892 21756 11060 21758
rect 10500 21644 10612 21700
rect 10444 21634 10500 21644
rect 10332 21422 10334 21474
rect 10386 21422 10388 21474
rect 10332 21410 10388 21422
rect 10108 21196 10500 21252
rect 9996 20850 10052 20860
rect 9548 20132 9604 20636
rect 9772 20244 9828 20254
rect 9660 20132 9716 20142
rect 9548 20130 9716 20132
rect 9548 20078 9662 20130
rect 9714 20078 9716 20130
rect 9548 20076 9716 20078
rect 9660 20066 9716 20076
rect 9772 20132 9828 20188
rect 9772 20130 10052 20132
rect 9772 20078 9774 20130
rect 9826 20078 10052 20130
rect 9772 20076 10052 20078
rect 9772 20066 9828 20076
rect 8652 20020 8708 20030
rect 6748 19458 6804 19740
rect 6748 19406 6750 19458
rect 6802 19406 6804 19458
rect 6748 19394 6804 19406
rect 7868 19906 7924 19918
rect 7868 19854 7870 19906
rect 7922 19854 7924 19906
rect 7868 19348 7924 19854
rect 7868 19282 7924 19292
rect 8316 19346 8372 19358
rect 8316 19294 8318 19346
rect 8370 19294 8372 19346
rect 7308 19236 7364 19246
rect 7308 19142 7364 19180
rect 8316 19236 8372 19294
rect 8316 19170 8372 19180
rect 8652 18676 8708 19964
rect 9772 19796 9828 19806
rect 9772 19702 9828 19740
rect 9548 19124 9604 19134
rect 8876 18676 8932 18686
rect 8652 18620 8876 18676
rect 8876 18582 8932 18620
rect 9548 17666 9604 19068
rect 9996 17778 10052 20076
rect 10444 20130 10500 21196
rect 10444 20078 10446 20130
rect 10498 20078 10500 20130
rect 10444 20066 10500 20078
rect 10556 20020 10612 21644
rect 10668 21698 10724 21710
rect 10668 21646 10670 21698
rect 10722 21646 10724 21698
rect 10668 21140 10724 21646
rect 10668 21074 10724 21084
rect 10780 21698 10836 21710
rect 10780 21646 10782 21698
rect 10834 21646 10836 21698
rect 10780 21028 10836 21646
rect 10780 20962 10836 20972
rect 10668 20914 10724 20926
rect 10668 20862 10670 20914
rect 10722 20862 10724 20914
rect 10668 20804 10724 20862
rect 10668 20738 10724 20748
rect 10668 20020 10724 20030
rect 10556 19964 10668 20020
rect 10668 19926 10724 19964
rect 10892 19684 10948 21756
rect 11116 21588 11172 21598
rect 11116 21494 11172 21532
rect 11116 21252 11172 21262
rect 11004 21196 11116 21252
rect 11004 20802 11060 21196
rect 11116 21186 11172 21196
rect 11004 20750 11006 20802
rect 11058 20750 11060 20802
rect 11004 20244 11060 20750
rect 11004 20178 11060 20188
rect 11340 19796 11396 23996
rect 11452 23604 11508 24670
rect 11564 23828 11620 26852
rect 11676 26516 11732 26526
rect 11676 26178 11732 26460
rect 11676 26126 11678 26178
rect 11730 26126 11732 26178
rect 11676 26114 11732 26126
rect 11788 25508 11844 25518
rect 11788 25414 11844 25452
rect 11564 23826 11732 23828
rect 11564 23774 11566 23826
rect 11618 23774 11732 23826
rect 11564 23772 11732 23774
rect 11564 23762 11620 23772
rect 11508 23548 11620 23604
rect 11452 23510 11508 23548
rect 11452 21588 11508 21598
rect 11452 21494 11508 21532
rect 11564 21476 11620 23548
rect 11676 22932 11732 23772
rect 12012 23714 12068 26852
rect 12124 24722 12180 27022
rect 13692 27074 13748 27086
rect 13692 27022 13694 27074
rect 13746 27022 13748 27074
rect 12124 24670 12126 24722
rect 12178 24670 12180 24722
rect 12124 23940 12180 24670
rect 12460 26962 12516 26974
rect 12460 26910 12462 26962
rect 12514 26910 12516 26962
rect 12124 23826 12180 23884
rect 12348 23940 12404 23950
rect 12348 23846 12404 23884
rect 12124 23774 12126 23826
rect 12178 23774 12180 23826
rect 12124 23762 12180 23774
rect 12012 23662 12014 23714
rect 12066 23662 12068 23714
rect 12012 23650 12068 23662
rect 11676 22866 11732 22876
rect 11788 23492 11844 23502
rect 11676 21700 11732 21710
rect 11676 21606 11732 21644
rect 11564 21420 11732 21476
rect 11452 21140 11508 21150
rect 11452 20020 11508 21084
rect 11564 20692 11620 20702
rect 11564 20598 11620 20636
rect 11676 20690 11732 21420
rect 11788 21474 11844 23436
rect 12124 23380 12180 23390
rect 12124 23154 12180 23324
rect 12124 23102 12126 23154
rect 12178 23102 12180 23154
rect 12124 23090 12180 23102
rect 12236 23268 12292 23278
rect 11788 21422 11790 21474
rect 11842 21422 11844 21474
rect 11788 21410 11844 21422
rect 11900 21586 11956 21598
rect 11900 21534 11902 21586
rect 11954 21534 11956 21586
rect 11900 20802 11956 21534
rect 12236 21586 12292 23212
rect 12460 22372 12516 26910
rect 12908 26962 12964 26974
rect 12908 26910 12910 26962
rect 12962 26910 12964 26962
rect 12908 26908 12964 26910
rect 13692 26908 13748 27022
rect 12908 26852 13188 26908
rect 12908 26404 12964 26414
rect 12796 25508 12852 25518
rect 12572 25506 12852 25508
rect 12572 25454 12798 25506
rect 12850 25454 12852 25506
rect 12572 25452 12852 25454
rect 12572 23380 12628 25452
rect 12796 25442 12852 25452
rect 12796 24164 12852 24174
rect 12796 24070 12852 24108
rect 12684 23938 12740 23950
rect 12684 23886 12686 23938
rect 12738 23886 12740 23938
rect 12684 23604 12740 23886
rect 12796 23828 12852 23838
rect 12908 23828 12964 26348
rect 12796 23826 12964 23828
rect 12796 23774 12798 23826
rect 12850 23774 12964 23826
rect 12796 23772 12964 23774
rect 13132 26292 13188 26852
rect 13132 24722 13188 26236
rect 13132 24670 13134 24722
rect 13186 24670 13188 24722
rect 12796 23762 12852 23772
rect 12684 23538 12740 23548
rect 12796 23380 12852 23390
rect 12572 23324 12740 23380
rect 12684 23266 12740 23324
rect 12684 23214 12686 23266
rect 12738 23214 12740 23266
rect 12572 23156 12628 23166
rect 12572 23062 12628 23100
rect 12684 23044 12740 23214
rect 12684 22978 12740 22988
rect 12684 22372 12740 22382
rect 12460 22370 12740 22372
rect 12460 22318 12686 22370
rect 12738 22318 12740 22370
rect 12460 22316 12740 22318
rect 12348 22260 12404 22270
rect 12348 22166 12404 22204
rect 12236 21534 12238 21586
rect 12290 21534 12292 21586
rect 12236 21522 12292 21534
rect 12572 21698 12628 21710
rect 12572 21646 12574 21698
rect 12626 21646 12628 21698
rect 12572 21588 12628 21646
rect 12572 21364 12628 21532
rect 11900 20750 11902 20802
rect 11954 20750 11956 20802
rect 11900 20738 11956 20750
rect 12236 21308 12628 21364
rect 11676 20638 11678 20690
rect 11730 20638 11732 20690
rect 11676 20626 11732 20638
rect 11676 20356 11732 20366
rect 11452 20018 11620 20020
rect 11452 19966 11454 20018
rect 11506 19966 11620 20018
rect 11452 19964 11620 19966
rect 11452 19954 11508 19964
rect 10892 19618 10948 19628
rect 11004 19740 11396 19796
rect 10220 19236 10276 19246
rect 10220 18450 10276 19180
rect 10556 19124 10612 19134
rect 10556 19122 10724 19124
rect 10556 19070 10558 19122
rect 10610 19070 10724 19122
rect 10556 19068 10724 19070
rect 10556 19058 10612 19068
rect 10220 18398 10222 18450
rect 10274 18398 10276 18450
rect 10220 18386 10276 18398
rect 9996 17726 9998 17778
rect 10050 17726 10052 17778
rect 9996 17714 10052 17726
rect 10668 17778 10724 19068
rect 10892 18452 10948 18462
rect 11004 18452 11060 19740
rect 11452 19684 11508 19694
rect 11340 19628 11452 19684
rect 10892 18450 11060 18452
rect 10892 18398 10894 18450
rect 10946 18398 11060 18450
rect 10892 18396 11060 18398
rect 11116 19012 11172 19022
rect 10892 18386 10948 18396
rect 10668 17726 10670 17778
rect 10722 17726 10724 17778
rect 10668 17714 10724 17726
rect 9548 17614 9550 17666
rect 9602 17614 9604 17666
rect 9548 17602 9604 17614
rect 10892 17668 10948 17678
rect 10892 17574 10948 17612
rect 11116 17666 11172 18956
rect 11340 17780 11396 19628
rect 11452 19618 11508 19628
rect 11452 19234 11508 19246
rect 11452 19182 11454 19234
rect 11506 19182 11508 19234
rect 11452 18676 11508 19182
rect 11564 19236 11620 19964
rect 11676 20018 11732 20300
rect 11900 20132 11956 20142
rect 11676 19966 11678 20018
rect 11730 19966 11732 20018
rect 11676 19954 11732 19966
rect 11788 20130 11956 20132
rect 11788 20078 11902 20130
rect 11954 20078 11956 20130
rect 11788 20076 11956 20078
rect 11676 19236 11732 19246
rect 11564 19234 11732 19236
rect 11564 19182 11678 19234
rect 11730 19182 11732 19234
rect 11564 19180 11732 19182
rect 11676 19170 11732 19180
rect 11452 18452 11508 18620
rect 11788 19124 11844 20076
rect 11900 20066 11956 20076
rect 12012 20132 12068 20142
rect 12012 20038 12068 20076
rect 12124 20020 12180 20030
rect 12236 20020 12292 21308
rect 12684 20804 12740 22316
rect 12796 22258 12852 23324
rect 12796 22206 12798 22258
rect 12850 22206 12852 22258
rect 12796 22194 12852 22206
rect 12908 22484 12964 22494
rect 12908 21810 12964 22428
rect 13132 22372 13188 24670
rect 13132 22306 13188 22316
rect 13244 26852 13748 26908
rect 13916 26964 13972 26974
rect 13020 22148 13076 22158
rect 13244 22148 13300 26852
rect 13692 25508 13748 25518
rect 13692 25414 13748 25452
rect 13804 25394 13860 25406
rect 13804 25342 13806 25394
rect 13858 25342 13860 25394
rect 13804 25284 13860 25342
rect 13804 25218 13860 25228
rect 13804 24612 13860 24622
rect 13804 24518 13860 24556
rect 13692 24276 13748 24286
rect 13692 24052 13748 24220
rect 13020 22146 13300 22148
rect 13020 22094 13022 22146
rect 13074 22094 13300 22146
rect 13020 22092 13300 22094
rect 13356 23996 13748 24052
rect 13020 22082 13076 22092
rect 13356 22036 13412 23996
rect 13692 23826 13748 23996
rect 13692 23774 13694 23826
rect 13746 23774 13748 23826
rect 13692 23762 13748 23774
rect 13916 23826 13972 26908
rect 14252 26404 14308 30046
rect 14476 29652 14532 33852
rect 15036 33796 15092 34750
rect 15036 33730 15092 33740
rect 15148 34690 15204 34702
rect 15148 34638 15150 34690
rect 15202 34638 15204 34690
rect 15148 33684 15204 34638
rect 15260 34580 15316 34972
rect 15372 34804 15428 34814
rect 15372 34710 15428 34748
rect 15260 34524 15428 34580
rect 15260 34132 15316 34142
rect 15260 34038 15316 34076
rect 15148 33618 15204 33628
rect 15260 33348 15316 33358
rect 15148 33122 15204 33134
rect 15148 33070 15150 33122
rect 15202 33070 15204 33122
rect 14700 32676 14756 32686
rect 14588 31780 14644 31790
rect 14588 31106 14644 31724
rect 14588 31054 14590 31106
rect 14642 31054 14644 31106
rect 14588 31042 14644 31054
rect 14700 30548 14756 32620
rect 14924 32562 14980 32574
rect 14924 32510 14926 32562
rect 14978 32510 14980 32562
rect 14924 31780 14980 32510
rect 15148 32564 15204 33070
rect 15148 32498 15204 32508
rect 15036 31780 15092 31790
rect 14924 31778 15092 31780
rect 14924 31726 15038 31778
rect 15090 31726 15092 31778
rect 14924 31724 15092 31726
rect 14924 31444 14980 31454
rect 14924 31108 14980 31388
rect 15036 31332 15092 31724
rect 15036 31266 15092 31276
rect 15036 31108 15092 31118
rect 14924 31106 15092 31108
rect 14924 31054 15038 31106
rect 15090 31054 15092 31106
rect 14924 31052 15092 31054
rect 14588 30492 14756 30548
rect 14588 30210 14644 30492
rect 14588 30158 14590 30210
rect 14642 30158 14644 30210
rect 14588 29988 14644 30158
rect 14588 29922 14644 29932
rect 14700 30324 14756 30334
rect 14588 29652 14644 29662
rect 14476 29650 14644 29652
rect 14476 29598 14590 29650
rect 14642 29598 14644 29650
rect 14476 29596 14644 29598
rect 14588 29586 14644 29596
rect 14700 29652 14756 30268
rect 14924 30100 14980 30110
rect 14924 30006 14980 30044
rect 14700 29428 14756 29596
rect 14700 29426 14868 29428
rect 14700 29374 14702 29426
rect 14754 29374 14868 29426
rect 14700 29372 14868 29374
rect 14700 29362 14756 29372
rect 14476 29092 14532 29102
rect 14476 27074 14532 29036
rect 14476 27022 14478 27074
rect 14530 27022 14532 27074
rect 14476 27010 14532 27022
rect 14700 28420 14756 28430
rect 14700 27074 14756 28364
rect 14700 27022 14702 27074
rect 14754 27022 14756 27074
rect 14700 27010 14756 27022
rect 14308 26348 14420 26404
rect 14252 26338 14308 26348
rect 14028 26180 14084 26190
rect 14364 26180 14420 26348
rect 14700 26292 14756 26302
rect 14700 26198 14756 26236
rect 14028 26178 14308 26180
rect 14028 26126 14030 26178
rect 14082 26126 14308 26178
rect 14028 26124 14308 26126
rect 14028 26114 14084 26124
rect 14028 25506 14084 25518
rect 14028 25454 14030 25506
rect 14082 25454 14084 25506
rect 14028 23940 14084 25454
rect 14140 24052 14196 24062
rect 14252 24052 14308 26124
rect 14364 26114 14420 26124
rect 14812 26068 14868 29372
rect 14924 29316 14980 29326
rect 14924 27858 14980 29260
rect 15036 28082 15092 31052
rect 15148 31106 15204 31118
rect 15148 31054 15150 31106
rect 15202 31054 15204 31106
rect 15148 30884 15204 31054
rect 15148 30818 15204 30828
rect 15260 29988 15316 33292
rect 15372 32338 15428 34524
rect 15372 32286 15374 32338
rect 15426 32286 15428 32338
rect 15372 32274 15428 32286
rect 15484 32228 15540 35420
rect 15708 34914 15764 35868
rect 15820 35698 15876 35710
rect 15820 35646 15822 35698
rect 15874 35646 15876 35698
rect 15820 35588 15876 35646
rect 15820 35522 15876 35532
rect 15708 34862 15710 34914
rect 15762 34862 15764 34914
rect 15708 34850 15764 34862
rect 16156 35252 16212 37436
rect 15596 34692 15652 34702
rect 15596 34242 15652 34636
rect 15596 34190 15598 34242
rect 15650 34190 15652 34242
rect 15596 34178 15652 34190
rect 15708 34356 15764 34366
rect 15708 34130 15764 34300
rect 16156 34356 16212 35196
rect 16156 34290 16212 34300
rect 16268 37266 16324 37278
rect 16268 37214 16270 37266
rect 16322 37214 16324 37266
rect 16268 34692 16324 37214
rect 16604 36932 16660 37996
rect 16716 37380 16772 37390
rect 16716 37154 16772 37324
rect 16716 37102 16718 37154
rect 16770 37102 16772 37154
rect 16716 37090 16772 37102
rect 16828 37044 16884 38892
rect 16828 36978 16884 36988
rect 16604 36866 16660 36876
rect 16940 36932 16996 46620
rect 17276 43092 17332 50372
rect 17500 49028 17556 49038
rect 17500 48914 17556 48972
rect 17500 48862 17502 48914
rect 17554 48862 17556 48914
rect 17500 48850 17556 48862
rect 17388 48802 17444 48814
rect 17388 48750 17390 48802
rect 17442 48750 17444 48802
rect 17388 47572 17444 48750
rect 17500 48244 17556 48254
rect 17612 48244 17668 50372
rect 18396 50370 18564 50372
rect 18396 50318 18510 50370
rect 18562 50318 18564 50370
rect 18396 50316 18564 50318
rect 18060 48916 18116 48926
rect 18060 48822 18116 48860
rect 18284 48914 18340 48926
rect 18284 48862 18286 48914
rect 18338 48862 18340 48914
rect 18284 48804 18340 48862
rect 18284 48738 18340 48748
rect 17500 48242 17668 48244
rect 17500 48190 17502 48242
rect 17554 48190 17668 48242
rect 17500 48188 17668 48190
rect 17500 48178 17556 48188
rect 17612 48020 17668 48188
rect 17612 47954 17668 47964
rect 18172 48130 18228 48142
rect 18172 48078 18174 48130
rect 18226 48078 18228 48130
rect 18172 47684 18228 48078
rect 18284 47684 18340 47694
rect 18172 47682 18340 47684
rect 18172 47630 18286 47682
rect 18338 47630 18340 47682
rect 18172 47628 18340 47630
rect 18284 47618 18340 47628
rect 17388 47506 17444 47516
rect 18284 47460 18340 47470
rect 18396 47460 18452 50316
rect 18508 50306 18564 50316
rect 18508 49140 18564 49150
rect 18620 49140 18676 53116
rect 19292 53106 19348 53116
rect 19628 55020 19908 55076
rect 22204 55074 22260 55086
rect 22204 55022 22206 55074
rect 22258 55022 22260 55074
rect 19628 52946 19684 55020
rect 19836 54908 20100 54918
rect 19892 54852 19940 54908
rect 19996 54852 20044 54908
rect 19836 54842 20100 54852
rect 22204 54516 22260 55022
rect 22316 54740 22372 55134
rect 22540 55076 22596 55086
rect 22540 54982 22596 55020
rect 22652 55076 22708 55086
rect 22988 55076 23044 55356
rect 23212 55300 23268 55356
rect 23884 55356 24052 55412
rect 25788 55412 25844 55422
rect 23436 55300 23492 55310
rect 23212 55298 23492 55300
rect 23212 55246 23438 55298
rect 23490 55246 23492 55298
rect 23212 55244 23492 55246
rect 22652 55074 23044 55076
rect 22652 55022 22654 55074
rect 22706 55022 23044 55074
rect 22652 55020 23044 55022
rect 23100 55186 23156 55198
rect 23100 55134 23102 55186
rect 23154 55134 23156 55186
rect 22652 55010 22708 55020
rect 22316 54684 22708 54740
rect 22092 54460 22260 54516
rect 22540 54514 22596 54526
rect 22540 54462 22542 54514
rect 22594 54462 22596 54514
rect 19852 54402 19908 54414
rect 19852 54350 19854 54402
rect 19906 54350 19908 54402
rect 19852 53956 19908 54350
rect 19852 53890 19908 53900
rect 21868 54404 21924 54414
rect 21868 53842 21924 54348
rect 21980 54402 22036 54414
rect 21980 54350 21982 54402
rect 22034 54350 22036 54402
rect 21980 54292 22036 54350
rect 22092 54292 22148 54460
rect 22540 54292 22596 54462
rect 21980 54236 22596 54292
rect 21868 53790 21870 53842
rect 21922 53790 21924 53842
rect 21868 53778 21924 53790
rect 22204 54068 22260 54078
rect 22204 53730 22260 54012
rect 22204 53678 22206 53730
rect 22258 53678 22260 53730
rect 22204 53666 22260 53678
rect 21644 53620 21700 53630
rect 20972 53508 21028 53518
rect 19836 53340 20100 53350
rect 19892 53284 19940 53340
rect 19996 53284 20044 53340
rect 19836 53274 20100 53284
rect 20524 53172 20580 53182
rect 20524 53078 20580 53116
rect 19628 52894 19630 52946
rect 19682 52894 19684 52946
rect 19628 52882 19684 52894
rect 19628 52220 20132 52276
rect 19628 52164 19684 52220
rect 19292 52108 19684 52164
rect 18732 51268 18788 51278
rect 18732 50818 18788 51212
rect 18732 50766 18734 50818
rect 18786 50766 18788 50818
rect 18732 50754 18788 50766
rect 19180 51044 19236 51054
rect 19180 50706 19236 50988
rect 19292 50818 19348 52108
rect 19628 52050 19684 52108
rect 20076 52162 20132 52220
rect 20076 52110 20078 52162
rect 20130 52110 20132 52162
rect 20076 52098 20132 52110
rect 19628 51998 19630 52050
rect 19682 51998 19684 52050
rect 19628 51986 19684 51998
rect 19740 52050 19796 52062
rect 19740 51998 19742 52050
rect 19794 51998 19796 52050
rect 19292 50766 19294 50818
rect 19346 50766 19348 50818
rect 19292 50754 19348 50766
rect 19404 51938 19460 51950
rect 19404 51886 19406 51938
rect 19458 51886 19460 51938
rect 19180 50654 19182 50706
rect 19234 50654 19236 50706
rect 19180 50642 19236 50654
rect 19404 50596 19460 51886
rect 19740 51940 19796 51998
rect 20412 52050 20468 52062
rect 20412 51998 20414 52050
rect 20466 51998 20468 52050
rect 19740 51874 19796 51884
rect 20300 51938 20356 51950
rect 20300 51886 20302 51938
rect 20354 51886 20356 51938
rect 19836 51772 20100 51782
rect 19892 51716 19940 51772
rect 19996 51716 20044 51772
rect 19836 51706 20100 51716
rect 20076 51492 20132 51502
rect 20300 51492 20356 51886
rect 20412 51940 20468 51998
rect 20412 51874 20468 51884
rect 20860 51492 20916 51502
rect 20300 51436 20580 51492
rect 19628 50596 19684 50606
rect 19404 50594 19684 50596
rect 19404 50542 19630 50594
rect 19682 50542 19684 50594
rect 19404 50540 19684 50542
rect 19628 50530 19684 50540
rect 20076 50482 20132 51436
rect 20300 51266 20356 51278
rect 20300 51214 20302 51266
rect 20354 51214 20356 51266
rect 20300 51044 20356 51214
rect 20300 50978 20356 50988
rect 20524 50594 20580 51436
rect 20860 51398 20916 51436
rect 20636 51268 20692 51278
rect 20636 51174 20692 51212
rect 20524 50542 20526 50594
rect 20578 50542 20580 50594
rect 20524 50530 20580 50542
rect 20076 50430 20078 50482
rect 20130 50430 20132 50482
rect 20076 50428 20132 50430
rect 18508 49138 18676 49140
rect 18508 49086 18510 49138
rect 18562 49086 18676 49138
rect 18508 49084 18676 49086
rect 18732 50372 18788 50382
rect 18508 49074 18564 49084
rect 18732 49028 18788 50316
rect 18732 48934 18788 48972
rect 19404 50372 20132 50428
rect 20524 50372 20580 50382
rect 18620 48132 18676 48142
rect 18620 47682 18676 48076
rect 18620 47630 18622 47682
rect 18674 47630 18676 47682
rect 18620 47618 18676 47630
rect 18284 47458 18452 47460
rect 18284 47406 18286 47458
rect 18338 47406 18452 47458
rect 18284 47404 18452 47406
rect 17388 47234 17444 47246
rect 17388 47182 17390 47234
rect 17442 47182 17444 47234
rect 17388 47124 17444 47182
rect 17388 46002 17444 47068
rect 17388 45950 17390 46002
rect 17442 45950 17444 46002
rect 17388 45938 17444 45950
rect 17724 46788 17780 46798
rect 18284 46788 18340 47404
rect 19404 47346 19460 50372
rect 20524 50278 20580 50316
rect 19836 50204 20100 50214
rect 19892 50148 19940 50204
rect 19996 50148 20044 50204
rect 19836 50138 20100 50148
rect 19628 49138 19684 49150
rect 19628 49086 19630 49138
rect 19682 49086 19684 49138
rect 19628 47570 19684 49086
rect 19964 48916 20020 48926
rect 20300 48916 20356 48926
rect 19964 48914 20300 48916
rect 19964 48862 19966 48914
rect 20018 48862 20300 48914
rect 19964 48860 20300 48862
rect 19964 48850 20020 48860
rect 19740 48804 19796 48842
rect 20300 48822 20356 48860
rect 19740 48738 19796 48748
rect 20412 48804 20468 48814
rect 20636 48804 20692 48814
rect 19836 48636 20100 48646
rect 19892 48580 19940 48636
rect 19996 48580 20044 48636
rect 19836 48570 20100 48580
rect 20300 48356 20356 48366
rect 20412 48356 20468 48748
rect 20356 48300 20468 48356
rect 20524 48802 20692 48804
rect 20524 48750 20638 48802
rect 20690 48750 20692 48802
rect 20524 48748 20692 48750
rect 20300 48130 20356 48300
rect 20300 48078 20302 48130
rect 20354 48078 20356 48130
rect 20300 48066 20356 48078
rect 19628 47518 19630 47570
rect 19682 47518 19684 47570
rect 19628 47506 19684 47518
rect 20076 47460 20132 47470
rect 20132 47404 20244 47460
rect 20076 47366 20132 47404
rect 19404 47294 19406 47346
rect 19458 47294 19460 47346
rect 19404 47282 19460 47294
rect 19836 47068 20100 47078
rect 19892 47012 19940 47068
rect 19996 47012 20044 47068
rect 19836 47002 20100 47012
rect 20188 46900 20244 47404
rect 20524 47458 20580 48748
rect 20636 48738 20692 48748
rect 20860 48354 20916 48366
rect 20860 48302 20862 48354
rect 20914 48302 20916 48354
rect 20636 48132 20692 48142
rect 20636 48038 20692 48076
rect 20524 47406 20526 47458
rect 20578 47406 20580 47458
rect 20524 47394 20580 47406
rect 20860 47460 20916 48302
rect 20860 47394 20916 47404
rect 20076 46844 20244 46900
rect 20972 46900 21028 53452
rect 21644 53506 21700 53564
rect 22092 53620 22148 53630
rect 22092 53526 22148 53564
rect 22428 53620 22484 53630
rect 22540 53620 22596 54236
rect 22428 53618 22596 53620
rect 22428 53566 22430 53618
rect 22482 53566 22596 53618
rect 22428 53564 22596 53566
rect 22652 54402 22708 54684
rect 22652 54350 22654 54402
rect 22706 54350 22708 54402
rect 22428 53554 22484 53564
rect 21644 53454 21646 53506
rect 21698 53454 21700 53506
rect 21644 52612 21700 53454
rect 22652 53506 22708 54350
rect 22988 53956 23044 53966
rect 22988 53862 23044 53900
rect 23100 53844 23156 55134
rect 23100 53732 23156 53788
rect 22652 53454 22654 53506
rect 22706 53454 22708 53506
rect 22540 53172 22596 53182
rect 22316 53170 22596 53172
rect 22316 53118 22542 53170
rect 22594 53118 22596 53170
rect 22316 53116 22596 53118
rect 21644 52546 21700 52556
rect 21756 52948 21812 52958
rect 21308 51940 21364 51950
rect 21308 51604 21364 51884
rect 21644 51940 21700 51950
rect 21644 51846 21700 51884
rect 21196 50820 21252 50830
rect 17724 46786 18340 46788
rect 17724 46734 17726 46786
rect 17778 46734 18340 46786
rect 17724 46732 18340 46734
rect 18396 46786 18452 46798
rect 18396 46734 18398 46786
rect 18450 46734 18452 46786
rect 17500 45106 17556 45118
rect 17500 45054 17502 45106
rect 17554 45054 17556 45106
rect 17500 44100 17556 45054
rect 17724 45108 17780 46732
rect 17836 46562 17892 46574
rect 17836 46510 17838 46562
rect 17890 46510 17892 46562
rect 17836 45668 17892 46510
rect 17948 46452 18004 46462
rect 17948 46450 18340 46452
rect 17948 46398 17950 46450
rect 18002 46398 18340 46450
rect 17948 46396 18340 46398
rect 17948 46386 18004 46396
rect 17836 45612 18228 45668
rect 18172 45218 18228 45612
rect 18172 45166 18174 45218
rect 18226 45166 18228 45218
rect 18172 45154 18228 45166
rect 17724 45052 18116 45108
rect 17500 44034 17556 44044
rect 17948 44436 18004 44446
rect 17948 43538 18004 44380
rect 17948 43486 17950 43538
rect 18002 43486 18004 43538
rect 17948 43474 18004 43486
rect 17052 43036 17332 43092
rect 17052 40852 17108 43036
rect 17164 42866 17220 42878
rect 17164 42814 17166 42866
rect 17218 42814 17220 42866
rect 17164 41972 17220 42814
rect 17836 42084 17892 42094
rect 17612 42028 17836 42084
rect 17612 41972 17668 42028
rect 17836 41990 17892 42028
rect 17164 41916 17668 41972
rect 18060 41972 18116 45052
rect 18284 43764 18340 46396
rect 18396 45780 18452 46734
rect 19180 46786 19236 46798
rect 19180 46734 19182 46786
rect 19234 46734 19236 46786
rect 18508 46676 18564 46686
rect 18956 46676 19012 46686
rect 18508 46674 19012 46676
rect 18508 46622 18510 46674
rect 18562 46622 18958 46674
rect 19010 46622 19012 46674
rect 18508 46620 19012 46622
rect 18508 46610 18564 46620
rect 18956 46610 19012 46620
rect 18620 46452 18676 46462
rect 18620 46358 18676 46396
rect 18396 45714 18452 45724
rect 19180 45108 19236 46734
rect 19292 46452 19348 46462
rect 19292 46450 19684 46452
rect 19292 46398 19294 46450
rect 19346 46398 19684 46450
rect 19292 46396 19684 46398
rect 19292 46386 19348 46396
rect 19292 45892 19348 45902
rect 19292 45798 19348 45836
rect 19628 45890 19684 46396
rect 20076 46002 20132 46844
rect 20972 46834 21028 46844
rect 21084 48020 21140 48030
rect 20412 46674 20468 46686
rect 20412 46622 20414 46674
rect 20466 46622 20468 46674
rect 20076 45950 20078 46002
rect 20130 45950 20132 46002
rect 20076 45938 20132 45950
rect 20188 46452 20244 46462
rect 19628 45838 19630 45890
rect 19682 45838 19684 45890
rect 19628 45826 19684 45838
rect 20188 45890 20244 46396
rect 20188 45838 20190 45890
rect 20242 45838 20244 45890
rect 20188 45668 20244 45838
rect 20412 45892 20468 46622
rect 20188 45602 20244 45612
rect 20300 45780 20356 45790
rect 19836 45500 20100 45510
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 19836 45434 20100 45444
rect 18620 44436 18676 44446
rect 18620 44322 18676 44380
rect 18620 44270 18622 44322
rect 18674 44270 18676 44322
rect 18620 44258 18676 44270
rect 19180 44212 19236 45052
rect 20300 44996 20356 45724
rect 20412 45444 20468 45836
rect 20412 45378 20468 45388
rect 21084 46562 21140 47964
rect 21084 46510 21086 46562
rect 21138 46510 21140 46562
rect 21084 45108 21140 46510
rect 21196 45668 21252 50764
rect 21308 50594 21364 51548
rect 21308 50542 21310 50594
rect 21362 50542 21364 50594
rect 21308 50530 21364 50542
rect 21420 51156 21476 51166
rect 21420 50482 21476 51100
rect 21420 50430 21422 50482
rect 21474 50430 21476 50482
rect 21420 50418 21476 50430
rect 21644 50484 21700 50494
rect 21756 50484 21812 52892
rect 22316 52164 22372 53116
rect 22540 53106 22596 53116
rect 22428 52948 22484 52958
rect 22428 52854 22484 52892
rect 22652 52836 22708 53454
rect 22988 53676 23156 53732
rect 22988 53060 23044 53676
rect 23100 53508 23156 53518
rect 23100 53414 23156 53452
rect 23212 53170 23268 55244
rect 23436 55234 23492 55244
rect 23772 55188 23828 55226
rect 23772 55122 23828 55132
rect 23660 55076 23716 55114
rect 23660 55010 23716 55020
rect 23884 54964 23940 55356
rect 24108 55300 24164 55310
rect 23772 54908 23940 54964
rect 23996 55298 24164 55300
rect 23996 55246 24110 55298
rect 24162 55246 24164 55298
rect 23996 55244 24164 55246
rect 23436 54516 23492 54526
rect 23324 54292 23380 54302
rect 23324 53954 23380 54236
rect 23324 53902 23326 53954
rect 23378 53902 23380 53954
rect 23324 53890 23380 53902
rect 23212 53118 23214 53170
rect 23266 53118 23268 53170
rect 23212 53106 23268 53118
rect 23436 53170 23492 54460
rect 23772 53618 23828 54908
rect 23884 54516 23940 54526
rect 23884 54422 23940 54460
rect 23772 53566 23774 53618
rect 23826 53566 23828 53618
rect 23772 53554 23828 53566
rect 23436 53118 23438 53170
rect 23490 53118 23492 53170
rect 23436 53106 23492 53118
rect 23100 53060 23156 53070
rect 22988 53058 23156 53060
rect 22988 53006 23102 53058
rect 23154 53006 23156 53058
rect 22988 53004 23156 53006
rect 23100 52994 23156 53004
rect 22652 52780 23044 52836
rect 22540 52724 22596 52734
rect 22540 52722 22708 52724
rect 22540 52670 22542 52722
rect 22594 52670 22708 52722
rect 22540 52668 22708 52670
rect 22540 52658 22596 52668
rect 22652 52164 22708 52668
rect 22316 52162 22484 52164
rect 22316 52110 22318 52162
rect 22370 52110 22484 52162
rect 22316 52108 22484 52110
rect 22316 52098 22372 52108
rect 22092 51940 22148 51950
rect 21980 51604 22036 51614
rect 21980 51378 22036 51548
rect 21980 51326 21982 51378
rect 22034 51326 22036 51378
rect 21980 51314 22036 51326
rect 21868 51156 21924 51166
rect 21868 50706 21924 51100
rect 21868 50654 21870 50706
rect 21922 50654 21924 50706
rect 21868 50642 21924 50654
rect 21980 50932 22036 50942
rect 21644 50482 21812 50484
rect 21644 50430 21646 50482
rect 21698 50430 21812 50482
rect 21644 50428 21812 50430
rect 21644 50418 21700 50428
rect 21644 47460 21700 47470
rect 21644 47366 21700 47404
rect 21308 47346 21364 47358
rect 21308 47294 21310 47346
rect 21362 47294 21364 47346
rect 21308 46564 21364 47294
rect 21420 47234 21476 47246
rect 21420 47182 21422 47234
rect 21474 47182 21476 47234
rect 21420 46676 21476 47182
rect 21420 46610 21476 46620
rect 21308 46004 21364 46508
rect 21308 45938 21364 45948
rect 21868 45890 21924 45902
rect 21868 45838 21870 45890
rect 21922 45838 21924 45890
rect 21868 45780 21924 45838
rect 21196 45612 21364 45668
rect 21084 45042 21140 45052
rect 21196 45444 21252 45454
rect 21196 45330 21252 45388
rect 21196 45278 21198 45330
rect 21250 45278 21252 45330
rect 20748 44996 20804 45006
rect 20188 44994 20356 44996
rect 20188 44942 20302 44994
rect 20354 44942 20356 44994
rect 20188 44940 20356 44942
rect 19852 44546 19908 44558
rect 19852 44494 19854 44546
rect 19906 44494 19908 44546
rect 19852 44436 19908 44494
rect 19852 44342 19908 44380
rect 19292 44212 19348 44222
rect 19180 44156 19292 44212
rect 19292 44146 19348 44156
rect 18284 43698 18340 43708
rect 19404 44100 19460 44110
rect 19404 43428 19460 44044
rect 19836 43932 20100 43942
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 19836 43866 20100 43876
rect 20188 43652 20244 44940
rect 20300 44930 20356 44940
rect 20636 44994 20804 44996
rect 20636 44942 20750 44994
rect 20802 44942 20804 44994
rect 20636 44940 20804 44942
rect 20300 44100 20356 44110
rect 20636 44100 20692 44940
rect 20748 44930 20804 44940
rect 21196 44660 21252 45278
rect 20748 44604 21252 44660
rect 20748 44546 20804 44604
rect 20748 44494 20750 44546
rect 20802 44494 20804 44546
rect 20748 44434 20804 44494
rect 20748 44382 20750 44434
rect 20802 44382 20804 44434
rect 20748 44370 20804 44382
rect 20356 44044 20692 44100
rect 20748 44212 20804 44222
rect 20300 44006 20356 44044
rect 20188 43586 20244 43596
rect 20300 43764 20356 43774
rect 20300 43650 20356 43708
rect 20300 43598 20302 43650
rect 20354 43598 20356 43650
rect 20300 43586 20356 43598
rect 20748 43538 20804 44156
rect 20748 43486 20750 43538
rect 20802 43486 20804 43538
rect 20748 43474 20804 43486
rect 19628 43428 19684 43438
rect 19404 43426 19684 43428
rect 19404 43374 19630 43426
rect 19682 43374 19684 43426
rect 19404 43372 19684 43374
rect 19628 42756 19684 43372
rect 19964 42756 20020 42766
rect 19628 42754 20020 42756
rect 19628 42702 19966 42754
rect 20018 42702 20020 42754
rect 19628 42700 20020 42702
rect 18508 42644 18564 42654
rect 18508 42194 18564 42588
rect 19292 42644 19348 42654
rect 19292 42550 19348 42588
rect 18508 42142 18510 42194
rect 18562 42142 18564 42194
rect 18508 42130 18564 42142
rect 19068 42084 19124 42094
rect 19068 41990 19124 42028
rect 18284 41972 18340 41982
rect 18060 41970 18340 41972
rect 18060 41918 18286 41970
rect 18338 41918 18340 41970
rect 18060 41916 18340 41918
rect 17388 41074 17444 41916
rect 17724 41858 17780 41870
rect 17724 41806 17726 41858
rect 17778 41806 17780 41858
rect 17612 41748 17668 41758
rect 17612 41186 17668 41692
rect 17612 41134 17614 41186
rect 17666 41134 17668 41186
rect 17612 41122 17668 41134
rect 17388 41022 17390 41074
rect 17442 41022 17444 41074
rect 17388 41010 17444 41022
rect 17052 40796 17444 40852
rect 17164 39394 17220 39406
rect 17164 39342 17166 39394
rect 17218 39342 17220 39394
rect 17164 39060 17220 39342
rect 17164 38994 17220 39004
rect 17388 38948 17444 40796
rect 17612 40516 17668 40526
rect 17612 40422 17668 40460
rect 17724 40402 17780 41806
rect 17948 41076 18004 41086
rect 17948 40404 18004 41020
rect 17724 40350 17726 40402
rect 17778 40350 17780 40402
rect 17724 40338 17780 40350
rect 17836 40402 18004 40404
rect 17836 40350 17950 40402
rect 18002 40350 18004 40402
rect 17836 40348 18004 40350
rect 17612 39396 17668 39406
rect 17612 39302 17668 39340
rect 17388 38834 17444 38892
rect 17388 38782 17390 38834
rect 17442 38782 17444 38834
rect 17388 38770 17444 38782
rect 17836 38274 17892 40348
rect 17948 40338 18004 40348
rect 17948 40068 18004 40078
rect 17948 39730 18004 40012
rect 17948 39678 17950 39730
rect 18002 39678 18004 39730
rect 17948 39284 18004 39678
rect 17948 39218 18004 39228
rect 17948 39060 18004 39070
rect 17948 38966 18004 39004
rect 18284 39058 18340 41916
rect 19180 41970 19236 41982
rect 19628 41972 19684 42700
rect 19964 42690 20020 42700
rect 20860 42756 20916 42766
rect 20860 42662 20916 42700
rect 20524 42644 20580 42654
rect 20524 42550 20580 42588
rect 20748 42644 20804 42654
rect 20636 42530 20692 42542
rect 20636 42478 20638 42530
rect 20690 42478 20692 42530
rect 19836 42364 20100 42374
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 19836 42298 20100 42308
rect 20524 42084 20580 42094
rect 19740 41972 19796 41982
rect 19180 41918 19182 41970
rect 19234 41918 19236 41970
rect 18620 41748 18676 41758
rect 18620 41746 18788 41748
rect 18620 41694 18622 41746
rect 18674 41694 18788 41746
rect 18620 41692 18788 41694
rect 18620 41682 18676 41692
rect 18396 41186 18452 41198
rect 18396 41134 18398 41186
rect 18450 41134 18452 41186
rect 18396 41076 18452 41134
rect 18396 41010 18452 41020
rect 18732 40962 18788 41692
rect 18732 40910 18734 40962
rect 18786 40910 18788 40962
rect 18732 40898 18788 40910
rect 19068 41746 19124 41758
rect 19068 41694 19070 41746
rect 19122 41694 19124 41746
rect 19068 40402 19124 41694
rect 19180 41748 19236 41918
rect 19180 40964 19236 41692
rect 19180 40898 19236 40908
rect 19404 41970 19796 41972
rect 19404 41918 19742 41970
rect 19794 41918 19796 41970
rect 19404 41916 19796 41918
rect 19068 40350 19070 40402
rect 19122 40350 19124 40402
rect 19068 40338 19124 40350
rect 19404 40404 19460 41916
rect 19740 41906 19796 41916
rect 20524 41970 20580 42028
rect 20524 41918 20526 41970
rect 20578 41918 20580 41970
rect 20524 41906 20580 41918
rect 20636 41972 20692 42478
rect 20636 41906 20692 41916
rect 19852 41188 19908 41198
rect 19516 41186 19908 41188
rect 19516 41134 19854 41186
rect 19906 41134 19908 41186
rect 19516 41132 19908 41134
rect 19516 40628 19572 41132
rect 19852 41122 19908 41132
rect 20524 41074 20580 41086
rect 20524 41022 20526 41074
rect 20578 41022 20580 41074
rect 19628 40964 19684 40974
rect 19628 40870 19684 40908
rect 20524 40964 20580 41022
rect 20636 41076 20692 41086
rect 20748 41076 20804 42588
rect 20636 41074 20804 41076
rect 20636 41022 20638 41074
rect 20690 41022 20804 41074
rect 20636 41020 20804 41022
rect 20636 41010 20692 41020
rect 20524 40898 20580 40908
rect 20860 40962 20916 40974
rect 20860 40910 20862 40962
rect 20914 40910 20916 40962
rect 19836 40796 20100 40806
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 19836 40730 20100 40740
rect 19516 40572 19684 40628
rect 19404 40338 19460 40348
rect 19516 40402 19572 40414
rect 19516 40350 19518 40402
rect 19570 40350 19572 40402
rect 19516 40068 19572 40350
rect 19516 40002 19572 40012
rect 19628 39844 19684 40572
rect 20860 40626 20916 40910
rect 21308 40628 21364 45612
rect 21756 45108 21812 45118
rect 21756 45014 21812 45052
rect 21868 44100 21924 45724
rect 21980 45556 22036 50876
rect 22092 50820 22148 51884
rect 22204 51490 22260 51502
rect 22204 51438 22206 51490
rect 22258 51438 22260 51490
rect 22204 51044 22260 51438
rect 22204 50978 22260 50988
rect 22092 50726 22148 50764
rect 22428 50818 22484 52108
rect 22652 52070 22708 52108
rect 22764 51938 22820 51950
rect 22764 51886 22766 51938
rect 22818 51886 22820 51938
rect 22540 51268 22596 51278
rect 22540 51044 22596 51212
rect 22764 51268 22820 51886
rect 22764 51202 22820 51212
rect 22876 51940 22932 51950
rect 22876 51044 22932 51884
rect 22540 50988 22932 51044
rect 22988 50932 23044 52780
rect 23772 52834 23828 52846
rect 23772 52782 23774 52834
rect 23826 52782 23828 52834
rect 23772 52722 23828 52782
rect 23772 52670 23774 52722
rect 23826 52670 23828 52722
rect 23324 52162 23380 52174
rect 23324 52110 23326 52162
rect 23378 52110 23380 52162
rect 23324 51940 23380 52110
rect 23548 52164 23604 52174
rect 23548 52070 23604 52108
rect 23324 51874 23380 51884
rect 23772 51380 23828 52670
rect 23996 52388 24052 55244
rect 24108 55234 24164 55244
rect 24892 55188 24948 55198
rect 25452 55188 25508 55198
rect 24892 55186 25172 55188
rect 24892 55134 24894 55186
rect 24946 55134 25172 55186
rect 24892 55132 25172 55134
rect 24892 55122 24948 55132
rect 24332 55076 24388 55086
rect 24108 54292 24164 54302
rect 24108 54198 24164 54236
rect 24220 53844 24276 53854
rect 24220 53750 24276 53788
rect 24332 53730 24388 55020
rect 25116 53842 25172 55132
rect 25116 53790 25118 53842
rect 25170 53790 25172 53842
rect 25116 53778 25172 53790
rect 25452 54402 25508 55132
rect 25788 55076 25844 55356
rect 27020 55412 27076 55422
rect 27020 55318 27076 55356
rect 27132 55300 27188 56030
rect 27188 55244 27412 55300
rect 27132 55234 27188 55244
rect 25788 54514 25844 55020
rect 27244 55074 27300 55086
rect 27244 55022 27246 55074
rect 27298 55022 27300 55074
rect 25788 54462 25790 54514
rect 25842 54462 25844 54514
rect 25788 54450 25844 54462
rect 27132 54516 27188 54526
rect 27132 54422 27188 54460
rect 25452 54350 25454 54402
rect 25506 54350 25508 54402
rect 24332 53678 24334 53730
rect 24386 53678 24388 53730
rect 24332 53666 24388 53678
rect 24780 53732 24836 53742
rect 24780 53638 24836 53676
rect 25340 53732 25396 53742
rect 25340 53638 25396 53676
rect 25004 53618 25060 53630
rect 25004 53566 25006 53618
rect 25058 53566 25060 53618
rect 24108 53506 24164 53518
rect 24108 53454 24110 53506
rect 24162 53454 24164 53506
rect 24108 52948 24164 53454
rect 24220 53508 24276 53518
rect 24220 53172 24276 53452
rect 25004 53508 25060 53566
rect 25004 53442 25060 53452
rect 24220 53078 24276 53116
rect 25228 53172 25284 53182
rect 24108 52722 24164 52892
rect 24108 52670 24110 52722
rect 24162 52670 24164 52722
rect 24108 52658 24164 52670
rect 25228 52500 25284 53116
rect 25340 52948 25396 52958
rect 25452 52948 25508 54350
rect 26236 54402 26292 54414
rect 26236 54350 26238 54402
rect 26290 54350 26292 54402
rect 25564 53732 25620 53742
rect 26012 53732 26068 53742
rect 25564 53730 26068 53732
rect 25564 53678 25566 53730
rect 25618 53678 26014 53730
rect 26066 53678 26068 53730
rect 25564 53676 26068 53678
rect 25564 53666 25620 53676
rect 26012 53666 26068 53676
rect 26124 53732 26180 53742
rect 26124 53638 26180 53676
rect 25900 53508 25956 53518
rect 25900 53284 25956 53452
rect 26236 53284 26292 54350
rect 26908 54402 26964 54414
rect 26908 54350 26910 54402
rect 26962 54350 26964 54402
rect 26908 53732 26964 54350
rect 27244 54068 27300 55022
rect 27244 54002 27300 54012
rect 26908 53676 27188 53732
rect 27132 53620 27188 53676
rect 25900 53228 26292 53284
rect 26348 53506 26404 53518
rect 27020 53508 27076 53518
rect 26348 53454 26350 53506
rect 26402 53454 26404 53506
rect 25788 53172 25844 53182
rect 25788 53078 25844 53116
rect 25396 52892 25508 52948
rect 25340 52854 25396 52892
rect 24780 52444 25396 52500
rect 23996 52332 24164 52388
rect 23548 51378 23828 51380
rect 23548 51326 23774 51378
rect 23826 51326 23828 51378
rect 23548 51324 23828 51326
rect 22428 50766 22430 50818
rect 22482 50766 22484 50818
rect 22428 50754 22484 50766
rect 22652 50876 23044 50932
rect 23324 51268 23380 51278
rect 23548 51268 23604 51324
rect 23772 51314 23828 51324
rect 23324 51266 23604 51268
rect 23324 51214 23326 51266
rect 23378 51214 23604 51266
rect 23324 51212 23604 51214
rect 23324 50932 23380 51212
rect 23660 51156 23716 51166
rect 23660 51062 23716 51100
rect 22652 49922 22708 50876
rect 23324 50866 23380 50876
rect 23100 50596 23156 50606
rect 23100 50502 23156 50540
rect 23660 50594 23716 50606
rect 23660 50542 23662 50594
rect 23714 50542 23716 50594
rect 23660 50428 23716 50542
rect 23772 50596 23828 50634
rect 23772 50530 23828 50540
rect 24108 50594 24164 52332
rect 24220 52164 24276 52174
rect 24220 52070 24276 52108
rect 24108 50542 24110 50594
rect 24162 50542 24164 50594
rect 23884 50484 23940 50494
rect 23660 50372 23828 50428
rect 22652 49870 22654 49922
rect 22706 49870 22708 49922
rect 22540 49812 22596 49822
rect 22092 49810 22596 49812
rect 22092 49758 22542 49810
rect 22594 49758 22596 49810
rect 22092 49756 22596 49758
rect 22092 48468 22148 49756
rect 22540 49746 22596 49756
rect 22540 48916 22596 48926
rect 22652 48916 22708 49870
rect 22876 49924 22932 49934
rect 23436 49924 23492 49934
rect 22876 49922 23492 49924
rect 22876 49870 22878 49922
rect 22930 49870 23438 49922
rect 23490 49870 23492 49922
rect 22876 49868 23492 49870
rect 22876 49858 22932 49868
rect 23436 49858 23492 49868
rect 23772 49924 23828 50372
rect 23772 49858 23828 49868
rect 23884 49922 23940 50428
rect 23884 49870 23886 49922
rect 23938 49870 23940 49922
rect 23884 49858 23940 49870
rect 23996 49924 24052 49934
rect 23996 49830 24052 49868
rect 23548 49810 23604 49822
rect 23548 49758 23550 49810
rect 23602 49758 23604 49810
rect 23436 49700 23492 49710
rect 23436 49586 23492 49644
rect 23436 49534 23438 49586
rect 23490 49534 23492 49586
rect 23436 49522 23492 49534
rect 23548 49588 23604 49758
rect 23996 49588 24052 49598
rect 23548 49586 24052 49588
rect 23548 49534 23998 49586
rect 24050 49534 24052 49586
rect 23548 49532 24052 49534
rect 23996 49522 24052 49532
rect 24108 49028 24164 50542
rect 22540 48914 22708 48916
rect 22540 48862 22542 48914
rect 22594 48862 22708 48914
rect 22540 48860 22708 48862
rect 23996 48972 24164 49028
rect 24220 49924 24276 49934
rect 22540 48850 22596 48860
rect 22092 47346 22148 48412
rect 22764 48804 22820 48814
rect 22204 48356 22260 48366
rect 22204 48262 22260 48300
rect 22092 47294 22094 47346
rect 22146 47294 22148 47346
rect 22092 47282 22148 47294
rect 22428 48132 22484 48142
rect 22428 47234 22484 48076
rect 22764 48130 22820 48748
rect 22876 48804 22932 48814
rect 23436 48804 23492 48814
rect 22876 48802 23604 48804
rect 22876 48750 22878 48802
rect 22930 48750 23438 48802
rect 23490 48750 23604 48802
rect 22876 48748 23604 48750
rect 22876 48738 22932 48748
rect 23436 48738 23492 48748
rect 23548 48244 23604 48748
rect 23772 48244 23828 48254
rect 23548 48242 23828 48244
rect 23548 48190 23774 48242
rect 23826 48190 23828 48242
rect 23548 48188 23828 48190
rect 22764 48078 22766 48130
rect 22818 48078 22820 48130
rect 22764 48066 22820 48078
rect 23324 48132 23380 48142
rect 23324 48038 23380 48076
rect 23772 47796 23828 48188
rect 23996 48020 24052 48972
rect 23996 47954 24052 47964
rect 24108 48802 24164 48814
rect 24108 48750 24110 48802
rect 24162 48750 24164 48802
rect 24108 47796 24164 48750
rect 24220 48354 24276 49868
rect 24556 49028 24612 49038
rect 24444 49026 24612 49028
rect 24444 48974 24558 49026
rect 24610 48974 24612 49026
rect 24444 48972 24612 48974
rect 24332 48804 24388 48814
rect 24332 48710 24388 48748
rect 24220 48302 24222 48354
rect 24274 48302 24276 48354
rect 24220 48290 24276 48302
rect 23772 47740 24164 47796
rect 24444 48244 24500 48972
rect 24556 48962 24612 48972
rect 23548 47460 23604 47470
rect 23548 47366 23604 47404
rect 22428 47182 22430 47234
rect 22482 47182 22484 47234
rect 21980 45490 22036 45500
rect 22092 46002 22148 46014
rect 22092 45950 22094 46002
rect 22146 45950 22148 46002
rect 22092 45892 22148 45950
rect 21980 44100 22036 44110
rect 21868 44044 21980 44100
rect 21980 44034 22036 44044
rect 21868 43652 21924 43662
rect 21868 43558 21924 43596
rect 21756 42868 21812 42878
rect 21756 42774 21812 42812
rect 21980 42756 22036 42766
rect 21980 42662 22036 42700
rect 21420 42644 21476 42654
rect 21420 41300 21476 42588
rect 21644 42530 21700 42542
rect 21644 42478 21646 42530
rect 21698 42478 21700 42530
rect 21644 41972 21700 42478
rect 21420 41298 21588 41300
rect 21420 41246 21422 41298
rect 21474 41246 21588 41298
rect 21420 41244 21588 41246
rect 21420 41234 21476 41244
rect 21532 40628 21588 41244
rect 21644 41074 21700 41916
rect 21644 41022 21646 41074
rect 21698 41022 21700 41074
rect 21644 41010 21700 41022
rect 21644 40628 21700 40638
rect 20860 40574 20862 40626
rect 20914 40574 20916 40626
rect 20860 40562 20916 40574
rect 20972 40572 21252 40628
rect 21308 40572 21476 40628
rect 21532 40626 21700 40628
rect 21532 40574 21646 40626
rect 21698 40574 21700 40626
rect 21532 40572 21700 40574
rect 20412 40404 20468 40414
rect 20972 40404 21028 40572
rect 21196 40516 21252 40572
rect 21196 40460 21364 40516
rect 20412 40402 21028 40404
rect 20412 40350 20414 40402
rect 20466 40350 21028 40402
rect 20412 40348 21028 40350
rect 21084 40402 21140 40414
rect 21084 40350 21086 40402
rect 21138 40350 21140 40402
rect 20412 40338 20468 40348
rect 19404 39788 19684 39844
rect 19740 40290 19796 40302
rect 19740 40238 19742 40290
rect 19794 40238 19796 40290
rect 18284 39006 18286 39058
rect 18338 39006 18340 39058
rect 18284 38994 18340 39006
rect 18396 39506 18452 39518
rect 18396 39454 18398 39506
rect 18450 39454 18452 39506
rect 18396 38948 18452 39454
rect 18396 38882 18452 38892
rect 18508 39396 18564 39406
rect 18508 39060 18564 39340
rect 18508 39004 19012 39060
rect 18508 38834 18564 39004
rect 18844 38836 18900 38846
rect 18508 38782 18510 38834
rect 18562 38782 18564 38834
rect 18508 38770 18564 38782
rect 18732 38834 18900 38836
rect 18732 38782 18846 38834
rect 18898 38782 18900 38834
rect 18732 38780 18900 38782
rect 18732 38668 18788 38780
rect 18844 38770 18900 38780
rect 18956 38668 19012 39004
rect 17836 38222 17838 38274
rect 17890 38222 17892 38274
rect 17836 38210 17892 38222
rect 18396 38612 18788 38668
rect 18844 38612 19012 38668
rect 19068 38946 19124 38958
rect 19068 38894 19070 38946
rect 19122 38894 19124 38946
rect 18396 38162 18452 38612
rect 18396 38110 18398 38162
rect 18450 38110 18452 38162
rect 18396 38098 18452 38110
rect 16940 36866 16996 36876
rect 17164 38050 17220 38062
rect 17164 37998 17166 38050
rect 17218 37998 17220 38050
rect 16492 36708 16548 36718
rect 16380 36036 16436 36046
rect 16380 35026 16436 35980
rect 16492 35922 16548 36652
rect 16492 35870 16494 35922
rect 16546 35870 16548 35922
rect 16492 35812 16548 35870
rect 16716 35812 16772 35822
rect 16492 35746 16548 35756
rect 16604 35810 16772 35812
rect 16604 35758 16718 35810
rect 16770 35758 16772 35810
rect 16604 35756 16772 35758
rect 16380 34974 16382 35026
rect 16434 34974 16436 35026
rect 16380 34962 16436 34974
rect 15708 34078 15710 34130
rect 15762 34078 15764 34130
rect 15708 34066 15764 34078
rect 15932 34242 15988 34254
rect 15932 34190 15934 34242
rect 15986 34190 15988 34242
rect 15932 34132 15988 34190
rect 15484 32162 15540 32172
rect 15708 32228 15764 32238
rect 15372 32004 15428 32014
rect 15708 32004 15764 32172
rect 15372 31218 15428 31948
rect 15372 31166 15374 31218
rect 15426 31166 15428 31218
rect 15372 31154 15428 31166
rect 15484 31948 15764 32004
rect 15484 30212 15540 31948
rect 15932 31780 15988 34076
rect 16044 33236 16100 33246
rect 16044 32228 16100 33180
rect 16044 32162 16100 32172
rect 15932 31714 15988 31724
rect 16044 32004 16100 32014
rect 15708 31556 15764 31566
rect 16044 31556 16100 31948
rect 16156 31892 16212 31902
rect 16268 31892 16324 34636
rect 16604 33908 16660 35756
rect 16716 35746 16772 35756
rect 16828 35700 16884 35710
rect 16828 35698 16996 35700
rect 16828 35646 16830 35698
rect 16882 35646 16996 35698
rect 16828 35644 16996 35646
rect 16828 35634 16884 35644
rect 16940 35140 16996 35644
rect 17164 35476 17220 37998
rect 18172 38050 18228 38062
rect 18172 37998 18174 38050
rect 18226 37998 18228 38050
rect 17612 37940 17668 37950
rect 17388 36596 17444 36606
rect 17276 36482 17332 36494
rect 17276 36430 17278 36482
rect 17330 36430 17332 36482
rect 17276 36148 17332 36430
rect 17276 36082 17332 36092
rect 17388 35698 17444 36540
rect 17612 36370 17668 37884
rect 18172 37492 18228 37998
rect 18844 37828 18900 38612
rect 18844 37734 18900 37772
rect 19068 37604 19124 38894
rect 19180 38836 19236 38846
rect 19180 38164 19236 38780
rect 19404 38500 19460 39788
rect 19516 39620 19572 39630
rect 19740 39620 19796 40238
rect 20748 40180 20804 40190
rect 20076 39844 20132 39854
rect 20076 39730 20132 39788
rect 20748 39732 20804 40124
rect 20076 39678 20078 39730
rect 20130 39678 20132 39730
rect 20076 39666 20132 39678
rect 20412 39730 20804 39732
rect 20412 39678 20750 39730
rect 20802 39678 20804 39730
rect 20412 39676 20804 39678
rect 19516 39618 19796 39620
rect 19516 39566 19518 39618
rect 19570 39566 19796 39618
rect 19516 39564 19796 39566
rect 19516 39172 19572 39564
rect 19836 39228 20100 39238
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 19836 39162 20100 39172
rect 19516 39106 19572 39116
rect 19628 38948 19684 38958
rect 19628 38722 19684 38892
rect 20412 38834 20468 39676
rect 20748 39666 20804 39676
rect 21084 38948 21140 40350
rect 21308 40402 21364 40460
rect 21308 40350 21310 40402
rect 21362 40350 21364 40402
rect 21308 40338 21364 40350
rect 21196 40292 21252 40302
rect 21196 40198 21252 40236
rect 21420 40068 21476 40572
rect 21644 40562 21700 40572
rect 21980 40402 22036 40414
rect 21980 40350 21982 40402
rect 22034 40350 22036 40402
rect 21980 40180 22036 40350
rect 21980 40114 22036 40124
rect 21084 38882 21140 38892
rect 21196 40012 21476 40068
rect 20412 38782 20414 38834
rect 20466 38782 20468 38834
rect 20412 38770 20468 38782
rect 19628 38670 19630 38722
rect 19682 38670 19684 38722
rect 19628 38658 19684 38670
rect 19740 38722 19796 38734
rect 19740 38670 19742 38722
rect 19794 38670 19796 38722
rect 19740 38500 19796 38670
rect 19404 38444 19796 38500
rect 20076 38500 20132 38510
rect 19180 38098 19236 38108
rect 19292 38276 19348 38286
rect 19180 37940 19236 37950
rect 19180 37846 19236 37884
rect 19292 37938 19348 38220
rect 19292 37886 19294 37938
rect 19346 37886 19348 37938
rect 19292 37874 19348 37886
rect 18172 37426 18228 37436
rect 18844 37548 19124 37604
rect 17948 37268 18004 37278
rect 18284 37268 18340 37278
rect 17948 37266 18228 37268
rect 17948 37214 17950 37266
rect 18002 37214 18228 37266
rect 17948 37212 18228 37214
rect 17948 37202 18004 37212
rect 18172 37156 18228 37212
rect 18284 37174 18340 37212
rect 18396 37268 18452 37278
rect 18732 37268 18788 37278
rect 18396 37266 18788 37268
rect 18396 37214 18398 37266
rect 18450 37214 18734 37266
rect 18786 37214 18788 37266
rect 18396 37212 18788 37214
rect 18396 37202 18452 37212
rect 17612 36318 17614 36370
rect 17666 36318 17668 36370
rect 17500 35812 17556 35822
rect 17612 35812 17668 36318
rect 18060 37044 18116 37054
rect 18060 36596 18116 36988
rect 18060 36370 18116 36540
rect 18060 36318 18062 36370
rect 18114 36318 18116 36370
rect 18060 35924 18116 36318
rect 18172 36036 18228 37100
rect 18396 37044 18452 37054
rect 18284 36820 18340 36830
rect 18284 36482 18340 36764
rect 18396 36594 18452 36988
rect 18396 36542 18398 36594
rect 18450 36542 18452 36594
rect 18396 36530 18452 36542
rect 18284 36430 18286 36482
rect 18338 36430 18340 36482
rect 18284 36418 18340 36430
rect 18508 36482 18564 37212
rect 18732 37202 18788 37212
rect 18844 37156 18900 37548
rect 19404 37492 19460 38444
rect 19628 38164 19684 38174
rect 19068 37436 19460 37492
rect 19516 37826 19572 37838
rect 19516 37774 19518 37826
rect 19570 37774 19572 37826
rect 18844 37090 18900 37100
rect 18956 37154 19012 37166
rect 18956 37102 18958 37154
rect 19010 37102 19012 37154
rect 18844 36932 18900 36942
rect 18844 36594 18900 36876
rect 18844 36542 18846 36594
rect 18898 36542 18900 36594
rect 18844 36530 18900 36542
rect 18508 36430 18510 36482
rect 18562 36430 18564 36482
rect 18508 36418 18564 36430
rect 18956 36036 19012 37102
rect 18172 35980 18564 36036
rect 18060 35868 18340 35924
rect 17612 35756 18116 35812
rect 17500 35718 17556 35756
rect 17388 35646 17390 35698
rect 17442 35646 17444 35698
rect 17388 35634 17444 35646
rect 17500 35586 17556 35598
rect 17500 35534 17502 35586
rect 17554 35534 17556 35586
rect 17500 35476 17556 35534
rect 17164 35420 17556 35476
rect 16940 35084 18004 35140
rect 17276 34916 17332 34926
rect 16604 33842 16660 33852
rect 16716 34244 16772 34254
rect 16716 33796 16772 34188
rect 17276 34242 17332 34860
rect 17276 34190 17278 34242
rect 17330 34190 17332 34242
rect 17276 34178 17332 34190
rect 17836 34242 17892 34254
rect 17836 34190 17838 34242
rect 17890 34190 17892 34242
rect 17500 34130 17556 34142
rect 17500 34078 17502 34130
rect 17554 34078 17556 34130
rect 16716 33740 16996 33796
rect 16604 32562 16660 32574
rect 16604 32510 16606 32562
rect 16658 32510 16660 32562
rect 16492 32452 16548 32462
rect 16492 32358 16548 32396
rect 16156 31890 16324 31892
rect 16156 31838 16158 31890
rect 16210 31838 16324 31890
rect 16156 31836 16324 31838
rect 16156 31826 16212 31836
rect 16604 31780 16660 32510
rect 16940 31890 16996 33740
rect 17052 33348 17108 33358
rect 17052 32452 17108 33292
rect 17388 33346 17444 33358
rect 17388 33294 17390 33346
rect 17442 33294 17444 33346
rect 17388 32676 17444 33294
rect 17388 32610 17444 32620
rect 17164 32452 17220 32462
rect 17052 32396 17164 32452
rect 16940 31838 16942 31890
rect 16994 31838 16996 31890
rect 16940 31826 16996 31838
rect 16268 31666 16324 31678
rect 16268 31614 16270 31666
rect 16322 31614 16324 31666
rect 15708 31554 15988 31556
rect 15708 31502 15710 31554
rect 15762 31502 15988 31554
rect 15708 31500 15988 31502
rect 15708 31490 15764 31500
rect 15484 30118 15540 30156
rect 15820 30770 15876 30782
rect 15820 30718 15822 30770
rect 15874 30718 15876 30770
rect 15820 29988 15876 30718
rect 15932 30212 15988 31500
rect 16044 31554 16212 31556
rect 16044 31502 16046 31554
rect 16098 31502 16212 31554
rect 16044 31500 16212 31502
rect 16044 31490 16100 31500
rect 16044 30212 16100 30222
rect 15932 30156 16044 30212
rect 16044 30118 16100 30156
rect 15260 29932 15876 29988
rect 15036 28030 15038 28082
rect 15090 28030 15092 28082
rect 15036 28018 15092 28030
rect 14924 27806 14926 27858
rect 14978 27806 14980 27858
rect 14924 26516 14980 27806
rect 15260 27860 15316 27870
rect 15484 27860 15540 29932
rect 15260 27858 15540 27860
rect 15260 27806 15262 27858
rect 15314 27806 15540 27858
rect 15260 27804 15540 27806
rect 15596 29764 15652 29774
rect 15260 27794 15316 27804
rect 14924 26450 14980 26460
rect 15484 26962 15540 26974
rect 15484 26910 15486 26962
rect 15538 26910 15540 26962
rect 14812 26002 14868 26012
rect 15148 26290 15204 26302
rect 15148 26238 15150 26290
rect 15202 26238 15204 26290
rect 15148 25844 15204 26238
rect 14364 25394 14420 25406
rect 14364 25342 14366 25394
rect 14418 25342 14420 25394
rect 14364 25284 14420 25342
rect 14924 25396 14980 25406
rect 14924 25394 15092 25396
rect 14924 25342 14926 25394
rect 14978 25342 15092 25394
rect 14924 25340 15092 25342
rect 14924 25330 14980 25340
rect 14364 25218 14420 25228
rect 14700 24612 14756 24622
rect 14756 24556 14868 24612
rect 14700 24546 14756 24556
rect 14140 24050 14308 24052
rect 14140 23998 14142 24050
rect 14194 23998 14308 24050
rect 14140 23996 14308 23998
rect 14812 24050 14868 24556
rect 14812 23998 14814 24050
rect 14866 23998 14868 24050
rect 14140 23986 14196 23996
rect 14812 23986 14868 23998
rect 14924 24164 14980 24174
rect 14028 23874 14084 23884
rect 13916 23774 13918 23826
rect 13970 23774 13972 23826
rect 13916 23762 13972 23774
rect 14140 23828 14196 23838
rect 13580 23716 13636 23726
rect 13580 23548 13636 23660
rect 13468 23492 13636 23548
rect 14028 23716 14084 23726
rect 14140 23716 14196 23772
rect 14252 23828 14308 23838
rect 14252 23826 14532 23828
rect 14252 23774 14254 23826
rect 14306 23774 14532 23826
rect 14252 23772 14532 23774
rect 14252 23762 14308 23772
rect 14028 23714 14196 23716
rect 14028 23662 14030 23714
rect 14082 23662 14196 23714
rect 14028 23660 14196 23662
rect 14476 23716 14532 23772
rect 14924 23826 14980 24108
rect 14924 23774 14926 23826
rect 14978 23774 14980 23826
rect 14924 23762 14980 23774
rect 14588 23716 14644 23726
rect 14476 23714 14644 23716
rect 14476 23662 14590 23714
rect 14642 23662 14644 23714
rect 14476 23660 14644 23662
rect 13468 23156 13524 23492
rect 13468 23062 13524 23100
rect 13916 23154 13972 23166
rect 13916 23102 13918 23154
rect 13970 23102 13972 23154
rect 13916 22596 13972 23102
rect 13916 22530 13972 22540
rect 13580 22370 13636 22382
rect 13580 22318 13582 22370
rect 13634 22318 13636 22370
rect 13580 22260 13636 22318
rect 14028 22372 14084 23660
rect 14588 23548 14644 23660
rect 14028 22306 14084 22316
rect 14476 23492 14644 23548
rect 14812 23714 14868 23726
rect 14812 23662 14814 23714
rect 14866 23662 14868 23714
rect 13580 22194 13636 22204
rect 14252 22258 14308 22270
rect 14252 22206 14254 22258
rect 14306 22206 14308 22258
rect 12908 21758 12910 21810
rect 12962 21758 12964 21810
rect 12908 21476 12964 21758
rect 12908 21410 12964 21420
rect 13244 21980 13412 22036
rect 14252 22036 14308 22206
rect 13244 21364 13300 21980
rect 14252 21970 14308 21980
rect 13916 21810 13972 21822
rect 13916 21758 13918 21810
rect 13970 21758 13972 21810
rect 13916 21700 13972 21758
rect 13916 21634 13972 21644
rect 14140 21700 14196 21738
rect 14140 21634 14196 21644
rect 14476 21700 14532 23492
rect 14812 22372 14868 23662
rect 15036 23380 15092 25340
rect 15148 25284 15204 25788
rect 15372 26292 15428 26302
rect 15372 25506 15428 26236
rect 15372 25454 15374 25506
rect 15426 25454 15428 25506
rect 15372 25442 15428 25454
rect 15148 25218 15204 25228
rect 15148 24164 15204 24174
rect 15148 23826 15204 24108
rect 15484 23940 15540 26910
rect 15596 26962 15652 29708
rect 16044 29428 16100 29438
rect 16044 29334 16100 29372
rect 16044 27748 16100 27758
rect 15596 26910 15598 26962
rect 15650 26910 15652 26962
rect 15596 26898 15652 26910
rect 15708 27188 15764 27198
rect 15596 26740 15652 26750
rect 15596 26514 15652 26684
rect 15596 26462 15598 26514
rect 15650 26462 15652 26514
rect 15596 26450 15652 26462
rect 15708 26516 15764 27132
rect 16044 27076 16100 27692
rect 16156 27300 16212 31500
rect 16268 29652 16324 31614
rect 16604 31444 16660 31724
rect 16604 31378 16660 31388
rect 16828 31778 16884 31790
rect 16828 31726 16830 31778
rect 16882 31726 16884 31778
rect 16604 30994 16660 31006
rect 16604 30942 16606 30994
rect 16658 30942 16660 30994
rect 16268 29586 16324 29596
rect 16492 30884 16548 30894
rect 16380 28756 16436 28766
rect 16380 28662 16436 28700
rect 16156 27234 16212 27244
rect 16268 28644 16324 28654
rect 16044 27010 16100 27020
rect 16268 27074 16324 28588
rect 16492 28532 16548 30828
rect 16268 27022 16270 27074
rect 16322 27022 16324 27074
rect 15820 26964 15876 27002
rect 15820 26898 15876 26908
rect 15820 26516 15876 26526
rect 15708 26514 15876 26516
rect 15708 26462 15822 26514
rect 15874 26462 15876 26514
rect 15708 26460 15876 26462
rect 15820 26450 15876 26460
rect 15932 26516 15988 26526
rect 15708 26292 15764 26302
rect 15932 26292 15988 26460
rect 15708 26290 15988 26292
rect 15708 26238 15710 26290
rect 15762 26238 15988 26290
rect 15708 26236 15988 26238
rect 16268 26292 16324 27022
rect 15708 26226 15764 26236
rect 16268 26226 16324 26236
rect 16380 28476 16548 28532
rect 16156 26180 16212 26190
rect 16156 26086 16212 26124
rect 15820 26068 15876 26078
rect 15148 23774 15150 23826
rect 15202 23774 15204 23826
rect 15148 23762 15204 23774
rect 15260 23884 15484 23940
rect 15036 23314 15092 23324
rect 15260 22596 15316 23884
rect 15484 23874 15540 23884
rect 15708 25284 15764 25294
rect 14812 22306 14868 22316
rect 14924 22540 15316 22596
rect 14588 22260 14644 22270
rect 14588 21810 14644 22204
rect 14924 22148 14980 22540
rect 14588 21758 14590 21810
rect 14642 21758 14644 21810
rect 14588 21746 14644 21758
rect 14812 22092 14980 22148
rect 13356 21588 13412 21598
rect 13692 21588 13748 21626
rect 13356 21586 13524 21588
rect 13356 21534 13358 21586
rect 13410 21534 13524 21586
rect 13356 21532 13524 21534
rect 13356 21522 13412 21532
rect 12684 20748 13076 20804
rect 12460 20692 12516 20702
rect 12460 20598 12516 20636
rect 12572 20690 12628 20702
rect 12572 20638 12574 20690
rect 12626 20638 12628 20690
rect 12460 20132 12516 20142
rect 12124 20018 12292 20020
rect 12124 19966 12126 20018
rect 12178 19966 12292 20018
rect 12124 19964 12292 19966
rect 12124 19954 12180 19964
rect 12012 19796 12068 19806
rect 12012 19234 12068 19740
rect 12124 19348 12180 19358
rect 12124 19254 12180 19292
rect 12012 19182 12014 19234
rect 12066 19182 12068 19234
rect 12012 19170 12068 19182
rect 12236 19236 12292 19964
rect 12348 20130 12516 20132
rect 12348 20078 12462 20130
rect 12514 20078 12516 20130
rect 12348 20076 12516 20078
rect 12348 20020 12404 20076
rect 12460 20066 12516 20076
rect 12572 20132 12628 20638
rect 12572 20066 12628 20076
rect 12684 20578 12740 20590
rect 12684 20526 12686 20578
rect 12738 20526 12740 20578
rect 12684 20244 12740 20526
rect 12348 19954 12404 19964
rect 12460 19236 12516 19246
rect 12236 19234 12516 19236
rect 12236 19182 12462 19234
rect 12514 19182 12516 19234
rect 12236 19180 12516 19182
rect 12460 19170 12516 19180
rect 11788 18564 11844 19068
rect 12236 19012 12292 19022
rect 12684 19012 12740 20188
rect 12236 19010 12740 19012
rect 12236 18958 12238 19010
rect 12290 18958 12740 19010
rect 12236 18956 12740 18958
rect 12796 20578 12852 20590
rect 12796 20526 12798 20578
rect 12850 20526 12852 20578
rect 12236 18946 12292 18956
rect 12796 18788 12852 20526
rect 12908 20580 12964 20590
rect 12908 20486 12964 20524
rect 13020 19908 13076 20748
rect 13244 20692 13300 21308
rect 13468 21140 13524 21532
rect 13692 21522 13748 21532
rect 14028 21474 14084 21486
rect 14028 21422 14030 21474
rect 14082 21422 14084 21474
rect 14028 21364 14084 21422
rect 14028 21298 14084 21308
rect 14364 21364 14420 21374
rect 13468 21074 13524 21084
rect 14252 21028 14308 21038
rect 14140 20916 14196 20926
rect 14140 20822 14196 20860
rect 12908 19684 12964 19694
rect 12908 19346 12964 19628
rect 12908 19294 12910 19346
rect 12962 19294 12964 19346
rect 12908 19282 12964 19294
rect 11788 18498 11844 18508
rect 12348 18732 12852 18788
rect 11676 18452 11732 18462
rect 11452 18450 11732 18452
rect 11452 18398 11678 18450
rect 11730 18398 11732 18450
rect 11452 18396 11732 18398
rect 11564 17780 11620 17790
rect 11340 17778 11620 17780
rect 11340 17726 11566 17778
rect 11618 17726 11620 17778
rect 11340 17724 11620 17726
rect 11564 17714 11620 17724
rect 11116 17614 11118 17666
rect 11170 17614 11172 17666
rect 11116 17602 11172 17614
rect 10556 17554 10612 17566
rect 10556 17502 10558 17554
rect 10610 17502 10612 17554
rect 10556 17108 10612 17502
rect 10556 17042 10612 17052
rect 11564 16884 11620 16894
rect 11676 16884 11732 18396
rect 12348 18450 12404 18732
rect 12348 18398 12350 18450
rect 12402 18398 12404 18450
rect 12348 18386 12404 18398
rect 12460 18564 12516 18574
rect 12460 17778 12516 18508
rect 12460 17726 12462 17778
rect 12514 17726 12516 17778
rect 12460 17714 12516 17726
rect 12796 17780 12852 17790
rect 12012 17108 12068 17118
rect 12012 17014 12068 17052
rect 12796 17106 12852 17724
rect 13020 17668 13076 19852
rect 13020 17602 13076 17612
rect 13132 20636 13244 20692
rect 13132 18452 13188 20636
rect 13244 20626 13300 20636
rect 13468 20692 13524 20702
rect 13468 20598 13524 20636
rect 13804 20578 13860 20590
rect 13804 20526 13806 20578
rect 13858 20526 13860 20578
rect 13244 20132 13300 20142
rect 13244 20038 13300 20076
rect 13804 20132 13860 20526
rect 13804 20066 13860 20076
rect 13580 20018 13636 20030
rect 13580 19966 13582 20018
rect 13634 19966 13636 20018
rect 13580 19236 13636 19966
rect 14028 19908 14084 19918
rect 13580 19170 13636 19180
rect 13916 19852 14028 19908
rect 13692 19124 13748 19134
rect 13916 19124 13972 19852
rect 14028 19814 14084 19852
rect 13692 19122 13972 19124
rect 13692 19070 13694 19122
rect 13746 19070 13972 19122
rect 13692 19068 13972 19070
rect 14140 19236 14196 19246
rect 13692 19058 13748 19068
rect 13020 17444 13076 17454
rect 13132 17444 13188 18396
rect 13468 19010 13524 19022
rect 13468 18958 13470 19010
rect 13522 18958 13524 19010
rect 13468 18004 13524 18958
rect 13580 19012 13636 19022
rect 13580 18918 13636 18956
rect 13692 18004 13748 18014
rect 13468 17948 13692 18004
rect 13580 17780 13636 17790
rect 13580 17686 13636 17724
rect 13020 17442 13188 17444
rect 13020 17390 13022 17442
rect 13074 17390 13188 17442
rect 13020 17388 13188 17390
rect 13020 17378 13076 17388
rect 12796 17054 12798 17106
rect 12850 17054 12852 17106
rect 12796 17042 12852 17054
rect 13580 17108 13636 17118
rect 13692 17108 13748 17948
rect 13636 17052 13748 17108
rect 14028 17666 14084 17678
rect 14028 17614 14030 17666
rect 14082 17614 14084 17666
rect 13580 17014 13636 17052
rect 11620 16828 11732 16884
rect 14028 16884 14084 17614
rect 11564 16790 11620 16828
rect 14028 16324 14084 16828
rect 14028 16258 14084 16268
rect 14140 16212 14196 19180
rect 14252 19234 14308 20972
rect 14252 19182 14254 19234
rect 14306 19182 14308 19234
rect 14252 19170 14308 19182
rect 14364 19124 14420 21308
rect 14476 20580 14532 21644
rect 14700 21588 14756 21598
rect 14812 21588 14868 22092
rect 15148 21924 15204 21934
rect 15148 21810 15204 21868
rect 15148 21758 15150 21810
rect 15202 21758 15204 21810
rect 15148 21746 15204 21758
rect 15596 21812 15652 21822
rect 15596 21718 15652 21756
rect 14700 21586 14868 21588
rect 14700 21534 14702 21586
rect 14754 21534 14868 21586
rect 14700 21532 14868 21534
rect 14924 21586 14980 21598
rect 14924 21534 14926 21586
rect 14978 21534 14980 21586
rect 14588 21476 14644 21486
rect 14588 21362 14644 21420
rect 14588 21310 14590 21362
rect 14642 21310 14644 21362
rect 14588 21298 14644 21310
rect 14700 21364 14756 21532
rect 14700 20692 14756 21308
rect 14700 20626 14756 20636
rect 14476 20242 14532 20524
rect 14476 20190 14478 20242
rect 14530 20190 14532 20242
rect 14476 20178 14532 20190
rect 14588 20468 14644 20478
rect 14588 19234 14644 20412
rect 14924 20356 14980 21534
rect 15260 21586 15316 21598
rect 15260 21534 15262 21586
rect 15314 21534 15316 21586
rect 15036 20468 15092 20478
rect 15260 20468 15316 21534
rect 15484 21588 15540 21598
rect 15092 20412 15316 20468
rect 15372 21364 15428 21374
rect 15036 20402 15092 20412
rect 14924 20290 14980 20300
rect 14700 20132 14756 20142
rect 14700 20018 14756 20076
rect 14700 19966 14702 20018
rect 14754 19966 14756 20018
rect 14700 19796 14756 19966
rect 15148 20132 15204 20142
rect 14924 19908 14980 19918
rect 14700 19730 14756 19740
rect 14812 19852 14924 19908
rect 14812 19236 14868 19852
rect 14924 19842 14980 19852
rect 15148 19796 15204 20076
rect 15260 20130 15316 20142
rect 15260 20078 15262 20130
rect 15314 20078 15316 20130
rect 15260 20020 15316 20078
rect 15372 20130 15428 21308
rect 15372 20078 15374 20130
rect 15426 20078 15428 20130
rect 15372 20066 15428 20078
rect 15484 20244 15540 21532
rect 15708 21476 15764 25228
rect 15820 23042 15876 26012
rect 16268 26068 16324 26078
rect 16156 25394 16212 25406
rect 16156 25342 16158 25394
rect 16210 25342 16212 25394
rect 16156 25172 16212 25342
rect 16156 25106 16212 25116
rect 16044 24948 16100 24958
rect 16268 24948 16324 26012
rect 16044 24946 16324 24948
rect 16044 24894 16046 24946
rect 16098 24894 16324 24946
rect 16044 24892 16324 24894
rect 16044 24882 16100 24892
rect 15932 24836 15988 24846
rect 15932 24050 15988 24780
rect 15932 23998 15934 24050
rect 15986 23998 15988 24050
rect 15932 23986 15988 23998
rect 16380 23380 16436 28476
rect 16492 27858 16548 27870
rect 16492 27806 16494 27858
rect 16546 27806 16548 27858
rect 16492 27524 16548 27806
rect 16492 27458 16548 27468
rect 16492 27300 16548 27310
rect 16492 25284 16548 27244
rect 16604 26290 16660 30942
rect 16828 30324 16884 31726
rect 17052 31780 17108 31790
rect 17052 31332 17108 31724
rect 17052 30436 17108 31276
rect 16828 30258 16884 30268
rect 16940 30380 17108 30436
rect 16828 30098 16884 30110
rect 16828 30046 16830 30098
rect 16882 30046 16884 30098
rect 16828 29988 16884 30046
rect 16828 29922 16884 29932
rect 16828 29652 16884 29662
rect 16940 29652 16996 30380
rect 16828 29650 16996 29652
rect 16828 29598 16830 29650
rect 16882 29598 16996 29650
rect 16828 29596 16996 29598
rect 17052 30212 17108 30222
rect 16828 29586 16884 29596
rect 17052 28644 17108 30156
rect 17052 28550 17108 28588
rect 17164 28420 17220 32396
rect 17500 31780 17556 34078
rect 17724 33684 17780 33694
rect 17724 32786 17780 33628
rect 17836 33460 17892 34190
rect 17836 33394 17892 33404
rect 17948 33236 18004 35084
rect 18060 33458 18116 35756
rect 18172 35588 18228 35598
rect 18172 35494 18228 35532
rect 18060 33406 18062 33458
rect 18114 33406 18116 33458
rect 18060 33394 18116 33406
rect 18172 34242 18228 34254
rect 18172 34190 18174 34242
rect 18226 34190 18228 34242
rect 18172 33348 18228 34190
rect 18172 33282 18228 33292
rect 17724 32734 17726 32786
rect 17778 32734 17780 32786
rect 17724 32722 17780 32734
rect 17836 33234 18004 33236
rect 17836 33182 17950 33234
rect 18002 33182 18004 33234
rect 17836 33180 18004 33182
rect 17500 31666 17556 31724
rect 17500 31614 17502 31666
rect 17554 31614 17556 31666
rect 17500 31602 17556 31614
rect 17500 31444 17556 31454
rect 17388 30996 17444 31006
rect 17388 30902 17444 30940
rect 17500 29650 17556 31388
rect 17836 30436 17892 33180
rect 17948 33170 18004 33180
rect 18284 33012 18340 35868
rect 18508 35026 18564 35980
rect 18956 35970 19012 35980
rect 18620 35698 18676 35710
rect 18620 35646 18622 35698
rect 18674 35646 18676 35698
rect 18620 35252 18676 35646
rect 18620 35186 18676 35196
rect 18844 35140 18900 35150
rect 19068 35140 19124 37436
rect 19180 37266 19236 37278
rect 19180 37214 19182 37266
rect 19234 37214 19236 37266
rect 19180 36932 19236 37214
rect 19292 37266 19348 37278
rect 19292 37214 19294 37266
rect 19346 37214 19348 37266
rect 19292 37044 19348 37214
rect 19292 36978 19348 36988
rect 19180 36866 19236 36876
rect 19404 36820 19460 36830
rect 19404 36482 19460 36764
rect 19404 36430 19406 36482
rect 19458 36430 19460 36482
rect 19404 36418 19460 36430
rect 19404 35924 19460 35934
rect 19404 35830 19460 35868
rect 19516 35812 19572 37774
rect 19628 37828 19684 38108
rect 20076 38050 20132 38444
rect 20076 37998 20078 38050
rect 20130 37998 20132 38050
rect 20076 37986 20132 37998
rect 20188 38164 20244 38174
rect 19740 37828 19796 37838
rect 19628 37826 19796 37828
rect 19628 37774 19742 37826
rect 19794 37774 19796 37826
rect 19628 37772 19796 37774
rect 19628 37268 19684 37772
rect 19740 37762 19796 37772
rect 19836 37660 20100 37670
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 19836 37594 20100 37604
rect 19852 37492 19908 37502
rect 20188 37492 20244 38108
rect 20524 38052 20580 38062
rect 20524 38050 20692 38052
rect 20524 37998 20526 38050
rect 20578 37998 20692 38050
rect 20524 37996 20692 37998
rect 20524 37986 20580 37996
rect 19852 37398 19908 37436
rect 20076 37490 20244 37492
rect 20076 37438 20190 37490
rect 20242 37438 20244 37490
rect 20076 37436 20244 37438
rect 19740 37268 19796 37278
rect 19628 37212 19740 37268
rect 19740 37174 19796 37212
rect 19964 37266 20020 37278
rect 19964 37214 19966 37266
rect 20018 37214 20020 37266
rect 19964 37156 20020 37214
rect 19964 37090 20020 37100
rect 20076 36932 20132 37436
rect 20188 37426 20244 37436
rect 20524 37268 20580 37278
rect 20076 36866 20132 36876
rect 20300 37266 20580 37268
rect 20300 37214 20526 37266
rect 20578 37214 20580 37266
rect 20300 37212 20580 37214
rect 20636 37268 20692 37996
rect 20748 37940 20804 37950
rect 20748 37846 20804 37884
rect 21196 37490 21252 40012
rect 21980 39620 22036 39630
rect 21756 39618 22036 39620
rect 21756 39566 21982 39618
rect 22034 39566 22036 39618
rect 21756 39564 22036 39566
rect 21420 39508 21476 39518
rect 21308 39506 21476 39508
rect 21308 39454 21422 39506
rect 21474 39454 21476 39506
rect 21308 39452 21476 39454
rect 21308 38724 21364 39452
rect 21420 39442 21476 39452
rect 21756 39506 21812 39564
rect 21980 39554 22036 39564
rect 21756 39454 21758 39506
rect 21810 39454 21812 39506
rect 21756 39442 21812 39454
rect 22092 39508 22148 45836
rect 22204 45556 22260 45566
rect 22204 43428 22260 45500
rect 22428 44660 22484 47182
rect 22764 47346 22820 47358
rect 22764 47294 22766 47346
rect 22818 47294 22820 47346
rect 22540 46676 22596 46686
rect 22540 46002 22596 46620
rect 22764 46116 22820 47294
rect 23436 47346 23492 47358
rect 23436 47294 23438 47346
rect 23490 47294 23492 47346
rect 22876 47236 22932 47246
rect 22876 47142 22932 47180
rect 23100 47236 23156 47246
rect 23436 47236 23492 47294
rect 23100 47234 23492 47236
rect 23100 47182 23102 47234
rect 23154 47182 23492 47234
rect 23100 47180 23492 47182
rect 23100 47170 23156 47180
rect 23100 46676 23156 46686
rect 23100 46582 23156 46620
rect 23212 46564 23268 46574
rect 23212 46470 23268 46508
rect 22764 46060 22932 46116
rect 22540 45950 22542 46002
rect 22594 45950 22596 46002
rect 22540 45938 22596 45950
rect 22876 45668 22932 46060
rect 22988 45892 23044 45902
rect 23212 45892 23268 45902
rect 23044 45890 23268 45892
rect 23044 45838 23214 45890
rect 23266 45838 23268 45890
rect 23044 45836 23268 45838
rect 22988 45826 23044 45836
rect 23212 45826 23268 45836
rect 22876 45574 22932 45612
rect 23436 45220 23492 45230
rect 22540 44996 22596 45006
rect 22540 44902 22596 44940
rect 22428 44604 22596 44660
rect 22316 43428 22372 43438
rect 22204 43426 22372 43428
rect 22204 43374 22318 43426
rect 22370 43374 22372 43426
rect 22204 43372 22372 43374
rect 22316 43362 22372 43372
rect 22428 40402 22484 40414
rect 22428 40350 22430 40402
rect 22482 40350 22484 40402
rect 22428 40180 22484 40350
rect 22204 39732 22260 39742
rect 22204 39638 22260 39676
rect 22316 39618 22372 39630
rect 22316 39566 22318 39618
rect 22370 39566 22372 39618
rect 22316 39508 22372 39566
rect 22092 39452 22260 39508
rect 21308 38658 21364 38668
rect 21756 38834 21812 38846
rect 21756 38782 21758 38834
rect 21810 38782 21812 38834
rect 21644 38052 21700 38062
rect 21196 37438 21198 37490
rect 21250 37438 21252 37490
rect 21196 37426 21252 37438
rect 21308 38050 21700 38052
rect 21308 37998 21646 38050
rect 21698 37998 21700 38050
rect 21308 37996 21700 37998
rect 20860 37380 20916 37390
rect 20636 37212 20804 37268
rect 20300 36706 20356 37212
rect 20524 37202 20580 37212
rect 20300 36654 20302 36706
rect 20354 36654 20356 36706
rect 20076 36482 20132 36494
rect 20076 36430 20078 36482
rect 20130 36430 20132 36482
rect 20076 36260 20132 36430
rect 20076 36204 20244 36260
rect 19836 36092 20100 36102
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 19836 36026 20100 36036
rect 19516 35746 19572 35756
rect 19964 35924 20020 35934
rect 20188 35924 20244 36204
rect 18844 35138 19124 35140
rect 18844 35086 18846 35138
rect 18898 35086 19124 35138
rect 18844 35084 19124 35086
rect 18844 35074 18900 35084
rect 18508 34974 18510 35026
rect 18562 34974 18564 35026
rect 18508 34962 18564 34974
rect 19404 35028 19460 35038
rect 19404 34914 19460 34972
rect 19404 34862 19406 34914
rect 19458 34862 19460 34914
rect 19404 34850 19460 34862
rect 19628 34916 19684 34926
rect 19964 34916 20020 35868
rect 20076 35868 20244 35924
rect 20076 35252 20132 35868
rect 20076 35186 20132 35196
rect 20300 34916 20356 36654
rect 20412 36484 20468 36494
rect 20412 35698 20468 36428
rect 20636 36258 20692 36270
rect 20636 36206 20638 36258
rect 20690 36206 20692 36258
rect 20636 36148 20692 36206
rect 20636 36082 20692 36092
rect 20412 35646 20414 35698
rect 20466 35646 20468 35698
rect 20412 35634 20468 35646
rect 20636 35698 20692 35710
rect 20636 35646 20638 35698
rect 20690 35646 20692 35698
rect 20636 35364 20692 35646
rect 20636 35298 20692 35308
rect 20748 35586 20804 37212
rect 20860 37044 20916 37324
rect 21084 37378 21140 37390
rect 21084 37326 21086 37378
rect 21138 37326 21140 37378
rect 20860 36978 20916 36988
rect 20972 37268 21028 37278
rect 20748 35534 20750 35586
rect 20802 35534 20804 35586
rect 20524 35252 20580 35262
rect 20524 35026 20580 35196
rect 20524 34974 20526 35026
rect 20578 34974 20580 35026
rect 20524 34962 20580 34974
rect 19964 34860 20132 34916
rect 19628 34822 19684 34860
rect 19292 34804 19348 34814
rect 19292 34710 19348 34748
rect 19964 34692 20020 34702
rect 19628 34690 20020 34692
rect 19628 34638 19966 34690
rect 20018 34638 20020 34690
rect 19628 34636 20020 34638
rect 20076 34692 20132 34860
rect 20076 34636 20244 34692
rect 17948 32956 18340 33012
rect 18508 34244 18564 34254
rect 18508 33572 18564 34188
rect 19404 34132 19460 34142
rect 19292 34130 19460 34132
rect 19292 34078 19406 34130
rect 19458 34078 19460 34130
rect 19292 34076 19460 34078
rect 19180 34018 19236 34030
rect 19180 33966 19182 34018
rect 19234 33966 19236 34018
rect 17948 30994 18004 32956
rect 18284 32450 18340 32462
rect 18284 32398 18286 32450
rect 18338 32398 18340 32450
rect 18060 32340 18116 32350
rect 18060 32246 18116 32284
rect 18284 32004 18340 32398
rect 18284 31938 18340 31948
rect 18284 31780 18340 31790
rect 18284 31686 18340 31724
rect 18508 31218 18564 33516
rect 19068 33908 19124 33918
rect 19068 33346 19124 33852
rect 19180 33796 19236 33966
rect 19180 33730 19236 33740
rect 19068 33294 19070 33346
rect 19122 33294 19124 33346
rect 18508 31166 18510 31218
rect 18562 31166 18564 31218
rect 18508 31154 18564 31166
rect 18620 32562 18676 32574
rect 18620 32510 18622 32562
rect 18674 32510 18676 32562
rect 18620 32340 18676 32510
rect 17948 30942 17950 30994
rect 18002 30942 18004 30994
rect 17948 30930 18004 30942
rect 18060 30996 18116 31006
rect 17500 29598 17502 29650
rect 17554 29598 17556 29650
rect 17500 29586 17556 29598
rect 17724 30380 17892 30436
rect 17388 29428 17444 29438
rect 17388 29334 17444 29372
rect 17724 28642 17780 30380
rect 17724 28590 17726 28642
rect 17778 28590 17780 28642
rect 16940 28364 17220 28420
rect 17388 28532 17444 28542
rect 16828 27970 16884 27982
rect 16828 27918 16830 27970
rect 16882 27918 16884 27970
rect 16828 27300 16884 27918
rect 16828 27234 16884 27244
rect 16604 26238 16606 26290
rect 16658 26238 16660 26290
rect 16604 26068 16660 26238
rect 16604 26002 16660 26012
rect 16492 25228 16772 25284
rect 16716 24836 16772 25228
rect 16716 24770 16772 24780
rect 16716 24610 16772 24622
rect 16716 24558 16718 24610
rect 16770 24558 16772 24610
rect 16716 23604 16772 24558
rect 16716 23538 16772 23548
rect 16828 24498 16884 24510
rect 16828 24446 16830 24498
rect 16882 24446 16884 24498
rect 16268 23324 16436 23380
rect 15820 22990 15822 23042
rect 15874 22990 15876 23042
rect 15820 22260 15876 22990
rect 16156 23156 16212 23166
rect 15820 22194 15876 22204
rect 15932 22708 15988 22718
rect 15260 19954 15316 19964
rect 15260 19796 15316 19806
rect 15148 19794 15316 19796
rect 15148 19742 15262 19794
rect 15314 19742 15316 19794
rect 15148 19740 15316 19742
rect 15260 19730 15316 19740
rect 14588 19182 14590 19234
rect 14642 19182 14644 19234
rect 14588 19170 14644 19182
rect 14700 19180 14868 19236
rect 14476 19124 14532 19134
rect 14364 19122 14532 19124
rect 14364 19070 14478 19122
rect 14530 19070 14532 19122
rect 14364 19068 14532 19070
rect 14476 19058 14532 19068
rect 14588 18676 14644 18686
rect 14700 18676 14756 19180
rect 15148 19124 15204 19134
rect 15148 19030 15204 19068
rect 14588 18674 14756 18676
rect 14588 18622 14590 18674
rect 14642 18622 14756 18674
rect 14588 18620 14756 18622
rect 14812 19012 14868 19022
rect 14588 18610 14644 18620
rect 14700 18340 14756 18350
rect 14700 16994 14756 18284
rect 14812 17778 14868 18956
rect 15484 18900 15540 20188
rect 15596 21420 15764 21476
rect 15932 21810 15988 22652
rect 15932 21758 15934 21810
rect 15986 21758 15988 21810
rect 15596 19236 15652 21420
rect 15820 20692 15876 20702
rect 15820 20242 15876 20636
rect 15820 20190 15822 20242
rect 15874 20190 15876 20242
rect 15820 20178 15876 20190
rect 15708 19908 15764 19918
rect 15708 19814 15764 19852
rect 15596 19170 15652 19180
rect 14812 17726 14814 17778
rect 14866 17726 14868 17778
rect 14812 17714 14868 17726
rect 15148 18844 15540 18900
rect 15708 19010 15764 19022
rect 15708 18958 15710 19010
rect 15762 18958 15764 19010
rect 15148 18450 15204 18844
rect 15148 18398 15150 18450
rect 15202 18398 15204 18450
rect 15148 17780 15204 18398
rect 15596 18452 15652 18462
rect 15596 18358 15652 18396
rect 15148 17714 15204 17724
rect 14700 16942 14702 16994
rect 14754 16942 14756 16994
rect 14700 16930 14756 16942
rect 14924 16324 14980 16334
rect 14588 16212 14644 16222
rect 14140 16210 14644 16212
rect 14140 16158 14590 16210
rect 14642 16158 14644 16210
rect 14140 16156 14644 16158
rect 14588 16146 14644 16156
rect 14924 16210 14980 16268
rect 14924 16158 14926 16210
rect 14978 16158 14980 16210
rect 14924 16146 14980 16158
rect 15708 16100 15764 18958
rect 15932 16212 15988 21758
rect 16156 21588 16212 23100
rect 16268 21812 16324 23324
rect 16380 23154 16436 23166
rect 16380 23102 16382 23154
rect 16434 23102 16436 23154
rect 16380 22482 16436 23102
rect 16828 22820 16884 24446
rect 16828 22754 16884 22764
rect 16380 22430 16382 22482
rect 16434 22430 16436 22482
rect 16380 22372 16436 22430
rect 16940 22482 16996 28364
rect 17388 28082 17444 28476
rect 17388 28030 17390 28082
rect 17442 28030 17444 28082
rect 17388 28018 17444 28030
rect 17500 28530 17556 28542
rect 17500 28478 17502 28530
rect 17554 28478 17556 28530
rect 17052 26962 17108 26974
rect 17052 26910 17054 26962
rect 17106 26910 17108 26962
rect 17052 26908 17108 26910
rect 17500 26908 17556 28478
rect 17724 27748 17780 28590
rect 17836 28756 17892 28766
rect 17836 28644 17892 28700
rect 17948 28644 18004 28654
rect 17836 28642 18004 28644
rect 17836 28590 17950 28642
rect 18002 28590 18004 28642
rect 17836 28588 18004 28590
rect 17948 28578 18004 28588
rect 17836 27748 17892 27758
rect 17780 27746 17892 27748
rect 17780 27694 17838 27746
rect 17890 27694 17892 27746
rect 17780 27692 17892 27694
rect 17724 27654 17780 27692
rect 17836 27682 17892 27692
rect 17052 26852 17332 26908
rect 17276 25732 17332 26852
rect 17388 26852 17556 26908
rect 17388 26516 17444 26852
rect 17388 26450 17444 26460
rect 17948 26516 18004 26526
rect 18060 26516 18116 30940
rect 18620 30884 18676 32284
rect 19068 31780 19124 33294
rect 19180 32676 19236 32686
rect 19292 32676 19348 34076
rect 19404 34066 19460 34076
rect 19628 33684 19684 34636
rect 19964 34626 20020 34636
rect 19836 34524 20100 34534
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 19836 34458 20100 34468
rect 20188 34356 20244 34636
rect 19964 34300 20244 34356
rect 19964 34244 20020 34300
rect 19628 33618 19684 33628
rect 19740 34242 20020 34244
rect 19740 34190 19966 34242
rect 20018 34190 20020 34242
rect 19740 34188 20020 34190
rect 19740 33460 19796 34188
rect 19964 34178 20020 34188
rect 19628 33404 19796 33460
rect 20300 33458 20356 34860
rect 20636 34242 20692 34254
rect 20636 34190 20638 34242
rect 20690 34190 20692 34242
rect 20524 34130 20580 34142
rect 20524 34078 20526 34130
rect 20578 34078 20580 34130
rect 20524 33796 20580 34078
rect 20524 33730 20580 33740
rect 20300 33406 20302 33458
rect 20354 33406 20356 33458
rect 19628 33236 19684 33404
rect 20300 33394 20356 33406
rect 20636 33348 20692 34190
rect 20748 33796 20804 35534
rect 20972 36372 21028 37212
rect 20860 34020 20916 34030
rect 20972 34020 21028 36316
rect 21084 35924 21140 37326
rect 21308 36260 21364 37996
rect 21644 37986 21700 37996
rect 21756 37940 21812 38782
rect 22092 38722 22148 38734
rect 22092 38670 22094 38722
rect 22146 38670 22148 38722
rect 22092 38668 22148 38670
rect 21980 38612 22148 38668
rect 21980 38500 22036 38612
rect 21756 37874 21812 37884
rect 21868 38276 21924 38286
rect 21420 37826 21476 37838
rect 21420 37774 21422 37826
rect 21474 37774 21476 37826
rect 21420 36820 21476 37774
rect 21532 37826 21588 37838
rect 21532 37774 21534 37826
rect 21586 37774 21588 37826
rect 21532 36932 21588 37774
rect 21644 37828 21700 37838
rect 21644 37490 21700 37772
rect 21644 37438 21646 37490
rect 21698 37438 21700 37490
rect 21644 37426 21700 37438
rect 21868 37716 21924 38220
rect 21868 37268 21924 37660
rect 21868 37174 21924 37212
rect 21756 37154 21812 37166
rect 21756 37102 21758 37154
rect 21810 37102 21812 37154
rect 21756 36932 21812 37102
rect 21756 36876 21924 36932
rect 21532 36866 21588 36876
rect 21420 36754 21476 36764
rect 21644 36820 21700 36830
rect 21700 36764 21812 36820
rect 21644 36754 21700 36764
rect 21308 36194 21364 36204
rect 21420 36482 21476 36494
rect 21420 36430 21422 36482
rect 21474 36430 21476 36482
rect 21084 35868 21252 35924
rect 21084 35700 21140 35710
rect 21084 35606 21140 35644
rect 21196 34580 21252 35868
rect 21420 35364 21476 36430
rect 21532 36484 21588 36494
rect 21532 36370 21588 36428
rect 21532 36318 21534 36370
rect 21586 36318 21588 36370
rect 21532 36306 21588 36318
rect 21532 35812 21588 35822
rect 21532 35718 21588 35756
rect 21420 35298 21476 35308
rect 21420 35028 21476 35038
rect 21420 34934 21476 34972
rect 21308 34804 21364 34814
rect 21308 34710 21364 34748
rect 21532 34692 21588 34702
rect 21420 34690 21588 34692
rect 21420 34638 21534 34690
rect 21586 34638 21588 34690
rect 21420 34636 21588 34638
rect 21420 34580 21476 34636
rect 21532 34626 21588 34636
rect 21756 34690 21812 36764
rect 21868 36372 21924 36876
rect 21980 36594 22036 38444
rect 22092 37938 22148 37950
rect 22092 37886 22094 37938
rect 22146 37886 22148 37938
rect 22092 37156 22148 37886
rect 22204 37492 22260 39452
rect 22316 39442 22372 39452
rect 22428 39172 22484 40124
rect 22428 39106 22484 39116
rect 22428 38276 22484 38286
rect 22540 38276 22596 44604
rect 23436 44322 23492 45164
rect 23548 44996 23604 45006
rect 23548 44434 23604 44940
rect 23548 44382 23550 44434
rect 23602 44382 23604 44434
rect 23548 44370 23604 44382
rect 23436 44270 23438 44322
rect 23490 44270 23492 44322
rect 23436 44258 23492 44270
rect 23660 44324 23716 44334
rect 22764 44100 22820 44110
rect 23660 44100 23716 44268
rect 22820 44044 22932 44100
rect 22764 44006 22820 44044
rect 22652 42868 22708 42878
rect 22652 42774 22708 42812
rect 22652 41972 22708 41982
rect 22652 41858 22708 41916
rect 22652 41806 22654 41858
rect 22706 41806 22708 41858
rect 22652 41794 22708 41806
rect 22652 39506 22708 39518
rect 22652 39454 22654 39506
rect 22706 39454 22708 39506
rect 22652 39058 22708 39454
rect 22652 39006 22654 39058
rect 22706 39006 22708 39058
rect 22652 38994 22708 39006
rect 22428 38274 22596 38276
rect 22428 38222 22430 38274
rect 22482 38222 22596 38274
rect 22428 38220 22596 38222
rect 22428 38210 22484 38220
rect 22316 37826 22372 37838
rect 22316 37774 22318 37826
rect 22370 37774 22372 37826
rect 22316 37716 22372 37774
rect 22652 37828 22708 37838
rect 22708 37772 22820 37828
rect 22652 37762 22708 37772
rect 22316 37650 22372 37660
rect 22764 37492 22820 37772
rect 22204 37436 22484 37492
rect 22316 37268 22372 37278
rect 22316 37174 22372 37212
rect 22204 37156 22260 37166
rect 22092 37100 22204 37156
rect 22204 37090 22260 37100
rect 21980 36542 21982 36594
rect 22034 36542 22036 36594
rect 21980 36530 22036 36542
rect 22316 36482 22372 36494
rect 22316 36430 22318 36482
rect 22370 36430 22372 36482
rect 21868 36316 22036 36372
rect 21868 36148 21924 36158
rect 21868 35698 21924 36092
rect 21868 35646 21870 35698
rect 21922 35646 21924 35698
rect 21868 35634 21924 35646
rect 21980 35700 22036 36316
rect 22316 36148 22372 36430
rect 22316 36082 22372 36092
rect 22428 35922 22484 37436
rect 22428 35870 22430 35922
rect 22482 35870 22484 35922
rect 22428 35858 22484 35870
rect 22540 37044 22596 37054
rect 22540 35810 22596 36988
rect 22540 35758 22542 35810
rect 22594 35758 22596 35810
rect 22540 35746 22596 35758
rect 22652 37042 22708 37054
rect 22652 36990 22654 37042
rect 22706 36990 22708 37042
rect 22204 35700 22260 35710
rect 21980 35698 22260 35700
rect 21980 35646 22206 35698
rect 22258 35646 22260 35698
rect 21980 35644 22260 35646
rect 22204 35634 22260 35644
rect 21756 34638 21758 34690
rect 21810 34638 21812 34690
rect 21196 34524 21476 34580
rect 20860 34018 21028 34020
rect 20860 33966 20862 34018
rect 20914 33966 21028 34018
rect 20860 33964 21028 33966
rect 21308 34018 21364 34030
rect 21308 33966 21310 34018
rect 21362 33966 21364 34018
rect 20860 33954 20916 33964
rect 20748 33740 20916 33796
rect 20412 33292 20692 33348
rect 19180 32674 19460 32676
rect 19180 32622 19182 32674
rect 19234 32622 19460 32674
rect 19180 32620 19460 32622
rect 19180 32610 19236 32620
rect 19068 31714 19124 31724
rect 18620 30790 18676 30828
rect 18732 31556 18788 31566
rect 18396 29652 18452 29662
rect 18396 29426 18452 29596
rect 18732 29650 18788 31500
rect 18732 29598 18734 29650
rect 18786 29598 18788 29650
rect 18732 29586 18788 29598
rect 18844 30994 18900 31006
rect 18844 30942 18846 30994
rect 18898 30942 18900 30994
rect 18844 29538 18900 30942
rect 18956 30324 19012 30334
rect 18956 30322 19348 30324
rect 18956 30270 18958 30322
rect 19010 30270 19348 30322
rect 18956 30268 19348 30270
rect 18956 30258 19012 30268
rect 18844 29486 18846 29538
rect 18898 29486 18900 29538
rect 18396 29374 18398 29426
rect 18450 29374 18452 29426
rect 18396 29362 18452 29374
rect 18620 29426 18676 29438
rect 18620 29374 18622 29426
rect 18674 29374 18676 29426
rect 18172 28868 18228 28878
rect 18228 28812 18340 28868
rect 18172 28802 18228 28812
rect 18172 28642 18228 28654
rect 18172 28590 18174 28642
rect 18226 28590 18228 28642
rect 18172 27188 18228 28590
rect 18284 28420 18340 28812
rect 18396 28644 18452 28654
rect 18452 28588 18564 28644
rect 18396 28578 18452 28588
rect 18396 28420 18452 28430
rect 18284 28418 18452 28420
rect 18284 28366 18398 28418
rect 18450 28366 18452 28418
rect 18284 28364 18452 28366
rect 18396 28354 18452 28364
rect 18508 27860 18564 28588
rect 18620 28084 18676 29374
rect 18620 28018 18676 28028
rect 18844 27972 18900 29486
rect 19180 30100 19236 30110
rect 19180 29428 19236 30044
rect 19068 29426 19236 29428
rect 19068 29374 19182 29426
rect 19234 29374 19236 29426
rect 19068 29372 19236 29374
rect 18956 28642 19012 28654
rect 18956 28590 18958 28642
rect 19010 28590 19012 28642
rect 18956 28420 19012 28590
rect 18956 28354 19012 28364
rect 18844 27916 19012 27972
rect 18620 27860 18676 27870
rect 18508 27858 18900 27860
rect 18508 27806 18622 27858
rect 18674 27806 18900 27858
rect 18508 27804 18900 27806
rect 18620 27794 18676 27804
rect 18732 27636 18788 27646
rect 18620 27300 18676 27310
rect 18228 27132 18452 27188
rect 18172 27094 18228 27132
rect 18396 27076 18452 27132
rect 18396 27020 18564 27076
rect 18396 26908 18452 26918
rect 18284 26516 18340 26526
rect 18060 26514 18340 26516
rect 18060 26462 18286 26514
rect 18338 26462 18340 26514
rect 18060 26460 18340 26462
rect 17948 26422 18004 26460
rect 18284 26450 18340 26460
rect 17388 26290 17444 26302
rect 17388 26238 17390 26290
rect 17442 26238 17444 26290
rect 17388 26068 17444 26238
rect 17388 26002 17444 26012
rect 17276 25676 17892 25732
rect 17724 25060 17780 25070
rect 17724 24724 17780 25004
rect 17612 24722 17780 24724
rect 17612 24670 17726 24722
rect 17778 24670 17780 24722
rect 17612 24668 17780 24670
rect 17612 23716 17668 24668
rect 17724 24658 17780 24668
rect 17836 24612 17892 25676
rect 18284 25620 18340 25630
rect 18396 25620 18452 26852
rect 18284 25618 18452 25620
rect 18284 25566 18286 25618
rect 18338 25566 18452 25618
rect 18284 25564 18452 25566
rect 18284 25554 18340 25564
rect 18172 25284 18228 25294
rect 18172 24834 18228 25228
rect 18508 24948 18564 27020
rect 18620 26404 18676 27244
rect 18620 26310 18676 26348
rect 18620 25732 18676 25742
rect 18732 25732 18788 27580
rect 18620 25730 18788 25732
rect 18620 25678 18622 25730
rect 18674 25678 18788 25730
rect 18620 25676 18788 25678
rect 18620 25666 18676 25676
rect 18620 25508 18676 25518
rect 18620 25172 18676 25452
rect 18732 25396 18788 25406
rect 18732 25302 18788 25340
rect 18620 25116 18788 25172
rect 18508 24892 18676 24948
rect 18172 24782 18174 24834
rect 18226 24782 18228 24834
rect 18172 24770 18228 24782
rect 18284 24834 18340 24846
rect 18284 24782 18286 24834
rect 18338 24782 18340 24834
rect 18172 24612 18228 24622
rect 17836 24610 18228 24612
rect 17836 24558 18174 24610
rect 18226 24558 18228 24610
rect 17836 24556 18228 24558
rect 18172 24546 18228 24556
rect 18284 24276 18340 24782
rect 17612 23268 17668 23660
rect 17948 23940 18004 23950
rect 17612 23154 17668 23212
rect 17612 23102 17614 23154
rect 17666 23102 17668 23154
rect 17612 23090 17668 23102
rect 17836 23604 17892 23614
rect 17724 22820 17780 22830
rect 16940 22430 16942 22482
rect 16994 22430 16996 22482
rect 16940 22418 16996 22430
rect 17612 22596 17668 22606
rect 16716 22372 16772 22382
rect 16380 22370 16772 22372
rect 16380 22318 16718 22370
rect 16770 22318 16772 22370
rect 16380 22316 16772 22318
rect 16716 22306 16772 22316
rect 17612 22372 17668 22540
rect 17612 22278 17668 22316
rect 16716 21924 16772 21934
rect 16268 21756 16436 21812
rect 16268 21588 16324 21598
rect 16212 21586 16324 21588
rect 16212 21534 16270 21586
rect 16322 21534 16324 21586
rect 16212 21532 16324 21534
rect 16156 21494 16212 21532
rect 16268 21522 16324 21532
rect 16268 20692 16324 20702
rect 16268 20598 16324 20636
rect 16380 20244 16436 21756
rect 16716 21476 16772 21868
rect 16268 20188 16436 20244
rect 16604 21474 16772 21476
rect 16604 21422 16718 21474
rect 16770 21422 16772 21474
rect 16604 21420 16772 21422
rect 16268 20020 16324 20188
rect 16492 20132 16548 20142
rect 16268 19954 16324 19964
rect 16380 20076 16492 20132
rect 16044 19348 16100 19358
rect 16044 19254 16100 19292
rect 16380 19234 16436 20076
rect 16492 20038 16548 20076
rect 16380 19182 16382 19234
rect 16434 19182 16436 19234
rect 16268 18564 16324 18574
rect 16380 18564 16436 19182
rect 16492 19012 16548 19022
rect 16492 18918 16548 18956
rect 16604 18788 16660 21420
rect 16716 21410 16772 21420
rect 16940 21588 16996 21598
rect 16828 20244 16884 20254
rect 16940 20244 16996 21532
rect 17724 21586 17780 22764
rect 17724 21534 17726 21586
rect 17778 21534 17780 21586
rect 17724 21522 17780 21534
rect 17724 21364 17780 21374
rect 16828 20242 16996 20244
rect 16828 20190 16830 20242
rect 16882 20190 16996 20242
rect 16828 20188 16996 20190
rect 16828 20178 16884 20188
rect 16940 20020 16996 20188
rect 16940 19954 16996 19964
rect 17052 20802 17108 20814
rect 17052 20750 17054 20802
rect 17106 20750 17108 20802
rect 16268 18562 16436 18564
rect 16268 18510 16270 18562
rect 16322 18510 16436 18562
rect 16268 18508 16436 18510
rect 16492 18732 16660 18788
rect 16716 19460 16772 19470
rect 16716 19234 16772 19404
rect 16716 19182 16718 19234
rect 16770 19182 16772 19234
rect 16268 18498 16324 18508
rect 16380 18340 16436 18350
rect 16380 18246 16436 18284
rect 16268 16212 16324 16222
rect 15932 16210 16324 16212
rect 15932 16158 16270 16210
rect 16322 16158 16324 16210
rect 15932 16156 16324 16158
rect 16268 16146 16324 16156
rect 15708 16044 16212 16100
rect 16156 15988 16212 16044
rect 16492 15988 16548 18732
rect 16604 18450 16660 18462
rect 16604 18398 16606 18450
rect 16658 18398 16660 18450
rect 16604 16212 16660 18398
rect 16604 16146 16660 16156
rect 16156 15932 16548 15988
rect 16044 15876 16100 15886
rect 14700 15204 14756 15214
rect 5852 15092 6020 15148
rect 4476 14924 4740 14934
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4476 14858 4740 14868
rect 4476 13356 4740 13366
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4476 13290 4740 13300
rect 4476 11788 4740 11798
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4476 11722 4740 11732
rect 4476 10220 4740 10230
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4476 10154 4740 10164
rect 5964 9940 6020 15092
rect 14700 13858 14756 15148
rect 16044 14642 16100 15820
rect 16268 15316 16324 15326
rect 16268 15222 16324 15260
rect 16380 15204 16436 15242
rect 16380 15138 16436 15148
rect 16492 15148 16548 15932
rect 16604 15428 16660 15438
rect 16716 15428 16772 19182
rect 16940 19122 16996 19134
rect 16940 19070 16942 19122
rect 16994 19070 16996 19122
rect 16940 19012 16996 19070
rect 16940 18946 16996 18956
rect 16828 18562 16884 18574
rect 16828 18510 16830 18562
rect 16882 18510 16884 18562
rect 16828 18452 16884 18510
rect 16940 18452 16996 18462
rect 16828 18396 16940 18452
rect 16940 18386 16996 18396
rect 16940 17778 16996 17790
rect 16940 17726 16942 17778
rect 16994 17726 16996 17778
rect 16940 17668 16996 17726
rect 16940 17602 16996 17612
rect 17052 17108 17108 20750
rect 17724 20804 17780 21308
rect 17836 20916 17892 23548
rect 17948 23154 18004 23884
rect 18060 23826 18116 23838
rect 18060 23774 18062 23826
rect 18114 23774 18116 23826
rect 18060 23492 18116 23774
rect 18284 23828 18340 24220
rect 18284 23762 18340 23772
rect 18508 24722 18564 24734
rect 18508 24670 18510 24722
rect 18562 24670 18564 24722
rect 18060 23436 18340 23492
rect 18284 23378 18340 23436
rect 18284 23326 18286 23378
rect 18338 23326 18340 23378
rect 18284 23314 18340 23326
rect 18396 23380 18452 23390
rect 18508 23380 18564 24670
rect 18620 24724 18676 24892
rect 18620 24658 18676 24668
rect 18452 23324 18564 23380
rect 18396 23286 18452 23324
rect 18172 23268 18228 23278
rect 17948 23102 17950 23154
rect 18002 23102 18004 23154
rect 17948 23090 18004 23102
rect 18060 23266 18228 23268
rect 18060 23214 18174 23266
rect 18226 23214 18228 23266
rect 18060 23212 18228 23214
rect 18060 23044 18116 23212
rect 18172 23202 18228 23212
rect 18060 21924 18116 22988
rect 18060 21858 18116 21868
rect 18172 22932 18228 22942
rect 18172 22370 18228 22876
rect 18508 22820 18564 22830
rect 18564 22764 18676 22820
rect 18508 22754 18564 22764
rect 18172 22318 18174 22370
rect 18226 22318 18228 22370
rect 17948 21812 18004 21822
rect 17948 21588 18004 21756
rect 17948 21586 18116 21588
rect 17948 21534 17950 21586
rect 18002 21534 18116 21586
rect 17948 21532 18116 21534
rect 17948 21522 18004 21532
rect 17948 20916 18004 20926
rect 17836 20860 17948 20916
rect 17948 20822 18004 20860
rect 17612 20244 17668 20254
rect 17724 20244 17780 20748
rect 17612 20242 17780 20244
rect 17612 20190 17614 20242
rect 17666 20190 17780 20242
rect 17612 20188 17780 20190
rect 18060 20188 18116 21532
rect 17612 20178 17668 20188
rect 17388 20132 17444 20142
rect 17164 19348 17220 19358
rect 17164 18788 17220 19292
rect 17276 19236 17332 19246
rect 17388 19236 17444 20076
rect 17836 20132 17892 20142
rect 17612 20020 17668 20030
rect 17500 19908 17556 19918
rect 17500 19814 17556 19852
rect 17276 19234 17444 19236
rect 17276 19182 17278 19234
rect 17330 19182 17444 19234
rect 17276 19180 17444 19182
rect 17276 19170 17332 19180
rect 17388 19012 17444 19022
rect 17388 18918 17444 18956
rect 17500 19010 17556 19022
rect 17500 18958 17502 19010
rect 17554 18958 17556 19010
rect 17164 18732 17444 18788
rect 17388 17780 17444 18732
rect 17500 18564 17556 18958
rect 17612 18674 17668 19964
rect 17836 20018 17892 20076
rect 17836 19966 17838 20018
rect 17890 19966 17892 20018
rect 17836 19954 17892 19966
rect 17948 20132 18116 20188
rect 17836 19346 17892 19358
rect 17836 19294 17838 19346
rect 17890 19294 17892 19346
rect 17836 19234 17892 19294
rect 17836 19182 17838 19234
rect 17890 19182 17892 19234
rect 17836 19170 17892 19182
rect 17612 18622 17614 18674
rect 17666 18622 17668 18674
rect 17612 18610 17668 18622
rect 17500 18498 17556 18508
rect 17724 18452 17780 18462
rect 17724 18358 17780 18396
rect 17836 18450 17892 18462
rect 17836 18398 17838 18450
rect 17890 18398 17892 18450
rect 17052 17042 17108 17052
rect 17164 17778 17444 17780
rect 17164 17726 17390 17778
rect 17442 17726 17444 17778
rect 17164 17724 17444 17726
rect 16828 16996 16884 17006
rect 16828 16770 16884 16940
rect 16828 16718 16830 16770
rect 16882 16718 16884 16770
rect 16828 16706 16884 16718
rect 17164 16324 17220 17724
rect 17388 17714 17444 17724
rect 17500 18340 17556 18350
rect 17500 17556 17556 18284
rect 16828 16268 17164 16324
rect 16828 16210 16884 16268
rect 17164 16230 17220 16268
rect 17388 17500 17556 17556
rect 17836 17556 17892 18398
rect 16828 16158 16830 16210
rect 16882 16158 16884 16210
rect 16828 16146 16884 16158
rect 16604 15426 16772 15428
rect 16604 15374 16606 15426
rect 16658 15374 16772 15426
rect 16604 15372 16772 15374
rect 16604 15362 16660 15372
rect 16716 15204 16772 15372
rect 17164 15986 17220 15998
rect 17164 15934 17166 15986
rect 17218 15934 17220 15986
rect 16492 15092 16660 15148
rect 16716 15138 16772 15148
rect 16828 15314 16884 15326
rect 16828 15262 16830 15314
rect 16882 15262 16884 15314
rect 16828 15148 16884 15262
rect 17164 15316 17220 15934
rect 17276 15876 17332 15886
rect 17276 15782 17332 15820
rect 16828 15092 16996 15148
rect 16044 14590 16046 14642
rect 16098 14590 16100 14642
rect 16044 14578 16100 14590
rect 14700 13806 14702 13858
rect 14754 13806 14756 13858
rect 14700 13794 14756 13806
rect 15260 14530 15316 14542
rect 15260 14478 15262 14530
rect 15314 14478 15316 14530
rect 14028 13746 14084 13758
rect 14028 13694 14030 13746
rect 14082 13694 14084 13746
rect 14028 13636 14084 13694
rect 14028 13570 14084 13580
rect 15260 13636 15316 14478
rect 15260 13570 15316 13580
rect 16604 12404 16660 15092
rect 16940 13860 16996 15092
rect 17164 15092 17220 15260
rect 17276 15092 17332 15102
rect 17164 15090 17332 15092
rect 17164 15038 17278 15090
rect 17330 15038 17332 15090
rect 17164 15036 17332 15038
rect 17276 15026 17332 15036
rect 17388 14532 17444 17500
rect 17836 17490 17892 17500
rect 17948 17778 18004 20132
rect 18060 20020 18116 20030
rect 18060 19926 18116 19964
rect 18172 19796 18228 22318
rect 18620 22370 18676 22764
rect 18620 22318 18622 22370
rect 18674 22318 18676 22370
rect 18620 22306 18676 22318
rect 18508 22258 18564 22270
rect 18508 22206 18510 22258
rect 18562 22206 18564 22258
rect 18284 21810 18340 21822
rect 18284 21758 18286 21810
rect 18338 21758 18340 21810
rect 18284 21588 18340 21758
rect 18284 21522 18340 21532
rect 18508 21364 18564 22206
rect 18732 22148 18788 25116
rect 18844 24948 18900 27804
rect 18956 27076 19012 27916
rect 18956 27010 19012 27020
rect 19068 26964 19124 29372
rect 19180 29362 19236 29372
rect 19292 28418 19348 30268
rect 19404 29652 19460 32620
rect 19628 32564 19684 33180
rect 20300 33236 20356 33246
rect 20412 33236 20468 33292
rect 20300 33234 20468 33236
rect 20300 33182 20302 33234
rect 20354 33182 20468 33234
rect 20300 33180 20468 33182
rect 20300 33170 20356 33180
rect 20524 33124 20580 33134
rect 19836 32956 20100 32966
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 19836 32890 20100 32900
rect 19628 32562 20020 32564
rect 19628 32510 19630 32562
rect 19682 32510 20020 32562
rect 19628 32508 20020 32510
rect 19628 32498 19684 32508
rect 19964 32002 20020 32508
rect 20188 32562 20244 32574
rect 20412 32564 20468 32574
rect 20188 32510 20190 32562
rect 20242 32510 20244 32562
rect 20188 32452 20244 32510
rect 20188 32228 20244 32396
rect 19964 31950 19966 32002
rect 20018 31950 20020 32002
rect 19964 31938 20020 31950
rect 20076 32172 20244 32228
rect 20300 32562 20468 32564
rect 20300 32510 20414 32562
rect 20466 32510 20468 32562
rect 20300 32508 20468 32510
rect 20076 31780 20132 32172
rect 20188 32004 20244 32014
rect 20300 32004 20356 32508
rect 20412 32498 20468 32508
rect 20188 32002 20356 32004
rect 20188 31950 20190 32002
rect 20242 31950 20356 32002
rect 20188 31948 20356 31950
rect 20188 31938 20244 31948
rect 20076 31724 20244 31780
rect 19836 31388 20100 31398
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 19836 31322 20100 31332
rect 20076 30994 20132 31006
rect 20076 30942 20078 30994
rect 20130 30942 20132 30994
rect 19628 30884 19684 30894
rect 19628 30790 19684 30828
rect 20076 30548 20132 30942
rect 20076 30482 20132 30492
rect 19404 29586 19460 29596
rect 19628 30212 19684 30222
rect 19292 28366 19294 28418
rect 19346 28366 19348 28418
rect 19180 28084 19236 28094
rect 19180 27412 19236 28028
rect 19180 27242 19236 27356
rect 19180 27190 19182 27242
rect 19234 27190 19236 27242
rect 19180 27178 19236 27190
rect 19292 27076 19348 28366
rect 19628 28084 19684 30156
rect 20076 30100 20132 30110
rect 20188 30100 20244 31724
rect 20076 30098 20244 30100
rect 20076 30046 20078 30098
rect 20130 30046 20244 30098
rect 20076 30044 20244 30046
rect 20076 30034 20132 30044
rect 19836 29820 20100 29830
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 19836 29754 20100 29764
rect 19740 29652 19796 29662
rect 19740 29538 19796 29596
rect 19740 29486 19742 29538
rect 19794 29486 19796 29538
rect 19740 29474 19796 29486
rect 20188 29428 20244 30044
rect 20300 29540 20356 31948
rect 20412 31892 20468 31902
rect 20412 31798 20468 31836
rect 20524 31220 20580 33068
rect 20636 31780 20692 33292
rect 20748 33234 20804 33246
rect 20748 33182 20750 33234
rect 20802 33182 20804 33234
rect 20748 32116 20804 33182
rect 20860 32786 20916 33740
rect 21308 33684 21364 33966
rect 21084 33628 21308 33684
rect 20860 32734 20862 32786
rect 20914 32734 20916 32786
rect 20860 32722 20916 32734
rect 20972 33572 21028 33582
rect 20972 32786 21028 33516
rect 20972 32734 20974 32786
rect 21026 32734 21028 32786
rect 20972 32722 21028 32734
rect 20748 32050 20804 32060
rect 20748 31892 20804 31902
rect 21084 31892 21140 33628
rect 21308 33618 21364 33628
rect 21308 33124 21364 33134
rect 21196 32674 21252 32686
rect 21196 32622 21198 32674
rect 21250 32622 21252 32674
rect 21196 32004 21252 32622
rect 21308 32674 21364 33068
rect 21308 32622 21310 32674
rect 21362 32622 21364 32674
rect 21308 32610 21364 32622
rect 21196 31938 21252 31948
rect 20748 31890 21140 31892
rect 20748 31838 20750 31890
rect 20802 31838 21140 31890
rect 20748 31836 21140 31838
rect 20748 31826 20804 31836
rect 20636 31686 20692 31724
rect 20748 31668 20804 31678
rect 20412 31164 20580 31220
rect 20636 31220 20692 31230
rect 20412 30212 20468 31164
rect 20524 30996 20580 31006
rect 20524 30902 20580 30940
rect 20636 30994 20692 31164
rect 20636 30942 20638 30994
rect 20690 30942 20692 30994
rect 20636 30930 20692 30942
rect 20748 30772 20804 31612
rect 20972 31668 21028 31678
rect 21308 31668 21364 31678
rect 20972 31106 21028 31612
rect 20972 31054 20974 31106
rect 21026 31054 21028 31106
rect 20972 31042 21028 31054
rect 21084 31666 21364 31668
rect 21084 31614 21310 31666
rect 21362 31614 21364 31666
rect 21084 31612 21364 31614
rect 20412 30118 20468 30156
rect 20636 30716 20804 30772
rect 20860 30882 20916 30894
rect 20860 30830 20862 30882
rect 20914 30830 20916 30882
rect 20300 29484 20580 29540
rect 20188 29372 20468 29428
rect 20300 29092 20356 29102
rect 19852 28756 19908 28766
rect 19852 28662 19908 28700
rect 20300 28754 20356 29036
rect 20300 28702 20302 28754
rect 20354 28702 20356 28754
rect 19836 28252 20100 28262
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 19836 28186 20100 28196
rect 19628 28028 19908 28084
rect 19068 26898 19124 26908
rect 19180 27020 19348 27076
rect 19404 27858 19460 27870
rect 19404 27806 19406 27858
rect 19458 27806 19460 27858
rect 19068 26740 19124 26750
rect 19068 26514 19124 26684
rect 19068 26462 19070 26514
rect 19122 26462 19124 26514
rect 19068 26450 19124 26462
rect 18956 26404 19012 26414
rect 18956 26310 19012 26348
rect 19068 25508 19124 25518
rect 19180 25508 19236 27020
rect 19404 26908 19460 27806
rect 19516 27412 19572 27422
rect 19516 27074 19572 27356
rect 19516 27022 19518 27074
rect 19570 27022 19572 27074
rect 19516 27010 19572 27022
rect 19292 26852 19460 26908
rect 19852 26962 19908 28028
rect 20188 27076 20244 27086
rect 20188 26982 20244 27020
rect 19852 26910 19854 26962
rect 19906 26910 19908 26962
rect 19852 26898 19908 26910
rect 19516 26852 19572 26862
rect 19292 25618 19348 26852
rect 19516 26514 19572 26796
rect 20300 26852 20356 28702
rect 20300 26786 20356 26796
rect 20188 26740 20244 26750
rect 19836 26684 20100 26694
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 19836 26618 20100 26628
rect 19516 26462 19518 26514
rect 19570 26462 19572 26514
rect 19516 26450 19572 26462
rect 20188 26402 20244 26684
rect 20300 26516 20356 26526
rect 20300 26422 20356 26460
rect 20188 26350 20190 26402
rect 20242 26350 20244 26402
rect 20188 26338 20244 26350
rect 19628 26292 19684 26302
rect 19628 26290 19908 26292
rect 19628 26238 19630 26290
rect 19682 26238 19908 26290
rect 19628 26236 19908 26238
rect 19628 26226 19684 26236
rect 19516 26068 19572 26078
rect 19740 26068 19796 26078
rect 19292 25566 19294 25618
rect 19346 25566 19348 25618
rect 19292 25554 19348 25566
rect 19404 26066 19572 26068
rect 19404 26014 19518 26066
rect 19570 26014 19572 26066
rect 19404 26012 19572 26014
rect 19124 25452 19236 25508
rect 19068 25442 19124 25452
rect 19292 25396 19348 25406
rect 19292 25302 19348 25340
rect 19404 25394 19460 26012
rect 19516 26002 19572 26012
rect 19628 26012 19740 26068
rect 19404 25342 19406 25394
rect 19458 25342 19460 25394
rect 19404 25330 19460 25342
rect 19516 25394 19572 25406
rect 19516 25342 19518 25394
rect 19570 25342 19572 25394
rect 19068 25284 19124 25294
rect 19068 25282 19236 25284
rect 19068 25230 19070 25282
rect 19122 25230 19236 25282
rect 19068 25228 19236 25230
rect 19068 25218 19124 25228
rect 18844 23938 18900 24892
rect 18956 24724 19012 24734
rect 18956 24630 19012 24668
rect 19180 24724 19236 25228
rect 19404 25172 19460 25182
rect 19404 24946 19460 25116
rect 19516 25060 19572 25342
rect 19516 24994 19572 25004
rect 19404 24894 19406 24946
rect 19458 24894 19460 24946
rect 19404 24882 19460 24894
rect 19516 24834 19572 24846
rect 19516 24782 19518 24834
rect 19570 24782 19572 24834
rect 19292 24724 19348 24734
rect 19180 24722 19348 24724
rect 19180 24670 19294 24722
rect 19346 24670 19348 24722
rect 19180 24668 19348 24670
rect 18844 23886 18846 23938
rect 18898 23886 18900 23938
rect 18844 23874 18900 23886
rect 18956 24052 19012 24062
rect 18508 21298 18564 21308
rect 18620 22092 18788 22148
rect 18844 22596 18900 22606
rect 18620 21140 18676 22092
rect 18732 21812 18788 21822
rect 18732 21718 18788 21756
rect 18508 21084 18676 21140
rect 18284 20578 18340 20590
rect 18284 20526 18286 20578
rect 18338 20526 18340 20578
rect 18284 20468 18340 20526
rect 18284 20402 18340 20412
rect 18060 19740 18228 19796
rect 18396 20020 18452 20030
rect 18060 18340 18116 19740
rect 18396 19572 18452 19964
rect 18396 19506 18452 19516
rect 18172 19346 18228 19358
rect 18172 19294 18174 19346
rect 18226 19294 18228 19346
rect 18172 19236 18228 19294
rect 18172 19180 18340 19236
rect 18060 18274 18116 18284
rect 18284 18450 18340 19180
rect 18284 18398 18286 18450
rect 18338 18398 18340 18450
rect 18284 17892 18340 18398
rect 17948 17726 17950 17778
rect 18002 17726 18004 17778
rect 17948 17444 18004 17726
rect 17948 17378 18004 17388
rect 18060 17836 18284 17892
rect 17500 17108 17556 17118
rect 17500 17014 17556 17052
rect 18060 17106 18116 17836
rect 18284 17826 18340 17836
rect 18060 17054 18062 17106
rect 18114 17054 18116 17106
rect 18060 17042 18116 17054
rect 18172 17442 18228 17454
rect 18172 17390 18174 17442
rect 18226 17390 18228 17442
rect 18172 16996 18228 17390
rect 18172 16930 18228 16940
rect 17612 16324 17668 16334
rect 17500 16212 17556 16222
rect 17500 16098 17556 16156
rect 17500 16046 17502 16098
rect 17554 16046 17556 16098
rect 17500 16034 17556 16046
rect 17612 15538 17668 16268
rect 17724 15988 17780 15998
rect 18508 15988 18564 21084
rect 18620 19906 18676 19918
rect 18620 19854 18622 19906
rect 18674 19854 18676 19906
rect 18620 18564 18676 19854
rect 18844 19908 18900 22540
rect 18956 21700 19012 23996
rect 19068 23380 19124 23390
rect 19180 23380 19236 24668
rect 19292 24658 19348 24668
rect 19516 24388 19572 24782
rect 19628 24834 19684 26012
rect 19740 26002 19796 26012
rect 19852 25396 19908 26236
rect 20300 26180 20356 26190
rect 20300 26066 20356 26124
rect 20300 26014 20302 26066
rect 20354 26014 20356 26066
rect 20300 26002 20356 26014
rect 20412 25844 20468 29372
rect 20524 26962 20580 29484
rect 20636 29204 20692 30716
rect 20860 30660 20916 30830
rect 20860 30594 20916 30604
rect 20748 30212 20804 30222
rect 20748 30118 20804 30156
rect 20748 29652 20804 29662
rect 20748 29558 20804 29596
rect 21084 29540 21140 31612
rect 21308 31602 21364 31612
rect 21420 31556 21476 34524
rect 21532 33908 21588 33918
rect 21532 33814 21588 33852
rect 21756 33796 21812 34638
rect 22204 35364 22260 35374
rect 21868 34356 21924 34366
rect 21868 34354 22148 34356
rect 21868 34302 21870 34354
rect 21922 34302 22148 34354
rect 21868 34300 22148 34302
rect 21868 34290 21924 34300
rect 22092 33796 22148 34300
rect 21756 33740 22036 33796
rect 21644 33348 21700 33358
rect 21980 33348 22036 33740
rect 22092 33730 22148 33740
rect 22092 33348 22148 33358
rect 21980 33292 22092 33348
rect 21420 31490 21476 31500
rect 21532 31890 21588 31902
rect 21532 31838 21534 31890
rect 21586 31838 21588 31890
rect 21532 31780 21588 31838
rect 21532 30994 21588 31724
rect 21532 30942 21534 30994
rect 21586 30942 21588 30994
rect 21532 30930 21588 30942
rect 21420 30210 21476 30222
rect 21420 30158 21422 30210
rect 21474 30158 21476 30210
rect 21420 30100 21476 30158
rect 21420 30034 21476 30044
rect 20972 29484 21588 29540
rect 20972 29428 21028 29484
rect 20636 29138 20692 29148
rect 20748 29426 21028 29428
rect 20748 29374 20974 29426
rect 21026 29374 21028 29426
rect 20748 29372 21028 29374
rect 20748 28642 20804 29372
rect 20972 29362 21028 29372
rect 21420 29204 21476 29214
rect 21420 28754 21476 29148
rect 21420 28702 21422 28754
rect 21474 28702 21476 28754
rect 21420 28690 21476 28702
rect 20748 28590 20750 28642
rect 20802 28590 20804 28642
rect 20748 28578 20804 28590
rect 21532 27746 21588 29484
rect 21644 29092 21700 33292
rect 22092 33254 22148 33292
rect 22092 32564 22148 32574
rect 21980 32450 22036 32462
rect 21980 32398 21982 32450
rect 22034 32398 22036 32450
rect 21644 29026 21700 29036
rect 21756 32116 21812 32126
rect 21980 32116 22036 32398
rect 21756 30100 21812 32060
rect 21868 32060 22036 32116
rect 21868 31892 21924 32060
rect 21868 31826 21924 31836
rect 21980 31780 22036 31790
rect 21980 31220 22036 31724
rect 21980 31154 22036 31164
rect 21868 30882 21924 30894
rect 21868 30830 21870 30882
rect 21922 30830 21924 30882
rect 21868 30212 21924 30830
rect 21868 30118 21924 30156
rect 21756 28756 21812 30044
rect 22092 29652 22148 32508
rect 22204 30434 22260 35308
rect 22652 35364 22708 36990
rect 22764 37044 22820 37436
rect 22876 37268 22932 44044
rect 23436 44044 23716 44100
rect 23100 42754 23156 42766
rect 23100 42702 23102 42754
rect 23154 42702 23156 42754
rect 23100 41076 23156 42702
rect 23436 42642 23492 44044
rect 23772 43652 23828 47740
rect 23996 47572 24052 47582
rect 23996 47478 24052 47516
rect 24108 47460 24164 47470
rect 24108 47068 24164 47404
rect 23996 47012 24164 47068
rect 24444 47124 24500 48188
rect 24668 48132 24724 48142
rect 24556 48020 24612 48030
rect 24556 47458 24612 47964
rect 24556 47406 24558 47458
rect 24610 47406 24612 47458
rect 24556 47394 24612 47406
rect 24668 47460 24724 48076
rect 24668 47394 24724 47404
rect 24444 47058 24500 47068
rect 24668 47236 24724 47246
rect 23884 46564 23940 46574
rect 23884 46470 23940 46508
rect 23996 46004 24052 47012
rect 24668 46898 24724 47180
rect 24668 46846 24670 46898
rect 24722 46846 24724 46898
rect 24668 46834 24724 46846
rect 24332 46676 24388 46686
rect 23884 45948 24052 46004
rect 24220 46674 24388 46676
rect 24220 46622 24334 46674
rect 24386 46622 24388 46674
rect 24220 46620 24388 46622
rect 23884 43876 23940 45948
rect 23996 45780 24052 45790
rect 24220 45780 24276 46620
rect 24332 46610 24388 46620
rect 24780 45892 24836 52444
rect 25228 52276 25284 52286
rect 24892 52274 25284 52276
rect 24892 52222 25230 52274
rect 25282 52222 25284 52274
rect 24892 52220 25284 52222
rect 24892 50706 24948 52220
rect 25228 52210 25284 52220
rect 25340 52050 25396 52444
rect 25788 52388 25844 52398
rect 25676 52332 25788 52388
rect 25340 51998 25342 52050
rect 25394 51998 25396 52050
rect 25340 51986 25396 51998
rect 25564 52050 25620 52062
rect 25564 51998 25566 52050
rect 25618 51998 25620 52050
rect 25564 51602 25620 51998
rect 25564 51550 25566 51602
rect 25618 51550 25620 51602
rect 25564 51538 25620 51550
rect 25676 51380 25732 52332
rect 25788 52322 25844 52332
rect 26348 52388 26404 53454
rect 26348 52322 26404 52332
rect 26908 53452 27020 53508
rect 26908 52388 26964 53452
rect 27020 53414 27076 53452
rect 26908 52322 26964 52332
rect 26796 52274 26852 52286
rect 26796 52222 26798 52274
rect 26850 52222 26852 52274
rect 26460 52164 26516 52174
rect 24892 50654 24894 50706
rect 24946 50654 24948 50706
rect 24892 50642 24948 50654
rect 25564 51324 25732 51380
rect 26012 52162 26516 52164
rect 26012 52110 26462 52162
rect 26514 52110 26516 52162
rect 26012 52108 26516 52110
rect 26012 51378 26068 52108
rect 26012 51326 26014 51378
rect 26066 51326 26068 51378
rect 25452 49698 25508 49710
rect 25452 49646 25454 49698
rect 25506 49646 25508 49698
rect 25340 49140 25396 49150
rect 25340 49046 25396 49084
rect 25452 48804 25508 49646
rect 25564 49028 25620 51324
rect 26012 51314 26068 51326
rect 25676 51156 25732 51166
rect 25676 49700 25732 51100
rect 26236 50484 26292 50494
rect 25676 49634 25732 49644
rect 25788 49698 25844 49710
rect 25788 49646 25790 49698
rect 25842 49646 25844 49698
rect 25564 48962 25620 48972
rect 25676 48804 25732 48814
rect 25452 48802 25732 48804
rect 25452 48750 25678 48802
rect 25730 48750 25732 48802
rect 25452 48748 25732 48750
rect 25340 48132 25396 48142
rect 25452 48132 25508 48748
rect 25676 48738 25732 48748
rect 25788 48580 25844 49646
rect 25900 49588 25956 49598
rect 25900 49494 25956 49532
rect 26236 49028 26292 50428
rect 26460 50428 26516 52108
rect 26796 51604 26852 52222
rect 27132 52164 27188 53564
rect 27244 53730 27300 53742
rect 27244 53678 27246 53730
rect 27298 53678 27300 53730
rect 27244 53284 27300 53678
rect 27356 53620 27412 55244
rect 27580 55186 27636 55198
rect 28028 55188 28084 55198
rect 27580 55134 27582 55186
rect 27634 55134 27636 55186
rect 27468 55074 27524 55086
rect 27468 55022 27470 55074
rect 27522 55022 27524 55074
rect 27468 54740 27524 55022
rect 27468 54674 27524 54684
rect 27468 54516 27524 54526
rect 27468 53732 27524 54460
rect 27580 53844 27636 55134
rect 27804 55186 28084 55188
rect 27804 55134 28030 55186
rect 28082 55134 28084 55186
rect 27804 55132 28084 55134
rect 27692 54404 27748 54414
rect 27804 54404 27860 55132
rect 28028 55122 28084 55132
rect 28364 55188 28420 55198
rect 28588 55188 28644 55198
rect 28364 55186 28532 55188
rect 28364 55134 28366 55186
rect 28418 55134 28532 55186
rect 28364 55132 28532 55134
rect 28364 55122 28420 55132
rect 28252 55076 28308 55086
rect 28252 54982 28308 55020
rect 27692 54402 27860 54404
rect 27692 54350 27694 54402
rect 27746 54350 27860 54402
rect 27692 54348 27860 54350
rect 27692 54338 27748 54348
rect 27692 53844 27748 53854
rect 27580 53842 27748 53844
rect 27580 53790 27694 53842
rect 27746 53790 27748 53842
rect 27580 53788 27748 53790
rect 27692 53778 27748 53788
rect 27804 53732 27860 54348
rect 27468 53676 27636 53732
rect 27356 53564 27524 53620
rect 27356 53284 27412 53294
rect 27244 53228 27356 53284
rect 27356 52386 27412 53228
rect 27468 53170 27524 53564
rect 27580 53618 27636 53676
rect 27916 54740 27972 54750
rect 27916 53732 27972 54684
rect 28028 54516 28084 54526
rect 28028 54404 28084 54460
rect 28028 54402 28308 54404
rect 28028 54350 28030 54402
rect 28082 54350 28308 54402
rect 28028 54348 28308 54350
rect 28028 54338 28084 54348
rect 28028 53732 28084 53742
rect 27916 53730 28084 53732
rect 27916 53678 28030 53730
rect 28082 53678 28084 53730
rect 27916 53676 28084 53678
rect 27804 53666 27860 53676
rect 28028 53666 28084 53676
rect 27580 53566 27582 53618
rect 27634 53566 27636 53618
rect 27580 53554 27636 53566
rect 27692 53620 27748 53630
rect 27692 53508 27748 53564
rect 28252 53618 28308 54348
rect 28252 53566 28254 53618
rect 28306 53566 28308 53618
rect 28252 53554 28308 53566
rect 28364 53618 28420 53630
rect 28364 53566 28366 53618
rect 28418 53566 28420 53618
rect 27804 53508 27860 53518
rect 27692 53506 28196 53508
rect 27692 53454 27806 53506
rect 27858 53454 28196 53506
rect 27692 53452 28196 53454
rect 27804 53442 27860 53452
rect 28140 53396 28196 53452
rect 28364 53396 28420 53566
rect 28140 53340 28420 53396
rect 28476 53284 28532 55132
rect 28588 55186 29092 55188
rect 28588 55134 28590 55186
rect 28642 55134 29092 55186
rect 28588 55132 29092 55134
rect 28588 55122 28644 55132
rect 29036 54292 29092 55132
rect 29148 55186 29204 57260
rect 30156 55972 30212 55982
rect 30268 55972 30324 59200
rect 30156 55970 30324 55972
rect 30156 55918 30158 55970
rect 30210 55918 30324 55970
rect 30156 55916 30324 55918
rect 31612 56082 31668 56094
rect 31612 56030 31614 56082
rect 31666 56030 31668 56082
rect 30156 55906 30212 55916
rect 29148 55134 29150 55186
rect 29202 55134 29204 55186
rect 29148 55122 29204 55134
rect 30044 55298 30100 55310
rect 30044 55246 30046 55298
rect 30098 55246 30100 55298
rect 30044 54404 30100 55246
rect 30716 55188 30772 55198
rect 30716 55094 30772 55132
rect 30156 55076 30212 55086
rect 30156 54626 30212 55020
rect 30156 54574 30158 54626
rect 30210 54574 30212 54626
rect 30156 54562 30212 54574
rect 30044 54338 30100 54348
rect 30940 54514 30996 54526
rect 30940 54462 30942 54514
rect 30994 54462 30996 54514
rect 30940 54404 30996 54462
rect 30940 54338 30996 54348
rect 31388 54404 31444 54414
rect 31612 54404 31668 56030
rect 31836 55412 31892 59200
rect 32172 55970 32228 55982
rect 32172 55918 32174 55970
rect 32226 55918 32228 55970
rect 32172 55524 32228 55918
rect 32172 55458 32228 55468
rect 31836 55346 31892 55356
rect 32844 55410 32900 55422
rect 32844 55358 32846 55410
rect 32898 55358 32900 55410
rect 32844 55300 32900 55358
rect 33180 55300 33236 55310
rect 32844 55298 33236 55300
rect 32844 55246 33182 55298
rect 33234 55246 33236 55298
rect 32844 55244 33236 55246
rect 33180 55234 33236 55244
rect 32508 55188 32564 55198
rect 31836 54404 31892 54414
rect 31612 54402 31892 54404
rect 31612 54350 31838 54402
rect 31890 54350 31892 54402
rect 31612 54348 31892 54350
rect 31388 54310 31444 54348
rect 29036 54236 29316 54292
rect 29260 53842 29316 54236
rect 31836 53956 31892 54348
rect 31836 53890 31892 53900
rect 32508 54402 32564 55132
rect 32508 54350 32510 54402
rect 32562 54350 32564 54402
rect 29260 53790 29262 53842
rect 29314 53790 29316 53842
rect 29260 53778 29316 53790
rect 32508 53844 32564 54350
rect 32508 53778 32564 53788
rect 33068 54402 33124 54414
rect 33068 54350 33070 54402
rect 33122 54350 33124 54402
rect 29148 53732 29204 53742
rect 29148 53638 29204 53676
rect 32956 53732 33012 53742
rect 32956 53638 33012 53676
rect 28476 53218 28532 53228
rect 28588 53620 28644 53630
rect 27468 53118 27470 53170
rect 27522 53118 27524 53170
rect 27468 53106 27524 53118
rect 27356 52334 27358 52386
rect 27410 52334 27412 52386
rect 27356 52322 27412 52334
rect 26796 51538 26852 51548
rect 26908 52108 27188 52164
rect 27244 52162 27300 52174
rect 27244 52110 27246 52162
rect 27298 52110 27300 52162
rect 26908 50820 26964 52108
rect 26796 50764 26964 50820
rect 27020 51492 27076 51502
rect 26796 50484 26852 50764
rect 27020 50708 27076 51436
rect 27244 50820 27300 52110
rect 28028 51604 28084 51614
rect 28028 51510 28084 51548
rect 28140 51492 28196 51502
rect 28140 51398 28196 51436
rect 27356 51268 27412 51278
rect 27916 51268 27972 51278
rect 27356 51266 27972 51268
rect 27356 51214 27358 51266
rect 27410 51214 27918 51266
rect 27970 51214 27972 51266
rect 27356 51212 27972 51214
rect 27356 51202 27412 51212
rect 27468 50820 27524 50830
rect 27244 50818 27524 50820
rect 27244 50766 27470 50818
rect 27522 50766 27524 50818
rect 27244 50764 27524 50766
rect 27468 50754 27524 50764
rect 27020 50706 27412 50708
rect 27020 50654 27022 50706
rect 27074 50654 27412 50706
rect 27020 50652 27412 50654
rect 27020 50642 27076 50652
rect 27356 50484 27412 50652
rect 27580 50596 27636 50606
rect 27804 50596 27860 51212
rect 27916 51202 27972 51212
rect 28028 51268 28084 51278
rect 28028 50708 28084 51212
rect 28588 50818 28644 53564
rect 30828 53620 30884 53630
rect 30828 53526 30884 53564
rect 31052 53618 31108 53630
rect 31052 53566 31054 53618
rect 31106 53566 31108 53618
rect 29372 53508 29428 53518
rect 29260 53506 29428 53508
rect 29260 53454 29374 53506
rect 29426 53454 29428 53506
rect 29260 53452 29428 53454
rect 29260 53284 29316 53452
rect 29372 53442 29428 53452
rect 29596 53508 29652 53518
rect 29596 53414 29652 53452
rect 30268 53508 30324 53518
rect 30268 53414 30324 53452
rect 29260 53218 29316 53228
rect 29372 53060 29428 53070
rect 29372 53058 29540 53060
rect 29372 53006 29374 53058
rect 29426 53006 29540 53058
rect 29372 53004 29540 53006
rect 29372 52994 29428 53004
rect 29260 52946 29316 52958
rect 29260 52894 29262 52946
rect 29314 52894 29316 52946
rect 29260 52164 29316 52894
rect 28924 51378 28980 51390
rect 28924 51326 28926 51378
rect 28978 51326 28980 51378
rect 28588 50766 28590 50818
rect 28642 50766 28644 50818
rect 28588 50754 28644 50766
rect 28700 51266 28756 51278
rect 28700 51214 28702 51266
rect 28754 51214 28756 51266
rect 28028 50614 28084 50652
rect 28700 50708 28756 51214
rect 28700 50642 28756 50652
rect 27580 50594 27860 50596
rect 27580 50542 27582 50594
rect 27634 50542 27860 50594
rect 27580 50540 27860 50542
rect 27580 50530 27636 50540
rect 27468 50484 27524 50494
rect 27356 50482 27524 50484
rect 27356 50430 27470 50482
rect 27522 50430 27524 50482
rect 27356 50428 27524 50430
rect 26460 50372 26628 50428
rect 26796 50418 26852 50428
rect 27468 50418 27524 50428
rect 26460 49812 26516 49822
rect 26460 49250 26516 49756
rect 26572 49698 26628 50372
rect 26572 49646 26574 49698
rect 26626 49646 26628 49698
rect 26572 49634 26628 49646
rect 26684 49922 26740 49934
rect 26684 49870 26686 49922
rect 26738 49870 26740 49922
rect 26460 49198 26462 49250
rect 26514 49198 26516 49250
rect 26460 49186 26516 49198
rect 26348 49028 26404 49038
rect 26012 49026 26404 49028
rect 26012 48974 26350 49026
rect 26402 48974 26404 49026
rect 26012 48972 26404 48974
rect 26012 48914 26068 48972
rect 26348 48962 26404 48972
rect 26460 49028 26516 49038
rect 26516 48972 26628 49028
rect 26460 48962 26516 48972
rect 26012 48862 26014 48914
rect 26066 48862 26068 48914
rect 26012 48850 26068 48862
rect 26460 48804 26516 48814
rect 26460 48710 26516 48748
rect 25788 48524 26292 48580
rect 26236 48354 26292 48524
rect 26236 48302 26238 48354
rect 26290 48302 26292 48354
rect 26236 48290 26292 48302
rect 25564 48244 25620 48254
rect 26572 48244 26628 48972
rect 25564 48150 25620 48188
rect 26460 48242 26628 48244
rect 26460 48190 26574 48242
rect 26626 48190 26628 48242
rect 26460 48188 26628 48190
rect 25396 48076 25508 48132
rect 25340 48038 25396 48076
rect 25004 47460 25060 47470
rect 24052 45724 24276 45780
rect 24668 45836 24836 45892
rect 24892 47404 25004 47460
rect 23996 45686 24052 45724
rect 24332 45666 24388 45678
rect 24332 45614 24334 45666
rect 24386 45614 24388 45666
rect 24332 45220 24388 45614
rect 24332 45154 24388 45164
rect 24444 45666 24500 45678
rect 24444 45614 24446 45666
rect 24498 45614 24500 45666
rect 24444 44996 24500 45614
rect 23996 44940 24500 44996
rect 24556 45668 24612 45678
rect 23996 44322 24052 44940
rect 23996 44270 23998 44322
rect 24050 44270 24052 44322
rect 23996 44258 24052 44270
rect 24556 44324 24612 45612
rect 24668 45220 24724 45836
rect 24668 45164 24836 45220
rect 24668 44996 24724 45006
rect 24668 44902 24724 44940
rect 24556 44258 24612 44268
rect 24668 44548 24724 44558
rect 24668 44434 24724 44492
rect 24668 44382 24670 44434
rect 24722 44382 24724 44434
rect 23884 43820 24164 43876
rect 23996 43652 24052 43662
rect 23772 43596 23996 43652
rect 23996 43586 24052 43596
rect 23996 42868 24052 42878
rect 23772 42644 23828 42654
rect 23436 42590 23438 42642
rect 23490 42590 23492 42642
rect 23436 42578 23492 42590
rect 23548 42642 23828 42644
rect 23548 42590 23774 42642
rect 23826 42590 23828 42642
rect 23548 42588 23828 42590
rect 23548 42084 23604 42588
rect 23772 42578 23828 42588
rect 23996 42642 24052 42812
rect 23996 42590 23998 42642
rect 24050 42590 24052 42642
rect 23996 42578 24052 42590
rect 23436 42028 23604 42084
rect 23884 42530 23940 42542
rect 23884 42478 23886 42530
rect 23938 42478 23940 42530
rect 23884 42084 23940 42478
rect 23324 41076 23380 41086
rect 23100 41074 23380 41076
rect 23100 41022 23326 41074
rect 23378 41022 23380 41074
rect 23100 41020 23380 41022
rect 23324 39396 23380 41020
rect 23436 40962 23492 42028
rect 23884 42018 23940 42028
rect 24108 41300 24164 43820
rect 24556 42978 24612 42990
rect 24556 42926 24558 42978
rect 24610 42926 24612 42978
rect 24556 42868 24612 42926
rect 24556 42774 24612 42812
rect 24220 41972 24276 41982
rect 24668 41972 24724 44382
rect 24780 42978 24836 45164
rect 24892 44546 24948 47404
rect 25004 47394 25060 47404
rect 25340 47348 25396 47358
rect 25340 47254 25396 47292
rect 25004 46900 25060 46910
rect 25004 45890 25060 46844
rect 25340 46900 25396 46910
rect 25340 46806 25396 46844
rect 26460 46900 26516 48188
rect 26572 48178 26628 48188
rect 26684 47796 26740 49870
rect 26796 49810 26852 49822
rect 26796 49758 26798 49810
rect 26850 49758 26852 49810
rect 26796 48020 26852 49758
rect 27356 49812 27412 49822
rect 27580 49812 27636 49822
rect 27356 49810 27524 49812
rect 27356 49758 27358 49810
rect 27410 49758 27524 49810
rect 27356 49756 27524 49758
rect 27356 49746 27412 49756
rect 27356 49140 27412 49150
rect 27356 49026 27412 49084
rect 27356 48974 27358 49026
rect 27410 48974 27412 49026
rect 27356 48962 27412 48974
rect 26796 47954 26852 47964
rect 26908 48242 26964 48254
rect 26908 48190 26910 48242
rect 26962 48190 26964 48242
rect 26908 47796 26964 48190
rect 27132 48244 27188 48254
rect 27356 48244 27412 48254
rect 27132 48242 27412 48244
rect 27132 48190 27134 48242
rect 27186 48190 27358 48242
rect 27410 48190 27412 48242
rect 27132 48188 27412 48190
rect 27132 48178 27188 48188
rect 27356 48178 27412 48188
rect 27020 48132 27076 48142
rect 27020 48038 27076 48076
rect 26684 47740 26964 47796
rect 26908 47460 26964 47740
rect 26908 47394 26964 47404
rect 27132 47796 27188 47806
rect 27468 47796 27524 49756
rect 27580 49718 27636 49756
rect 27580 48244 27636 48254
rect 27580 48242 27748 48244
rect 27580 48190 27582 48242
rect 27634 48190 27748 48242
rect 27580 48188 27748 48190
rect 27580 48178 27636 48188
rect 27132 47236 27188 47740
rect 27132 47170 27188 47180
rect 27244 47740 27524 47796
rect 26460 46898 26740 46900
rect 26460 46846 26462 46898
rect 26514 46846 26740 46898
rect 26460 46844 26740 46846
rect 26460 46834 26516 46844
rect 25788 46562 25844 46574
rect 25788 46510 25790 46562
rect 25842 46510 25844 46562
rect 25340 46116 25396 46126
rect 25004 45838 25006 45890
rect 25058 45838 25060 45890
rect 25004 45556 25060 45838
rect 25004 45490 25060 45500
rect 25228 46114 25396 46116
rect 25228 46062 25342 46114
rect 25394 46062 25396 46114
rect 25228 46060 25396 46062
rect 25004 45220 25060 45230
rect 25228 45220 25284 46060
rect 25340 46050 25396 46060
rect 25452 45780 25508 45790
rect 25676 45780 25732 45790
rect 25452 45778 25732 45780
rect 25452 45726 25454 45778
rect 25506 45726 25678 45778
rect 25730 45726 25732 45778
rect 25452 45724 25732 45726
rect 25452 45714 25508 45724
rect 25676 45714 25732 45724
rect 25340 45668 25396 45678
rect 25340 45574 25396 45612
rect 25452 45556 25508 45566
rect 25508 45500 25620 45556
rect 25452 45490 25508 45500
rect 25060 45164 25172 45220
rect 25228 45164 25396 45220
rect 25004 45154 25060 45164
rect 24892 44494 24894 44546
rect 24946 44494 24948 44546
rect 24892 44482 24948 44494
rect 25004 44996 25060 45006
rect 25116 44996 25172 45164
rect 25228 44996 25284 45006
rect 25116 44994 25284 44996
rect 25116 44942 25230 44994
rect 25282 44942 25284 44994
rect 25116 44940 25284 44942
rect 24892 44324 24948 44334
rect 24892 44230 24948 44268
rect 25004 43708 25060 44940
rect 25228 44930 25284 44940
rect 25340 44322 25396 45164
rect 25452 45108 25508 45118
rect 25452 44548 25508 45052
rect 25452 44482 25508 44492
rect 25340 44270 25342 44322
rect 25394 44270 25396 44322
rect 25340 44258 25396 44270
rect 25452 44324 25508 44334
rect 25340 43764 25396 43774
rect 25452 43764 25508 44268
rect 25340 43762 25508 43764
rect 25340 43710 25342 43762
rect 25394 43710 25508 43762
rect 25340 43708 25508 43710
rect 24780 42926 24782 42978
rect 24834 42926 24836 42978
rect 24780 42914 24836 42926
rect 24892 43652 24948 43662
rect 25004 43652 25284 43708
rect 25340 43698 25396 43708
rect 24220 41970 24388 41972
rect 24220 41918 24222 41970
rect 24274 41918 24388 41970
rect 24220 41916 24388 41918
rect 24220 41906 24276 41916
rect 23436 40910 23438 40962
rect 23490 40910 23492 40962
rect 23436 40898 23492 40910
rect 23996 41244 24164 41300
rect 24332 41300 24388 41916
rect 24668 41878 24724 41916
rect 24556 41300 24612 41310
rect 24332 41298 24612 41300
rect 24332 41246 24558 41298
rect 24610 41246 24612 41298
rect 24332 41244 24612 41246
rect 23884 40516 23940 40526
rect 23772 40460 23884 40516
rect 23772 40292 23828 40460
rect 23884 40422 23940 40460
rect 23996 40292 24052 41244
rect 24444 40404 24500 40414
rect 24444 40310 24500 40348
rect 23660 40236 23828 40292
rect 23884 40236 24052 40292
rect 23548 39508 23604 39518
rect 23548 39414 23604 39452
rect 23324 39330 23380 39340
rect 22988 38836 23044 38846
rect 22988 38742 23044 38780
rect 23212 38836 23268 38846
rect 23100 38050 23156 38062
rect 23100 37998 23102 38050
rect 23154 37998 23156 38050
rect 23100 37940 23156 37998
rect 23212 37940 23268 38780
rect 23324 37940 23380 37950
rect 23212 37938 23380 37940
rect 23212 37886 23326 37938
rect 23378 37886 23380 37938
rect 23212 37884 23380 37886
rect 23100 37874 23156 37884
rect 23324 37874 23380 37884
rect 22988 37492 23044 37502
rect 23548 37492 23604 37502
rect 23660 37492 23716 40236
rect 23772 39618 23828 39630
rect 23772 39566 23774 39618
rect 23826 39566 23828 39618
rect 23772 38836 23828 39566
rect 23772 38770 23828 38780
rect 22988 37490 23380 37492
rect 22988 37438 22990 37490
rect 23042 37438 23380 37490
rect 22988 37436 23380 37438
rect 22988 37426 23044 37436
rect 22876 37212 23156 37268
rect 22876 37044 22932 37054
rect 22764 37042 22932 37044
rect 22764 36990 22878 37042
rect 22930 36990 22932 37042
rect 22764 36988 22932 36990
rect 22876 36978 22932 36988
rect 22988 37044 23044 37054
rect 22652 35298 22708 35308
rect 22876 36482 22932 36494
rect 22876 36430 22878 36482
rect 22930 36430 22932 36482
rect 22876 35700 22932 36430
rect 22764 35252 22820 35262
rect 22764 34914 22820 35196
rect 22764 34862 22766 34914
rect 22818 34862 22820 34914
rect 22764 34850 22820 34862
rect 22316 34130 22372 34142
rect 22316 34078 22318 34130
rect 22370 34078 22372 34130
rect 22316 33572 22372 34078
rect 22876 34132 22932 35644
rect 22988 35698 23044 36988
rect 23100 36372 23156 37212
rect 23324 36594 23380 37436
rect 23548 37490 23716 37492
rect 23548 37438 23550 37490
rect 23602 37438 23716 37490
rect 23548 37436 23716 37438
rect 23772 37492 23828 37502
rect 23548 37426 23604 37436
rect 23324 36542 23326 36594
rect 23378 36542 23380 36594
rect 23324 36530 23380 36542
rect 23436 37266 23492 37278
rect 23436 37214 23438 37266
rect 23490 37214 23492 37266
rect 23436 37156 23492 37214
rect 23660 37268 23716 37278
rect 23772 37268 23828 37436
rect 23660 37266 23828 37268
rect 23660 37214 23662 37266
rect 23714 37214 23828 37266
rect 23660 37212 23828 37214
rect 23660 37202 23716 37212
rect 23100 36316 23380 36372
rect 22988 35646 22990 35698
rect 23042 35646 23044 35698
rect 22988 35634 23044 35646
rect 23212 34914 23268 34926
rect 23212 34862 23214 34914
rect 23266 34862 23268 34914
rect 23212 34804 23268 34862
rect 23212 34244 23268 34748
rect 23212 34178 23268 34188
rect 23100 34132 23156 34142
rect 22876 34130 23156 34132
rect 22876 34078 23102 34130
rect 23154 34078 23156 34130
rect 22876 34076 23156 34078
rect 23100 34066 23156 34076
rect 22540 34020 22596 34030
rect 22540 33926 22596 33964
rect 23212 34018 23268 34030
rect 23212 33966 23214 34018
rect 23266 33966 23268 34018
rect 23212 33796 23268 33966
rect 22316 33506 22372 33516
rect 22652 33572 22708 33582
rect 22316 33346 22372 33358
rect 22316 33294 22318 33346
rect 22370 33294 22372 33346
rect 22316 32788 22372 33294
rect 22316 32722 22372 32732
rect 22652 32564 22708 33516
rect 22876 33236 22932 33246
rect 22876 33142 22932 33180
rect 22316 32562 22708 32564
rect 22316 32510 22654 32562
rect 22706 32510 22708 32562
rect 22316 32508 22708 32510
rect 22316 30770 22372 32508
rect 22652 32498 22708 32508
rect 22988 32562 23044 32574
rect 22988 32510 22990 32562
rect 23042 32510 23044 32562
rect 22988 32452 23044 32510
rect 23212 32562 23268 33740
rect 23212 32510 23214 32562
rect 23266 32510 23268 32562
rect 23212 32498 23268 32510
rect 22988 32386 23044 32396
rect 23324 32228 23380 36316
rect 23436 35140 23492 37100
rect 23548 36482 23604 36494
rect 23548 36430 23550 36482
rect 23602 36430 23604 36482
rect 23548 35252 23604 36430
rect 23548 35186 23604 35196
rect 23660 35586 23716 35598
rect 23660 35534 23662 35586
rect 23714 35534 23716 35586
rect 23436 35074 23492 35084
rect 23548 35028 23604 35038
rect 23660 35028 23716 35534
rect 23548 35026 23716 35028
rect 23548 34974 23550 35026
rect 23602 34974 23716 35026
rect 23548 34972 23716 34974
rect 23772 35252 23828 35262
rect 23548 33684 23604 34972
rect 23548 33618 23604 33628
rect 23436 33236 23492 33246
rect 23436 32338 23492 33180
rect 23772 33124 23828 35196
rect 23772 33030 23828 33068
rect 23436 32286 23438 32338
rect 23490 32286 23492 32338
rect 23436 32274 23492 32286
rect 23100 32172 23380 32228
rect 22988 31778 23044 31790
rect 22988 31726 22990 31778
rect 23042 31726 23044 31778
rect 22428 31668 22484 31678
rect 22764 31668 22820 31678
rect 22428 31666 22708 31668
rect 22428 31614 22430 31666
rect 22482 31614 22708 31666
rect 22428 31612 22708 31614
rect 22428 31602 22484 31612
rect 22316 30718 22318 30770
rect 22370 30718 22372 30770
rect 22316 30706 22372 30718
rect 22204 30382 22206 30434
rect 22258 30382 22260 30434
rect 22204 30370 22260 30382
rect 22316 30210 22372 30222
rect 22316 30158 22318 30210
rect 22370 30158 22372 30210
rect 22316 30100 22372 30158
rect 22316 30034 22372 30044
rect 22092 29586 22148 29596
rect 22652 28868 22708 31612
rect 22764 31666 22932 31668
rect 22764 31614 22766 31666
rect 22818 31614 22932 31666
rect 22764 31612 22932 31614
rect 22764 31602 22820 31612
rect 22764 31220 22820 31230
rect 22764 29092 22820 31164
rect 22876 30212 22932 31612
rect 22988 30436 23044 31726
rect 22988 30370 23044 30380
rect 22988 30212 23044 30222
rect 22876 30210 23044 30212
rect 22876 30158 22990 30210
rect 23042 30158 23044 30210
rect 22876 30156 23044 30158
rect 22988 30146 23044 30156
rect 23100 29986 23156 32172
rect 23884 32004 23940 40236
rect 24556 40068 24612 41244
rect 24668 41186 24724 41198
rect 24668 41134 24670 41186
rect 24722 41134 24724 41186
rect 24668 40516 24724 41134
rect 24892 40964 24948 43596
rect 25228 43650 25284 43652
rect 25228 43598 25230 43650
rect 25282 43598 25284 43650
rect 25228 43586 25284 43598
rect 25564 42196 25620 45500
rect 25788 45444 25844 46510
rect 26684 46452 26740 46844
rect 27020 46562 27076 46574
rect 27020 46510 27022 46562
rect 27074 46510 27076 46562
rect 26684 46396 26964 46452
rect 26012 45778 26068 45790
rect 26012 45726 26014 45778
rect 26066 45726 26068 45778
rect 25452 42140 25620 42196
rect 25676 42754 25732 42766
rect 25676 42702 25678 42754
rect 25730 42702 25732 42754
rect 25340 41972 25396 41982
rect 25340 41878 25396 41916
rect 25228 41860 25284 41870
rect 25116 41300 25172 41310
rect 25116 41186 25172 41244
rect 25116 41134 25118 41186
rect 25170 41134 25172 41186
rect 25116 41122 25172 41134
rect 24892 40908 25172 40964
rect 24668 40450 24724 40460
rect 24444 40012 24612 40068
rect 24108 39730 24164 39742
rect 24108 39678 24110 39730
rect 24162 39678 24164 39730
rect 24108 39620 24164 39678
rect 24108 39554 24164 39564
rect 23996 39508 24052 39518
rect 23996 38834 24052 39452
rect 23996 38782 23998 38834
rect 24050 38782 24052 38834
rect 23996 38668 24052 38782
rect 24332 38724 24388 38734
rect 23996 38612 24388 38668
rect 24332 38162 24388 38612
rect 24332 38110 24334 38162
rect 24386 38110 24388 38162
rect 24332 38098 24388 38110
rect 23996 38052 24052 38062
rect 23996 37940 24052 37996
rect 24220 38052 24276 38062
rect 24108 37940 24164 37950
rect 23996 37938 24164 37940
rect 23996 37886 24110 37938
rect 24162 37886 24164 37938
rect 23996 37884 24164 37886
rect 24108 37492 24164 37884
rect 24108 37426 24164 37436
rect 23996 37266 24052 37278
rect 23996 37214 23998 37266
rect 24050 37214 24052 37266
rect 23996 35028 24052 37214
rect 24220 36594 24276 37996
rect 24220 36542 24222 36594
rect 24274 36542 24276 36594
rect 24220 36530 24276 36542
rect 24444 36484 24500 40012
rect 24668 39620 24724 39630
rect 25004 39620 25060 39630
rect 24668 39618 24836 39620
rect 24668 39566 24670 39618
rect 24722 39566 24836 39618
rect 24668 39564 24836 39566
rect 24668 39554 24724 39564
rect 24556 39396 24612 39406
rect 24556 39302 24612 39340
rect 24668 38948 24724 38958
rect 24668 38854 24724 38892
rect 24556 38836 24612 38846
rect 24556 38274 24612 38780
rect 24780 38668 24836 39564
rect 25004 39526 25060 39564
rect 24780 38612 24948 38668
rect 24556 38222 24558 38274
rect 24610 38222 24612 38274
rect 24556 38210 24612 38222
rect 24780 38388 24836 38398
rect 24780 37490 24836 38332
rect 24892 38274 24948 38612
rect 24892 38222 24894 38274
rect 24946 38222 24948 38274
rect 24892 38210 24948 38222
rect 24780 37438 24782 37490
rect 24834 37438 24836 37490
rect 24556 37268 24612 37278
rect 24780 37268 24836 37438
rect 24612 37212 24724 37268
rect 24556 37202 24612 37212
rect 24668 36706 24724 37212
rect 24780 37202 24836 37212
rect 24668 36654 24670 36706
rect 24722 36654 24724 36706
rect 24668 36642 24724 36654
rect 25116 36596 25172 40908
rect 25228 40404 25284 41804
rect 25452 41636 25508 42140
rect 25564 41970 25620 41982
rect 25564 41918 25566 41970
rect 25618 41918 25620 41970
rect 25564 41860 25620 41918
rect 25564 41794 25620 41804
rect 25676 41636 25732 42702
rect 25228 40338 25284 40348
rect 25340 41580 25508 41636
rect 25564 41580 25732 41636
rect 25228 38724 25284 38762
rect 25228 38658 25284 38668
rect 25340 38668 25396 41580
rect 25452 41300 25508 41310
rect 25564 41300 25620 41580
rect 25676 41412 25732 41422
rect 25676 41318 25732 41356
rect 25508 41244 25620 41300
rect 25788 41300 25844 45388
rect 25900 45666 25956 45678
rect 25900 45614 25902 45666
rect 25954 45614 25956 45666
rect 25900 45106 25956 45614
rect 25900 45054 25902 45106
rect 25954 45054 25956 45106
rect 25900 44324 25956 45054
rect 26012 45108 26068 45726
rect 26012 45042 26068 45052
rect 26124 45332 26180 45342
rect 26124 45108 26180 45276
rect 26572 45218 26628 45230
rect 26572 45166 26574 45218
rect 26626 45166 26628 45218
rect 26572 45108 26628 45166
rect 26124 45052 26628 45108
rect 26796 45106 26852 45118
rect 26796 45054 26798 45106
rect 26850 45054 26852 45106
rect 26012 44436 26068 44446
rect 26124 44436 26180 45052
rect 26236 44548 26292 44558
rect 26236 44454 26292 44492
rect 26012 44434 26180 44436
rect 26012 44382 26014 44434
rect 26066 44382 26180 44434
rect 26012 44380 26180 44382
rect 26012 44370 26068 44380
rect 26796 44324 26852 45054
rect 25900 44258 25956 44268
rect 26460 44268 26852 44324
rect 26348 43540 26404 43550
rect 26460 43540 26516 44268
rect 26348 43538 26516 43540
rect 26348 43486 26350 43538
rect 26402 43486 26516 43538
rect 26348 43484 26516 43486
rect 26572 44098 26628 44110
rect 26572 44046 26574 44098
rect 26626 44046 26628 44098
rect 26572 43540 26628 44046
rect 26908 43876 26964 46396
rect 27020 45892 27076 46510
rect 27244 46116 27300 47740
rect 27468 47570 27524 47582
rect 27468 47518 27470 47570
rect 27522 47518 27524 47570
rect 27356 46676 27412 46686
rect 27468 46676 27524 47518
rect 27692 47460 27748 48188
rect 27804 47796 27860 50540
rect 28252 50596 28308 50606
rect 28252 50502 28308 50540
rect 28924 50596 28980 51326
rect 29260 50818 29316 52108
rect 29260 50766 29262 50818
rect 29314 50766 29316 50818
rect 29260 50754 29316 50766
rect 29484 52162 29540 53004
rect 29484 52110 29486 52162
rect 29538 52110 29540 52162
rect 28924 50530 28980 50540
rect 28476 50484 28532 50494
rect 28476 49922 28532 50428
rect 29484 50484 29540 52110
rect 29596 52946 29652 52958
rect 29596 52894 29598 52946
rect 29650 52894 29652 52946
rect 29596 52052 29652 52894
rect 31052 52946 31108 53566
rect 31388 53618 31444 53630
rect 31388 53566 31390 53618
rect 31442 53566 31444 53618
rect 31276 53508 31332 53518
rect 31276 53414 31332 53452
rect 31052 52894 31054 52946
rect 31106 52894 31108 52946
rect 29596 51986 29652 51996
rect 29708 52836 29764 52846
rect 29596 51492 29652 51502
rect 29708 51492 29764 52780
rect 30828 52836 30884 52846
rect 30828 52742 30884 52780
rect 30156 52164 30212 52174
rect 30156 52070 30212 52108
rect 30828 52162 30884 52174
rect 30828 52110 30830 52162
rect 30882 52110 30884 52162
rect 29596 51490 29764 51492
rect 29596 51438 29598 51490
rect 29650 51438 29764 51490
rect 29596 51436 29764 51438
rect 30604 52052 30660 52062
rect 29596 51426 29652 51436
rect 30268 51380 30324 51390
rect 29596 50820 29652 50830
rect 29596 50726 29652 50764
rect 30156 50708 30212 50718
rect 30156 50614 30212 50652
rect 29484 50418 29540 50428
rect 29596 50596 29652 50606
rect 28476 49870 28478 49922
rect 28530 49870 28532 49922
rect 28476 49858 28532 49870
rect 29372 49922 29428 49934
rect 29372 49870 29374 49922
rect 29426 49870 29428 49922
rect 28700 49812 28756 49822
rect 28700 49718 28756 49756
rect 29372 49812 29428 49870
rect 29372 49746 29428 49756
rect 28252 49700 28308 49710
rect 27916 49698 28308 49700
rect 27916 49646 28254 49698
rect 28306 49646 28308 49698
rect 27916 49644 28308 49646
rect 27916 49588 27972 49644
rect 28252 49634 28308 49644
rect 27916 49026 27972 49532
rect 29596 49250 29652 50540
rect 30268 50596 30324 51324
rect 30604 51378 30660 51996
rect 30604 51326 30606 51378
rect 30658 51326 30660 51378
rect 30604 51314 30660 51326
rect 30828 52052 30884 52110
rect 30828 50932 30884 51996
rect 31052 51490 31108 52894
rect 31388 52836 31444 53566
rect 32060 53508 32116 53518
rect 31948 53452 32060 53508
rect 31724 53284 31780 53294
rect 31724 53058 31780 53228
rect 31724 53006 31726 53058
rect 31778 53006 31780 53058
rect 31724 52994 31780 53006
rect 31388 52770 31444 52780
rect 31612 52274 31668 52286
rect 31612 52222 31614 52274
rect 31666 52222 31668 52274
rect 31388 52164 31444 52174
rect 31052 51438 31054 51490
rect 31106 51438 31108 51490
rect 31052 51426 31108 51438
rect 31276 52162 31444 52164
rect 31276 52110 31390 52162
rect 31442 52110 31444 52162
rect 31276 52108 31444 52110
rect 30828 50866 30884 50876
rect 31164 51378 31220 51390
rect 31164 51326 31166 51378
rect 31218 51326 31220 51378
rect 31164 50820 31220 51326
rect 31276 51044 31332 52108
rect 31388 52098 31444 52108
rect 31612 52052 31668 52222
rect 31612 51986 31668 51996
rect 31500 51378 31556 51390
rect 31500 51326 31502 51378
rect 31554 51326 31556 51378
rect 31276 50978 31332 50988
rect 31388 51156 31444 51166
rect 31164 50754 31220 50764
rect 29932 50484 29988 50522
rect 30268 50502 30324 50540
rect 29932 50418 29988 50428
rect 30380 50484 30436 50494
rect 29596 49198 29598 49250
rect 29650 49198 29652 49250
rect 29596 49186 29652 49198
rect 29708 49810 29764 49822
rect 29708 49758 29710 49810
rect 29762 49758 29764 49810
rect 29708 49700 29764 49758
rect 30156 49700 30212 49710
rect 29708 49698 30212 49700
rect 29708 49646 30158 49698
rect 30210 49646 30212 49698
rect 29708 49644 30212 49646
rect 29708 49140 29764 49644
rect 30156 49634 30212 49644
rect 29708 49074 29764 49084
rect 30044 49138 30100 49150
rect 30044 49086 30046 49138
rect 30098 49086 30100 49138
rect 27916 48974 27918 49026
rect 27970 48974 27972 49026
rect 27916 48962 27972 48974
rect 28028 49028 28084 49038
rect 27804 47730 27860 47740
rect 27916 48356 27972 48366
rect 27916 47572 27972 48300
rect 28028 48242 28084 48972
rect 28588 49028 28644 49038
rect 28588 48914 28644 48972
rect 29260 49028 29316 49038
rect 29260 48934 29316 48972
rect 28588 48862 28590 48914
rect 28642 48862 28644 48914
rect 28588 48850 28644 48862
rect 29484 48804 29540 48814
rect 30044 48804 30100 49086
rect 29484 48802 30100 48804
rect 29484 48750 29486 48802
rect 29538 48750 30100 48802
rect 29484 48748 30100 48750
rect 30268 48914 30324 48926
rect 30268 48862 30270 48914
rect 30322 48862 30324 48914
rect 29484 48356 29540 48748
rect 29484 48290 29540 48300
rect 28028 48190 28030 48242
rect 28082 48190 28084 48242
rect 28028 48178 28084 48190
rect 29932 48242 29988 48254
rect 29932 48190 29934 48242
rect 29986 48190 29988 48242
rect 27916 47506 27972 47516
rect 28364 48132 28420 48142
rect 28028 47460 28084 47470
rect 27692 47458 27860 47460
rect 27692 47406 27694 47458
rect 27746 47406 27860 47458
rect 27692 47404 27860 47406
rect 27692 47394 27748 47404
rect 27804 46786 27860 47404
rect 28028 47366 28084 47404
rect 28364 47458 28420 48076
rect 28364 47406 28366 47458
rect 28418 47406 28420 47458
rect 28364 47394 28420 47406
rect 28700 48020 28756 48030
rect 27916 47348 27972 47358
rect 27916 47254 27972 47292
rect 28700 46898 28756 47964
rect 29484 47684 29540 47694
rect 28700 46846 28702 46898
rect 28754 46846 28756 46898
rect 28700 46834 28756 46846
rect 29372 47460 29428 47470
rect 27804 46734 27806 46786
rect 27858 46734 27860 46786
rect 27804 46722 27860 46734
rect 29260 46788 29316 46798
rect 29148 46676 29204 46686
rect 29260 46676 29316 46732
rect 27356 46674 27748 46676
rect 27356 46622 27358 46674
rect 27410 46622 27748 46674
rect 27356 46620 27748 46622
rect 27356 46610 27412 46620
rect 27692 46564 27748 46620
rect 29148 46674 29316 46676
rect 29148 46622 29150 46674
rect 29202 46622 29316 46674
rect 29148 46620 29316 46622
rect 29372 46674 29428 47404
rect 29372 46622 29374 46674
rect 29426 46622 29428 46674
rect 29148 46610 29204 46620
rect 29372 46610 29428 46622
rect 29484 46674 29540 47628
rect 29708 47570 29764 47582
rect 29708 47518 29710 47570
rect 29762 47518 29764 47570
rect 29708 47124 29764 47518
rect 29484 46622 29486 46674
rect 29538 46622 29540 46674
rect 29484 46610 29540 46622
rect 29596 47068 29764 47124
rect 29820 47458 29876 47470
rect 29820 47406 29822 47458
rect 29874 47406 29876 47458
rect 29820 47124 29876 47406
rect 28140 46564 28196 46574
rect 27692 46562 28196 46564
rect 27692 46510 28142 46562
rect 28194 46510 28196 46562
rect 27692 46508 28196 46510
rect 27356 46116 27412 46126
rect 27244 46114 27412 46116
rect 27244 46062 27358 46114
rect 27410 46062 27412 46114
rect 27244 46060 27412 46062
rect 27356 46050 27412 46060
rect 27916 46002 27972 46508
rect 28140 46498 28196 46508
rect 29596 46564 29652 47068
rect 29820 47058 29876 47068
rect 29932 46788 29988 48190
rect 30268 47684 30324 48862
rect 30380 48466 30436 50428
rect 31052 50484 31108 50522
rect 31052 50418 31108 50428
rect 30380 48414 30382 48466
rect 30434 48414 30436 48466
rect 30380 48402 30436 48414
rect 30492 48244 30548 48254
rect 30492 48242 30772 48244
rect 30492 48190 30494 48242
rect 30546 48190 30772 48242
rect 30492 48188 30772 48190
rect 30492 48178 30548 48188
rect 30268 47618 30324 47628
rect 30716 47570 30772 48188
rect 30716 47518 30718 47570
rect 30770 47518 30772 47570
rect 30716 47460 30772 47518
rect 30716 47394 30772 47404
rect 31276 48242 31332 48254
rect 31276 48190 31278 48242
rect 31330 48190 31332 48242
rect 31276 47458 31332 48190
rect 31276 47406 31278 47458
rect 31330 47406 31332 47458
rect 29932 46694 29988 46732
rect 30380 47012 30436 47022
rect 27916 45950 27918 46002
rect 27970 45950 27972 46002
rect 27916 45938 27972 45950
rect 28364 46450 28420 46462
rect 28364 46398 28366 46450
rect 28418 46398 28420 46450
rect 27692 45892 27748 45902
rect 27020 45890 27748 45892
rect 27020 45838 27694 45890
rect 27746 45838 27748 45890
rect 27020 45836 27748 45838
rect 27692 45780 27748 45836
rect 28364 45780 28420 46398
rect 29596 45890 29652 46508
rect 29596 45838 29598 45890
rect 29650 45838 29652 45890
rect 29596 45826 29652 45838
rect 29708 46676 29764 46686
rect 27692 45724 28420 45780
rect 27580 45220 27636 45230
rect 27692 45220 27748 45724
rect 27580 45218 27748 45220
rect 27580 45166 27582 45218
rect 27634 45166 27748 45218
rect 27580 45164 27748 45166
rect 28140 45556 28196 45566
rect 29708 45556 29764 46620
rect 30268 46674 30324 46686
rect 30268 46622 30270 46674
rect 30322 46622 30324 46674
rect 29932 45780 29988 45790
rect 30268 45780 30324 46622
rect 29932 45778 30324 45780
rect 29932 45726 29934 45778
rect 29986 45726 30324 45778
rect 29932 45724 30324 45726
rect 30380 46562 30436 46956
rect 30380 46510 30382 46562
rect 30434 46510 30436 46562
rect 29932 45714 29988 45724
rect 30380 45556 30436 46510
rect 30940 46900 30996 46910
rect 30940 45890 30996 46844
rect 31276 46676 31332 47406
rect 31276 46610 31332 46620
rect 30940 45838 30942 45890
rect 30994 45838 30996 45890
rect 30940 45826 30996 45838
rect 29708 45500 29988 45556
rect 27244 45108 27300 45118
rect 27244 45106 27412 45108
rect 27244 45054 27246 45106
rect 27298 45054 27412 45106
rect 27244 45052 27412 45054
rect 27244 45042 27300 45052
rect 26908 43810 26964 43820
rect 27244 44322 27300 44334
rect 27244 44270 27246 44322
rect 27298 44270 27300 44322
rect 27244 43708 27300 44270
rect 25900 42866 25956 42878
rect 25900 42814 25902 42866
rect 25954 42814 25956 42866
rect 25900 41412 25956 42814
rect 26236 42756 26292 42766
rect 26236 42662 26292 42700
rect 26236 41972 26292 41982
rect 25900 41346 25956 41356
rect 26012 41970 26292 41972
rect 26012 41918 26238 41970
rect 26290 41918 26292 41970
rect 26012 41916 26292 41918
rect 26012 41410 26068 41916
rect 26236 41906 26292 41916
rect 26348 41636 26404 43484
rect 26572 43474 26628 43484
rect 26684 43652 26740 43662
rect 26684 43538 26740 43596
rect 26796 43652 27300 43708
rect 26796 43650 26852 43652
rect 26796 43598 26798 43650
rect 26850 43598 26852 43650
rect 26796 43586 26852 43598
rect 27244 43650 27300 43652
rect 27244 43598 27246 43650
rect 27298 43598 27300 43650
rect 27244 43586 27300 43598
rect 27356 43652 27412 45052
rect 27580 44548 27636 45164
rect 27580 44482 27636 44492
rect 27356 43586 27412 43596
rect 27692 44322 27748 44334
rect 27692 44270 27694 44322
rect 27746 44270 27748 44322
rect 26684 43486 26686 43538
rect 26738 43486 26740 43538
rect 26460 43204 26516 43214
rect 26460 41858 26516 43148
rect 26460 41806 26462 41858
rect 26514 41806 26516 41858
rect 26460 41794 26516 41806
rect 26348 41580 26628 41636
rect 26012 41358 26014 41410
rect 26066 41358 26068 41410
rect 26012 41346 26068 41358
rect 25452 41206 25508 41244
rect 25788 41234 25844 41244
rect 25564 39788 26180 39844
rect 25564 39506 25620 39788
rect 25564 39454 25566 39506
rect 25618 39454 25620 39506
rect 25564 39442 25620 39454
rect 25340 38612 25732 38668
rect 25676 37828 25732 38612
rect 25900 37828 25956 39788
rect 26012 39618 26068 39630
rect 26012 39566 26014 39618
rect 26066 39566 26068 39618
rect 26012 38162 26068 39566
rect 26124 39618 26180 39788
rect 26124 39566 26126 39618
rect 26178 39566 26180 39618
rect 26124 39554 26180 39566
rect 26460 39506 26516 39518
rect 26460 39454 26462 39506
rect 26514 39454 26516 39506
rect 26348 39396 26404 39406
rect 26348 39302 26404 39340
rect 26012 38110 26014 38162
rect 26066 38110 26068 38162
rect 26012 38098 26068 38110
rect 26124 38948 26180 38958
rect 26460 38948 26516 39454
rect 26180 38892 26516 38948
rect 26124 38050 26180 38892
rect 26124 37998 26126 38050
rect 26178 37998 26180 38050
rect 26124 37986 26180 37998
rect 26572 38052 26628 41580
rect 26572 37986 26628 37996
rect 25676 37826 25844 37828
rect 25676 37774 25678 37826
rect 25730 37774 25844 37826
rect 25676 37772 25844 37774
rect 25676 37762 25732 37772
rect 25452 37492 25508 37502
rect 25340 37380 25396 37390
rect 25340 37286 25396 37324
rect 25228 37268 25284 37278
rect 25228 37174 25284 37212
rect 25452 36820 25508 37436
rect 24332 36428 24500 36484
rect 24892 36540 25172 36596
rect 25228 36764 25508 36820
rect 25564 37268 25620 37278
rect 24108 35700 24164 35710
rect 24108 35698 24276 35700
rect 24108 35646 24110 35698
rect 24162 35646 24276 35698
rect 24108 35644 24276 35646
rect 24108 35634 24164 35644
rect 24108 35476 24164 35486
rect 24108 35382 24164 35420
rect 24220 35252 24276 35644
rect 23996 34962 24052 34972
rect 24108 35196 24276 35252
rect 24108 34356 24164 35196
rect 23996 34300 24164 34356
rect 24220 34356 24276 34366
rect 24332 34356 24388 36428
rect 24668 36372 24724 36382
rect 24668 36278 24724 36316
rect 24780 36370 24836 36382
rect 24780 36318 24782 36370
rect 24834 36318 24836 36370
rect 24780 34804 24836 36318
rect 24780 34738 24836 34748
rect 24220 34354 24388 34356
rect 24220 34302 24222 34354
rect 24274 34302 24388 34354
rect 24220 34300 24388 34302
rect 23996 33908 24052 34300
rect 24220 34290 24276 34300
rect 23996 33842 24052 33852
rect 24108 34130 24164 34142
rect 24108 34078 24110 34130
rect 24162 34078 24164 34130
rect 24108 32676 24164 34078
rect 24332 34132 24388 34142
rect 24332 34038 24388 34076
rect 24668 34132 24724 34142
rect 24668 34038 24724 34076
rect 24780 33348 24836 33358
rect 24556 33346 24836 33348
rect 24556 33294 24782 33346
rect 24834 33294 24836 33346
rect 24556 33292 24836 33294
rect 24444 33124 24500 33134
rect 23996 32620 24164 32676
rect 24332 33122 24500 33124
rect 24332 33070 24446 33122
rect 24498 33070 24500 33122
rect 24332 33068 24500 33070
rect 23996 32452 24052 32620
rect 23996 32386 24052 32396
rect 24220 32340 24276 32350
rect 24220 32246 24276 32284
rect 23996 32004 24052 32014
rect 23884 32002 24052 32004
rect 23884 31950 23998 32002
rect 24050 31950 24052 32002
rect 23884 31948 24052 31950
rect 23996 31938 24052 31948
rect 23548 31892 23604 31902
rect 23436 31780 23492 31790
rect 23548 31780 23604 31836
rect 23436 31778 23716 31780
rect 23436 31726 23438 31778
rect 23490 31726 23716 31778
rect 23436 31724 23716 31726
rect 23436 31714 23492 31724
rect 23660 30996 23716 31724
rect 23100 29934 23102 29986
rect 23154 29934 23156 29986
rect 23100 29922 23156 29934
rect 23548 30210 23604 30222
rect 23548 30158 23550 30210
rect 23602 30158 23604 30210
rect 22876 29316 22932 29326
rect 22876 29314 23380 29316
rect 22876 29262 22878 29314
rect 22930 29262 23380 29314
rect 22876 29260 23380 29262
rect 22876 29250 22932 29260
rect 22764 29036 23156 29092
rect 21756 28642 21812 28700
rect 21756 28590 21758 28642
rect 21810 28590 21812 28642
rect 21756 28578 21812 28590
rect 21980 28812 22708 28868
rect 21980 28082 22036 28812
rect 22652 28756 22708 28812
rect 22988 28756 23044 28766
rect 22652 28700 22932 28756
rect 22428 28644 22484 28654
rect 21980 28030 21982 28082
rect 22034 28030 22036 28082
rect 21532 27694 21534 27746
rect 21586 27694 21588 27746
rect 21532 27682 21588 27694
rect 21868 27858 21924 27870
rect 21868 27806 21870 27858
rect 21922 27806 21924 27858
rect 20524 26910 20526 26962
rect 20578 26910 20580 26962
rect 20524 26404 20580 26910
rect 21420 27074 21476 27086
rect 21420 27022 21422 27074
rect 21474 27022 21476 27074
rect 21196 26516 21252 26526
rect 20524 26338 20580 26348
rect 20860 26404 20916 26414
rect 20860 26310 20916 26348
rect 20972 26290 21028 26302
rect 20972 26238 20974 26290
rect 21026 26238 21028 26290
rect 20860 26068 20916 26078
rect 20860 25974 20916 26012
rect 20300 25788 20468 25844
rect 20188 25508 20244 25518
rect 19964 25396 20020 25406
rect 19852 25340 19964 25396
rect 19964 25330 20020 25340
rect 20076 25284 20132 25322
rect 20076 25218 20132 25228
rect 20188 25172 20244 25452
rect 20300 25394 20356 25788
rect 20300 25342 20302 25394
rect 20354 25342 20356 25394
rect 20300 25330 20356 25342
rect 20412 25396 20468 25406
rect 20412 25284 20468 25340
rect 20972 25284 21028 26238
rect 20412 25228 21028 25284
rect 21196 25508 21252 26460
rect 21420 26180 21476 27022
rect 21868 26852 21924 27806
rect 21868 26786 21924 26796
rect 21980 26516 22036 28030
rect 22204 28642 22484 28644
rect 22204 28590 22430 28642
rect 22482 28590 22484 28642
rect 22204 28588 22484 28590
rect 22204 28082 22260 28588
rect 22428 28578 22484 28588
rect 22876 28530 22932 28700
rect 22988 28662 23044 28700
rect 23100 28532 23156 29036
rect 22876 28478 22878 28530
rect 22930 28478 22932 28530
rect 22876 28466 22932 28478
rect 22988 28530 23156 28532
rect 22988 28478 23102 28530
rect 23154 28478 23156 28530
rect 22988 28476 23156 28478
rect 22204 28030 22206 28082
rect 22258 28030 22260 28082
rect 22204 28018 22260 28030
rect 22316 28420 22372 28430
rect 21980 26450 22036 26460
rect 22092 26962 22148 26974
rect 22092 26910 22094 26962
rect 22146 26910 22148 26962
rect 21420 26114 21476 26124
rect 21756 26178 21812 26190
rect 21756 26126 21758 26178
rect 21810 26126 21812 26178
rect 19836 25116 20100 25126
rect 20188 25116 20468 25172
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 19836 25050 20100 25060
rect 19628 24782 19630 24834
rect 19682 24782 19684 24834
rect 19628 24770 19684 24782
rect 20076 24724 20132 24734
rect 20076 24630 20132 24668
rect 20300 24722 20356 24734
rect 20300 24670 20302 24722
rect 20354 24670 20356 24722
rect 19516 24052 19572 24332
rect 19516 23986 19572 23996
rect 20188 24052 20244 24062
rect 19292 23938 19348 23950
rect 19292 23886 19294 23938
rect 19346 23886 19348 23938
rect 19292 23548 19348 23886
rect 20188 23938 20244 23996
rect 20188 23886 20190 23938
rect 20242 23886 20244 23938
rect 20188 23874 20244 23886
rect 20300 23940 20356 24670
rect 20300 23874 20356 23884
rect 19516 23828 19572 23838
rect 19516 23734 19572 23772
rect 19964 23716 20020 23754
rect 19964 23650 20020 23660
rect 19836 23548 20100 23558
rect 19292 23492 19460 23548
rect 19124 23324 19236 23380
rect 19068 23286 19124 23324
rect 18956 21634 19012 21644
rect 19068 23156 19124 23166
rect 19068 21476 19124 23100
rect 19404 23154 19460 23492
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 19836 23482 20100 23492
rect 19404 23102 19406 23154
rect 19458 23102 19460 23154
rect 19404 22372 19460 23102
rect 19740 23156 19796 23166
rect 19740 23062 19796 23100
rect 20300 23042 20356 23054
rect 20300 22990 20302 23042
rect 20354 22990 20356 23042
rect 19852 22932 19908 22942
rect 19852 22930 20132 22932
rect 19852 22878 19854 22930
rect 19906 22878 20132 22930
rect 19852 22876 20132 22878
rect 19852 22866 19908 22876
rect 19628 22372 19684 22382
rect 19964 22372 20020 22382
rect 19404 22370 19684 22372
rect 19404 22318 19630 22370
rect 19682 22318 19684 22370
rect 19404 22316 19684 22318
rect 19628 22306 19684 22316
rect 19740 22370 20020 22372
rect 19740 22318 19966 22370
rect 20018 22318 20020 22370
rect 19740 22316 20020 22318
rect 19180 22258 19236 22270
rect 19180 22206 19182 22258
rect 19234 22206 19236 22258
rect 19180 21700 19236 22206
rect 19740 22148 19796 22316
rect 19964 22306 20020 22316
rect 19180 21634 19236 21644
rect 19628 22092 19796 22148
rect 19852 22148 19908 22186
rect 20076 22148 20132 22876
rect 20188 22372 20244 22382
rect 20188 22278 20244 22316
rect 19908 22092 20132 22148
rect 19292 21476 19348 21486
rect 19068 21474 19348 21476
rect 19068 21422 19294 21474
rect 19346 21422 19348 21474
rect 19068 21420 19348 21422
rect 19180 21140 19236 21150
rect 18956 20578 19012 20590
rect 18956 20526 18958 20578
rect 19010 20526 19012 20578
rect 18956 20020 19012 20526
rect 19068 20580 19124 20590
rect 19068 20486 19124 20524
rect 19180 20578 19236 21084
rect 19180 20526 19182 20578
rect 19234 20526 19236 20578
rect 19180 20468 19236 20526
rect 19180 20188 19236 20412
rect 18956 19954 19012 19964
rect 19068 20132 19236 20188
rect 18732 19236 18788 19246
rect 18732 19142 18788 19180
rect 18844 19124 18900 19852
rect 18844 19058 18900 19068
rect 18732 18676 18788 18686
rect 18732 18674 19012 18676
rect 18732 18622 18734 18674
rect 18786 18622 19012 18674
rect 18732 18620 19012 18622
rect 18732 18610 18788 18620
rect 18620 18498 18676 18508
rect 18844 17892 18900 17902
rect 18732 17556 18788 17566
rect 18732 17462 18788 17500
rect 18620 16996 18676 17006
rect 18620 16902 18676 16940
rect 18732 16884 18788 16894
rect 18732 16790 18788 16828
rect 18844 16100 18900 17836
rect 17724 15986 18116 15988
rect 17724 15934 17726 15986
rect 17778 15934 18116 15986
rect 17724 15932 18116 15934
rect 17724 15922 17780 15932
rect 17612 15486 17614 15538
rect 17666 15486 17668 15538
rect 17612 15474 17668 15486
rect 18060 15538 18116 15932
rect 18508 15894 18564 15932
rect 18732 16044 18900 16100
rect 18060 15486 18062 15538
rect 18114 15486 18116 15538
rect 18060 15474 18116 15486
rect 18396 15876 18452 15886
rect 17948 15316 18004 15326
rect 17724 15314 18004 15316
rect 17724 15262 17950 15314
rect 18002 15262 18004 15314
rect 17724 15260 18004 15262
rect 16940 13794 16996 13804
rect 17164 14476 17444 14532
rect 17612 15090 17668 15102
rect 17612 15038 17614 15090
rect 17666 15038 17668 15090
rect 16828 13748 16884 13758
rect 16716 13636 16772 13646
rect 16716 13412 16772 13580
rect 16828 13634 16884 13692
rect 16828 13582 16830 13634
rect 16882 13582 16884 13634
rect 16828 13570 16884 13582
rect 16716 13356 17108 13412
rect 16268 12292 16324 12302
rect 16268 12290 16548 12292
rect 16268 12238 16270 12290
rect 16322 12238 16548 12290
rect 16268 12236 16548 12238
rect 16268 12226 16324 12236
rect 16380 12066 16436 12078
rect 16380 12014 16382 12066
rect 16434 12014 16436 12066
rect 16380 11620 16436 12014
rect 15596 11564 16436 11620
rect 15596 11506 15652 11564
rect 15596 11454 15598 11506
rect 15650 11454 15652 11506
rect 15596 11442 15652 11454
rect 14924 11394 14980 11406
rect 14924 11342 14926 11394
rect 14978 11342 14980 11394
rect 14924 10836 14980 11342
rect 16492 11172 16548 12236
rect 16604 12290 16660 12348
rect 17052 13074 17108 13356
rect 17052 13022 17054 13074
rect 17106 13022 17108 13074
rect 16604 12238 16606 12290
rect 16658 12238 16660 12290
rect 16604 12226 16660 12238
rect 16828 12290 16884 12302
rect 16828 12238 16830 12290
rect 16882 12238 16884 12290
rect 16828 12180 16884 12238
rect 16940 12180 16996 12190
rect 16828 12124 16940 12180
rect 16940 12114 16996 12124
rect 16044 10948 16100 10958
rect 15036 10836 15092 10846
rect 14924 10780 15036 10836
rect 5964 9874 6020 9884
rect 15036 9826 15092 10780
rect 16044 10834 16100 10892
rect 16044 10782 16046 10834
rect 16098 10782 16100 10834
rect 16044 10770 16100 10782
rect 16268 10724 16324 10734
rect 16492 10724 16548 11116
rect 16268 10722 16548 10724
rect 16268 10670 16270 10722
rect 16322 10670 16548 10722
rect 16268 10668 16548 10670
rect 16268 10658 16324 10668
rect 16380 10498 16436 10510
rect 16380 10446 16382 10498
rect 16434 10446 16436 10498
rect 16380 10052 16436 10446
rect 15708 9996 16436 10052
rect 15708 9938 15764 9996
rect 15708 9886 15710 9938
rect 15762 9886 15764 9938
rect 15708 9874 15764 9886
rect 15036 9774 15038 9826
rect 15090 9774 15092 9826
rect 4476 8652 4740 8662
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4476 8586 4740 8596
rect 15036 8428 15092 9774
rect 16492 9156 16548 10668
rect 16604 10948 16660 10958
rect 16604 10722 16660 10892
rect 17052 10836 17108 13022
rect 17164 10948 17220 14476
rect 17612 12740 17668 15038
rect 17724 13970 17780 15260
rect 17948 15250 18004 15260
rect 18172 15314 18228 15326
rect 18172 15262 18174 15314
rect 18226 15262 18228 15314
rect 18172 14642 18228 15262
rect 18172 14590 18174 14642
rect 18226 14590 18228 14642
rect 17724 13918 17726 13970
rect 17778 13918 17780 13970
rect 17724 13076 17780 13918
rect 18060 14532 18116 14542
rect 17836 13860 17892 13870
rect 17836 13766 17892 13804
rect 17948 13748 18004 13758
rect 18060 13748 18116 14476
rect 18172 13972 18228 14590
rect 18172 13906 18228 13916
rect 18004 13692 18116 13748
rect 18396 13746 18452 15820
rect 18620 15316 18676 15326
rect 18732 15316 18788 16044
rect 18844 15876 18900 15886
rect 18844 15782 18900 15820
rect 18508 15314 18788 15316
rect 18508 15262 18622 15314
rect 18674 15262 18788 15314
rect 18508 15260 18788 15262
rect 18844 15652 18900 15662
rect 18508 15148 18564 15260
rect 18620 15250 18676 15260
rect 18508 15092 18788 15148
rect 18732 14644 18788 15092
rect 18844 14868 18900 15596
rect 18956 15148 19012 18620
rect 19068 18564 19124 20132
rect 19180 20018 19236 20030
rect 19180 19966 19182 20018
rect 19234 19966 19236 20018
rect 19180 19684 19236 19966
rect 19180 19618 19236 19628
rect 19068 18562 19236 18564
rect 19068 18510 19070 18562
rect 19122 18510 19236 18562
rect 19068 18508 19236 18510
rect 19068 18498 19124 18508
rect 19068 17890 19124 17902
rect 19068 17838 19070 17890
rect 19122 17838 19124 17890
rect 19068 16882 19124 17838
rect 19180 17668 19236 18508
rect 19292 17890 19348 21420
rect 19404 21028 19460 21038
rect 19628 21028 19684 22092
rect 19852 22082 19908 22092
rect 19836 21980 20100 21990
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 19836 21914 20100 21924
rect 20076 21812 20132 21822
rect 20076 21718 20132 21756
rect 19740 21700 19796 21710
rect 19796 21644 19908 21700
rect 19740 21634 19796 21644
rect 19852 21028 19908 21644
rect 19964 21588 20020 21598
rect 19964 21586 20132 21588
rect 19964 21534 19966 21586
rect 20018 21534 20132 21586
rect 19964 21532 20132 21534
rect 19964 21522 20020 21532
rect 19964 21028 20020 21038
rect 19628 20972 19796 21028
rect 19852 21026 20020 21028
rect 19852 20974 19966 21026
rect 20018 20974 20020 21026
rect 19852 20972 20020 20974
rect 19404 20914 19460 20972
rect 19404 20862 19406 20914
rect 19458 20862 19460 20914
rect 19404 20850 19460 20862
rect 19516 20804 19572 20814
rect 19292 17838 19294 17890
rect 19346 17838 19348 17890
rect 19292 17826 19348 17838
rect 19404 20692 19460 20702
rect 19404 17780 19460 20636
rect 19404 17714 19460 17724
rect 19180 17612 19348 17668
rect 19180 17444 19236 17454
rect 19180 17350 19236 17388
rect 19068 16830 19070 16882
rect 19122 16830 19124 16882
rect 19068 15314 19124 16830
rect 19180 15876 19236 15886
rect 19180 15782 19236 15820
rect 19180 15428 19236 15438
rect 19292 15428 19348 17612
rect 19404 17556 19460 17566
rect 19404 16100 19460 17500
rect 19516 16324 19572 20748
rect 19628 20802 19684 20814
rect 19628 20750 19630 20802
rect 19682 20750 19684 20802
rect 19628 20244 19684 20750
rect 19740 20692 19796 20972
rect 19740 20626 19796 20636
rect 19964 20580 20020 20972
rect 20076 20804 20132 21532
rect 20188 21586 20244 21598
rect 20188 21534 20190 21586
rect 20242 21534 20244 21586
rect 20188 21140 20244 21534
rect 20188 21074 20244 21084
rect 20188 20804 20244 20814
rect 20076 20748 20188 20804
rect 20188 20710 20244 20748
rect 19964 20524 20244 20580
rect 19836 20412 20100 20422
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 19836 20346 20100 20356
rect 20188 20188 20244 20524
rect 19628 20178 19684 20188
rect 19964 20132 20244 20188
rect 19964 20018 20020 20132
rect 19964 19966 19966 20018
rect 20018 19966 20020 20018
rect 19628 19908 19684 19918
rect 19628 19814 19684 19852
rect 19964 19012 20020 19966
rect 20188 20020 20244 20030
rect 20188 19926 20244 19964
rect 19628 18956 20020 19012
rect 20188 19572 20244 19582
rect 19628 16994 19684 18956
rect 19836 18844 20100 18854
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 19836 18778 20100 18788
rect 20076 18450 20132 18462
rect 20076 18398 20078 18450
rect 20130 18398 20132 18450
rect 20076 17890 20132 18398
rect 20076 17838 20078 17890
rect 20130 17838 20132 17890
rect 20076 17826 20132 17838
rect 19740 17780 19796 17790
rect 19740 17686 19796 17724
rect 20188 17778 20244 19516
rect 20300 19348 20356 22990
rect 20412 22932 20468 25116
rect 20524 24836 20580 24846
rect 20524 24742 20580 24780
rect 20636 24722 20692 25228
rect 20636 24670 20638 24722
rect 20690 24670 20692 24722
rect 20636 23828 20692 24670
rect 20972 24612 21028 24622
rect 20636 23762 20692 23772
rect 20860 24276 20916 24286
rect 20748 23714 20804 23726
rect 20748 23662 20750 23714
rect 20802 23662 20804 23714
rect 20748 23268 20804 23662
rect 20636 23212 20804 23268
rect 20524 22932 20580 22942
rect 20636 22932 20692 23212
rect 20748 23044 20804 23054
rect 20860 23044 20916 24220
rect 20748 23042 20916 23044
rect 20748 22990 20750 23042
rect 20802 22990 20916 23042
rect 20748 22988 20916 22990
rect 20748 22978 20804 22988
rect 20412 22876 20524 22932
rect 20580 22876 20692 22932
rect 20524 22866 20580 22876
rect 20860 22484 20916 22988
rect 20860 22418 20916 22428
rect 20524 22258 20580 22270
rect 20524 22206 20526 22258
rect 20578 22206 20580 22258
rect 20412 22148 20468 22158
rect 20412 22054 20468 22092
rect 20524 21812 20580 22206
rect 20972 21924 21028 24556
rect 21196 24610 21252 25452
rect 21756 26066 21812 26126
rect 22092 26068 22148 26910
rect 22316 26908 22372 28364
rect 22988 28308 23044 28476
rect 23100 28466 23156 28476
rect 22428 28252 23044 28308
rect 22428 28082 22484 28252
rect 23324 28196 23380 29260
rect 23436 28868 23492 28878
rect 23436 28774 23492 28812
rect 23548 28756 23604 30158
rect 23660 30098 23716 30940
rect 23660 30046 23662 30098
rect 23714 30046 23716 30098
rect 23660 30034 23716 30046
rect 23772 31778 23828 31790
rect 23772 31726 23774 31778
rect 23826 31726 23828 31778
rect 23772 28868 23828 31726
rect 24332 31108 24388 33068
rect 24444 33058 24500 33068
rect 24556 32788 24612 33292
rect 24780 33282 24836 33292
rect 24444 32732 24612 32788
rect 24444 31668 24500 32732
rect 24556 32564 24612 32602
rect 24556 32498 24612 32508
rect 24556 32340 24612 32350
rect 24892 32340 24948 36540
rect 25228 36370 25284 36764
rect 25564 36594 25620 37212
rect 25788 37042 25844 37772
rect 25900 37734 25956 37772
rect 26572 37826 26628 37838
rect 26572 37774 26574 37826
rect 26626 37774 26628 37826
rect 26012 37492 26068 37502
rect 26012 37398 26068 37436
rect 26460 37268 26516 37278
rect 26460 37174 26516 37212
rect 25788 36990 25790 37042
rect 25842 36990 25844 37042
rect 25788 36978 25844 36990
rect 26572 37042 26628 37774
rect 26572 36990 26574 37042
rect 26626 36990 26628 37042
rect 26572 36932 26628 36990
rect 26460 36876 26628 36932
rect 25564 36542 25566 36594
rect 25618 36542 25620 36594
rect 25564 36530 25620 36542
rect 25676 36706 25732 36718
rect 25676 36654 25678 36706
rect 25730 36654 25732 36706
rect 25228 36318 25230 36370
rect 25282 36318 25284 36370
rect 25228 36306 25284 36318
rect 25340 35476 25396 35486
rect 25396 35420 25508 35476
rect 25340 35410 25396 35420
rect 25340 35140 25396 35150
rect 25116 35028 25172 35038
rect 25116 34934 25172 34972
rect 25340 34914 25396 35084
rect 25340 34862 25342 34914
rect 25394 34862 25396 34914
rect 25340 34850 25396 34862
rect 25452 34354 25508 35420
rect 25452 34302 25454 34354
rect 25506 34302 25508 34354
rect 25452 34290 25508 34302
rect 25564 35028 25620 35038
rect 25564 34354 25620 34972
rect 25564 34302 25566 34354
rect 25618 34302 25620 34354
rect 25564 34290 25620 34302
rect 25676 34354 25732 36654
rect 26012 35810 26068 35822
rect 26012 35758 26014 35810
rect 26066 35758 26068 35810
rect 25676 34302 25678 34354
rect 25730 34302 25732 34354
rect 25676 34290 25732 34302
rect 25788 35698 25844 35710
rect 25788 35646 25790 35698
rect 25842 35646 25844 35698
rect 25788 34356 25844 35646
rect 25788 34354 25956 34356
rect 25788 34302 25790 34354
rect 25842 34302 25956 34354
rect 25788 34300 25956 34302
rect 25788 34290 25844 34300
rect 25900 34132 25956 34300
rect 26012 34244 26068 35758
rect 26012 34150 26068 34188
rect 25900 34020 25956 34076
rect 26348 34020 26404 34030
rect 25900 34018 26404 34020
rect 25900 33966 26350 34018
rect 26402 33966 26404 34018
rect 25900 33964 26404 33966
rect 25788 33460 25844 33470
rect 25676 33404 25788 33460
rect 25228 33348 25284 33358
rect 25228 33346 25396 33348
rect 25228 33294 25230 33346
rect 25282 33294 25396 33346
rect 25228 33292 25396 33294
rect 25228 33282 25284 33292
rect 25340 32452 25396 33292
rect 25676 33346 25732 33404
rect 25788 33394 25844 33404
rect 25676 33294 25678 33346
rect 25730 33294 25732 33346
rect 25676 33282 25732 33294
rect 24556 32338 24948 32340
rect 24556 32286 24558 32338
rect 24610 32286 24948 32338
rect 24556 32284 24948 32286
rect 25116 32340 25172 32350
rect 24556 32274 24612 32284
rect 24444 31602 24500 31612
rect 25116 31892 25172 32284
rect 25228 31892 25284 31902
rect 25116 31890 25284 31892
rect 25116 31838 25230 31890
rect 25282 31838 25284 31890
rect 25116 31836 25284 31838
rect 24668 31220 24724 31230
rect 24444 31108 24500 31118
rect 24332 31052 24444 31108
rect 24444 31042 24500 31052
rect 24556 31106 24612 31118
rect 24556 31054 24558 31106
rect 24610 31054 24612 31106
rect 23884 30994 23940 31006
rect 23884 30942 23886 30994
rect 23938 30942 23940 30994
rect 23884 30100 23940 30942
rect 24332 30772 24388 30782
rect 23884 30034 23940 30044
rect 24108 30770 24388 30772
rect 24108 30718 24334 30770
rect 24386 30718 24388 30770
rect 24108 30716 24388 30718
rect 23548 28690 23604 28700
rect 23660 28812 23828 28868
rect 23996 29540 24052 29550
rect 23660 28420 23716 28812
rect 23996 28754 24052 29484
rect 23996 28702 23998 28754
rect 24050 28702 24052 28754
rect 23996 28690 24052 28702
rect 24108 29538 24164 30716
rect 24332 30706 24388 30716
rect 24220 30548 24276 30558
rect 24220 30100 24276 30492
rect 24556 30436 24612 31054
rect 24668 30882 24724 31164
rect 24668 30830 24670 30882
rect 24722 30830 24724 30882
rect 24668 30818 24724 30830
rect 25116 30884 25172 31836
rect 25228 31826 25284 31836
rect 25228 31108 25284 31118
rect 25228 30994 25284 31052
rect 25228 30942 25230 30994
rect 25282 30942 25284 30994
rect 25228 30930 25284 30942
rect 24556 30380 24948 30436
rect 24220 29764 24276 30044
rect 24556 30212 24612 30222
rect 24220 29708 24500 29764
rect 24108 29486 24110 29538
rect 24162 29486 24164 29538
rect 24108 28756 24164 29486
rect 24108 28690 24164 28700
rect 23772 28644 23828 28654
rect 23772 28550 23828 28588
rect 24444 28642 24500 29708
rect 24556 29650 24612 30156
rect 24556 29598 24558 29650
rect 24610 29598 24612 29650
rect 24556 29316 24612 29598
rect 24780 30210 24836 30222
rect 24780 30158 24782 30210
rect 24834 30158 24836 30210
rect 24780 29540 24836 30158
rect 24780 29474 24836 29484
rect 24556 29250 24612 29260
rect 24668 29426 24724 29438
rect 24668 29374 24670 29426
rect 24722 29374 24724 29426
rect 24444 28590 24446 28642
rect 24498 28590 24500 28642
rect 24444 28578 24500 28590
rect 24332 28532 24388 28542
rect 23660 28354 23716 28364
rect 24108 28530 24388 28532
rect 24108 28478 24334 28530
rect 24386 28478 24388 28530
rect 24108 28476 24388 28478
rect 24108 28196 24164 28476
rect 24332 28466 24388 28476
rect 24668 28420 24724 29374
rect 24668 28354 24724 28364
rect 23324 28130 23380 28140
rect 23660 28140 24164 28196
rect 24332 28196 24388 28206
rect 22428 28030 22430 28082
rect 22482 28030 22484 28082
rect 22428 28018 22484 28030
rect 22764 28084 22820 28094
rect 22764 27990 22820 28028
rect 23660 28082 23716 28140
rect 23660 28030 23662 28082
rect 23714 28030 23716 28082
rect 23660 28018 23716 28030
rect 23324 27972 23380 27982
rect 23324 27878 23380 27916
rect 23436 27970 23492 27982
rect 23436 27918 23438 27970
rect 23490 27918 23492 27970
rect 23436 27860 23492 27918
rect 23436 27804 23604 27860
rect 23548 27412 23604 27804
rect 24332 27858 24388 28140
rect 24332 27806 24334 27858
rect 24386 27806 24388 27858
rect 22204 26852 22372 26908
rect 23436 27356 23604 27412
rect 23884 27746 23940 27758
rect 23884 27694 23886 27746
rect 23938 27694 23940 27746
rect 22204 26292 22260 26852
rect 22204 26226 22260 26236
rect 22540 26348 22820 26404
rect 21756 26014 21758 26066
rect 21810 26014 21812 26066
rect 21644 25394 21700 25406
rect 21644 25342 21646 25394
rect 21698 25342 21700 25394
rect 21644 25172 21700 25342
rect 21196 24558 21198 24610
rect 21250 24558 21252 24610
rect 21196 24546 21252 24558
rect 21308 25116 21644 25172
rect 21308 24724 21364 25116
rect 21644 25106 21700 25116
rect 21308 23826 21364 24668
rect 21308 23774 21310 23826
rect 21362 23774 21364 23826
rect 21308 23762 21364 23774
rect 21420 24948 21476 24958
rect 21308 23156 21364 23166
rect 20972 21858 21028 21868
rect 21084 22148 21140 22158
rect 20524 21746 20580 21756
rect 21084 21700 21140 22092
rect 21308 21810 21364 23100
rect 21420 22482 21476 24892
rect 21756 24948 21812 26014
rect 21868 26012 22148 26068
rect 22316 26180 22372 26190
rect 22540 26180 22596 26348
rect 22316 26178 22596 26180
rect 22316 26126 22318 26178
rect 22370 26126 22596 26178
rect 22316 26124 22596 26126
rect 22652 26178 22708 26190
rect 22652 26126 22654 26178
rect 22706 26126 22708 26178
rect 21868 25618 21924 26012
rect 22316 25844 22372 26124
rect 22092 25788 22372 25844
rect 21868 25566 21870 25618
rect 21922 25566 21924 25618
rect 21868 25554 21924 25566
rect 21980 25620 22036 25630
rect 21868 25396 21924 25406
rect 21868 25302 21924 25340
rect 21980 25394 22036 25564
rect 21980 25342 21982 25394
rect 22034 25342 22036 25394
rect 21980 25330 22036 25342
rect 21756 24882 21812 24892
rect 21644 24052 21700 24062
rect 21644 23938 21700 23996
rect 21644 23886 21646 23938
rect 21698 23886 21700 23938
rect 21644 23874 21700 23886
rect 21532 23716 21588 23726
rect 21532 23378 21588 23660
rect 21532 23326 21534 23378
rect 21586 23326 21588 23378
rect 21532 23314 21588 23326
rect 21868 23156 21924 23166
rect 21868 23062 21924 23100
rect 21980 23044 22036 23054
rect 22092 23044 22148 25788
rect 22652 25620 22708 26126
rect 22652 25554 22708 25564
rect 22764 25394 22820 26348
rect 23100 26178 23156 26190
rect 23100 26126 23102 26178
rect 23154 26126 23156 26178
rect 23100 26066 23156 26126
rect 23100 26014 23102 26066
rect 23154 26014 23156 26066
rect 23100 26002 23156 26014
rect 23212 25956 23268 25966
rect 22764 25342 22766 25394
rect 22818 25342 22820 25394
rect 22764 25330 22820 25342
rect 22876 25394 22932 25406
rect 22876 25342 22878 25394
rect 22930 25342 22932 25394
rect 22204 25284 22260 25294
rect 22540 25284 22596 25294
rect 22204 25282 22596 25284
rect 22204 25230 22206 25282
rect 22258 25230 22542 25282
rect 22594 25230 22596 25282
rect 22204 25228 22596 25230
rect 22204 23716 22260 25228
rect 22540 25218 22596 25228
rect 22652 25172 22708 25182
rect 22316 24276 22372 24286
rect 22316 24050 22372 24220
rect 22316 23998 22318 24050
rect 22370 23998 22372 24050
rect 22316 23986 22372 23998
rect 22652 23938 22708 25116
rect 22652 23886 22654 23938
rect 22706 23886 22708 23938
rect 22652 23874 22708 23886
rect 22764 24836 22820 24846
rect 22204 23650 22260 23660
rect 22316 23604 22372 23614
rect 22204 23380 22260 23390
rect 22316 23380 22372 23548
rect 22764 23604 22820 24780
rect 22876 24052 22932 25342
rect 22988 25394 23044 25406
rect 22988 25342 22990 25394
rect 23042 25342 23044 25394
rect 22988 25172 23044 25342
rect 22988 25106 23044 25116
rect 23100 25284 23156 25294
rect 22876 23996 23044 24052
rect 22764 23538 22820 23548
rect 22876 23828 22932 23838
rect 22204 23378 22372 23380
rect 22204 23326 22206 23378
rect 22258 23326 22372 23378
rect 22204 23324 22372 23326
rect 22204 23314 22260 23324
rect 22652 23044 22708 23054
rect 22876 23044 22932 23772
rect 22988 23378 23044 23996
rect 23100 23826 23156 25228
rect 23212 24500 23268 25900
rect 23324 25618 23380 25630
rect 23324 25566 23326 25618
rect 23378 25566 23380 25618
rect 23324 24834 23380 25566
rect 23436 25172 23492 27356
rect 23884 26964 23940 27694
rect 24332 27188 24388 27806
rect 24332 27094 24388 27132
rect 23548 26516 23604 26526
rect 23604 26460 23828 26516
rect 23548 26422 23604 26460
rect 23548 25396 23604 25406
rect 23548 25302 23604 25340
rect 23772 25394 23828 26460
rect 23884 26514 23940 26908
rect 23884 26462 23886 26514
rect 23938 26462 23940 26514
rect 23884 26450 23940 26462
rect 24668 26180 24724 26190
rect 23772 25342 23774 25394
rect 23826 25342 23828 25394
rect 23772 25330 23828 25342
rect 23884 25396 23940 25406
rect 24444 25396 24500 25406
rect 23884 25394 24500 25396
rect 23884 25342 23886 25394
rect 23938 25342 24446 25394
rect 24498 25342 24500 25394
rect 23884 25340 24500 25342
rect 23436 25106 23492 25116
rect 23324 24782 23326 24834
rect 23378 24782 23380 24834
rect 23324 24770 23380 24782
rect 23884 24836 23940 25340
rect 24444 25330 24500 25340
rect 24556 25396 24612 25406
rect 24556 25302 24612 25340
rect 24668 25060 24724 26124
rect 24892 26180 24948 30380
rect 25116 30098 25172 30828
rect 25340 30772 25396 32396
rect 25564 32562 25620 32574
rect 25564 32510 25566 32562
rect 25618 32510 25620 32562
rect 25116 30046 25118 30098
rect 25170 30046 25172 30098
rect 25116 30034 25172 30046
rect 25228 30716 25396 30772
rect 25452 32004 25508 32014
rect 25116 26852 25172 26862
rect 25228 26852 25284 30716
rect 25116 26850 25284 26852
rect 25116 26798 25118 26850
rect 25170 26798 25284 26850
rect 25116 26796 25284 26798
rect 25116 26786 25172 26796
rect 25228 26740 25284 26796
rect 25228 26674 25284 26684
rect 25340 27188 25396 27198
rect 25340 26290 25396 27132
rect 25340 26238 25342 26290
rect 25394 26238 25396 26290
rect 25340 26226 25396 26238
rect 24892 25508 24948 26124
rect 24892 25442 24948 25452
rect 24780 25284 24836 25294
rect 25452 25284 25508 31948
rect 25564 30100 25620 32510
rect 25900 32450 25956 33964
rect 26348 33954 26404 33964
rect 25900 32398 25902 32450
rect 25954 32398 25956 32450
rect 25900 32386 25956 32398
rect 26348 33346 26404 33358
rect 26348 33294 26350 33346
rect 26402 33294 26404 33346
rect 26348 32004 26404 33294
rect 26460 33348 26516 36876
rect 26572 34244 26628 34254
rect 26572 34130 26628 34188
rect 26572 34078 26574 34130
rect 26626 34078 26628 34130
rect 26572 33570 26628 34078
rect 26572 33518 26574 33570
rect 26626 33518 26628 33570
rect 26572 33506 26628 33518
rect 26684 33460 26740 43486
rect 27692 43538 27748 44270
rect 27916 44324 27972 44334
rect 27916 44230 27972 44268
rect 28140 43762 28196 45500
rect 29372 45218 29428 45230
rect 29372 45166 29374 45218
rect 29426 45166 29428 45218
rect 28140 43710 28142 43762
rect 28194 43710 28196 43762
rect 28140 43698 28196 43710
rect 29260 45106 29316 45118
rect 29260 45054 29262 45106
rect 29314 45054 29316 45106
rect 27692 43486 27694 43538
rect 27746 43486 27748 43538
rect 27692 43316 27748 43486
rect 28028 43540 28084 43550
rect 28028 43446 28084 43484
rect 29148 43540 29204 43550
rect 29260 43540 29316 45054
rect 29148 43538 29316 43540
rect 29148 43486 29150 43538
rect 29202 43486 29316 43538
rect 29148 43484 29316 43486
rect 29372 44434 29428 45166
rect 29596 45108 29652 45118
rect 29596 45014 29652 45052
rect 29820 44996 29876 45006
rect 29372 44382 29374 44434
rect 29426 44382 29428 44434
rect 29372 44324 29428 44382
rect 29708 44994 29876 44996
rect 29708 44942 29822 44994
rect 29874 44942 29876 44994
rect 29708 44940 29876 44942
rect 27692 43250 27748 43260
rect 29148 43204 29204 43484
rect 29372 43426 29428 44268
rect 29596 44322 29652 44334
rect 29596 44270 29598 44322
rect 29650 44270 29652 44322
rect 29372 43374 29374 43426
rect 29426 43374 29428 43426
rect 29372 43362 29428 43374
rect 29484 43764 29540 43774
rect 29148 43138 29204 43148
rect 27132 42754 27188 42766
rect 27132 42702 27134 42754
rect 27186 42702 27188 42754
rect 27132 41972 27188 42702
rect 27356 42756 27412 42766
rect 27412 42700 27524 42756
rect 27356 42662 27412 42700
rect 27356 41972 27412 41982
rect 27132 41970 27412 41972
rect 27132 41918 27358 41970
rect 27410 41918 27412 41970
rect 27132 41916 27412 41918
rect 27244 41074 27300 41086
rect 27244 41022 27246 41074
rect 27298 41022 27300 41074
rect 27132 40404 27188 40414
rect 27244 40404 27300 41022
rect 27132 40402 27300 40404
rect 27132 40350 27134 40402
rect 27186 40350 27300 40402
rect 27132 40348 27300 40350
rect 27132 39732 27188 40348
rect 27356 40292 27412 41916
rect 27468 41858 27524 42700
rect 27692 42530 27748 42542
rect 27692 42478 27694 42530
rect 27746 42478 27748 42530
rect 27692 41972 27748 42478
rect 27692 41906 27748 41916
rect 28364 42532 28420 42542
rect 27468 41806 27470 41858
rect 27522 41806 27524 41858
rect 27468 41794 27524 41806
rect 27804 41298 27860 41310
rect 27804 41246 27806 41298
rect 27858 41246 27860 41298
rect 27356 40226 27412 40236
rect 27468 41186 27524 41198
rect 27468 41134 27470 41186
rect 27522 41134 27524 41186
rect 27468 40290 27524 41134
rect 27804 41188 27860 41246
rect 27804 41122 27860 41132
rect 27468 40238 27470 40290
rect 27522 40238 27524 40290
rect 27468 39844 27524 40238
rect 27916 40516 27972 40526
rect 27916 40290 27972 40460
rect 27916 40238 27918 40290
rect 27970 40238 27972 40290
rect 27916 40226 27972 40238
rect 28028 40404 28084 40414
rect 27468 39778 27524 39788
rect 27132 39666 27188 39676
rect 28028 39618 28084 40348
rect 28364 40068 28420 42476
rect 29484 42194 29540 43708
rect 29596 43204 29652 44270
rect 29708 43650 29764 44940
rect 29820 44930 29876 44940
rect 29932 44882 29988 45500
rect 30380 45490 30436 45500
rect 29932 44830 29934 44882
rect 29986 44830 29988 44882
rect 29932 44818 29988 44830
rect 30268 45106 30324 45118
rect 30268 45054 30270 45106
rect 30322 45054 30324 45106
rect 30268 44548 30324 45054
rect 30268 44492 30772 44548
rect 30156 44324 30212 44334
rect 30604 44324 30660 44334
rect 30156 44322 30660 44324
rect 30156 44270 30158 44322
rect 30210 44270 30606 44322
rect 30658 44270 30660 44322
rect 30156 44268 30660 44270
rect 30716 44324 30772 44492
rect 30828 44324 30884 44334
rect 30716 44322 30884 44324
rect 30716 44270 30830 44322
rect 30882 44270 30884 44322
rect 30716 44268 30884 44270
rect 30156 44258 30212 44268
rect 30604 44258 30660 44268
rect 29708 43598 29710 43650
rect 29762 43598 29764 43650
rect 29708 43586 29764 43598
rect 30604 43876 30660 43886
rect 29596 43138 29652 43148
rect 30380 43538 30436 43550
rect 30380 43486 30382 43538
rect 30434 43486 30436 43538
rect 29484 42142 29486 42194
rect 29538 42142 29540 42194
rect 29484 42130 29540 42142
rect 30044 42868 30100 42878
rect 30380 42868 30436 43486
rect 30044 42866 30436 42868
rect 30044 42814 30046 42866
rect 30098 42814 30436 42866
rect 30044 42812 30436 42814
rect 30492 43316 30548 43326
rect 30044 42084 30100 42812
rect 30492 42642 30548 43260
rect 30492 42590 30494 42642
rect 30546 42590 30548 42642
rect 30492 42578 30548 42590
rect 30156 42084 30212 42094
rect 30044 42082 30212 42084
rect 30044 42030 30158 42082
rect 30210 42030 30212 42082
rect 30044 42028 30212 42030
rect 29260 41972 29316 41982
rect 29260 41878 29316 41916
rect 29820 41970 29876 41982
rect 29820 41918 29822 41970
rect 29874 41918 29876 41970
rect 28588 41860 28644 41870
rect 28588 41766 28644 41804
rect 29820 41860 29876 41918
rect 29820 41794 29876 41804
rect 30156 41410 30212 42028
rect 30156 41358 30158 41410
rect 30210 41358 30212 41410
rect 30156 41346 30212 41358
rect 28700 41300 28756 41310
rect 28364 40002 28420 40012
rect 28476 40628 28532 40638
rect 28028 39566 28030 39618
rect 28082 39566 28084 39618
rect 28028 39554 28084 39566
rect 27916 39508 27972 39518
rect 27916 39414 27972 39452
rect 27356 39396 27412 39406
rect 27356 38946 27412 39340
rect 28476 39394 28532 40572
rect 28588 39620 28644 39630
rect 28588 39526 28644 39564
rect 28476 39342 28478 39394
rect 28530 39342 28532 39394
rect 28476 39330 28532 39342
rect 27356 38894 27358 38946
rect 27410 38894 27412 38946
rect 27356 38882 27412 38894
rect 28028 39172 28084 39182
rect 28028 38668 28084 39116
rect 28140 38836 28196 38846
rect 28140 38834 28420 38836
rect 28140 38782 28142 38834
rect 28194 38782 28420 38834
rect 28140 38780 28420 38782
rect 28140 38770 28196 38780
rect 27356 38612 28084 38668
rect 28364 38612 28420 38780
rect 26908 37940 26964 37950
rect 26796 37268 26852 37278
rect 26796 36706 26852 37212
rect 26796 36654 26798 36706
rect 26850 36654 26852 36706
rect 26796 36642 26852 36654
rect 26908 34132 26964 37884
rect 27020 36482 27076 36494
rect 27020 36430 27022 36482
rect 27074 36430 27076 36482
rect 27020 36148 27076 36430
rect 27020 36082 27076 36092
rect 27132 35810 27188 35822
rect 27132 35758 27134 35810
rect 27186 35758 27188 35810
rect 27132 35028 27188 35758
rect 27132 34962 27188 34972
rect 26908 34076 27076 34132
rect 26908 33906 26964 33918
rect 26908 33854 26910 33906
rect 26962 33854 26964 33906
rect 26908 33684 26964 33854
rect 26908 33618 26964 33628
rect 26684 33394 26740 33404
rect 26796 33458 26852 33470
rect 26796 33406 26798 33458
rect 26850 33406 26852 33458
rect 26572 33348 26628 33358
rect 26460 33292 26572 33348
rect 26572 33282 26628 33292
rect 26796 32676 26852 33406
rect 26796 32610 26852 32620
rect 26572 32562 26628 32574
rect 26572 32510 26574 32562
rect 26626 32510 26628 32562
rect 26572 32452 26628 32510
rect 26572 32386 26628 32396
rect 26348 31938 26404 31948
rect 26796 31780 26852 31790
rect 26796 31686 26852 31724
rect 25676 31666 25732 31678
rect 25676 31614 25678 31666
rect 25730 31614 25732 31666
rect 25676 30212 25732 31614
rect 27020 30322 27076 34076
rect 27020 30270 27022 30322
rect 27074 30270 27076 30322
rect 27020 30258 27076 30270
rect 26684 30212 26740 30222
rect 25676 30210 26740 30212
rect 25676 30158 26686 30210
rect 26738 30158 26740 30210
rect 25676 30156 26740 30158
rect 25564 30034 25620 30044
rect 26684 29650 26740 30156
rect 27244 30100 27300 30110
rect 26684 29598 26686 29650
rect 26738 29598 26740 29650
rect 26684 29586 26740 29598
rect 27020 30044 27244 30100
rect 25788 29540 25844 29550
rect 25788 29538 25956 29540
rect 25788 29486 25790 29538
rect 25842 29486 25956 29538
rect 25788 29484 25956 29486
rect 25788 29474 25844 29484
rect 25564 28644 25620 28654
rect 25564 27970 25620 28588
rect 25564 27918 25566 27970
rect 25618 27918 25620 27970
rect 25564 27906 25620 27918
rect 25900 28084 25956 29484
rect 26796 29428 26852 29438
rect 26796 29334 26852 29372
rect 27020 29426 27076 30044
rect 27244 30034 27300 30044
rect 27020 29374 27022 29426
rect 27074 29374 27076 29426
rect 27020 29362 27076 29374
rect 26012 29316 26068 29326
rect 26012 28642 26068 29260
rect 27356 29204 27412 38612
rect 28252 38164 28308 38174
rect 28028 38052 28084 38062
rect 28028 37490 28084 37996
rect 28028 37438 28030 37490
rect 28082 37438 28084 37490
rect 28028 37426 28084 37438
rect 27804 37380 27860 37390
rect 27692 37268 27748 37278
rect 27580 37266 27748 37268
rect 27580 37214 27694 37266
rect 27746 37214 27748 37266
rect 27580 37212 27748 37214
rect 27468 37156 27524 37166
rect 27468 37062 27524 37100
rect 27580 36594 27636 37212
rect 27692 37202 27748 37212
rect 27580 36542 27582 36594
rect 27634 36542 27636 36594
rect 27580 36148 27636 36542
rect 27804 36482 27860 37324
rect 27804 36430 27806 36482
rect 27858 36430 27860 36482
rect 27804 36418 27860 36430
rect 27580 36092 28084 36148
rect 28028 35026 28084 36092
rect 28028 34974 28030 35026
rect 28082 34974 28084 35026
rect 28028 34962 28084 34974
rect 27580 34916 27636 34926
rect 27580 34822 27636 34860
rect 27916 34914 27972 34926
rect 27916 34862 27918 34914
rect 27970 34862 27972 34914
rect 27916 33684 27972 34862
rect 28252 33908 28308 38108
rect 28364 38162 28420 38556
rect 28364 38110 28366 38162
rect 28418 38110 28420 38162
rect 28364 38098 28420 38110
rect 28364 37044 28420 37054
rect 28364 36594 28420 36988
rect 28364 36542 28366 36594
rect 28418 36542 28420 36594
rect 28364 36530 28420 36542
rect 28364 36148 28420 36158
rect 28364 35586 28420 36092
rect 28588 35700 28644 35710
rect 28588 35606 28644 35644
rect 28364 35534 28366 35586
rect 28418 35534 28420 35586
rect 28364 35522 28420 35534
rect 28700 34916 28756 41244
rect 29708 41298 29764 41310
rect 29708 41246 29710 41298
rect 29762 41246 29764 41298
rect 29036 41188 29092 41198
rect 29036 41094 29092 41132
rect 28924 40628 28980 40638
rect 28924 40402 28980 40572
rect 28924 40350 28926 40402
rect 28978 40350 28980 40402
rect 28924 40338 28980 40350
rect 29036 40516 29092 40526
rect 29036 40290 29092 40460
rect 29708 40516 29764 41246
rect 29820 41186 29876 41198
rect 29820 41134 29822 41186
rect 29874 41134 29876 41186
rect 29820 40628 29876 41134
rect 29820 40562 29876 40572
rect 29932 41076 29988 41086
rect 29708 40450 29764 40460
rect 29820 40404 29876 40414
rect 29932 40404 29988 41020
rect 30268 40516 30324 40526
rect 30156 40514 30324 40516
rect 30156 40462 30270 40514
rect 30322 40462 30324 40514
rect 30156 40460 30324 40462
rect 29820 40402 29988 40404
rect 29820 40350 29822 40402
rect 29874 40350 29988 40402
rect 29820 40348 29988 40350
rect 30044 40404 30100 40414
rect 29820 40338 29876 40348
rect 30044 40310 30100 40348
rect 29036 40238 29038 40290
rect 29090 40238 29092 40290
rect 29036 40226 29092 40238
rect 28812 39956 28868 39966
rect 28812 38946 28868 39900
rect 29260 39956 29316 39966
rect 29260 39730 29316 39900
rect 30156 39844 30212 40460
rect 30268 40450 30324 40460
rect 30380 40402 30436 40414
rect 30380 40350 30382 40402
rect 30434 40350 30436 40402
rect 30380 39956 30436 40350
rect 30380 39890 30436 39900
rect 29260 39678 29262 39730
rect 29314 39678 29316 39730
rect 29260 39666 29316 39678
rect 29708 39788 30212 39844
rect 28924 39620 28980 39630
rect 28924 39058 28980 39564
rect 28924 39006 28926 39058
rect 28978 39006 28980 39058
rect 28924 38994 28980 39006
rect 29036 39508 29092 39518
rect 28812 38894 28814 38946
rect 28866 38894 28868 38946
rect 28812 38882 28868 38894
rect 29036 38668 29092 39452
rect 29708 39506 29764 39788
rect 29708 39454 29710 39506
rect 29762 39454 29764 39506
rect 29148 38836 29204 38846
rect 29708 38836 29764 39454
rect 30380 39060 30436 39070
rect 30380 38966 30436 39004
rect 29148 38834 29764 38836
rect 29148 38782 29150 38834
rect 29202 38782 29764 38834
rect 29148 38780 29764 38782
rect 29148 38770 29204 38780
rect 29036 38612 29316 38668
rect 29260 38162 29316 38612
rect 29260 38110 29262 38162
rect 29314 38110 29316 38162
rect 29260 38098 29316 38110
rect 29148 38052 29204 38062
rect 29148 37958 29204 37996
rect 29260 37938 29316 37950
rect 29260 37886 29262 37938
rect 29314 37886 29316 37938
rect 28588 34860 28756 34916
rect 28812 37378 28868 37390
rect 28812 37326 28814 37378
rect 28866 37326 28868 37378
rect 28812 35812 28868 37326
rect 29260 36148 29316 37886
rect 29372 37268 29428 37278
rect 29372 37266 29540 37268
rect 29372 37214 29374 37266
rect 29426 37214 29540 37266
rect 29372 37212 29540 37214
rect 29372 37202 29428 37212
rect 29260 36082 29316 36092
rect 29484 37156 29540 37212
rect 29484 36594 29540 37100
rect 29484 36542 29486 36594
rect 29538 36542 29540 36594
rect 29484 36260 29540 36542
rect 28252 33842 28308 33852
rect 28364 34130 28420 34142
rect 28364 34078 28366 34130
rect 28418 34078 28420 34130
rect 27916 33618 27972 33628
rect 27804 33572 27860 33582
rect 27468 33346 27524 33358
rect 27468 33294 27470 33346
rect 27522 33294 27524 33346
rect 27468 31892 27524 33294
rect 27804 33346 27860 33516
rect 27804 33294 27806 33346
rect 27858 33294 27860 33346
rect 27804 33282 27860 33294
rect 28252 33346 28308 33358
rect 28252 33294 28254 33346
rect 28306 33294 28308 33346
rect 27916 33234 27972 33246
rect 27916 33182 27918 33234
rect 27970 33182 27972 33234
rect 27468 31826 27524 31836
rect 27692 32564 27748 32574
rect 26908 29148 27412 29204
rect 27580 29428 27636 29438
rect 26908 28754 26964 29148
rect 26908 28702 26910 28754
rect 26962 28702 26964 28754
rect 26908 28690 26964 28702
rect 27132 28756 27188 28766
rect 26012 28590 26014 28642
rect 26066 28590 26068 28642
rect 26012 28578 26068 28590
rect 27020 28642 27076 28654
rect 27020 28590 27022 28642
rect 27074 28590 27076 28642
rect 27020 28084 27076 28590
rect 25788 26964 25844 26974
rect 25564 26404 25620 26414
rect 25564 26310 25620 26348
rect 25676 25620 25732 25630
rect 25676 25506 25732 25564
rect 25676 25454 25678 25506
rect 25730 25454 25732 25506
rect 25676 25442 25732 25454
rect 25788 25506 25844 26908
rect 25788 25454 25790 25506
rect 25842 25454 25844 25506
rect 25788 25442 25844 25454
rect 25564 25284 25620 25294
rect 25452 25282 25620 25284
rect 25452 25230 25566 25282
rect 25618 25230 25620 25282
rect 25452 25228 25620 25230
rect 24780 25190 24836 25228
rect 25564 25218 25620 25228
rect 23884 24770 23940 24780
rect 24108 25004 24724 25060
rect 24108 24722 24164 25004
rect 24444 24836 24500 24846
rect 24444 24742 24500 24780
rect 24556 24834 24612 24846
rect 24556 24782 24558 24834
rect 24610 24782 24612 24834
rect 24108 24670 24110 24722
rect 24162 24670 24164 24722
rect 24108 24658 24164 24670
rect 24556 24724 24612 24782
rect 24556 24658 24612 24668
rect 24556 24500 24612 24510
rect 23212 24444 23380 24500
rect 23100 23774 23102 23826
rect 23154 23774 23156 23826
rect 23100 23762 23156 23774
rect 23212 24276 23268 24286
rect 23212 23826 23268 24220
rect 23324 23940 23380 24444
rect 24108 24498 24612 24500
rect 24108 24446 24558 24498
rect 24610 24446 24612 24498
rect 24108 24444 24612 24446
rect 23324 23874 23380 23884
rect 23996 24388 24052 24398
rect 23996 23828 24052 24332
rect 23212 23774 23214 23826
rect 23266 23774 23268 23826
rect 23212 23762 23268 23774
rect 23884 23826 24052 23828
rect 23884 23774 23998 23826
rect 24050 23774 24052 23826
rect 23884 23772 24052 23774
rect 23324 23714 23380 23726
rect 23324 23662 23326 23714
rect 23378 23662 23380 23714
rect 22988 23326 22990 23378
rect 23042 23326 23044 23378
rect 22988 23314 23044 23326
rect 23100 23604 23156 23614
rect 23100 23156 23156 23548
rect 23212 23492 23268 23502
rect 23212 23378 23268 23436
rect 23212 23326 23214 23378
rect 23266 23326 23268 23378
rect 23212 23314 23268 23326
rect 23324 23380 23380 23662
rect 23436 23716 23492 23726
rect 23772 23716 23828 23726
rect 23492 23714 23828 23716
rect 23492 23662 23774 23714
rect 23826 23662 23828 23714
rect 23492 23660 23828 23662
rect 23436 23622 23492 23660
rect 23772 23650 23828 23660
rect 23324 23324 23716 23380
rect 23324 23156 23380 23166
rect 23100 23154 23380 23156
rect 23100 23102 23326 23154
rect 23378 23102 23380 23154
rect 23100 23100 23380 23102
rect 23324 23090 23380 23100
rect 22036 22988 22148 23044
rect 22428 23042 22932 23044
rect 22428 22990 22654 23042
rect 22706 22990 22932 23042
rect 22428 22988 22932 22990
rect 21980 22978 22036 22988
rect 22428 22484 22484 22988
rect 22652 22978 22708 22988
rect 21420 22430 21422 22482
rect 21474 22430 21476 22482
rect 21420 22418 21476 22430
rect 22204 22482 22484 22484
rect 22204 22430 22430 22482
rect 22482 22430 22484 22482
rect 22204 22428 22484 22430
rect 21980 22146 22036 22158
rect 21980 22094 21982 22146
rect 22034 22094 22036 22146
rect 21980 22036 22036 22094
rect 21868 21980 21980 22036
rect 21308 21758 21310 21810
rect 21362 21758 21364 21810
rect 21308 21746 21364 21758
rect 21644 21812 21700 21822
rect 21868 21812 21924 21980
rect 21980 21970 22036 21980
rect 22204 21812 22260 22428
rect 22428 22418 22484 22428
rect 23660 22482 23716 23324
rect 23884 23268 23940 23772
rect 23996 23762 24052 23772
rect 24108 23826 24164 24444
rect 24556 24434 24612 24444
rect 24556 24050 24612 24062
rect 24556 23998 24558 24050
rect 24610 23998 24612 24050
rect 24108 23774 24110 23826
rect 24162 23774 24164 23826
rect 24108 23762 24164 23774
rect 24220 23826 24276 23838
rect 24220 23774 24222 23826
rect 24274 23774 24276 23826
rect 24220 23604 24276 23774
rect 24556 23828 24612 23998
rect 24668 23940 24724 25004
rect 25788 25172 25844 25182
rect 25788 24722 25844 25116
rect 25900 24948 25956 28028
rect 26796 28028 27076 28084
rect 26124 27860 26180 27870
rect 26124 27766 26180 27804
rect 26236 27748 26292 27758
rect 26236 27654 26292 27692
rect 26124 27076 26180 27086
rect 26012 26964 26068 26974
rect 26124 26964 26180 27020
rect 26012 26962 26180 26964
rect 26012 26910 26014 26962
rect 26066 26910 26180 26962
rect 26012 26908 26180 26910
rect 26012 26898 26068 26908
rect 26012 26516 26068 26526
rect 26012 25844 26068 26460
rect 26012 25778 26068 25788
rect 26124 25620 26180 26908
rect 26572 27074 26628 27086
rect 26572 27022 26574 27074
rect 26626 27022 26628 27074
rect 26572 26628 26628 27022
rect 26796 27074 26852 28028
rect 26796 27022 26798 27074
rect 26850 27022 26852 27074
rect 26796 26964 26852 27022
rect 26796 26898 26852 26908
rect 26908 27746 26964 27758
rect 26908 27694 26910 27746
rect 26962 27694 26964 27746
rect 26684 26852 26740 26862
rect 26684 26740 26740 26796
rect 26908 26740 26964 27694
rect 27132 26908 27188 28700
rect 27356 28308 27412 28318
rect 27356 27858 27412 28252
rect 27356 27806 27358 27858
rect 27410 27806 27412 27858
rect 27356 26908 27412 27806
rect 26684 26684 26964 26740
rect 27020 26852 27188 26908
rect 27244 26852 27412 26908
rect 27468 28084 27524 28094
rect 26572 26562 26628 26572
rect 26796 25844 26852 26684
rect 27020 26290 27076 26852
rect 27020 26238 27022 26290
rect 27074 26238 27076 26290
rect 27020 26226 27076 26238
rect 27132 26628 27188 26638
rect 27132 25844 27188 26572
rect 26796 25778 26852 25788
rect 27020 25788 27188 25844
rect 26124 25618 26292 25620
rect 26124 25566 26126 25618
rect 26178 25566 26292 25618
rect 26124 25564 26292 25566
rect 26124 25554 26180 25564
rect 26012 24948 26068 24958
rect 25900 24946 26068 24948
rect 25900 24894 26014 24946
rect 26066 24894 26068 24946
rect 25900 24892 26068 24894
rect 26012 24882 26068 24892
rect 25788 24670 25790 24722
rect 25842 24670 25844 24722
rect 24892 23940 24948 23950
rect 24668 23938 24948 23940
rect 24668 23886 24894 23938
rect 24946 23886 24948 23938
rect 24668 23884 24948 23886
rect 24556 23762 24612 23772
rect 24220 23538 24276 23548
rect 23660 22430 23662 22482
rect 23714 22430 23716 22482
rect 23660 22418 23716 22430
rect 23772 23212 23940 23268
rect 22988 22370 23044 22382
rect 22988 22318 22990 22370
rect 23042 22318 23044 22370
rect 22988 22148 23044 22318
rect 22988 22082 23044 22092
rect 22876 22036 22932 22046
rect 22876 21812 22932 21980
rect 23436 22036 23492 22046
rect 23436 21812 23492 21980
rect 21644 21810 21924 21812
rect 21644 21758 21646 21810
rect 21698 21758 21924 21810
rect 21644 21756 21924 21758
rect 21980 21810 22260 21812
rect 21980 21758 22206 21810
rect 22258 21758 22260 21810
rect 21980 21756 22260 21758
rect 21644 21746 21700 21756
rect 21980 21700 22036 21756
rect 22204 21746 22260 21756
rect 22652 21810 22932 21812
rect 22652 21758 22878 21810
rect 22930 21758 22932 21810
rect 22652 21756 22932 21758
rect 21084 21606 21140 21644
rect 21756 21644 22036 21700
rect 20972 21588 21028 21598
rect 21756 21588 21812 21644
rect 20524 21586 21028 21588
rect 20524 21534 20974 21586
rect 21026 21534 21028 21586
rect 20524 21532 21028 21534
rect 20412 21474 20468 21486
rect 20412 21422 20414 21474
rect 20466 21422 20468 21474
rect 20412 21028 20468 21422
rect 20412 20962 20468 20972
rect 20524 20914 20580 21532
rect 20972 21522 21028 21532
rect 21532 21586 21812 21588
rect 21532 21534 21758 21586
rect 21810 21534 21812 21586
rect 21532 21532 21812 21534
rect 20636 21364 20692 21374
rect 20636 21270 20692 21308
rect 21308 21364 21364 21374
rect 20524 20862 20526 20914
rect 20578 20862 20580 20914
rect 20524 20850 20580 20862
rect 20636 21140 20692 21150
rect 20412 20804 20468 20814
rect 20412 20710 20468 20748
rect 20636 20802 20692 21084
rect 20636 20750 20638 20802
rect 20690 20750 20692 20802
rect 20636 20580 20692 20750
rect 21308 20804 21364 21308
rect 21420 21028 21476 21038
rect 21420 20934 21476 20972
rect 21308 20738 21364 20748
rect 21532 20916 21588 21532
rect 21756 21522 21812 21532
rect 21644 21362 21700 21374
rect 21644 21310 21646 21362
rect 21698 21310 21700 21362
rect 21644 21140 21700 21310
rect 21644 21074 21700 21084
rect 22540 20916 22596 20926
rect 21532 20802 21588 20860
rect 21532 20750 21534 20802
rect 21586 20750 21588 20802
rect 21532 20738 21588 20750
rect 22092 20914 22596 20916
rect 22092 20862 22542 20914
rect 22594 20862 22596 20914
rect 22092 20860 22596 20862
rect 20412 20524 20692 20580
rect 20748 20692 20804 20702
rect 20412 20242 20468 20524
rect 20748 20244 20804 20636
rect 21420 20692 21476 20702
rect 21420 20598 21476 20636
rect 22092 20692 22148 20860
rect 22540 20850 22596 20860
rect 22652 20914 22708 21756
rect 22876 21746 22932 21756
rect 23324 21810 23492 21812
rect 23324 21758 23438 21810
rect 23490 21758 23492 21810
rect 23324 21756 23492 21758
rect 23100 21700 23156 21710
rect 23100 21606 23156 21644
rect 22652 20862 22654 20914
rect 22706 20862 22708 20914
rect 22652 20850 22708 20862
rect 22764 21588 22820 21598
rect 22092 20598 22148 20636
rect 22204 20692 22260 20702
rect 22764 20692 22820 21532
rect 22204 20690 22820 20692
rect 22204 20638 22206 20690
rect 22258 20638 22820 20690
rect 22204 20636 22820 20638
rect 22204 20626 22260 20636
rect 21868 20578 21924 20590
rect 23100 20580 23156 20590
rect 21868 20526 21870 20578
rect 21922 20526 21924 20578
rect 21868 20356 21924 20526
rect 22988 20578 23156 20580
rect 22988 20526 23102 20578
rect 23154 20526 23156 20578
rect 22988 20524 23156 20526
rect 20972 20244 21028 20254
rect 20412 20190 20414 20242
rect 20466 20190 20468 20242
rect 20412 20178 20468 20190
rect 20524 20188 20804 20244
rect 20860 20188 20972 20244
rect 20524 20130 20580 20188
rect 20524 20078 20526 20130
rect 20578 20078 20580 20130
rect 20524 20066 20580 20078
rect 20636 20020 20692 20030
rect 20860 20020 20916 20188
rect 20972 20178 21028 20188
rect 21308 20242 21364 20254
rect 21308 20190 21310 20242
rect 21362 20190 21364 20242
rect 21308 20188 21364 20190
rect 21308 20132 21700 20188
rect 21532 20020 21588 20030
rect 20636 20018 20916 20020
rect 20636 19966 20638 20018
rect 20690 19966 20916 20018
rect 20636 19964 20916 19966
rect 21196 20018 21588 20020
rect 21196 19966 21534 20018
rect 21586 19966 21588 20018
rect 21196 19964 21588 19966
rect 20636 19954 20692 19964
rect 20300 19254 20356 19292
rect 20188 17726 20190 17778
rect 20242 17726 20244 17778
rect 20188 17714 20244 17726
rect 20524 17780 20580 17790
rect 20524 17686 20580 17724
rect 19836 17276 20100 17286
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 19836 17210 20100 17220
rect 19628 16942 19630 16994
rect 19682 16942 19684 16994
rect 19628 16930 19684 16942
rect 20076 17108 20132 17118
rect 19740 16324 19796 16334
rect 19516 16322 19796 16324
rect 19516 16270 19742 16322
rect 19794 16270 19796 16322
rect 19516 16268 19796 16270
rect 19740 16258 19796 16268
rect 19404 16044 19796 16100
rect 19740 15986 19796 16044
rect 19628 15932 19684 15942
rect 19516 15930 19684 15932
rect 19516 15878 19630 15930
rect 19682 15878 19684 15930
rect 19740 15934 19742 15986
rect 19794 15934 19796 15986
rect 19740 15922 19796 15934
rect 19516 15876 19684 15878
rect 19516 15764 19572 15876
rect 19628 15866 19684 15876
rect 20076 15876 20132 17052
rect 20412 16100 20468 16110
rect 20412 15986 20468 16044
rect 21196 16100 21252 19964
rect 21532 19954 21588 19964
rect 21420 19236 21476 19246
rect 21308 19180 21420 19236
rect 21308 17780 21364 19180
rect 21420 19170 21476 19180
rect 21532 19234 21588 19246
rect 21532 19182 21534 19234
rect 21586 19182 21588 19234
rect 21532 18340 21588 19182
rect 21644 18900 21700 20132
rect 21868 20132 21924 20300
rect 22764 20468 22820 20478
rect 21868 20066 21924 20076
rect 22092 20130 22148 20142
rect 22316 20132 22372 20142
rect 22092 20078 22094 20130
rect 22146 20078 22148 20130
rect 21980 20018 22036 20030
rect 21980 19966 21982 20018
rect 22034 19966 22036 20018
rect 21980 19684 22036 19966
rect 21980 19618 22036 19628
rect 22092 19460 22148 20078
rect 22204 20130 22372 20132
rect 22204 20078 22318 20130
rect 22370 20078 22372 20130
rect 22204 20076 22372 20078
rect 22204 20020 22260 20076
rect 22316 20066 22372 20076
rect 22652 20132 22708 20142
rect 22652 20038 22708 20076
rect 22764 20130 22820 20412
rect 22764 20078 22766 20130
rect 22818 20078 22820 20130
rect 22764 20066 22820 20078
rect 22204 19954 22260 19964
rect 22652 19796 22708 19806
rect 22652 19702 22708 19740
rect 22092 19404 22372 19460
rect 21756 19348 21812 19358
rect 21756 19122 21812 19292
rect 22092 19236 22148 19246
rect 22092 19142 22148 19180
rect 21756 19070 21758 19122
rect 21810 19070 21812 19122
rect 21756 19058 21812 19070
rect 21644 18844 21812 18900
rect 21420 17780 21476 17790
rect 21308 17778 21476 17780
rect 21308 17726 21422 17778
rect 21474 17726 21476 17778
rect 21308 17724 21476 17726
rect 21420 17714 21476 17724
rect 21532 17106 21588 18284
rect 21532 17054 21534 17106
rect 21586 17054 21588 17106
rect 21532 17042 21588 17054
rect 21644 18562 21700 18574
rect 21644 18510 21646 18562
rect 21698 18510 21700 18562
rect 21644 17556 21700 18510
rect 21644 16994 21700 17500
rect 21644 16942 21646 16994
rect 21698 16942 21700 16994
rect 21644 16930 21700 16942
rect 21756 17892 21812 18844
rect 21196 16034 21252 16044
rect 21644 16772 21700 16782
rect 21644 16212 21700 16716
rect 21644 16098 21700 16156
rect 21644 16046 21646 16098
rect 21698 16046 21700 16098
rect 21644 16034 21700 16046
rect 20412 15934 20414 15986
rect 20466 15934 20468 15986
rect 20412 15876 20468 15934
rect 20748 15988 20804 15998
rect 20748 15894 20804 15932
rect 21308 15986 21364 15998
rect 21308 15934 21310 15986
rect 21362 15934 21364 15986
rect 20076 15820 20244 15876
rect 19628 15764 19684 15774
rect 19516 15708 19628 15764
rect 19628 15698 19684 15708
rect 19836 15708 20100 15718
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 19836 15642 20100 15652
rect 20188 15540 20244 15820
rect 20412 15810 20468 15820
rect 19180 15426 19348 15428
rect 19180 15374 19182 15426
rect 19234 15374 19348 15426
rect 19180 15372 19348 15374
rect 20076 15484 20244 15540
rect 20524 15538 20580 15550
rect 20524 15486 20526 15538
rect 20578 15486 20580 15538
rect 19180 15362 19236 15372
rect 19068 15262 19070 15314
rect 19122 15262 19124 15314
rect 19068 15250 19124 15262
rect 19740 15316 19796 15326
rect 19292 15204 19348 15214
rect 18956 15092 19124 15148
rect 18844 14812 19012 14868
rect 18844 14644 18900 14654
rect 18732 14642 18900 14644
rect 18732 14590 18846 14642
rect 18898 14590 18900 14642
rect 18732 14588 18900 14590
rect 18844 14578 18900 14588
rect 18956 13972 19012 14812
rect 18396 13694 18398 13746
rect 18450 13694 18452 13746
rect 17948 13654 18004 13692
rect 17724 13020 18004 13076
rect 17836 12740 17892 12750
rect 17612 12738 17892 12740
rect 17612 12686 17838 12738
rect 17890 12686 17892 12738
rect 17612 12684 17892 12686
rect 17500 12404 17556 12414
rect 17500 12310 17556 12348
rect 17724 11788 17780 12684
rect 17836 12674 17892 12684
rect 17612 11732 17780 11788
rect 17836 12404 17892 12414
rect 17948 12404 18004 13020
rect 18172 12852 18228 12862
rect 18228 12796 18340 12852
rect 18172 12758 18228 12796
rect 17836 12402 17948 12404
rect 17836 12350 17838 12402
rect 17890 12350 17948 12402
rect 17836 12348 17948 12350
rect 17612 11060 17668 11732
rect 17724 11508 17780 11518
rect 17724 11414 17780 11452
rect 17612 11004 17780 11060
rect 17164 10882 17220 10892
rect 17052 10770 17108 10780
rect 17612 10836 17668 10846
rect 17612 10742 17668 10780
rect 16604 10670 16606 10722
rect 16658 10670 16660 10722
rect 16604 10658 16660 10670
rect 16828 10722 16884 10734
rect 16828 10670 16830 10722
rect 16882 10670 16884 10722
rect 16828 10612 16884 10670
rect 16940 10612 16996 10622
rect 16828 10556 16940 10612
rect 16940 10546 16996 10556
rect 15036 8372 15204 8428
rect 15148 8260 15204 8372
rect 15372 8260 15428 8270
rect 15148 8258 15428 8260
rect 15148 8206 15374 8258
rect 15426 8206 15428 8258
rect 15148 8204 15428 8206
rect 4476 7084 4740 7094
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4476 7018 4740 7028
rect 15372 6692 15428 8204
rect 16044 8148 16100 8158
rect 16044 8146 16436 8148
rect 16044 8094 16046 8146
rect 16098 8094 16436 8146
rect 16044 8092 16436 8094
rect 16044 8082 16100 8092
rect 16380 7698 16436 8092
rect 16380 7646 16382 7698
rect 16434 7646 16436 7698
rect 16380 7634 16436 7646
rect 16268 7476 16324 7486
rect 16492 7476 16548 9100
rect 17724 8820 17780 11004
rect 17836 10836 17892 12348
rect 17948 12338 18004 12348
rect 17948 12180 18004 12190
rect 17948 12086 18004 12124
rect 18060 12178 18116 12190
rect 18060 12126 18062 12178
rect 18114 12126 18116 12178
rect 18060 11508 18116 12126
rect 18060 11442 18116 11452
rect 18284 11394 18340 12796
rect 18396 12178 18452 13694
rect 18844 13916 19012 13972
rect 18732 13636 18788 13646
rect 18732 13542 18788 13580
rect 18732 12964 18788 12974
rect 18844 12964 18900 13916
rect 18732 12962 18900 12964
rect 18732 12910 18734 12962
rect 18786 12910 18900 12962
rect 18732 12908 18900 12910
rect 18956 13746 19012 13758
rect 18956 13694 18958 13746
rect 19010 13694 19012 13746
rect 18956 13636 19012 13694
rect 18732 12898 18788 12908
rect 18956 12738 19012 13580
rect 18956 12686 18958 12738
rect 19010 12686 19012 12738
rect 18956 12628 19012 12686
rect 18396 12126 18398 12178
rect 18450 12126 18452 12178
rect 18396 11732 18452 12126
rect 18620 12572 19012 12628
rect 19068 12852 19124 15092
rect 19180 14530 19236 14542
rect 19180 14478 19182 14530
rect 19234 14478 19236 14530
rect 19180 14084 19236 14478
rect 19292 14530 19348 15148
rect 19292 14478 19294 14530
rect 19346 14478 19348 14530
rect 19292 14466 19348 14478
rect 19740 14530 19796 15260
rect 19740 14478 19742 14530
rect 19794 14478 19796 14530
rect 19740 14466 19796 14478
rect 19516 14306 19572 14318
rect 19516 14254 19518 14306
rect 19570 14254 19572 14306
rect 19516 14196 19572 14254
rect 20076 14308 20132 15484
rect 20524 15148 20580 15486
rect 20748 15540 20804 15550
rect 20748 15148 20804 15484
rect 21308 15316 21364 15934
rect 21308 15250 21364 15260
rect 21420 15874 21476 15886
rect 21420 15822 21422 15874
rect 21474 15822 21476 15874
rect 21420 15148 21476 15822
rect 21756 15148 21812 17836
rect 22204 18452 22260 18462
rect 21868 17666 21924 17678
rect 21868 17614 21870 17666
rect 21922 17614 21924 17666
rect 21868 17108 21924 17614
rect 22204 17668 22260 18396
rect 22204 17602 22260 17612
rect 21868 17042 21924 17052
rect 22316 16884 22372 19404
rect 22652 19348 22708 19358
rect 22652 18450 22708 19292
rect 22652 18398 22654 18450
rect 22706 18398 22708 18450
rect 22652 18386 22708 18398
rect 22988 18450 23044 20524
rect 23100 20514 23156 20524
rect 23324 20242 23380 21756
rect 23436 21746 23492 21756
rect 23548 21924 23604 21934
rect 23772 21924 23828 23212
rect 23884 23044 23940 23054
rect 24332 23044 24388 23054
rect 24892 23044 24948 23884
rect 25676 23828 25732 23838
rect 25676 23734 25732 23772
rect 25452 23716 25508 23726
rect 23884 23042 24948 23044
rect 23884 22990 23886 23042
rect 23938 22990 24334 23042
rect 24386 22990 24948 23042
rect 23884 22988 24948 22990
rect 25340 23604 25396 23614
rect 25340 23044 25396 23548
rect 23884 22148 23940 22988
rect 24332 22978 24388 22988
rect 25340 22950 25396 22988
rect 25228 22932 25284 22942
rect 23884 22082 23940 22092
rect 24444 22260 24500 22270
rect 23772 21868 24388 21924
rect 23548 21028 23604 21868
rect 24332 21810 24388 21868
rect 24332 21758 24334 21810
rect 24386 21758 24388 21810
rect 24332 21746 24388 21758
rect 23884 21698 23940 21710
rect 23884 21646 23886 21698
rect 23938 21646 23940 21698
rect 23660 21586 23716 21598
rect 23660 21534 23662 21586
rect 23714 21534 23716 21586
rect 23660 21364 23716 21534
rect 23660 21298 23716 21308
rect 23884 21140 23940 21646
rect 23884 21074 23940 21084
rect 23996 21586 24052 21598
rect 23996 21534 23998 21586
rect 24050 21534 24052 21586
rect 23996 21476 24052 21534
rect 23548 20972 23828 21028
rect 23436 20692 23492 20702
rect 23436 20598 23492 20636
rect 23324 20190 23326 20242
rect 23378 20190 23380 20242
rect 23324 20178 23380 20190
rect 23660 20578 23716 20590
rect 23660 20526 23662 20578
rect 23714 20526 23716 20578
rect 23660 20244 23716 20526
rect 23660 20178 23716 20188
rect 23548 20018 23604 20030
rect 23548 19966 23550 20018
rect 23602 19966 23604 20018
rect 22988 18398 22990 18450
rect 23042 18398 23044 18450
rect 22764 18338 22820 18350
rect 22764 18286 22766 18338
rect 22818 18286 22820 18338
rect 22764 17892 22820 18286
rect 22540 17836 22820 17892
rect 22540 17778 22596 17836
rect 22540 17726 22542 17778
rect 22594 17726 22596 17778
rect 22540 17714 22596 17726
rect 22764 17668 22820 17678
rect 21980 16660 22036 16670
rect 21868 15986 21924 15998
rect 21868 15934 21870 15986
rect 21922 15934 21924 15986
rect 21868 15540 21924 15934
rect 21868 15474 21924 15484
rect 20412 15092 20580 15148
rect 20636 15092 20804 15148
rect 20860 15092 21476 15148
rect 21644 15092 21812 15148
rect 20076 14252 20244 14308
rect 19516 14140 19684 14196
rect 19180 14028 19572 14084
rect 19516 13970 19572 14028
rect 19516 13918 19518 13970
rect 19570 13918 19572 13970
rect 19516 13906 19572 13918
rect 19628 13972 19684 14140
rect 19836 14140 20100 14150
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 19836 14074 20100 14084
rect 20188 13972 20244 14252
rect 19628 13916 19796 13972
rect 19404 13746 19460 13758
rect 19404 13694 19406 13746
rect 19458 13694 19460 13746
rect 19404 13524 19460 13694
rect 19628 13748 19684 13758
rect 19628 13654 19684 13692
rect 19404 13458 19460 13468
rect 18620 12180 18676 12572
rect 18732 12404 18788 12414
rect 18732 12310 18788 12348
rect 19068 12402 19124 12796
rect 19740 12852 19796 13916
rect 20076 13916 20244 13972
rect 20300 14306 20356 14318
rect 20300 14254 20302 14306
rect 20354 14254 20356 14306
rect 20076 13746 20132 13916
rect 20076 13694 20078 13746
rect 20130 13694 20132 13746
rect 20076 13682 20132 13694
rect 20188 13636 20244 13646
rect 20300 13636 20356 14254
rect 20244 13580 20356 13636
rect 20188 13570 20244 13580
rect 19740 12786 19796 12796
rect 20188 13412 20244 13422
rect 19836 12572 20100 12582
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 19836 12506 20100 12516
rect 19068 12350 19070 12402
rect 19122 12350 19124 12402
rect 19068 12338 19124 12350
rect 19740 12292 19796 12302
rect 18844 12180 18900 12190
rect 18620 12124 18788 12180
rect 18396 11676 18564 11732
rect 18284 11342 18286 11394
rect 18338 11342 18340 11394
rect 18284 11330 18340 11342
rect 18060 11172 18116 11182
rect 18060 11078 18116 11116
rect 17948 10836 18004 10846
rect 17836 10834 18004 10836
rect 17836 10782 17950 10834
rect 18002 10782 18004 10834
rect 17836 10780 18004 10782
rect 17948 10770 18004 10780
rect 18284 10836 18340 10846
rect 18060 10612 18116 10622
rect 18060 10518 18116 10556
rect 18172 10610 18228 10622
rect 18172 10558 18174 10610
rect 18226 10558 18228 10610
rect 17836 9940 17892 9950
rect 18172 9940 18228 10558
rect 17836 9938 18228 9940
rect 17836 9886 17838 9938
rect 17890 9886 18228 9938
rect 17836 9884 18228 9886
rect 18284 9938 18340 10780
rect 18284 9886 18286 9938
rect 18338 9886 18340 9938
rect 17836 9044 17892 9884
rect 18284 9874 18340 9886
rect 18508 10610 18564 11676
rect 18732 11396 18788 12124
rect 18508 10558 18510 10610
rect 18562 10558 18564 10610
rect 18284 9266 18340 9278
rect 18284 9214 18286 9266
rect 18338 9214 18340 9266
rect 17836 8978 17892 8988
rect 17948 9156 18004 9166
rect 17948 9042 18004 9100
rect 17948 8990 17950 9042
rect 18002 8990 18004 9042
rect 17948 8978 18004 8990
rect 17724 8764 18004 8820
rect 17948 8260 18004 8764
rect 17052 7700 17108 7710
rect 16828 7644 17052 7700
rect 16828 7586 16884 7644
rect 17052 7634 17108 7644
rect 17948 7698 18004 8204
rect 18172 8370 18228 8382
rect 18172 8318 18174 8370
rect 18226 8318 18228 8370
rect 17948 7646 17950 7698
rect 18002 7646 18004 7698
rect 17948 7634 18004 7646
rect 18060 7700 18116 7710
rect 18060 7606 18116 7644
rect 16828 7534 16830 7586
rect 16882 7534 16884 7586
rect 16828 7522 16884 7534
rect 16268 7474 16548 7476
rect 16268 7422 16270 7474
rect 16322 7422 16548 7474
rect 16268 7420 16548 7422
rect 16604 7474 16660 7486
rect 16604 7422 16606 7474
rect 16658 7422 16660 7474
rect 16268 7410 16324 7420
rect 16604 7364 16660 7422
rect 18172 7476 18228 8318
rect 18172 7382 18228 7420
rect 16604 7298 16660 7308
rect 17500 7364 17556 7374
rect 17500 7270 17556 7308
rect 18284 7140 18340 9214
rect 18396 9156 18452 9166
rect 18396 9062 18452 9100
rect 18508 7474 18564 10558
rect 18620 10948 18676 10958
rect 18620 9268 18676 10892
rect 18732 10388 18788 11340
rect 18844 11394 18900 12124
rect 19740 11956 19796 12236
rect 19740 11890 19796 11900
rect 20188 11788 20244 13356
rect 20300 12180 20356 12218
rect 20412 12180 20468 15092
rect 20636 14642 20692 15092
rect 20636 14590 20638 14642
rect 20690 14590 20692 14642
rect 20636 14578 20692 14590
rect 20524 14420 20580 14430
rect 20524 14326 20580 14364
rect 20748 14308 20804 14318
rect 20636 14306 20804 14308
rect 20636 14254 20750 14306
rect 20802 14254 20804 14306
rect 20636 14252 20804 14254
rect 20636 13748 20692 14252
rect 20748 14242 20804 14252
rect 20748 13860 20804 13870
rect 20860 13860 20916 15092
rect 20748 13858 20916 13860
rect 20748 13806 20750 13858
rect 20802 13806 20916 13858
rect 20748 13804 20916 13806
rect 20748 13794 20804 13804
rect 20524 12404 20580 12414
rect 20636 12404 20692 13692
rect 21308 13076 21364 13086
rect 21308 12964 21364 13020
rect 20580 12348 20692 12404
rect 21196 12962 21364 12964
rect 21196 12910 21310 12962
rect 21362 12910 21364 12962
rect 21196 12908 21364 12910
rect 20524 12310 20580 12348
rect 20356 12124 20468 12180
rect 20300 12114 20356 12124
rect 20300 11956 20356 11966
rect 20356 11900 20468 11956
rect 20300 11890 20356 11900
rect 20076 11732 20244 11788
rect 19964 11396 20020 11406
rect 18844 11342 18846 11394
rect 18898 11342 18900 11394
rect 18844 11172 18900 11342
rect 19292 11394 20020 11396
rect 19292 11342 19966 11394
rect 20018 11342 20020 11394
rect 19292 11340 20020 11342
rect 18844 11106 18900 11116
rect 19068 11172 19124 11182
rect 19292 11172 19348 11340
rect 19068 11170 19348 11172
rect 19068 11118 19070 11170
rect 19122 11118 19348 11170
rect 19068 11116 19348 11118
rect 19404 11172 19460 11182
rect 19068 11106 19124 11116
rect 19404 11078 19460 11116
rect 19180 10836 19236 10846
rect 19180 10612 19236 10780
rect 19628 10724 19684 11340
rect 19964 11330 20020 11340
rect 20076 11396 20132 11732
rect 20076 11340 20356 11396
rect 19740 11172 19796 11182
rect 20076 11172 20132 11340
rect 19740 11170 20132 11172
rect 19740 11118 19742 11170
rect 19794 11118 20132 11170
rect 19740 11116 20132 11118
rect 20188 11170 20244 11182
rect 20188 11118 20190 11170
rect 20242 11118 20244 11170
rect 19740 11106 19796 11116
rect 19836 11004 20100 11014
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 19836 10938 20100 10948
rect 20188 10836 20244 11118
rect 19964 10780 20244 10836
rect 19628 10668 19908 10724
rect 19180 10610 19684 10612
rect 19180 10558 19182 10610
rect 19234 10558 19684 10610
rect 19180 10556 19684 10558
rect 19180 10546 19236 10556
rect 18732 10332 19236 10388
rect 18620 9202 18676 9212
rect 19068 9604 19124 9614
rect 19068 9266 19124 9548
rect 19068 9214 19070 9266
rect 19122 9214 19124 9266
rect 19068 9156 19124 9214
rect 18620 9044 18676 9054
rect 18620 9042 18900 9044
rect 18620 8990 18622 9042
rect 18674 8990 18900 9042
rect 18620 8988 18900 8990
rect 18620 8978 18676 8988
rect 18844 8370 18900 8988
rect 19068 8596 19124 9100
rect 19068 8530 19124 8540
rect 18844 8318 18846 8370
rect 18898 8318 18900 8370
rect 18844 8306 18900 8318
rect 18732 8260 18788 8270
rect 18732 8166 18788 8204
rect 18956 8260 19012 8270
rect 19012 8204 19124 8260
rect 18956 8166 19012 8204
rect 18508 7422 18510 7474
rect 18562 7422 18564 7474
rect 18508 7410 18564 7422
rect 17164 7084 18340 7140
rect 18396 7364 18452 7374
rect 15372 6626 15428 6636
rect 16492 6692 16548 6702
rect 4476 5516 4740 5526
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4476 5450 4740 5460
rect 16492 5124 16548 6636
rect 17164 6690 17220 7084
rect 17164 6638 17166 6690
rect 17218 6638 17220 6690
rect 17164 6626 17220 6638
rect 18396 6130 18452 7308
rect 19068 6804 19124 8204
rect 19180 8146 19236 10332
rect 19628 10164 19684 10556
rect 19628 8372 19684 10108
rect 19852 9604 19908 10668
rect 19964 10722 20020 10780
rect 19964 10670 19966 10722
rect 20018 10670 20020 10722
rect 19964 10658 20020 10670
rect 19852 9548 20244 9604
rect 19836 9436 20100 9446
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 19836 9370 20100 9380
rect 19852 9268 19908 9278
rect 19852 9174 19908 9212
rect 20076 9156 20132 9166
rect 20188 9156 20244 9548
rect 20076 9154 20244 9156
rect 20076 9102 20078 9154
rect 20130 9102 20244 9154
rect 20076 9100 20244 9102
rect 19740 8372 19796 8382
rect 19180 8094 19182 8146
rect 19234 8094 19236 8146
rect 19180 8082 19236 8094
rect 19292 8370 19796 8372
rect 19292 8318 19742 8370
rect 19794 8318 19796 8370
rect 19292 8316 19796 8318
rect 19292 7476 19348 8316
rect 19740 8306 19796 8316
rect 20076 8036 20132 9100
rect 19516 7980 20132 8036
rect 20188 8930 20244 8942
rect 20188 8878 20190 8930
rect 20242 8878 20244 8930
rect 19292 7474 19460 7476
rect 19292 7422 19294 7474
rect 19346 7422 19460 7474
rect 19292 7420 19460 7422
rect 19292 7410 19348 7420
rect 19292 6804 19348 6814
rect 19068 6802 19348 6804
rect 19068 6750 19294 6802
rect 19346 6750 19348 6802
rect 19068 6748 19348 6750
rect 19292 6738 19348 6748
rect 19404 6692 19460 7420
rect 19404 6626 19460 6636
rect 18396 6078 18398 6130
rect 18450 6078 18452 6130
rect 18396 5908 18452 6078
rect 19516 6020 19572 7980
rect 19836 7868 20100 7878
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 19836 7802 20100 7812
rect 20188 7700 20244 8878
rect 20300 8932 20356 11340
rect 20412 11394 20468 11900
rect 20412 11342 20414 11394
rect 20466 11342 20468 11394
rect 20412 11330 20468 11342
rect 20636 11284 20692 11294
rect 20636 11190 20692 11228
rect 20972 10164 21028 10174
rect 21196 10164 21252 12908
rect 21308 12898 21364 12908
rect 21308 12404 21364 12414
rect 21308 11170 21364 12348
rect 21420 11284 21476 11294
rect 21420 11190 21476 11228
rect 21308 11118 21310 11170
rect 21362 11118 21364 11170
rect 21308 11060 21364 11118
rect 21532 11170 21588 11182
rect 21532 11118 21534 11170
rect 21586 11118 21588 11170
rect 21308 11004 21476 11060
rect 21028 10108 21364 10164
rect 20972 10098 21028 10108
rect 21308 9826 21364 10108
rect 21308 9774 21310 9826
rect 21362 9774 21364 9826
rect 21308 9762 21364 9774
rect 20412 9268 20468 9278
rect 21196 9268 21252 9278
rect 20412 9154 20468 9212
rect 20412 9102 20414 9154
rect 20466 9102 20468 9154
rect 20412 9090 20468 9102
rect 20636 9266 21252 9268
rect 20636 9214 21198 9266
rect 21250 9214 21252 9266
rect 20636 9212 21252 9214
rect 20636 9154 20692 9212
rect 21196 9202 21252 9212
rect 20636 9102 20638 9154
rect 20690 9102 20692 9154
rect 20636 9090 20692 9102
rect 21308 9156 21364 9166
rect 21308 9062 21364 9100
rect 21084 9044 21140 9054
rect 21084 9042 21252 9044
rect 21084 8990 21086 9042
rect 21138 8990 21252 9042
rect 21084 8988 21252 8990
rect 21084 8978 21140 8988
rect 20300 8876 20468 8932
rect 19964 7644 20244 7700
rect 20300 8596 20356 8606
rect 19964 7586 20020 7644
rect 19964 7534 19966 7586
rect 20018 7534 20020 7586
rect 19964 7522 20020 7534
rect 19740 6692 19796 6702
rect 20300 6692 20356 8540
rect 19740 6598 19796 6636
rect 20188 6690 20356 6692
rect 20188 6638 20302 6690
rect 20354 6638 20356 6690
rect 20188 6636 20356 6638
rect 19836 6300 20100 6310
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 19836 6234 20100 6244
rect 20188 6132 20244 6636
rect 20300 6626 20356 6636
rect 18956 5964 19236 6020
rect 18396 5842 18452 5852
rect 18620 5906 18676 5918
rect 18620 5854 18622 5906
rect 18674 5854 18676 5906
rect 18620 5460 18676 5854
rect 18844 5908 18900 5918
rect 18844 5814 18900 5852
rect 18620 5394 18676 5404
rect 18956 5348 19012 5964
rect 18732 5292 19012 5348
rect 19068 5794 19124 5806
rect 19068 5742 19070 5794
rect 19122 5742 19124 5794
rect 18620 5236 18676 5246
rect 18732 5236 18788 5292
rect 18620 5234 18788 5236
rect 18620 5182 18622 5234
rect 18674 5182 18788 5234
rect 18620 5180 18788 5182
rect 18620 5170 18676 5180
rect 16492 5058 16548 5068
rect 17948 5124 18004 5134
rect 17948 4340 18004 5068
rect 19068 4450 19124 5742
rect 19180 5684 19236 5964
rect 19292 6018 19572 6020
rect 19292 5966 19518 6018
rect 19570 5966 19572 6018
rect 19292 5964 19572 5966
rect 19292 5906 19348 5964
rect 19516 5954 19572 5964
rect 19852 6076 20244 6132
rect 19852 6018 19908 6076
rect 19852 5966 19854 6018
rect 19906 5966 19908 6018
rect 19852 5954 19908 5966
rect 19292 5854 19294 5906
rect 19346 5854 19348 5906
rect 19292 5842 19348 5854
rect 19964 5908 20020 5918
rect 19964 5814 20020 5852
rect 20412 5906 20468 8876
rect 21196 8820 21252 8988
rect 21420 8820 21476 11004
rect 21532 10276 21588 11118
rect 21532 10210 21588 10220
rect 21196 8764 21476 8820
rect 21644 9042 21700 15092
rect 21756 12066 21812 12078
rect 21756 12014 21758 12066
rect 21810 12014 21812 12066
rect 21756 11844 21812 12014
rect 21756 11778 21812 11788
rect 21868 11396 21924 11406
rect 21868 11302 21924 11340
rect 21980 9604 22036 16604
rect 22204 16100 22260 16110
rect 22204 16006 22260 16044
rect 22204 15428 22260 15438
rect 22316 15428 22372 16828
rect 22540 17444 22596 17454
rect 22540 15986 22596 17388
rect 22540 15934 22542 15986
rect 22594 15934 22596 15986
rect 22540 15922 22596 15934
rect 22764 16882 22820 17612
rect 22764 16830 22766 16882
rect 22818 16830 22820 16882
rect 22204 15426 22372 15428
rect 22204 15374 22206 15426
rect 22258 15374 22372 15426
rect 22204 15372 22372 15374
rect 22204 15362 22260 15372
rect 22764 15314 22820 16830
rect 22988 16772 23044 18398
rect 23212 18452 23268 18462
rect 23212 18358 23268 18396
rect 23436 18450 23492 18462
rect 23436 18398 23438 18450
rect 23490 18398 23492 18450
rect 23436 18116 23492 18398
rect 23548 18340 23604 19966
rect 23548 18274 23604 18284
rect 23660 19346 23716 19358
rect 23660 19294 23662 19346
rect 23714 19294 23716 19346
rect 23660 18676 23716 19294
rect 23436 18060 23604 18116
rect 23548 17892 23604 18060
rect 23548 17826 23604 17836
rect 22988 16706 23044 16716
rect 23100 17108 23156 17118
rect 23100 16210 23156 17052
rect 23660 17108 23716 18620
rect 23660 17042 23716 17052
rect 23772 16884 23828 20972
rect 23996 20802 24052 21420
rect 24444 20916 24500 22204
rect 24668 21588 24724 21598
rect 24668 21494 24724 21532
rect 23996 20750 23998 20802
rect 24050 20750 24052 20802
rect 23996 20738 24052 20750
rect 24220 20860 24500 20916
rect 24892 20916 24948 20926
rect 23884 20692 23940 20702
rect 23884 20598 23940 20636
rect 23884 20132 23940 20142
rect 23884 20130 24164 20132
rect 23884 20078 23886 20130
rect 23938 20078 24164 20130
rect 23884 20076 24164 20078
rect 23884 20066 23940 20076
rect 24108 18674 24164 20076
rect 24220 19572 24276 20860
rect 24332 20692 24388 20702
rect 24332 20598 24388 20636
rect 24444 20692 24500 20702
rect 24444 20690 24724 20692
rect 24444 20638 24446 20690
rect 24498 20638 24724 20690
rect 24444 20636 24724 20638
rect 24444 20626 24500 20636
rect 24668 20244 24724 20636
rect 24892 20690 24948 20860
rect 25116 20804 25172 20814
rect 25228 20804 25284 22876
rect 25452 22708 25508 23660
rect 25452 22642 25508 22652
rect 25788 22482 25844 24670
rect 26124 24724 26180 24734
rect 26124 24630 26180 24668
rect 26236 24610 26292 25564
rect 26908 25508 26964 25518
rect 26796 25506 26964 25508
rect 26796 25454 26910 25506
rect 26962 25454 26964 25506
rect 26796 25452 26964 25454
rect 26796 25172 26852 25452
rect 26908 25442 26964 25452
rect 27020 25396 27076 25788
rect 27132 25620 27188 25630
rect 27244 25620 27300 26852
rect 27468 26514 27524 28028
rect 27580 27076 27636 29372
rect 27692 28084 27748 32508
rect 27916 31780 27972 33182
rect 28140 33234 28196 33246
rect 28140 33182 28142 33234
rect 28194 33182 28196 33234
rect 28140 32004 28196 33182
rect 28252 32228 28308 33294
rect 28364 33236 28420 34078
rect 28364 33170 28420 33180
rect 28476 34018 28532 34030
rect 28476 33966 28478 34018
rect 28530 33966 28532 34018
rect 28476 33348 28532 33966
rect 28364 32564 28420 32574
rect 28364 32470 28420 32508
rect 28252 32172 28420 32228
rect 28140 31948 28308 32004
rect 27916 31714 27972 31724
rect 28252 31778 28308 31948
rect 28252 31726 28254 31778
rect 28306 31726 28308 31778
rect 28028 31668 28084 31678
rect 28028 30772 28084 31612
rect 28028 30706 28084 30716
rect 27916 30660 27972 30670
rect 27916 29204 27972 30604
rect 28252 30324 28308 31726
rect 28364 31668 28420 32172
rect 28476 32002 28532 33292
rect 28476 31950 28478 32002
rect 28530 31950 28532 32002
rect 28476 31938 28532 31950
rect 28364 31602 28420 31612
rect 28588 31108 28644 34860
rect 28700 34692 28756 34702
rect 28700 34598 28756 34636
rect 28812 34018 28868 35756
rect 28812 33966 28814 34018
rect 28866 33966 28868 34018
rect 28812 33954 28868 33966
rect 28924 35698 28980 35710
rect 28924 35646 28926 35698
rect 28978 35646 28980 35698
rect 28700 33572 28756 33582
rect 28924 33572 28980 35646
rect 29372 35700 29428 35710
rect 29372 35138 29428 35644
rect 29372 35086 29374 35138
rect 29426 35086 29428 35138
rect 29372 35074 29428 35086
rect 29484 35698 29540 36204
rect 29596 36482 29652 36494
rect 29596 36430 29598 36482
rect 29650 36430 29652 36482
rect 29596 35812 29652 36430
rect 29596 35718 29652 35756
rect 29484 35646 29486 35698
rect 29538 35646 29540 35698
rect 29148 35028 29204 35038
rect 29148 34934 29204 34972
rect 29484 34804 29540 35646
rect 29708 35586 29764 38780
rect 30604 38668 30660 43820
rect 30828 43764 30884 44268
rect 30828 43698 30884 43708
rect 31052 44100 31108 44110
rect 31052 43650 31108 44044
rect 31052 43598 31054 43650
rect 31106 43598 31108 43650
rect 31052 43586 31108 43598
rect 30716 43426 30772 43438
rect 30716 43374 30718 43426
rect 30770 43374 30772 43426
rect 30716 42756 30772 43374
rect 31388 42980 31444 51100
rect 31500 50820 31556 51326
rect 31612 50820 31668 50830
rect 31500 50818 31668 50820
rect 31500 50766 31614 50818
rect 31666 50766 31668 50818
rect 31500 50764 31668 50766
rect 31612 50754 31668 50764
rect 31948 50428 32004 53452
rect 32060 53442 32116 53452
rect 32956 53508 33012 53518
rect 32284 52164 32340 52174
rect 32732 52164 32788 52174
rect 32284 52162 32788 52164
rect 32284 52110 32286 52162
rect 32338 52110 32734 52162
rect 32786 52110 32788 52162
rect 32284 52108 32788 52110
rect 32284 50428 32340 52108
rect 32732 52098 32788 52108
rect 32956 52162 33012 53452
rect 33068 53060 33124 54350
rect 33068 52994 33124 53004
rect 33292 54404 33348 54414
rect 33292 53506 33348 54348
rect 33292 53454 33294 53506
rect 33346 53454 33348 53506
rect 32956 52110 32958 52162
rect 33010 52110 33012 52162
rect 32956 52098 33012 52110
rect 32508 51380 32564 51390
rect 32508 51286 32564 51324
rect 33180 51266 33236 51278
rect 33180 51214 33182 51266
rect 33234 51214 33236 51266
rect 32732 51044 32788 51054
rect 32620 50932 32676 50942
rect 31948 50372 32116 50428
rect 32060 49924 32116 50372
rect 32172 50372 32340 50428
rect 32508 50596 32564 50606
rect 32172 50260 32228 50372
rect 32172 50204 32452 50260
rect 32396 50034 32452 50204
rect 32396 49982 32398 50034
rect 32450 49982 32452 50034
rect 32396 49970 32452 49982
rect 32172 49924 32228 49934
rect 32060 49922 32228 49924
rect 32060 49870 32174 49922
rect 32226 49870 32228 49922
rect 32060 49868 32228 49870
rect 32172 49858 32228 49868
rect 32508 49698 32564 50540
rect 32620 50594 32676 50876
rect 32620 50542 32622 50594
rect 32674 50542 32676 50594
rect 32620 50530 32676 50542
rect 32732 50482 32788 50988
rect 33180 50932 33236 51214
rect 33180 50866 33236 50876
rect 32732 50430 32734 50482
rect 32786 50430 32788 50482
rect 32732 50418 32788 50430
rect 33292 50428 33348 53454
rect 33404 53508 33460 59200
rect 34300 55972 34356 55982
rect 34300 55970 34804 55972
rect 34300 55918 34302 55970
rect 34354 55918 34804 55970
rect 34300 55916 34804 55918
rect 34300 55906 34356 55916
rect 33628 55524 33684 55534
rect 33404 53442 33460 53452
rect 33516 53844 33572 53854
rect 33516 53284 33572 53788
rect 33628 53730 33684 55468
rect 34188 55412 34244 55422
rect 34188 55318 34244 55356
rect 33628 53678 33630 53730
rect 33682 53678 33684 53730
rect 33628 53666 33684 53678
rect 33740 53956 33796 53966
rect 33180 50372 33348 50428
rect 33404 53228 33572 53284
rect 33180 49812 33236 50372
rect 33180 49810 33348 49812
rect 33180 49758 33182 49810
rect 33234 49758 33348 49810
rect 33180 49756 33348 49758
rect 33180 49746 33236 49756
rect 32508 49646 32510 49698
rect 32562 49646 32564 49698
rect 32508 49634 32564 49646
rect 32844 49140 32900 49150
rect 32844 49046 32900 49084
rect 31500 49028 31556 49038
rect 31500 48934 31556 48972
rect 31500 47460 31556 47470
rect 31500 47366 31556 47404
rect 32172 47460 32228 47470
rect 32172 47366 32228 47404
rect 32732 47404 33124 47460
rect 32732 47234 32788 47404
rect 32732 47182 32734 47234
rect 32786 47182 32788 47234
rect 32732 47124 32788 47182
rect 32060 47068 32788 47124
rect 32844 47234 32900 47246
rect 32844 47182 32846 47234
rect 32898 47182 32900 47234
rect 31948 46788 32004 46798
rect 32060 46788 32116 47068
rect 32844 47012 32900 47182
rect 31948 46786 32116 46788
rect 31948 46734 31950 46786
rect 32002 46734 32116 46786
rect 31948 46732 32116 46734
rect 32508 46956 32900 47012
rect 32956 47234 33012 47246
rect 32956 47182 32958 47234
rect 33010 47182 33012 47234
rect 32508 46786 32564 46956
rect 32508 46734 32510 46786
rect 32562 46734 32564 46786
rect 31948 46722 32004 46732
rect 32508 46722 32564 46734
rect 32284 46674 32340 46686
rect 32284 46622 32286 46674
rect 32338 46622 32340 46674
rect 32060 46562 32116 46574
rect 32060 46510 32062 46562
rect 32114 46510 32116 46562
rect 32060 46228 32116 46510
rect 32284 46564 32340 46622
rect 32956 46564 33012 47182
rect 33068 46900 33124 47404
rect 33292 46900 33348 49756
rect 33404 48804 33460 53228
rect 33628 52052 33684 52062
rect 33628 51958 33684 51996
rect 33516 50596 33572 50606
rect 33740 50596 33796 53900
rect 34636 53508 34692 53518
rect 34636 53414 34692 53452
rect 34300 53060 34356 53070
rect 34300 52966 34356 53004
rect 33852 52836 33908 52846
rect 33852 52834 34020 52836
rect 33852 52782 33854 52834
rect 33906 52782 34020 52834
rect 33852 52780 34020 52782
rect 33852 52770 33908 52780
rect 33964 51378 34020 52780
rect 33964 51326 33966 51378
rect 34018 51326 34020 51378
rect 33964 50708 34020 51326
rect 34300 52724 34356 52734
rect 34300 52164 34356 52668
rect 34748 52276 34804 55916
rect 34972 54628 35028 59200
rect 36540 56308 36596 59200
rect 38108 57092 38164 59200
rect 39676 57428 39732 59200
rect 39676 57372 39956 57428
rect 38108 57026 38164 57036
rect 36540 56242 36596 56252
rect 35084 56084 35140 56094
rect 35084 55990 35140 56028
rect 35868 56084 35924 56094
rect 35196 55692 35460 55702
rect 35252 55636 35300 55692
rect 35356 55636 35404 55692
rect 35196 55626 35460 55636
rect 34972 54562 35028 54572
rect 35868 54516 35924 56028
rect 38780 56084 38836 56094
rect 39788 56084 39844 56094
rect 38780 55990 38836 56028
rect 39004 56082 39844 56084
rect 39004 56030 39790 56082
rect 39842 56030 39844 56082
rect 39004 56028 39844 56030
rect 35980 55970 36036 55982
rect 35980 55918 35982 55970
rect 36034 55918 36036 55970
rect 35980 55524 36036 55918
rect 38108 55972 38164 55982
rect 38108 55878 38164 55916
rect 37548 55524 37604 55534
rect 35980 55458 36036 55468
rect 37436 55468 37548 55524
rect 36876 55300 36932 55310
rect 37212 55300 37268 55310
rect 36316 55298 36932 55300
rect 36316 55246 36878 55298
rect 36930 55246 36932 55298
rect 36316 55244 36932 55246
rect 36204 55188 36260 55198
rect 35868 54422 35924 54460
rect 36092 55186 36260 55188
rect 36092 55134 36206 55186
rect 36258 55134 36260 55186
rect 36092 55132 36260 55134
rect 35196 54404 35252 54414
rect 35084 54402 35252 54404
rect 35084 54350 35198 54402
rect 35250 54350 35252 54402
rect 35084 54348 35252 54350
rect 35084 53172 35140 54348
rect 35196 54338 35252 54348
rect 35196 54124 35460 54134
rect 35252 54068 35300 54124
rect 35356 54068 35404 54124
rect 35196 54058 35460 54068
rect 35084 53106 35140 53116
rect 34972 52948 35028 52958
rect 34748 52182 34804 52220
rect 34860 52892 34972 52948
rect 34300 51266 34356 52108
rect 34860 52052 34916 52892
rect 34972 52882 35028 52892
rect 35196 52946 35252 52958
rect 35196 52894 35198 52946
rect 35250 52894 35252 52946
rect 35084 52836 35140 52846
rect 35084 52162 35140 52780
rect 35196 52724 35252 52894
rect 35868 52836 35924 52846
rect 35868 52742 35924 52780
rect 35196 52658 35252 52668
rect 35196 52556 35460 52566
rect 35252 52500 35300 52556
rect 35356 52500 35404 52556
rect 35196 52490 35460 52500
rect 35532 52276 35588 52286
rect 36092 52276 36148 55132
rect 36204 55122 36260 55132
rect 36316 55186 36372 55244
rect 36876 55234 36932 55244
rect 36988 55298 37268 55300
rect 36988 55246 37214 55298
rect 37266 55246 37268 55298
rect 36988 55244 37268 55246
rect 36316 55134 36318 55186
rect 36370 55134 36372 55186
rect 36316 55122 36372 55134
rect 36540 55074 36596 55086
rect 36540 55022 36542 55074
rect 36594 55022 36596 55074
rect 36540 54404 36596 55022
rect 36540 54338 36596 54348
rect 36988 53508 37044 55244
rect 37212 55234 37268 55244
rect 37100 55074 37156 55086
rect 37100 55022 37102 55074
rect 37154 55022 37156 55074
rect 37100 54852 37156 55022
rect 37100 54796 37268 54852
rect 37100 54628 37156 54638
rect 37100 54534 37156 54572
rect 37212 53730 37268 54796
rect 37436 54740 37492 55468
rect 37548 55458 37604 55468
rect 37996 55524 38052 55534
rect 37996 55298 38052 55468
rect 38556 55524 38612 55534
rect 37996 55246 37998 55298
rect 38050 55246 38052 55298
rect 37996 55234 38052 55246
rect 38444 55298 38500 55310
rect 38444 55246 38446 55298
rect 38498 55246 38500 55298
rect 37548 55188 37604 55198
rect 37548 55186 37828 55188
rect 37548 55134 37550 55186
rect 37602 55134 37828 55186
rect 37548 55132 37828 55134
rect 37548 55122 37604 55132
rect 37436 54684 37716 54740
rect 37436 53844 37492 53854
rect 37212 53678 37214 53730
rect 37266 53678 37268 53730
rect 37100 53508 37156 53518
rect 36764 53452 37100 53508
rect 36204 52948 36260 52958
rect 36204 52854 36260 52892
rect 36764 52946 36820 53452
rect 37100 53414 37156 53452
rect 37212 53060 37268 53678
rect 37324 53788 37436 53844
rect 37324 53730 37380 53788
rect 37436 53778 37492 53788
rect 37324 53678 37326 53730
rect 37378 53678 37380 53730
rect 37324 53666 37380 53678
rect 37660 53730 37716 54684
rect 37660 53678 37662 53730
rect 37714 53678 37716 53730
rect 37660 53666 37716 53678
rect 37772 54628 37828 55132
rect 38444 54740 38500 55246
rect 38444 54674 38500 54684
rect 37436 53618 37492 53630
rect 37436 53566 37438 53618
rect 37490 53566 37492 53618
rect 37436 53508 37492 53566
rect 37324 53452 37492 53508
rect 37324 53284 37380 53452
rect 37772 53396 37828 54572
rect 37324 53218 37380 53228
rect 37436 53340 37828 53396
rect 37884 54516 37940 54526
rect 37436 53170 37492 53340
rect 37436 53118 37438 53170
rect 37490 53118 37492 53170
rect 37436 53106 37492 53118
rect 37884 53060 37940 54460
rect 38332 54404 38388 54414
rect 37212 52994 37268 53004
rect 37772 53004 37940 53060
rect 37996 53844 38052 53854
rect 36988 52948 37044 52958
rect 36764 52894 36766 52946
rect 36818 52894 36820 52946
rect 36764 52882 36820 52894
rect 36876 52946 37044 52948
rect 36876 52894 36990 52946
rect 37042 52894 37044 52946
rect 36876 52892 37044 52894
rect 36876 52388 36932 52892
rect 36988 52882 37044 52892
rect 37324 52948 37380 52958
rect 36428 52332 36932 52388
rect 36204 52276 36260 52286
rect 36092 52220 36204 52276
rect 35532 52182 35588 52220
rect 36204 52210 36260 52220
rect 36428 52274 36484 52332
rect 36428 52222 36430 52274
rect 36482 52222 36484 52274
rect 36428 52210 36484 52222
rect 35084 52110 35086 52162
rect 35138 52110 35140 52162
rect 35084 52098 35140 52110
rect 35644 52164 35700 52174
rect 35980 52164 36036 52174
rect 35644 52162 35924 52164
rect 35644 52110 35646 52162
rect 35698 52110 35924 52162
rect 35644 52108 35924 52110
rect 35644 52098 35700 52108
rect 34636 51996 34916 52052
rect 34636 51490 34692 51996
rect 35420 51940 35476 51950
rect 35420 51846 35476 51884
rect 35532 51604 35588 51614
rect 35532 51510 35588 51548
rect 34636 51438 34638 51490
rect 34690 51438 34692 51490
rect 34636 51426 34692 51438
rect 34300 51214 34302 51266
rect 34354 51214 34356 51266
rect 34300 51202 34356 51214
rect 35868 51154 35924 52108
rect 35980 51602 36036 52108
rect 35980 51550 35982 51602
rect 36034 51550 36036 51602
rect 35980 51538 36036 51550
rect 36092 51940 36148 51950
rect 36092 51602 36148 51884
rect 36092 51550 36094 51602
rect 36146 51550 36148 51602
rect 35868 51102 35870 51154
rect 35922 51102 35924 51154
rect 35196 50988 35460 50998
rect 35252 50932 35300 50988
rect 35356 50932 35404 50988
rect 35196 50922 35460 50932
rect 33964 50642 34020 50652
rect 35756 50708 35812 50718
rect 33852 50596 33908 50606
rect 33740 50540 33852 50596
rect 33516 50502 33572 50540
rect 33852 50530 33908 50540
rect 34076 50596 34132 50606
rect 34636 50596 34692 50606
rect 35084 50596 35140 50606
rect 34076 50594 34356 50596
rect 34076 50542 34078 50594
rect 34130 50542 34356 50594
rect 34076 50540 34356 50542
rect 34076 50530 34132 50540
rect 33516 50370 33572 50382
rect 34188 50372 34244 50382
rect 33516 50318 33518 50370
rect 33570 50318 33572 50370
rect 33516 49924 33572 50318
rect 33516 49858 33572 49868
rect 33852 50370 34244 50372
rect 33852 50318 34190 50370
rect 34242 50318 34244 50370
rect 33852 50316 34244 50318
rect 33852 49922 33908 50316
rect 34188 50306 34244 50316
rect 34300 50260 34356 50540
rect 34636 50594 35140 50596
rect 34636 50542 34638 50594
rect 34690 50542 35086 50594
rect 35138 50542 35140 50594
rect 34636 50540 35140 50542
rect 34636 50530 34692 50540
rect 35084 50530 35140 50540
rect 35644 50596 35700 50606
rect 35756 50596 35812 50652
rect 35644 50594 35812 50596
rect 35644 50542 35646 50594
rect 35698 50542 35812 50594
rect 35644 50540 35812 50542
rect 35644 50530 35700 50540
rect 34412 50484 34468 50522
rect 35196 50482 35252 50494
rect 35196 50430 35198 50482
rect 35250 50430 35252 50482
rect 35196 50428 35252 50430
rect 34412 50418 34468 50428
rect 34972 50370 35028 50382
rect 34972 50318 34974 50370
rect 35026 50318 35028 50370
rect 34300 50194 34356 50204
rect 34636 50260 34692 50270
rect 33852 49870 33854 49922
rect 33906 49870 33908 49922
rect 33852 49858 33908 49870
rect 33740 49140 33796 49150
rect 33740 49046 33796 49084
rect 34636 49138 34692 50204
rect 34972 50260 35028 50318
rect 34972 50194 35028 50204
rect 35084 50372 35252 50428
rect 34636 49086 34638 49138
rect 34690 49086 34692 49138
rect 34636 49074 34692 49086
rect 34188 49028 34244 49038
rect 35084 49028 35140 50316
rect 35532 49812 35588 49822
rect 35196 49420 35460 49430
rect 35252 49364 35300 49420
rect 35356 49364 35404 49420
rect 35196 49354 35460 49364
rect 35420 49252 35476 49262
rect 35196 49028 35252 49038
rect 35084 49026 35252 49028
rect 35084 48974 35198 49026
rect 35250 48974 35252 49026
rect 35084 48972 35252 48974
rect 34188 48934 34244 48972
rect 35196 48962 35252 48972
rect 35420 48914 35476 49196
rect 35420 48862 35422 48914
rect 35474 48862 35476 48914
rect 35420 48850 35476 48862
rect 35532 48914 35588 49756
rect 35532 48862 35534 48914
rect 35586 48862 35588 48914
rect 33404 48738 33460 48748
rect 35532 48692 35588 48862
rect 35084 48636 35588 48692
rect 35084 47570 35140 48636
rect 35532 48242 35588 48254
rect 35532 48190 35534 48242
rect 35586 48190 35588 48242
rect 35196 47852 35460 47862
rect 35252 47796 35300 47852
rect 35356 47796 35404 47852
rect 35196 47786 35460 47796
rect 35084 47518 35086 47570
rect 35138 47518 35140 47570
rect 35084 47506 35140 47518
rect 33404 47458 33460 47470
rect 33404 47406 33406 47458
rect 33458 47406 33460 47458
rect 33404 47236 33460 47406
rect 34972 47460 35028 47470
rect 34972 47366 35028 47404
rect 35420 47458 35476 47470
rect 35420 47406 35422 47458
rect 35474 47406 35476 47458
rect 33740 47348 33796 47358
rect 33740 47236 33796 47292
rect 34524 47348 34580 47358
rect 34524 47346 34692 47348
rect 34524 47294 34526 47346
rect 34578 47294 34692 47346
rect 34524 47292 34692 47294
rect 34524 47282 34580 47292
rect 33404 47234 33796 47236
rect 33404 47182 33742 47234
rect 33794 47182 33796 47234
rect 33404 47180 33796 47182
rect 33068 46844 33236 46900
rect 33180 46676 33236 46844
rect 33292 46834 33348 46844
rect 33292 46676 33348 46686
rect 33180 46674 33348 46676
rect 33180 46622 33294 46674
rect 33346 46622 33348 46674
rect 33180 46620 33348 46622
rect 33292 46610 33348 46620
rect 32284 46508 33012 46564
rect 31612 46172 32116 46228
rect 31612 46002 31668 46172
rect 31612 45950 31614 46002
rect 31666 45950 31668 46002
rect 31612 45938 31668 45950
rect 32396 45220 32452 45230
rect 31948 45108 32004 45118
rect 31948 45014 32004 45052
rect 31500 44436 31556 44446
rect 31500 44342 31556 44380
rect 32396 44434 32452 45164
rect 32396 44382 32398 44434
rect 32450 44382 32452 44434
rect 32396 44370 32452 44382
rect 32956 44324 33012 46508
rect 33404 45220 33460 45230
rect 33404 45126 33460 45164
rect 33516 45218 33572 45230
rect 33516 45166 33518 45218
rect 33570 45166 33572 45218
rect 32956 44258 33012 44268
rect 31836 44100 31892 44110
rect 31836 44006 31892 44044
rect 33068 43428 33124 43438
rect 33516 43428 33572 45166
rect 33628 45108 33684 47180
rect 33740 47170 33796 47180
rect 34412 47234 34468 47246
rect 34412 47182 34414 47234
rect 34466 47182 34468 47234
rect 33740 46674 33796 46686
rect 33740 46622 33742 46674
rect 33794 46622 33796 46674
rect 33740 46002 33796 46622
rect 34188 46676 34244 46686
rect 34412 46676 34468 47182
rect 34636 47124 34692 47292
rect 35196 47234 35252 47246
rect 35196 47182 35198 47234
rect 35250 47182 35252 47234
rect 35196 47124 35252 47182
rect 34636 47068 35140 47124
rect 34188 46674 34412 46676
rect 34188 46622 34190 46674
rect 34242 46622 34412 46674
rect 34188 46620 34412 46622
rect 34188 46610 34244 46620
rect 34412 46610 34468 46620
rect 34524 47012 34580 47022
rect 33740 45950 33742 46002
rect 33794 45950 33796 46002
rect 33740 45780 33796 45950
rect 33740 45724 34244 45780
rect 33740 45332 33796 45342
rect 33740 45238 33796 45276
rect 33964 45332 34020 45342
rect 33628 45052 33796 45108
rect 33068 43426 33572 43428
rect 33068 43374 33070 43426
rect 33122 43374 33572 43426
rect 33068 43372 33572 43374
rect 33068 43316 33124 43372
rect 33068 43250 33124 43260
rect 31388 42924 31556 42980
rect 31388 42756 31444 42766
rect 30716 42754 31444 42756
rect 30716 42702 31390 42754
rect 31442 42702 31444 42754
rect 30716 42700 31444 42702
rect 30716 41860 30772 42700
rect 31388 42690 31444 42700
rect 30716 41794 30772 41804
rect 31500 41412 31556 42924
rect 32060 42756 32116 42766
rect 32060 42662 32116 42700
rect 32956 42754 33012 42766
rect 32956 42702 32958 42754
rect 33010 42702 33012 42754
rect 32956 42532 33012 42702
rect 33068 42756 33124 42766
rect 33292 42756 33348 42766
rect 33068 42662 33124 42700
rect 33180 42700 33292 42756
rect 33012 42476 33124 42532
rect 32956 42466 33012 42476
rect 31500 41346 31556 41356
rect 31836 42196 31892 42206
rect 31724 40740 31780 40750
rect 30940 40068 30996 40078
rect 30716 39618 30772 39630
rect 30716 39566 30718 39618
rect 30770 39566 30772 39618
rect 30716 39508 30772 39566
rect 30716 39442 30772 39452
rect 30940 38834 30996 40012
rect 31724 39732 31780 40684
rect 31836 40628 31892 42140
rect 33068 41972 33124 42476
rect 33180 42194 33236 42700
rect 33292 42662 33348 42700
rect 33628 42754 33684 42766
rect 33628 42702 33630 42754
rect 33682 42702 33684 42754
rect 33180 42142 33182 42194
rect 33234 42142 33236 42194
rect 33180 42130 33236 42142
rect 33404 42642 33460 42654
rect 33404 42590 33406 42642
rect 33458 42590 33460 42642
rect 33292 42082 33348 42094
rect 33292 42030 33294 42082
rect 33346 42030 33348 42082
rect 33068 41916 33236 41972
rect 33068 41748 33124 41758
rect 32508 41300 32564 41310
rect 32508 41206 32564 41244
rect 32844 41188 32900 41198
rect 32844 41094 32900 41132
rect 33068 41076 33124 41692
rect 33180 41298 33236 41916
rect 33180 41246 33182 41298
rect 33234 41246 33236 41298
rect 33180 41234 33236 41246
rect 33292 41188 33348 42030
rect 33404 41972 33460 42590
rect 33628 42644 33684 42702
rect 33628 42578 33684 42588
rect 33404 41906 33460 41916
rect 33404 41188 33460 41198
rect 33292 41132 33404 41188
rect 33404 41122 33460 41132
rect 33516 41186 33572 41198
rect 33516 41134 33518 41186
rect 33570 41134 33572 41186
rect 33068 40982 33124 41020
rect 33292 40962 33348 40974
rect 33292 40910 33294 40962
rect 33346 40910 33348 40962
rect 33180 40740 33236 40750
rect 33292 40740 33348 40910
rect 33292 40684 33460 40740
rect 32172 40628 32228 40638
rect 31836 40572 32004 40628
rect 31500 39730 31780 39732
rect 31500 39678 31726 39730
rect 31778 39678 31780 39730
rect 31500 39676 31780 39678
rect 30940 38782 30942 38834
rect 30994 38782 30996 38834
rect 30940 38668 30996 38782
rect 30604 38612 30772 38668
rect 30156 38050 30212 38062
rect 30156 37998 30158 38050
rect 30210 37998 30212 38050
rect 30156 37940 30212 37998
rect 30604 37940 30660 37950
rect 30156 37938 30660 37940
rect 30156 37886 30606 37938
rect 30658 37886 30660 37938
rect 30156 37884 30660 37886
rect 30044 37268 30100 37278
rect 30044 37174 30100 37212
rect 30156 36706 30212 37884
rect 30604 37874 30660 37884
rect 30716 37380 30772 38612
rect 30156 36654 30158 36706
rect 30210 36654 30212 36706
rect 30156 36642 30212 36654
rect 30492 37324 30772 37380
rect 30828 38612 30996 38668
rect 31276 39508 31332 39518
rect 31276 39060 31332 39452
rect 31164 38612 31220 38622
rect 29708 35534 29710 35586
rect 29762 35534 29764 35586
rect 29708 35522 29764 35534
rect 30380 36484 30436 36494
rect 29708 34916 29764 34926
rect 29708 34822 29764 34860
rect 30380 34914 30436 36428
rect 30380 34862 30382 34914
rect 30434 34862 30436 34914
rect 30380 34850 30436 34862
rect 29484 34738 29540 34748
rect 29372 34356 29428 34366
rect 29372 34354 30100 34356
rect 29372 34302 29374 34354
rect 29426 34302 30100 34354
rect 29372 34300 30100 34302
rect 29372 34290 29428 34300
rect 30044 34242 30100 34300
rect 30044 34190 30046 34242
rect 30098 34190 30100 34242
rect 28700 33570 28980 33572
rect 28700 33518 28702 33570
rect 28754 33518 28980 33570
rect 28700 33516 28980 33518
rect 29260 34130 29316 34142
rect 29260 34078 29262 34130
rect 29314 34078 29316 34130
rect 29260 33572 29316 34078
rect 29596 34130 29652 34142
rect 29596 34078 29598 34130
rect 29650 34078 29652 34130
rect 29484 33572 29540 33582
rect 29260 33516 29484 33572
rect 28700 33506 28756 33516
rect 29148 33236 29204 33246
rect 29148 33142 29204 33180
rect 29484 33122 29540 33516
rect 29596 33348 29652 34078
rect 29820 33906 29876 33918
rect 29820 33854 29822 33906
rect 29874 33854 29876 33906
rect 29820 33572 29876 33854
rect 29820 33506 29876 33516
rect 29932 33348 29988 33358
rect 29596 33346 29988 33348
rect 29596 33294 29934 33346
rect 29986 33294 29988 33346
rect 29596 33292 29988 33294
rect 29932 33282 29988 33292
rect 29484 33070 29486 33122
rect 29538 33070 29540 33122
rect 29036 32564 29092 32574
rect 29036 31444 29092 32508
rect 29372 32452 29428 32462
rect 29484 32452 29540 33070
rect 30044 32676 30100 34190
rect 30156 33906 30212 33918
rect 30156 33854 30158 33906
rect 30210 33854 30212 33906
rect 30156 33572 30212 33854
rect 30156 33506 30212 33516
rect 30156 32676 30212 32686
rect 30044 32674 30212 32676
rect 30044 32622 30158 32674
rect 30210 32622 30212 32674
rect 30044 32620 30212 32622
rect 29596 32452 29652 32462
rect 29484 32450 29652 32452
rect 29484 32398 29598 32450
rect 29650 32398 29652 32450
rect 29484 32396 29652 32398
rect 29148 31892 29204 31902
rect 29148 31798 29204 31836
rect 29372 31556 29428 32396
rect 29596 32386 29652 32396
rect 30156 31890 30212 32620
rect 30156 31838 30158 31890
rect 30210 31838 30212 31890
rect 30156 31826 30212 31838
rect 29596 31778 29652 31790
rect 29596 31726 29598 31778
rect 29650 31726 29652 31778
rect 29484 31556 29540 31566
rect 29372 31500 29484 31556
rect 29036 31388 29204 31444
rect 28588 31106 28980 31108
rect 28588 31054 28590 31106
rect 28642 31054 28980 31106
rect 28588 31052 28980 31054
rect 28588 31042 28644 31052
rect 28252 30258 28308 30268
rect 28588 30212 28644 30222
rect 28588 30118 28644 30156
rect 28476 30100 28532 30110
rect 28476 30006 28532 30044
rect 27916 29138 27972 29148
rect 28588 29652 28644 29662
rect 28588 29426 28644 29596
rect 28588 29374 28590 29426
rect 28642 29374 28644 29426
rect 27804 28644 27860 28654
rect 27804 28550 27860 28588
rect 27692 28018 27748 28028
rect 27916 28532 27972 28542
rect 27804 27972 27860 27982
rect 27804 27858 27860 27916
rect 27804 27806 27806 27858
rect 27858 27806 27860 27858
rect 27804 27794 27860 27806
rect 27916 27860 27972 28476
rect 27916 27748 27972 27804
rect 28364 27860 28420 27870
rect 27916 27746 28196 27748
rect 27916 27694 27918 27746
rect 27970 27694 28196 27746
rect 27916 27692 28196 27694
rect 27916 27682 27972 27692
rect 27580 27020 27972 27076
rect 27916 26962 27972 27020
rect 28140 27074 28196 27692
rect 28140 27022 28142 27074
rect 28194 27022 28196 27074
rect 28140 27010 28196 27022
rect 27916 26910 27918 26962
rect 27970 26910 27972 26962
rect 27916 26898 27972 26910
rect 28364 26908 28420 27804
rect 27468 26462 27470 26514
rect 27522 26462 27524 26514
rect 27468 26450 27524 26462
rect 28252 26852 28420 26908
rect 28476 27748 28532 27758
rect 28476 27076 28532 27692
rect 27356 26292 27412 26302
rect 28140 26292 28196 26302
rect 28252 26292 28308 26852
rect 28476 26514 28532 27020
rect 28588 26908 28644 29374
rect 28812 29314 28868 29326
rect 28812 29262 28814 29314
rect 28866 29262 28868 29314
rect 28812 28308 28868 29262
rect 28812 28242 28868 28252
rect 28588 26852 28756 26908
rect 28476 26462 28478 26514
rect 28530 26462 28532 26514
rect 28476 26450 28532 26462
rect 28588 26740 28644 26750
rect 27356 26290 27748 26292
rect 27356 26238 27358 26290
rect 27410 26238 27748 26290
rect 27356 26236 27748 26238
rect 27356 26226 27412 26236
rect 27132 25618 27300 25620
rect 27132 25566 27134 25618
rect 27186 25566 27300 25618
rect 27132 25564 27300 25566
rect 27468 25620 27524 25630
rect 27132 25554 27188 25564
rect 27468 25526 27524 25564
rect 27692 25506 27748 26236
rect 28140 26290 28308 26292
rect 28140 26238 28142 26290
rect 28194 26238 28308 26290
rect 28140 26236 28308 26238
rect 28140 26226 28196 26236
rect 27916 26180 27972 26190
rect 27916 26086 27972 26124
rect 28252 25618 28308 26236
rect 28252 25566 28254 25618
rect 28306 25566 28308 25618
rect 28252 25554 28308 25566
rect 28588 25618 28644 26684
rect 28700 26404 28756 26852
rect 28700 26338 28756 26348
rect 28588 25566 28590 25618
rect 28642 25566 28644 25618
rect 28588 25554 28644 25566
rect 27692 25454 27694 25506
rect 27746 25454 27748 25506
rect 27076 25340 27300 25396
rect 27020 25330 27076 25340
rect 26796 24946 26852 25116
rect 26796 24894 26798 24946
rect 26850 24894 26852 24946
rect 26796 24882 26852 24894
rect 26236 24558 26238 24610
rect 26290 24558 26292 24610
rect 26236 24546 26292 24558
rect 27244 24610 27300 25340
rect 27692 24948 27748 25454
rect 28588 24948 28644 24958
rect 27748 24892 27860 24948
rect 27692 24882 27748 24892
rect 27244 24558 27246 24610
rect 27298 24558 27300 24610
rect 27244 24546 27300 24558
rect 27692 24610 27748 24622
rect 27692 24558 27694 24610
rect 27746 24558 27748 24610
rect 26236 23380 26292 23390
rect 25788 22430 25790 22482
rect 25842 22430 25844 22482
rect 25788 22418 25844 22430
rect 25900 22484 25956 22494
rect 25340 21588 25396 21598
rect 25340 21028 25396 21532
rect 25340 20962 25396 20972
rect 25676 21474 25732 21486
rect 25676 21422 25678 21474
rect 25730 21422 25732 21474
rect 25676 21140 25732 21422
rect 24892 20638 24894 20690
rect 24946 20638 24948 20690
rect 24892 20626 24948 20638
rect 25004 20802 25620 20804
rect 25004 20750 25118 20802
rect 25170 20750 25620 20802
rect 25004 20748 25620 20750
rect 24780 20244 24836 20254
rect 25004 20244 25060 20748
rect 25116 20738 25172 20748
rect 24668 20242 25060 20244
rect 24668 20190 24782 20242
rect 24834 20190 25060 20242
rect 24668 20188 25060 20190
rect 24780 20178 24836 20188
rect 25564 20130 25620 20748
rect 25564 20078 25566 20130
rect 25618 20078 25620 20130
rect 25564 20066 25620 20078
rect 24220 19506 24276 19516
rect 25564 19460 25620 19470
rect 25452 19404 25564 19460
rect 25116 19348 25172 19358
rect 24108 18622 24110 18674
rect 24162 18622 24164 18674
rect 23884 18450 23940 18462
rect 23884 18398 23886 18450
rect 23938 18398 23940 18450
rect 23884 18340 23940 18398
rect 23996 18452 24052 18462
rect 23996 18358 24052 18396
rect 23884 18274 23940 18284
rect 24108 17668 24164 18622
rect 24108 17602 24164 17612
rect 24220 19236 24276 19246
rect 23100 16158 23102 16210
rect 23154 16158 23156 16210
rect 23100 16146 23156 16158
rect 23548 16828 23828 16884
rect 23548 15540 23604 16828
rect 22764 15262 22766 15314
rect 22818 15262 22820 15314
rect 22764 15250 22820 15262
rect 22988 15428 23044 15438
rect 22988 15148 23044 15372
rect 22876 15092 23044 15148
rect 22092 14418 22148 14430
rect 22092 14366 22094 14418
rect 22146 14366 22148 14418
rect 22092 13076 22148 14366
rect 22876 14420 22932 15092
rect 22876 13634 22932 14364
rect 22876 13582 22878 13634
rect 22930 13582 22932 13634
rect 22876 13570 22932 13582
rect 23548 13970 23604 15484
rect 23660 16098 23716 16110
rect 23660 16046 23662 16098
rect 23714 16046 23716 16098
rect 23660 14196 23716 16046
rect 24108 15316 24164 15326
rect 24108 15222 24164 15260
rect 23884 15204 23940 15214
rect 23884 15110 23940 15148
rect 23884 14530 23940 14542
rect 23884 14478 23886 14530
rect 23938 14478 23940 14530
rect 23884 14308 23940 14478
rect 24220 14308 24276 19180
rect 25116 19234 25172 19292
rect 25116 19182 25118 19234
rect 25170 19182 25172 19234
rect 25116 19170 25172 19182
rect 25452 19234 25508 19404
rect 25564 19394 25620 19404
rect 25452 19182 25454 19234
rect 25506 19182 25508 19234
rect 25452 19170 25508 19182
rect 25340 19124 25396 19134
rect 24668 18676 24724 18714
rect 24668 18610 24724 18620
rect 25228 18676 25284 18686
rect 24668 18452 24724 18462
rect 24668 17778 24724 18396
rect 25228 18450 25284 18620
rect 25228 18398 25230 18450
rect 25282 18398 25284 18450
rect 24668 17726 24670 17778
rect 24722 17726 24724 17778
rect 24668 17714 24724 17726
rect 25004 18228 25060 18238
rect 25004 17666 25060 18172
rect 25004 17614 25006 17666
rect 25058 17614 25060 17666
rect 25004 17602 25060 17614
rect 25228 17108 25284 18398
rect 25340 17554 25396 19068
rect 25452 19010 25508 19022
rect 25452 18958 25454 19010
rect 25506 18958 25508 19010
rect 25452 18564 25508 18958
rect 25452 18498 25508 18508
rect 25340 17502 25342 17554
rect 25394 17502 25396 17554
rect 25340 17490 25396 17502
rect 25340 17108 25396 17118
rect 25228 17106 25396 17108
rect 25228 17054 25342 17106
rect 25394 17054 25396 17106
rect 25228 17052 25396 17054
rect 25340 17042 25396 17052
rect 25676 16660 25732 21084
rect 25788 20578 25844 20590
rect 25788 20526 25790 20578
rect 25842 20526 25844 20578
rect 25788 19460 25844 20526
rect 25900 19684 25956 22428
rect 26236 22148 26292 23324
rect 27692 23044 27748 24558
rect 27804 24050 27860 24892
rect 28588 24854 28644 24892
rect 27804 23998 27806 24050
rect 27858 23998 27860 24050
rect 27804 23986 27860 23998
rect 28140 24722 28196 24734
rect 28140 24670 28142 24722
rect 28194 24670 28196 24722
rect 28140 24052 28196 24670
rect 28140 23986 28196 23996
rect 28476 24164 28532 24174
rect 28476 23826 28532 24108
rect 28476 23774 28478 23826
rect 28530 23774 28532 23826
rect 28476 23762 28532 23774
rect 28140 23716 28196 23726
rect 28140 23622 28196 23660
rect 27916 23380 27972 23390
rect 27972 23324 28308 23380
rect 27916 23286 27972 23324
rect 28252 23154 28308 23324
rect 28252 23102 28254 23154
rect 28306 23102 28308 23154
rect 28252 23090 28308 23102
rect 27804 23044 27860 23054
rect 27692 22988 27804 23044
rect 27804 22978 27860 22988
rect 28140 23044 28196 23054
rect 28140 22932 28196 22988
rect 28140 22876 28308 22932
rect 28028 22596 28084 22606
rect 26124 21924 26180 21934
rect 26124 20802 26180 21868
rect 26124 20750 26126 20802
rect 26178 20750 26180 20802
rect 26124 20738 26180 20750
rect 26236 20188 26292 22092
rect 27020 22372 27076 22382
rect 27580 22372 27636 22382
rect 27020 22370 27636 22372
rect 27020 22318 27022 22370
rect 27074 22318 27582 22370
rect 27634 22318 27636 22370
rect 27020 22316 27636 22318
rect 27020 21924 27076 22316
rect 27580 22306 27636 22316
rect 28028 22370 28084 22540
rect 28028 22318 28030 22370
rect 28082 22318 28084 22370
rect 28028 22306 28084 22318
rect 27692 22260 27748 22270
rect 27692 22258 27860 22260
rect 27692 22206 27694 22258
rect 27746 22206 27860 22258
rect 27692 22204 27860 22206
rect 27692 22194 27748 22204
rect 27020 21858 27076 21868
rect 27132 22146 27188 22158
rect 27132 22094 27134 22146
rect 27186 22094 27188 22146
rect 26348 21812 26404 21822
rect 27132 21812 27188 22094
rect 27356 22148 27412 22158
rect 27356 22146 27636 22148
rect 27356 22094 27358 22146
rect 27410 22094 27636 22146
rect 27356 22092 27636 22094
rect 27356 22082 27412 22092
rect 27580 21924 27636 22092
rect 27580 21868 27748 21924
rect 26348 21810 26852 21812
rect 26348 21758 26350 21810
rect 26402 21758 26852 21810
rect 26348 21756 26852 21758
rect 27132 21756 27524 21812
rect 26348 21476 26404 21756
rect 26684 21588 26740 21598
rect 26796 21588 26852 21756
rect 27356 21588 27412 21598
rect 26796 21532 26964 21588
rect 26684 21494 26740 21532
rect 26348 21410 26404 21420
rect 26460 21028 26516 21038
rect 26908 21028 26964 21532
rect 27244 21586 27412 21588
rect 27244 21534 27358 21586
rect 27410 21534 27412 21586
rect 27244 21532 27412 21534
rect 27468 21588 27524 21756
rect 27580 21588 27636 21598
rect 27468 21586 27636 21588
rect 27468 21534 27582 21586
rect 27634 21534 27636 21586
rect 27468 21532 27636 21534
rect 27132 21028 27188 21038
rect 27244 21028 27300 21532
rect 27356 21522 27412 21532
rect 26908 21026 27300 21028
rect 26908 20974 27134 21026
rect 27186 20974 27300 21026
rect 26908 20972 27300 20974
rect 26460 20934 26516 20972
rect 27132 20962 27188 20972
rect 27356 20916 27412 20926
rect 27580 20916 27636 21532
rect 27692 21588 27748 21868
rect 27692 21522 27748 21532
rect 27804 21028 27860 22204
rect 28028 21812 28084 21822
rect 28028 21474 28084 21756
rect 28028 21422 28030 21474
rect 28082 21422 28084 21474
rect 28028 21410 28084 21422
rect 28140 21364 28196 21374
rect 28140 21270 28196 21308
rect 28028 21028 28084 21038
rect 27804 21026 28084 21028
rect 27804 20974 28030 21026
rect 28082 20974 28084 21026
rect 27804 20972 28084 20974
rect 27412 20860 27636 20916
rect 28028 20914 28084 20972
rect 28028 20862 28030 20914
rect 28082 20862 28084 20914
rect 27356 20822 27412 20860
rect 28028 20850 28084 20862
rect 26908 20802 26964 20814
rect 26908 20750 26910 20802
rect 26962 20750 26964 20802
rect 26572 20692 26628 20702
rect 26572 20598 26628 20636
rect 26908 20356 26964 20750
rect 26908 20290 26964 20300
rect 27468 20690 27524 20702
rect 27468 20638 27470 20690
rect 27522 20638 27524 20690
rect 26236 20132 26404 20188
rect 25900 19618 25956 19628
rect 26236 19908 26292 19918
rect 26348 19908 26404 20132
rect 26796 20076 26964 20132
rect 26572 19908 26628 19918
rect 26796 19908 26852 20076
rect 26908 20018 26964 20076
rect 26908 19966 26910 20018
rect 26962 19966 26964 20018
rect 26908 19954 26964 19966
rect 26348 19906 26852 19908
rect 26348 19854 26574 19906
rect 26626 19854 26852 19906
rect 26348 19852 26852 19854
rect 25788 19394 25844 19404
rect 26236 19236 26292 19852
rect 26236 19142 26292 19180
rect 25788 19124 25844 19134
rect 25788 19122 26180 19124
rect 25788 19070 25790 19122
rect 25842 19070 26180 19122
rect 25788 19068 26180 19070
rect 25788 19058 25844 19068
rect 25900 18564 25956 18574
rect 25956 18508 26068 18564
rect 25900 18498 25956 18508
rect 26012 18450 26068 18508
rect 26012 18398 26014 18450
rect 26066 18398 26068 18450
rect 26012 18386 26068 18398
rect 26124 17778 26180 19068
rect 26572 18676 26628 19852
rect 26572 18610 26628 18620
rect 26796 19684 26852 19694
rect 26796 18676 26852 19628
rect 26796 18610 26852 18620
rect 27468 17892 27524 20638
rect 28252 20356 28308 22876
rect 28588 22596 28644 22606
rect 28476 22540 28588 22596
rect 28476 22482 28532 22540
rect 28588 22530 28644 22540
rect 28476 22430 28478 22482
rect 28530 22430 28532 22482
rect 28476 22418 28532 22430
rect 28476 21924 28532 21934
rect 28364 20580 28420 20590
rect 28364 20486 28420 20524
rect 28252 20300 28420 20356
rect 27692 19908 27748 19918
rect 27692 19906 28196 19908
rect 27692 19854 27694 19906
rect 27746 19854 28196 19906
rect 27692 19852 28196 19854
rect 27692 19842 27748 19852
rect 27916 19684 27972 19694
rect 27916 19234 27972 19628
rect 28140 19346 28196 19852
rect 28140 19294 28142 19346
rect 28194 19294 28196 19346
rect 28140 19282 28196 19294
rect 27916 19182 27918 19234
rect 27970 19182 27972 19234
rect 27916 19124 27972 19182
rect 27916 19058 27972 19068
rect 28252 19234 28308 19246
rect 28252 19182 28254 19234
rect 28306 19182 28308 19234
rect 27804 19010 27860 19022
rect 27804 18958 27806 19010
rect 27858 18958 27860 19010
rect 27804 18900 27860 18958
rect 28252 18900 28308 19182
rect 27804 18844 28308 18900
rect 28140 18338 28196 18350
rect 28140 18286 28142 18338
rect 28194 18286 28196 18338
rect 27468 17836 28084 17892
rect 26124 17726 26126 17778
rect 26178 17726 26180 17778
rect 26124 17714 26180 17726
rect 26012 17668 26068 17678
rect 26012 17574 26068 17612
rect 26236 17668 26292 17678
rect 26236 17574 26292 17612
rect 27132 17666 27188 17678
rect 27132 17614 27134 17666
rect 27186 17614 27188 17666
rect 26460 17444 26516 17454
rect 26460 17350 26516 17388
rect 26908 17442 26964 17454
rect 26908 17390 26910 17442
rect 26962 17390 26964 17442
rect 26908 17220 26964 17390
rect 26908 17154 26964 17164
rect 27132 17444 27188 17614
rect 27692 17444 27748 17454
rect 27132 17442 27748 17444
rect 27132 17390 27694 17442
rect 27746 17390 27748 17442
rect 27132 17388 27748 17390
rect 26908 16994 26964 17006
rect 26908 16942 26910 16994
rect 26962 16942 26964 16994
rect 25676 16594 25732 16604
rect 26572 16882 26628 16894
rect 26572 16830 26574 16882
rect 26626 16830 26628 16882
rect 26460 16210 26516 16222
rect 26460 16158 26462 16210
rect 26514 16158 26516 16210
rect 24332 15988 24388 15998
rect 25788 15988 25844 15998
rect 24332 15986 24724 15988
rect 24332 15934 24334 15986
rect 24386 15934 24724 15986
rect 24332 15932 24724 15934
rect 24332 15922 24388 15932
rect 24556 15090 24612 15102
rect 24556 15038 24558 15090
rect 24610 15038 24612 15090
rect 24332 14308 24388 14318
rect 23884 14306 24500 14308
rect 23884 14254 24334 14306
rect 24386 14254 24500 14306
rect 23884 14252 24500 14254
rect 24332 14242 24388 14252
rect 23660 14140 24164 14196
rect 23548 13918 23550 13970
rect 23602 13918 23604 13970
rect 23548 13636 23604 13918
rect 23996 13972 24052 13982
rect 23884 13860 23940 13870
rect 23884 13766 23940 13804
rect 23660 13746 23716 13758
rect 23660 13694 23662 13746
rect 23714 13694 23716 13746
rect 23660 13636 23716 13694
rect 23996 13746 24052 13916
rect 23996 13694 23998 13746
rect 24050 13694 24052 13746
rect 23996 13682 24052 13694
rect 23548 13580 23716 13636
rect 22092 13010 22148 13020
rect 22876 13300 22932 13310
rect 22092 12852 22148 12862
rect 22092 12758 22148 12796
rect 22092 10498 22148 10510
rect 22092 10446 22094 10498
rect 22146 10446 22148 10498
rect 22092 10276 22148 10446
rect 22652 10498 22708 10510
rect 22652 10446 22654 10498
rect 22706 10446 22708 10498
rect 22540 10388 22596 10398
rect 22092 10210 22148 10220
rect 22204 10386 22596 10388
rect 22204 10334 22542 10386
rect 22594 10334 22596 10386
rect 22204 10332 22596 10334
rect 22092 9940 22148 9950
rect 22204 9940 22260 10332
rect 22540 10322 22596 10332
rect 22092 9938 22260 9940
rect 22092 9886 22094 9938
rect 22146 9886 22260 9938
rect 22092 9884 22260 9886
rect 22652 9940 22708 10446
rect 22092 9874 22148 9884
rect 22652 9874 22708 9884
rect 21980 9538 22036 9548
rect 21644 8990 21646 9042
rect 21698 8990 21700 9042
rect 21308 6692 21364 6702
rect 20636 6244 20692 6254
rect 20636 6132 20692 6188
rect 20972 6132 21028 6142
rect 20636 6130 20804 6132
rect 20636 6078 20638 6130
rect 20690 6078 20804 6130
rect 20636 6076 20804 6078
rect 20636 6066 20692 6076
rect 20412 5854 20414 5906
rect 20466 5854 20468 5906
rect 19628 5794 19684 5806
rect 19628 5742 19630 5794
rect 19682 5742 19684 5794
rect 19628 5684 19684 5742
rect 19180 5628 19684 5684
rect 20412 5012 20468 5854
rect 20524 5908 20580 5918
rect 20524 5814 20580 5852
rect 20748 5234 20804 6076
rect 20972 5906 21028 6076
rect 20972 5854 20974 5906
rect 21026 5854 21028 5906
rect 20972 5842 21028 5854
rect 21308 5908 21364 6636
rect 21532 6466 21588 6478
rect 21532 6414 21534 6466
rect 21586 6414 21588 6466
rect 21532 6244 21588 6414
rect 21532 6178 21588 6188
rect 21644 6132 21700 8990
rect 22092 9156 22148 9166
rect 22092 7812 22148 9100
rect 22092 7362 22148 7756
rect 22764 8036 22820 8046
rect 22092 7310 22094 7362
rect 22146 7310 22148 7362
rect 22092 7298 22148 7310
rect 22540 7362 22596 7374
rect 22540 7310 22542 7362
rect 22594 7310 22596 7362
rect 22204 7252 22260 7262
rect 21980 6804 22036 6814
rect 21980 6690 22036 6748
rect 21980 6638 21982 6690
rect 22034 6638 22036 6690
rect 21980 6626 22036 6638
rect 22092 6466 22148 6478
rect 22092 6414 22094 6466
rect 22146 6414 22148 6466
rect 21700 6076 21924 6132
rect 21644 6066 21700 6076
rect 21308 5906 21700 5908
rect 21308 5854 21310 5906
rect 21362 5854 21700 5906
rect 21308 5852 21700 5854
rect 21308 5842 21364 5852
rect 20748 5182 20750 5234
rect 20802 5182 20804 5234
rect 20748 5170 20804 5182
rect 21420 5460 21476 5470
rect 21420 5234 21476 5404
rect 21420 5182 21422 5234
rect 21474 5182 21476 5234
rect 21420 5170 21476 5182
rect 21308 5012 21364 5022
rect 21532 5012 21588 5022
rect 20412 5010 21364 5012
rect 20412 4958 21310 5010
rect 21362 4958 21364 5010
rect 20412 4956 21364 4958
rect 21308 4946 21364 4956
rect 21420 4956 21532 5012
rect 21420 4788 21476 4956
rect 21532 4918 21588 4956
rect 19836 4732 20100 4742
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 19836 4666 20100 4676
rect 21196 4732 21476 4788
rect 19068 4398 19070 4450
rect 19122 4398 19124 4450
rect 19068 4386 19124 4398
rect 18284 4340 18340 4350
rect 17948 4338 18340 4340
rect 17948 4286 18286 4338
rect 18338 4286 18340 4338
rect 17948 4284 18340 4286
rect 18284 4274 18340 4284
rect 21196 4226 21252 4732
rect 21644 4340 21700 5852
rect 21868 5122 21924 6076
rect 22092 6018 22148 6414
rect 22092 5966 22094 6018
rect 22146 5966 22148 6018
rect 22092 5954 22148 5966
rect 21868 5070 21870 5122
rect 21922 5070 21924 5122
rect 21868 5058 21924 5070
rect 22204 5012 22260 7196
rect 22540 6692 22596 7310
rect 22764 6916 22820 7980
rect 22876 7364 22932 13244
rect 24108 12292 24164 14140
rect 24332 13748 24388 13758
rect 24332 13654 24388 13692
rect 24220 13524 24276 13534
rect 24220 13074 24276 13468
rect 24444 13188 24500 14252
rect 24556 13412 24612 15038
rect 24668 13524 24724 15932
rect 25228 15540 25284 15550
rect 25228 15446 25284 15484
rect 25788 15314 25844 15932
rect 25788 15262 25790 15314
rect 25842 15262 25844 15314
rect 25788 15250 25844 15262
rect 26012 15314 26068 15326
rect 26012 15262 26014 15314
rect 26066 15262 26068 15314
rect 24780 15204 24836 15214
rect 24780 14532 24836 15148
rect 25564 15204 25620 15242
rect 25564 15138 25620 15148
rect 25676 14642 25732 14654
rect 25676 14590 25678 14642
rect 25730 14590 25732 14642
rect 25004 14532 25060 14570
rect 24780 14530 24948 14532
rect 24780 14478 24782 14530
rect 24834 14478 24948 14530
rect 24780 14476 24948 14478
rect 24780 14466 24836 14476
rect 24668 13468 24836 13524
rect 24556 13356 24724 13412
rect 24556 13188 24612 13198
rect 24444 13132 24556 13188
rect 24556 13122 24612 13132
rect 24220 13022 24222 13074
rect 24274 13022 24276 13074
rect 24220 13010 24276 13022
rect 24668 12964 24724 13356
rect 24108 12226 24164 12236
rect 24444 12908 24724 12964
rect 23772 12068 23828 12078
rect 23436 11620 23492 11630
rect 23660 11620 23716 11630
rect 23436 11618 23660 11620
rect 23436 11566 23438 11618
rect 23490 11566 23660 11618
rect 23436 11564 23660 11566
rect 23212 11508 23268 11518
rect 23212 11414 23268 11452
rect 22988 11396 23044 11406
rect 22988 11302 23044 11340
rect 23100 10498 23156 10510
rect 23100 10446 23102 10498
rect 23154 10446 23156 10498
rect 23100 10164 23156 10446
rect 23100 10098 23156 10108
rect 23212 9268 23268 9278
rect 23436 9268 23492 11564
rect 23660 11554 23716 11564
rect 23772 11618 23828 12012
rect 23772 11566 23774 11618
rect 23826 11566 23828 11618
rect 23772 11554 23828 11566
rect 23884 12066 23940 12078
rect 23884 12014 23886 12066
rect 23938 12014 23940 12066
rect 23884 11172 23940 12014
rect 24444 11618 24500 12908
rect 24556 12292 24612 12302
rect 24556 12178 24612 12236
rect 24556 12126 24558 12178
rect 24610 12126 24612 12178
rect 24556 12114 24612 12126
rect 24780 11732 24836 13468
rect 24444 11566 24446 11618
rect 24498 11566 24500 11618
rect 24444 11554 24500 11566
rect 24556 11676 24836 11732
rect 24220 11508 24276 11518
rect 24220 11282 24276 11452
rect 24332 11396 24388 11406
rect 24556 11396 24612 11676
rect 24892 11620 24948 14476
rect 25004 14466 25060 14476
rect 25340 14420 25396 14430
rect 25676 14420 25732 14590
rect 25340 14418 25732 14420
rect 25340 14366 25342 14418
rect 25394 14366 25732 14418
rect 25340 14364 25732 14366
rect 25340 14354 25396 14364
rect 25004 14308 25060 14318
rect 25004 14214 25060 14252
rect 25564 13972 25620 13982
rect 25228 13746 25284 13758
rect 25228 13694 25230 13746
rect 25282 13694 25284 13746
rect 25116 13188 25172 13198
rect 25116 12962 25172 13132
rect 25116 12910 25118 12962
rect 25170 12910 25172 12962
rect 25116 12898 25172 12910
rect 25228 12516 25284 13694
rect 25452 13746 25508 13758
rect 25452 13694 25454 13746
rect 25506 13694 25508 13746
rect 25116 12460 25284 12516
rect 25340 13634 25396 13646
rect 25340 13582 25342 13634
rect 25394 13582 25396 13634
rect 25116 12068 25172 12460
rect 25340 12404 25396 13582
rect 25452 13636 25508 13694
rect 25452 13570 25508 13580
rect 25564 13412 25620 13916
rect 25676 13524 25732 14364
rect 26012 14308 26068 15262
rect 26236 15316 26292 15326
rect 26236 15202 26292 15260
rect 26236 15150 26238 15202
rect 26290 15150 26292 15202
rect 26236 15092 26292 15150
rect 26236 15026 26292 15036
rect 26348 15314 26404 15326
rect 26348 15262 26350 15314
rect 26402 15262 26404 15314
rect 25676 13458 25732 13468
rect 25900 13746 25956 13758
rect 25900 13694 25902 13746
rect 25954 13694 25956 13746
rect 25116 12002 25172 12012
rect 25228 12348 25396 12404
rect 25452 13356 25620 13412
rect 25788 13412 25844 13422
rect 24892 11554 24948 11564
rect 25116 11844 25172 11854
rect 24332 11394 24612 11396
rect 24332 11342 24334 11394
rect 24386 11342 24612 11394
rect 24332 11340 24612 11342
rect 24332 11330 24388 11340
rect 24220 11230 24222 11282
rect 24274 11230 24276 11282
rect 24220 11218 24276 11230
rect 23884 11106 23940 11116
rect 24892 11170 24948 11182
rect 24892 11118 24894 11170
rect 24946 11118 24948 11170
rect 23660 10836 23716 10846
rect 23660 10834 24052 10836
rect 23660 10782 23662 10834
rect 23714 10782 24052 10834
rect 23660 10780 24052 10782
rect 23660 10770 23716 10780
rect 23996 10724 24052 10780
rect 24332 10724 24388 10734
rect 23996 10722 24388 10724
rect 23996 10670 24334 10722
rect 24386 10670 24388 10722
rect 23996 10668 24388 10670
rect 23212 9266 23492 9268
rect 23212 9214 23214 9266
rect 23266 9214 23492 9266
rect 23212 9212 23492 9214
rect 23548 10610 23604 10622
rect 23548 10558 23550 10610
rect 23602 10558 23604 10610
rect 23548 10164 23604 10558
rect 23884 10612 23940 10622
rect 23884 10518 23940 10556
rect 24108 10386 24164 10398
rect 24108 10334 24110 10386
rect 24162 10334 24164 10386
rect 24108 10164 24164 10334
rect 23548 10108 24164 10164
rect 23548 9268 23604 10108
rect 24220 9938 24276 9950
rect 24220 9886 24222 9938
rect 24274 9886 24276 9938
rect 23660 9268 23716 9278
rect 23548 9266 23716 9268
rect 23548 9214 23662 9266
rect 23714 9214 23716 9266
rect 23548 9212 23716 9214
rect 23212 9202 23268 9212
rect 22988 9042 23044 9054
rect 22988 8990 22990 9042
rect 23042 8990 23044 9042
rect 22988 8372 23044 8990
rect 23436 9042 23492 9212
rect 23660 9202 23716 9212
rect 23436 8990 23438 9042
rect 23490 8990 23492 9042
rect 23436 8978 23492 8990
rect 23772 9044 23828 9054
rect 23772 8950 23828 8988
rect 24108 9044 24164 9054
rect 24220 9044 24276 9886
rect 24108 9042 24276 9044
rect 24108 8990 24110 9042
rect 24162 8990 24276 9042
rect 24108 8988 24276 8990
rect 24108 8978 24164 8988
rect 24220 8818 24276 8988
rect 24220 8766 24222 8818
rect 24274 8766 24276 8818
rect 24220 8754 24276 8766
rect 24332 8596 24388 10668
rect 24444 10386 24500 10398
rect 24444 10334 24446 10386
rect 24498 10334 24500 10386
rect 24444 10052 24500 10334
rect 24444 9986 24500 9996
rect 24556 10164 24612 10174
rect 24892 10164 24948 11118
rect 24612 10108 24948 10164
rect 24556 9266 24612 10108
rect 24668 9940 24724 9950
rect 24668 9846 24724 9884
rect 24556 9214 24558 9266
rect 24610 9214 24612 9266
rect 24556 9202 24612 9214
rect 24668 9714 24724 9726
rect 24668 9662 24670 9714
rect 24722 9662 24724 9714
rect 24668 8820 24724 9662
rect 24892 9714 24948 9726
rect 24892 9662 24894 9714
rect 24946 9662 24948 9714
rect 24892 8932 24948 9662
rect 24892 8866 24948 8876
rect 24780 8820 24836 8830
rect 24668 8818 24836 8820
rect 24668 8766 24782 8818
rect 24834 8766 24836 8818
rect 24668 8764 24836 8766
rect 24108 8540 24388 8596
rect 22988 8306 23044 8316
rect 23772 8372 23828 8382
rect 23772 8260 23828 8316
rect 23660 8258 23828 8260
rect 23660 8206 23774 8258
rect 23826 8206 23828 8258
rect 23660 8204 23828 8206
rect 23660 7586 23716 8204
rect 23772 8194 23828 8204
rect 23996 8260 24052 8270
rect 23996 8166 24052 8204
rect 23884 8036 23940 8046
rect 23884 7942 23940 7980
rect 23660 7534 23662 7586
rect 23714 7534 23716 7586
rect 23660 7522 23716 7534
rect 23884 7476 23940 7486
rect 23884 7382 23940 7420
rect 22876 7298 22932 7308
rect 23772 7362 23828 7374
rect 23772 7310 23774 7362
rect 23826 7310 23828 7362
rect 23772 6916 23828 7310
rect 24108 7252 24164 8540
rect 24780 8484 24836 8764
rect 25004 8484 25060 8494
rect 24780 8482 25060 8484
rect 24780 8430 25006 8482
rect 25058 8430 25060 8482
rect 24780 8428 25060 8430
rect 25004 8418 25060 8428
rect 24332 8260 24388 8270
rect 24332 8166 24388 8204
rect 24780 8260 24836 8270
rect 25116 8260 25172 11788
rect 25228 11394 25284 12348
rect 25340 12068 25396 12078
rect 25340 11974 25396 12012
rect 25228 11342 25230 11394
rect 25282 11342 25284 11394
rect 25228 11330 25284 11342
rect 25340 10836 25396 10846
rect 25452 10836 25508 13356
rect 25676 13076 25732 13086
rect 25676 12292 25732 13020
rect 25676 12226 25732 12236
rect 25788 12178 25844 13356
rect 25900 12516 25956 13694
rect 26012 13636 26068 14252
rect 26012 13570 26068 13580
rect 26124 13634 26180 13646
rect 26124 13582 26126 13634
rect 26178 13582 26180 13634
rect 26124 13412 26180 13582
rect 26124 13346 26180 13356
rect 26236 13522 26292 13534
rect 26236 13470 26238 13522
rect 26290 13470 26292 13522
rect 25900 12460 26068 12516
rect 25788 12126 25790 12178
rect 25842 12126 25844 12178
rect 25676 11956 25732 11966
rect 25676 11394 25732 11900
rect 25788 11844 25844 12126
rect 25788 11778 25844 11788
rect 25900 12292 25956 12302
rect 25676 11342 25678 11394
rect 25730 11342 25732 11394
rect 25676 11330 25732 11342
rect 25788 11396 25844 11434
rect 25788 11330 25844 11340
rect 25676 11172 25732 11182
rect 25676 11078 25732 11116
rect 25340 10834 25844 10836
rect 25340 10782 25342 10834
rect 25394 10782 25844 10834
rect 25340 10780 25844 10782
rect 25340 10770 25396 10780
rect 25452 10612 25508 10622
rect 25452 10518 25508 10556
rect 25340 10388 25396 10398
rect 25788 10388 25844 10780
rect 25900 10612 25956 12236
rect 26012 12180 26068 12460
rect 26124 12180 26180 12190
rect 26012 12178 26180 12180
rect 26012 12126 26126 12178
rect 26178 12126 26180 12178
rect 26012 12124 26180 12126
rect 26012 11396 26068 11406
rect 26012 11302 26068 11340
rect 26012 10836 26068 10846
rect 26124 10836 26180 12124
rect 26236 11394 26292 13470
rect 26348 13412 26404 15262
rect 26460 13748 26516 16158
rect 26572 15988 26628 16830
rect 26908 16772 26964 16942
rect 26572 15922 26628 15932
rect 26796 16716 26964 16772
rect 26572 15540 26628 15550
rect 26796 15540 26852 16716
rect 26908 16660 26964 16716
rect 26908 16594 26964 16604
rect 27132 16100 27188 17388
rect 27692 17378 27748 17388
rect 27244 16996 27300 17006
rect 27244 16770 27300 16940
rect 27244 16718 27246 16770
rect 27298 16718 27300 16770
rect 27244 16706 27300 16718
rect 27132 16034 27188 16044
rect 26572 15538 26852 15540
rect 26572 15486 26574 15538
rect 26626 15486 26852 15538
rect 26572 15484 26852 15486
rect 27132 15540 27188 15550
rect 27132 15538 27860 15540
rect 27132 15486 27134 15538
rect 27186 15486 27860 15538
rect 27132 15484 27860 15486
rect 26572 15474 26628 15484
rect 27132 15474 27188 15484
rect 26796 15314 26852 15326
rect 26796 15262 26798 15314
rect 26850 15262 26852 15314
rect 26572 15204 26628 15214
rect 26572 13972 26628 15148
rect 26572 13906 26628 13916
rect 26796 13970 26852 15262
rect 27244 15314 27300 15326
rect 27244 15262 27246 15314
rect 27298 15262 27300 15314
rect 27132 15092 27188 15102
rect 27244 15092 27300 15262
rect 27468 15314 27524 15326
rect 27468 15262 27470 15314
rect 27522 15262 27524 15314
rect 27468 15204 27524 15262
rect 27468 15138 27524 15148
rect 27188 15036 27300 15092
rect 27132 15026 27188 15036
rect 26796 13918 26798 13970
rect 26850 13918 26852 13970
rect 26796 13906 26852 13918
rect 26908 14980 26964 14990
rect 26460 13682 26516 13692
rect 26684 13748 26740 13758
rect 26684 13746 26852 13748
rect 26684 13694 26686 13746
rect 26738 13694 26852 13746
rect 26684 13692 26852 13694
rect 26684 13682 26740 13692
rect 26572 13412 26628 13422
rect 26348 13356 26572 13412
rect 26572 12402 26628 13356
rect 26572 12350 26574 12402
rect 26626 12350 26628 12402
rect 26572 12338 26628 12350
rect 26796 12404 26852 13692
rect 26796 12178 26852 12348
rect 26796 12126 26798 12178
rect 26850 12126 26852 12178
rect 26796 12114 26852 12126
rect 26796 11956 26852 11966
rect 26796 11862 26852 11900
rect 26236 11342 26238 11394
rect 26290 11342 26292 11394
rect 26236 11330 26292 11342
rect 26684 11396 26740 11406
rect 26684 11060 26740 11340
rect 26684 10994 26740 11004
rect 26068 10780 26180 10836
rect 26012 10770 26068 10780
rect 26684 10724 26740 10734
rect 26684 10630 26740 10668
rect 25900 10610 26516 10612
rect 25900 10558 25902 10610
rect 25954 10558 26516 10610
rect 25900 10556 26516 10558
rect 25900 10546 25956 10556
rect 25340 10386 25620 10388
rect 25340 10334 25342 10386
rect 25394 10334 25620 10386
rect 25340 10332 25620 10334
rect 25788 10332 26180 10388
rect 25340 10322 25396 10332
rect 25452 10052 25508 10062
rect 25452 9958 25508 9996
rect 25564 10050 25620 10332
rect 25564 9998 25566 10050
rect 25618 9998 25620 10050
rect 25564 9986 25620 9998
rect 26124 9938 26180 10332
rect 26124 9886 26126 9938
rect 26178 9886 26180 9938
rect 26124 9874 26180 9886
rect 25228 9716 25284 9726
rect 25452 9716 25508 9726
rect 25228 9714 25452 9716
rect 25228 9662 25230 9714
rect 25282 9662 25452 9714
rect 25228 9660 25452 9662
rect 25228 9650 25284 9660
rect 25452 9650 25508 9660
rect 26012 9716 26068 9726
rect 25788 8932 25844 8942
rect 24780 8258 25172 8260
rect 24780 8206 24782 8258
rect 24834 8206 25172 8258
rect 24780 8204 25172 8206
rect 25228 8258 25284 8270
rect 25228 8206 25230 8258
rect 25282 8206 25284 8258
rect 24780 8194 24836 8204
rect 25004 8036 25060 8046
rect 24220 7476 24276 7486
rect 24276 7420 24500 7476
rect 24220 7382 24276 7420
rect 24108 7196 24388 7252
rect 22764 6914 23268 6916
rect 22764 6862 22766 6914
rect 22818 6862 23268 6914
rect 22764 6860 23268 6862
rect 22764 6850 22820 6860
rect 22428 6466 22484 6478
rect 22428 6414 22430 6466
rect 22482 6414 22484 6466
rect 22428 6356 22484 6414
rect 22428 6290 22484 6300
rect 22540 6132 22596 6636
rect 22988 6692 23044 6702
rect 22988 6598 23044 6636
rect 22316 5236 22372 5246
rect 22540 5236 22596 6076
rect 22316 5234 22596 5236
rect 22316 5182 22318 5234
rect 22370 5182 22596 5234
rect 22316 5180 22596 5182
rect 22876 5236 22932 5246
rect 22316 5170 22372 5180
rect 22204 4946 22260 4956
rect 21196 4174 21198 4226
rect 21250 4174 21252 4226
rect 21196 4162 21252 4174
rect 21532 4338 21700 4340
rect 21532 4286 21646 4338
rect 21698 4286 21700 4338
rect 21532 4284 21700 4286
rect 4476 3948 4740 3958
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4476 3882 4740 3892
rect 21532 3666 21588 4284
rect 21644 4274 21700 4284
rect 22316 4228 22372 4238
rect 22316 4226 22820 4228
rect 22316 4174 22318 4226
rect 22370 4174 22820 4226
rect 22316 4172 22820 4174
rect 22316 4162 22372 4172
rect 22764 3778 22820 4172
rect 22764 3726 22766 3778
rect 22818 3726 22820 3778
rect 22764 3714 22820 3726
rect 21532 3614 21534 3666
rect 21586 3614 21588 3666
rect 21532 3602 21588 3614
rect 22876 3666 22932 5180
rect 23212 5010 23268 6860
rect 23324 6692 23380 6702
rect 23772 6692 23828 6860
rect 24332 6802 24388 7196
rect 24332 6750 24334 6802
rect 24386 6750 24388 6802
rect 23884 6692 23940 6702
rect 24220 6692 24276 6702
rect 23772 6690 23940 6692
rect 23772 6638 23886 6690
rect 23938 6638 23940 6690
rect 23772 6636 23940 6638
rect 23324 5796 23380 6636
rect 23884 6626 23940 6636
rect 24108 6690 24276 6692
rect 24108 6638 24222 6690
rect 24274 6638 24276 6690
rect 24108 6636 24276 6638
rect 23436 6468 23492 6478
rect 23492 6412 23604 6468
rect 23436 6374 23492 6412
rect 23548 5908 23604 6412
rect 23660 6466 23716 6478
rect 23660 6414 23662 6466
rect 23714 6414 23716 6466
rect 23660 6356 23716 6414
rect 23772 6468 23828 6478
rect 24108 6468 24164 6636
rect 24220 6626 24276 6636
rect 24332 6692 24388 6750
rect 24332 6626 24388 6636
rect 24444 6468 24500 7420
rect 24892 7364 24948 7374
rect 24892 6690 24948 7308
rect 24892 6638 24894 6690
rect 24946 6638 24948 6690
rect 24892 6626 24948 6638
rect 24668 6580 24724 6590
rect 23772 6466 24164 6468
rect 23772 6414 23774 6466
rect 23826 6414 24164 6466
rect 23772 6412 24164 6414
rect 24220 6412 24500 6468
rect 24556 6524 24668 6580
rect 23772 6402 23828 6412
rect 23660 6020 23716 6300
rect 23660 5964 24164 6020
rect 23548 5852 23828 5908
rect 23324 5684 23380 5740
rect 23324 5628 23492 5684
rect 23324 5124 23380 5134
rect 23324 5030 23380 5068
rect 23436 5122 23492 5628
rect 23436 5070 23438 5122
rect 23490 5070 23492 5122
rect 23436 5058 23492 5070
rect 23772 5122 23828 5852
rect 24108 5348 24164 5964
rect 24220 5794 24276 6412
rect 24220 5742 24222 5794
rect 24274 5742 24276 5794
rect 24220 5730 24276 5742
rect 24220 5348 24276 5358
rect 24108 5346 24276 5348
rect 24108 5294 24222 5346
rect 24274 5294 24276 5346
rect 24108 5292 24276 5294
rect 24220 5282 24276 5292
rect 23772 5070 23774 5122
rect 23826 5070 23828 5122
rect 23772 5058 23828 5070
rect 24108 5124 24164 5134
rect 24108 5030 24164 5068
rect 23212 4958 23214 5010
rect 23266 4958 23268 5010
rect 23212 4946 23268 4958
rect 24556 5010 24612 6524
rect 24668 6486 24724 6524
rect 25004 6356 25060 7980
rect 25228 7476 25284 8206
rect 25452 8260 25508 8270
rect 25452 8166 25508 8204
rect 25116 6804 25172 6814
rect 25116 6710 25172 6748
rect 25228 6690 25284 7420
rect 25452 7476 25508 7486
rect 25788 7476 25844 8876
rect 25900 8034 25956 8046
rect 25900 7982 25902 8034
rect 25954 7982 25956 8034
rect 25900 7588 25956 7982
rect 25900 7522 25956 7532
rect 25452 7474 25844 7476
rect 25452 7422 25454 7474
rect 25506 7422 25844 7474
rect 25452 7420 25844 7422
rect 25340 7364 25396 7374
rect 25452 7364 25508 7420
rect 25396 7308 25508 7364
rect 25340 7298 25396 7308
rect 25788 6916 25844 6926
rect 25788 6822 25844 6860
rect 25228 6638 25230 6690
rect 25282 6638 25284 6690
rect 25228 6626 25284 6638
rect 25564 6690 25620 6702
rect 25564 6638 25566 6690
rect 25618 6638 25620 6690
rect 25564 6356 25620 6638
rect 26012 6580 26068 9660
rect 26460 9044 26516 10556
rect 26908 9940 26964 14924
rect 27804 14642 27860 15484
rect 27916 15204 27972 15242
rect 27916 15138 27972 15148
rect 27804 14590 27806 14642
rect 27858 14590 27860 14642
rect 27804 14578 27860 14590
rect 27692 13970 27748 13982
rect 27692 13918 27694 13970
rect 27746 13918 27748 13970
rect 27244 13860 27300 13870
rect 27692 13860 27748 13918
rect 27244 13858 27748 13860
rect 27244 13806 27246 13858
rect 27298 13806 27748 13858
rect 27244 13804 27748 13806
rect 27244 13794 27300 13804
rect 27020 13746 27076 13758
rect 28028 13748 28084 17836
rect 28140 17668 28196 18286
rect 28140 17602 28196 17612
rect 28140 17444 28196 17454
rect 28140 17350 28196 17388
rect 28252 15148 28308 18844
rect 28364 18340 28420 20300
rect 28364 18274 28420 18284
rect 28476 17892 28532 21868
rect 28700 21476 28756 21486
rect 28700 21026 28756 21420
rect 28700 20974 28702 21026
rect 28754 20974 28756 21026
rect 28700 20962 28756 20974
rect 28924 19908 28980 31052
rect 29036 30324 29092 30334
rect 29036 30230 29092 30268
rect 29148 29988 29204 31388
rect 29484 30098 29540 31500
rect 29596 31220 29652 31726
rect 29596 31154 29652 31164
rect 30380 31332 30436 31342
rect 29484 30046 29486 30098
rect 29538 30046 29540 30098
rect 29484 30034 29540 30046
rect 29820 30212 29876 30222
rect 29708 29988 29764 29998
rect 29148 29932 29316 29988
rect 29148 29764 29204 29774
rect 29148 29426 29204 29708
rect 29148 29374 29150 29426
rect 29202 29374 29204 29426
rect 29148 29362 29204 29374
rect 29260 29314 29316 29932
rect 29596 29932 29708 29988
rect 29372 29428 29428 29438
rect 29428 29372 29540 29428
rect 29372 29362 29428 29372
rect 29260 29262 29262 29314
rect 29314 29262 29316 29314
rect 29260 29250 29316 29262
rect 29148 29204 29204 29214
rect 29148 28530 29204 29148
rect 29148 28478 29150 28530
rect 29202 28478 29204 28530
rect 29148 28466 29204 28478
rect 29372 28644 29428 28654
rect 29036 27748 29092 27758
rect 29036 24724 29092 27692
rect 29372 27746 29428 28588
rect 29484 28642 29540 29372
rect 29484 28590 29486 28642
rect 29538 28590 29540 28642
rect 29484 28578 29540 28590
rect 29372 27694 29374 27746
rect 29426 27694 29428 27746
rect 29372 27300 29428 27694
rect 29596 27300 29652 29932
rect 29708 29922 29764 29932
rect 29708 29540 29764 29550
rect 29708 29446 29764 29484
rect 29820 28530 29876 30156
rect 30156 30210 30212 30222
rect 30156 30158 30158 30210
rect 30210 30158 30212 30210
rect 29932 30098 29988 30110
rect 29932 30046 29934 30098
rect 29986 30046 29988 30098
rect 29932 29988 29988 30046
rect 29932 29922 29988 29932
rect 29932 29764 29988 29774
rect 29932 29540 29988 29708
rect 30044 29540 30100 29550
rect 29932 29484 30044 29540
rect 29932 29426 29988 29484
rect 30044 29474 30100 29484
rect 29932 29374 29934 29426
rect 29986 29374 29988 29426
rect 29932 29362 29988 29374
rect 30156 28980 30212 30158
rect 30380 29652 30436 31276
rect 30492 30212 30548 37324
rect 30716 37156 30772 37166
rect 30716 37062 30772 37100
rect 30716 36260 30772 36270
rect 30716 36166 30772 36204
rect 30828 35812 30884 38612
rect 30940 38052 30996 38062
rect 30940 37938 30996 37996
rect 30940 37886 30942 37938
rect 30994 37886 30996 37938
rect 30940 37874 30996 37886
rect 30716 35756 30884 35812
rect 30940 36596 30996 36606
rect 30604 33572 30660 33582
rect 30604 33458 30660 33516
rect 30604 33406 30606 33458
rect 30658 33406 30660 33458
rect 30604 33394 30660 33406
rect 30492 30118 30548 30156
rect 30604 31108 30660 31118
rect 30716 31108 30772 35756
rect 30940 35700 30996 36540
rect 31164 36484 31220 38556
rect 31276 38164 31332 39004
rect 31500 38722 31556 39676
rect 31724 39666 31780 39676
rect 31836 40402 31892 40414
rect 31836 40350 31838 40402
rect 31890 40350 31892 40402
rect 31724 39284 31780 39294
rect 31724 38834 31780 39228
rect 31836 39060 31892 40350
rect 31836 38994 31892 39004
rect 31724 38782 31726 38834
rect 31778 38782 31780 38834
rect 31724 38770 31780 38782
rect 31948 38836 32004 40572
rect 32172 40626 33124 40628
rect 32172 40574 32174 40626
rect 32226 40574 33124 40626
rect 32172 40572 33124 40574
rect 32172 40562 32228 40572
rect 32060 40516 32116 40526
rect 32060 40402 32116 40460
rect 32060 40350 32062 40402
rect 32114 40350 32116 40402
rect 32060 40338 32116 40350
rect 32284 40402 32340 40414
rect 32284 40350 32286 40402
rect 32338 40350 32340 40402
rect 32172 40180 32228 40190
rect 31948 38770 32004 38780
rect 32060 39396 32116 39406
rect 31500 38670 31502 38722
rect 31554 38670 31556 38722
rect 31500 38658 31556 38670
rect 32060 38668 32116 39340
rect 31836 38612 32116 38668
rect 31836 38546 31892 38556
rect 32172 38276 32228 40124
rect 32284 39060 32340 40350
rect 32396 40292 32452 40302
rect 32396 39618 32452 40236
rect 33068 39732 33124 40572
rect 33180 40514 33236 40684
rect 33180 40462 33182 40514
rect 33234 40462 33236 40514
rect 33180 40450 33236 40462
rect 33292 40514 33348 40526
rect 33292 40462 33294 40514
rect 33346 40462 33348 40514
rect 33180 39732 33236 39742
rect 33068 39730 33236 39732
rect 33068 39678 33182 39730
rect 33234 39678 33236 39730
rect 33068 39676 33236 39678
rect 33180 39666 33236 39676
rect 33292 39732 33348 40462
rect 33404 40404 33460 40684
rect 33516 40628 33572 41134
rect 33740 40964 33796 45052
rect 33852 44324 33908 44334
rect 33852 44230 33908 44268
rect 33964 44100 34020 45276
rect 34076 45106 34132 45118
rect 34076 45054 34078 45106
rect 34130 45054 34132 45106
rect 34076 44324 34132 45054
rect 34188 44436 34244 45724
rect 34524 45778 34580 46956
rect 34748 46900 34804 46910
rect 34524 45726 34526 45778
rect 34578 45726 34580 45778
rect 34524 45714 34580 45726
rect 34636 46788 34692 46798
rect 34300 45444 34356 45454
rect 34300 45330 34356 45388
rect 34300 45278 34302 45330
rect 34354 45278 34356 45330
rect 34300 45266 34356 45278
rect 34412 45332 34468 45342
rect 34412 45238 34468 45276
rect 34524 45332 34580 45342
rect 34636 45332 34692 46732
rect 34748 46004 34804 46844
rect 35084 46450 35140 47068
rect 35196 47058 35252 47068
rect 35308 46788 35364 46798
rect 35308 46694 35364 46732
rect 35084 46398 35086 46450
rect 35138 46398 35140 46450
rect 34748 45938 34804 45948
rect 34860 46116 34916 46126
rect 34860 45890 34916 46060
rect 34860 45838 34862 45890
rect 34914 45838 34916 45890
rect 34860 45826 34916 45838
rect 34524 45330 34692 45332
rect 34524 45278 34526 45330
rect 34578 45278 34692 45330
rect 34524 45276 34692 45278
rect 34524 44884 34580 45276
rect 34748 45108 34804 45118
rect 35084 45108 35140 46398
rect 35420 46452 35476 47406
rect 35532 47460 35588 48190
rect 35532 47394 35588 47404
rect 35644 47458 35700 47470
rect 35644 47406 35646 47458
rect 35698 47406 35700 47458
rect 35644 46452 35700 47406
rect 35756 47348 35812 50540
rect 35868 50036 35924 51102
rect 36092 50706 36148 51550
rect 36092 50654 36094 50706
rect 36146 50654 36148 50706
rect 36092 50642 36148 50654
rect 36876 50708 36932 52332
rect 37100 52836 37156 52846
rect 37100 52162 37156 52780
rect 37100 52110 37102 52162
rect 37154 52110 37156 52162
rect 37100 52098 37156 52110
rect 36988 52050 37044 52062
rect 36988 51998 36990 52050
rect 37042 51998 37044 52050
rect 36988 51716 37044 51998
rect 36988 51660 37268 51716
rect 36988 51492 37044 51502
rect 36988 51398 37044 51436
rect 37212 51490 37268 51660
rect 37212 51438 37214 51490
rect 37266 51438 37268 51490
rect 37212 51426 37268 51438
rect 37100 51268 37156 51278
rect 37324 51268 37380 52892
rect 37660 52948 37716 52958
rect 37660 52854 37716 52892
rect 37548 52834 37604 52846
rect 37548 52782 37550 52834
rect 37602 52782 37604 52834
rect 37548 52724 37604 52782
rect 37772 52724 37828 53004
rect 37996 52946 38052 53788
rect 37996 52894 37998 52946
rect 38050 52894 38052 52946
rect 37996 52882 38052 52894
rect 38108 53506 38164 53518
rect 38108 53454 38110 53506
rect 38162 53454 38164 53506
rect 37548 52668 37828 52724
rect 37436 52164 37492 52174
rect 37436 52070 37492 52108
rect 38108 52164 38164 53454
rect 38220 53058 38276 53070
rect 38220 53006 38222 53058
rect 38274 53006 38276 53058
rect 38220 52276 38276 53006
rect 38332 52948 38388 54348
rect 38444 53732 38500 53742
rect 38444 53638 38500 53676
rect 38556 53508 38612 55468
rect 38892 54740 38948 54750
rect 38668 54514 38724 54526
rect 38668 54462 38670 54514
rect 38722 54462 38724 54514
rect 38668 53844 38724 54462
rect 38668 53778 38724 53788
rect 38332 52882 38388 52892
rect 38444 53452 38612 53508
rect 38220 52210 38276 52220
rect 38108 51940 38164 52108
rect 38332 52164 38388 52174
rect 38444 52164 38500 53452
rect 38892 53396 38948 54684
rect 39004 53508 39060 56028
rect 39788 56018 39844 56028
rect 39340 55748 39396 55758
rect 39116 55298 39172 55310
rect 39116 55246 39118 55298
rect 39170 55246 39172 55298
rect 39116 53732 39172 55246
rect 39340 54738 39396 55692
rect 39900 55468 39956 57372
rect 40796 56308 40852 56318
rect 40796 56214 40852 56252
rect 39340 54686 39342 54738
rect 39394 54686 39396 54738
rect 39340 54674 39396 54686
rect 39788 55412 39956 55468
rect 41132 56084 41188 56094
rect 39452 54628 39508 54638
rect 39228 54514 39284 54526
rect 39228 54462 39230 54514
rect 39282 54462 39284 54514
rect 39228 54404 39284 54462
rect 39452 54514 39508 54572
rect 39452 54462 39454 54514
rect 39506 54462 39508 54514
rect 39452 54450 39508 54462
rect 39676 54516 39732 54526
rect 39676 54422 39732 54460
rect 39228 54338 39284 54348
rect 39116 53666 39172 53676
rect 39228 53732 39284 53742
rect 39228 53730 39732 53732
rect 39228 53678 39230 53730
rect 39282 53678 39732 53730
rect 39228 53676 39732 53678
rect 39228 53666 39284 53676
rect 39004 53452 39284 53508
rect 38892 53340 39172 53396
rect 39004 53170 39060 53182
rect 39004 53118 39006 53170
rect 39058 53118 39060 53170
rect 38892 52948 38948 52958
rect 38556 52946 38948 52948
rect 38556 52894 38894 52946
rect 38946 52894 38948 52946
rect 38556 52892 38948 52894
rect 38556 52274 38612 52892
rect 38892 52882 38948 52892
rect 39004 52612 39060 53118
rect 39004 52546 39060 52556
rect 38668 52388 38724 52398
rect 39116 52388 39172 53340
rect 38668 52386 39172 52388
rect 38668 52334 38670 52386
rect 38722 52334 39172 52386
rect 38668 52332 39172 52334
rect 38668 52322 38724 52332
rect 38556 52222 38558 52274
rect 38610 52222 38612 52274
rect 38556 52210 38612 52222
rect 38332 52162 38500 52164
rect 38332 52110 38334 52162
rect 38386 52110 38500 52162
rect 38332 52108 38500 52110
rect 39116 52164 39172 52174
rect 38332 52098 38388 52108
rect 39116 52070 39172 52108
rect 37996 51884 38164 51940
rect 38556 52052 38612 52062
rect 37660 51604 37716 51614
rect 37996 51604 38052 51884
rect 37716 51548 38052 51604
rect 37660 51510 37716 51548
rect 37100 51266 37380 51268
rect 37100 51214 37102 51266
rect 37154 51214 37380 51266
rect 37100 51212 37380 51214
rect 37100 51202 37156 51212
rect 37100 50820 37156 50830
rect 37100 50726 37156 50764
rect 36876 50642 36932 50652
rect 37548 50708 37604 50718
rect 37548 50614 37604 50652
rect 35980 50594 36036 50606
rect 37884 50596 37940 51548
rect 35980 50542 35982 50594
rect 36034 50542 36036 50594
rect 35980 50260 36036 50542
rect 37660 50594 37940 50596
rect 37660 50542 37886 50594
rect 37938 50542 37940 50594
rect 37660 50540 37940 50542
rect 36316 50484 36372 50522
rect 36316 50418 36372 50428
rect 36988 50484 37044 50522
rect 37660 50484 37716 50540
rect 37884 50530 37940 50540
rect 38108 51492 38164 51502
rect 35980 50194 36036 50204
rect 36764 50260 36820 50270
rect 35868 49970 35924 49980
rect 36652 50036 36708 50046
rect 36652 49942 36708 49980
rect 36316 49812 36372 49822
rect 36540 49812 36596 49822
rect 36316 49718 36372 49756
rect 36428 49810 36596 49812
rect 36428 49758 36542 49810
rect 36594 49758 36596 49810
rect 36428 49756 36596 49758
rect 35980 49700 36036 49710
rect 35980 49606 36036 49644
rect 36428 49364 36484 49756
rect 36540 49746 36596 49756
rect 36764 49810 36820 50204
rect 36764 49758 36766 49810
rect 36818 49758 36820 49810
rect 35980 49308 36484 49364
rect 35980 49252 36036 49308
rect 35980 49158 36036 49196
rect 36764 49028 36820 49758
rect 36988 49810 37044 50428
rect 36988 49758 36990 49810
rect 37042 49758 37044 49810
rect 36988 49140 37044 49758
rect 37436 50428 37716 50484
rect 38108 50428 38164 51436
rect 37436 50034 37492 50428
rect 37436 49982 37438 50034
rect 37490 49982 37492 50034
rect 36988 49074 37044 49084
rect 37100 49588 37156 49598
rect 37100 49138 37156 49532
rect 37436 49476 37492 49982
rect 37436 49410 37492 49420
rect 37996 50372 38164 50428
rect 37100 49086 37102 49138
rect 37154 49086 37156 49138
rect 35756 47282 35812 47292
rect 35868 48972 36148 49028
rect 35868 48130 35924 48972
rect 36092 48916 36148 48972
rect 36764 48962 36820 48972
rect 36092 48822 36148 48860
rect 37100 48916 37156 49086
rect 37100 48850 37156 48860
rect 37772 49140 37828 49150
rect 37996 49140 38052 50372
rect 38108 50260 38164 50270
rect 38108 50034 38164 50204
rect 38108 49982 38110 50034
rect 38162 49982 38164 50034
rect 38108 49970 38164 49982
rect 38220 49700 38276 49710
rect 38220 49606 38276 49644
rect 37828 49084 38052 49140
rect 35868 48078 35870 48130
rect 35922 48078 35924 48130
rect 35644 46396 35812 46452
rect 35420 46386 35476 46396
rect 35196 46284 35460 46294
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35196 46218 35460 46228
rect 35196 46004 35252 46014
rect 35252 45948 35364 46004
rect 35196 45938 35252 45948
rect 34748 45106 35140 45108
rect 34748 45054 34750 45106
rect 34802 45054 35140 45106
rect 34748 45052 35140 45054
rect 35308 45108 35364 45948
rect 35756 45332 35812 46396
rect 35868 46116 35924 48078
rect 35980 48802 36036 48814
rect 35980 48750 35982 48802
rect 36034 48750 36036 48802
rect 35980 48132 36036 48750
rect 37212 48804 37268 48814
rect 37268 48748 37380 48804
rect 37212 48738 37268 48748
rect 36316 48132 36372 48142
rect 35980 48130 36372 48132
rect 35980 48078 36318 48130
rect 36370 48078 36372 48130
rect 35980 48076 36372 48078
rect 36204 47234 36260 47246
rect 36204 47182 36206 47234
rect 36258 47182 36260 47234
rect 36204 46676 36260 47182
rect 36316 47124 36372 48076
rect 36316 47058 36372 47068
rect 36428 47348 36484 47358
rect 36316 46676 36372 46686
rect 36204 46674 36372 46676
rect 36204 46622 36318 46674
rect 36370 46622 36372 46674
rect 36204 46620 36372 46622
rect 35868 46050 35924 46060
rect 36092 46452 36148 46462
rect 35308 45106 35700 45108
rect 35308 45054 35310 45106
rect 35362 45054 35700 45106
rect 35308 45052 35700 45054
rect 34524 44828 34692 44884
rect 34636 44546 34692 44828
rect 34636 44494 34638 44546
rect 34690 44494 34692 44546
rect 34636 44482 34692 44494
rect 34524 44436 34580 44446
rect 34188 44434 34580 44436
rect 34188 44382 34526 44434
rect 34578 44382 34580 44434
rect 34188 44380 34580 44382
rect 34524 44370 34580 44380
rect 34748 44436 34804 45052
rect 35308 45042 35364 45052
rect 35196 44716 35460 44726
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35196 44650 35460 44660
rect 34748 44370 34804 44380
rect 34076 44268 34244 44324
rect 34188 44210 34244 44268
rect 34188 44158 34190 44210
rect 34242 44158 34244 44210
rect 34076 44100 34132 44110
rect 33964 44098 34132 44100
rect 33964 44046 34078 44098
rect 34130 44046 34132 44098
rect 33964 44044 34132 44046
rect 34076 44034 34132 44044
rect 34188 42868 34244 44158
rect 35644 43540 35700 45052
rect 35756 44546 35812 45276
rect 35756 44494 35758 44546
rect 35810 44494 35812 44546
rect 35756 44482 35812 44494
rect 35868 45890 35924 45902
rect 35868 45838 35870 45890
rect 35922 45838 35924 45890
rect 35868 44434 35924 45838
rect 35868 44382 35870 44434
rect 35922 44382 35924 44434
rect 35868 44370 35924 44382
rect 35980 44994 36036 45006
rect 35980 44942 35982 44994
rect 36034 44942 36036 44994
rect 35980 44100 36036 44942
rect 36092 44322 36148 46396
rect 36316 45892 36372 46620
rect 36428 46002 36484 47292
rect 37212 47348 37268 47358
rect 37212 47254 37268 47292
rect 37100 47012 37156 47022
rect 36988 46564 37044 46574
rect 36428 45950 36430 46002
rect 36482 45950 36484 46002
rect 36428 45938 36484 45950
rect 36876 46508 36988 46564
rect 36876 46004 36932 46508
rect 36988 46470 37044 46508
rect 36876 45938 36932 45948
rect 36316 45826 36372 45836
rect 36764 45892 36820 45902
rect 36092 44270 36094 44322
rect 36146 44270 36148 44322
rect 36092 44258 36148 44270
rect 35980 44044 36484 44100
rect 36428 43762 36484 44044
rect 36428 43710 36430 43762
rect 36482 43710 36484 43762
rect 36428 43698 36484 43710
rect 36316 43652 36372 43662
rect 36316 43558 36372 43596
rect 35868 43540 35924 43550
rect 35644 43538 36260 43540
rect 35644 43486 35870 43538
rect 35922 43486 36260 43538
rect 35644 43484 36260 43486
rect 35868 43474 35924 43484
rect 35196 43428 35252 43438
rect 35084 43426 35252 43428
rect 35084 43374 35198 43426
rect 35250 43374 35252 43426
rect 35084 43372 35252 43374
rect 34188 42866 34692 42868
rect 34188 42814 34190 42866
rect 34242 42814 34692 42866
rect 34188 42812 34692 42814
rect 34188 42802 34244 42812
rect 34076 42756 34132 42766
rect 34076 42662 34132 42700
rect 34636 42754 34692 42812
rect 34636 42702 34638 42754
rect 34690 42702 34692 42754
rect 34636 42690 34692 42702
rect 34300 42532 34356 42542
rect 34300 42438 34356 42476
rect 34748 42530 34804 42542
rect 34972 42532 35028 42542
rect 34748 42478 34750 42530
rect 34802 42478 34804 42530
rect 34524 42308 34580 42318
rect 34524 42196 34580 42252
rect 34524 42194 34692 42196
rect 34524 42142 34526 42194
rect 34578 42142 34692 42194
rect 34524 42140 34692 42142
rect 34524 42130 34580 42140
rect 34300 42082 34356 42094
rect 34300 42030 34302 42082
rect 34354 42030 34356 42082
rect 33964 41970 34020 41982
rect 33964 41918 33966 41970
rect 34018 41918 34020 41970
rect 33852 41860 33908 41870
rect 33852 41300 33908 41804
rect 33852 41186 33908 41244
rect 33852 41134 33854 41186
rect 33906 41134 33908 41186
rect 33852 41122 33908 41134
rect 33852 40964 33908 40974
rect 33740 40908 33852 40964
rect 33852 40898 33908 40908
rect 33516 40562 33572 40572
rect 33628 40516 33684 40526
rect 33516 40404 33572 40414
rect 33404 40402 33572 40404
rect 33404 40350 33518 40402
rect 33570 40350 33572 40402
rect 33404 40348 33572 40350
rect 32396 39566 32398 39618
rect 32450 39566 32452 39618
rect 32396 39396 32452 39566
rect 32396 39330 32452 39340
rect 33292 39284 33348 39676
rect 33292 39218 33348 39228
rect 33516 39284 33572 40348
rect 33516 39218 33572 39228
rect 33068 39060 33124 39070
rect 32284 39058 33124 39060
rect 32284 39006 33070 39058
rect 33122 39006 33124 39058
rect 32284 39004 33124 39006
rect 32284 38946 32340 39004
rect 33068 38994 33124 39004
rect 33180 39060 33236 39070
rect 33180 38966 33236 39004
rect 33292 39060 33348 39070
rect 33628 39060 33684 40460
rect 33964 40516 34020 41918
rect 34300 40852 34356 42030
rect 33292 39058 33684 39060
rect 33292 39006 33294 39058
rect 33346 39006 33684 39058
rect 33292 39004 33684 39006
rect 33740 39396 33796 39406
rect 33292 38994 33348 39004
rect 32284 38894 32286 38946
rect 32338 38894 32340 38946
rect 32284 38882 32340 38894
rect 31948 38220 32228 38276
rect 33068 38836 33124 38846
rect 31388 38164 31444 38174
rect 31276 38162 31444 38164
rect 31276 38110 31390 38162
rect 31442 38110 31444 38162
rect 31276 38108 31444 38110
rect 31388 38098 31444 38108
rect 31276 36484 31332 36494
rect 31220 36482 31332 36484
rect 31220 36430 31278 36482
rect 31330 36430 31332 36482
rect 31220 36428 31332 36430
rect 31164 36390 31220 36428
rect 31276 36418 31332 36428
rect 31948 36260 32004 38220
rect 33068 38162 33124 38780
rect 33740 38834 33796 39340
rect 33964 39172 34020 40460
rect 34076 40796 34356 40852
rect 34412 41858 34468 41870
rect 34412 41806 34414 41858
rect 34466 41806 34468 41858
rect 34076 39732 34132 40796
rect 34188 40626 34244 40638
rect 34188 40574 34190 40626
rect 34242 40574 34244 40626
rect 34188 39844 34244 40574
rect 34412 40628 34468 41806
rect 34412 40562 34468 40572
rect 34524 41748 34580 41758
rect 34524 40402 34580 41692
rect 34636 40740 34692 42140
rect 34748 42084 34804 42478
rect 34748 42018 34804 42028
rect 34860 42530 35028 42532
rect 34860 42478 34974 42530
rect 35026 42478 35028 42530
rect 34860 42476 35028 42478
rect 34860 42082 34916 42476
rect 34972 42466 35028 42476
rect 35084 42308 35140 43372
rect 35196 43362 35252 43372
rect 35196 43148 35460 43158
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35196 43082 35460 43092
rect 36204 42868 36260 43484
rect 36540 43538 36596 43550
rect 36540 43486 36542 43538
rect 36594 43486 36596 43538
rect 36316 42868 36372 42878
rect 36204 42866 36372 42868
rect 36204 42814 36318 42866
rect 36370 42814 36372 42866
rect 36204 42812 36372 42814
rect 36316 42802 36372 42812
rect 34972 42252 35140 42308
rect 36316 42532 36372 42542
rect 34972 42194 35028 42252
rect 34972 42142 34974 42194
rect 35026 42142 35028 42194
rect 34972 42130 35028 42142
rect 34860 42030 34862 42082
rect 34914 42030 34916 42082
rect 34860 42018 34916 42030
rect 35196 41972 35252 41982
rect 35196 41878 35252 41916
rect 35532 41970 35588 41982
rect 35532 41918 35534 41970
rect 35586 41918 35588 41970
rect 35196 41580 35460 41590
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35196 41514 35460 41524
rect 35308 41300 35364 41310
rect 35532 41300 35588 41918
rect 36316 41970 36372 42476
rect 36316 41918 36318 41970
rect 36370 41918 36372 41970
rect 36316 41906 36372 41918
rect 36540 41748 36596 43486
rect 36764 41860 36820 45836
rect 37100 45890 37156 46956
rect 37100 45838 37102 45890
rect 37154 45838 37156 45890
rect 37100 45826 37156 45838
rect 37212 46116 37268 46126
rect 37212 44434 37268 46060
rect 37212 44382 37214 44434
rect 37266 44382 37268 44434
rect 37212 44370 37268 44382
rect 36988 43652 37044 43662
rect 36876 43540 36932 43550
rect 36876 43446 36932 43484
rect 36988 42754 37044 43596
rect 37324 43652 37380 48748
rect 37772 48802 37828 49084
rect 37772 48750 37774 48802
rect 37826 48750 37828 48802
rect 37548 47684 37604 47694
rect 37548 47590 37604 47628
rect 37548 47460 37604 47470
rect 37772 47460 37828 48750
rect 38332 49028 38388 49038
rect 37548 47458 37828 47460
rect 37548 47406 37550 47458
rect 37602 47406 37828 47458
rect 37548 47404 37828 47406
rect 38220 47460 38276 47470
rect 38332 47460 38388 48972
rect 38444 48130 38500 48142
rect 38444 48078 38446 48130
rect 38498 48078 38500 48130
rect 38444 47684 38500 48078
rect 38444 47618 38500 47628
rect 38220 47458 38388 47460
rect 38220 47406 38222 47458
rect 38274 47406 38388 47458
rect 38220 47404 38388 47406
rect 37548 47394 37604 47404
rect 38220 47012 38276 47404
rect 38220 46946 38276 46956
rect 38556 46788 38612 51996
rect 39228 51828 39284 53452
rect 39452 53284 39508 53294
rect 39452 53170 39508 53228
rect 39452 53118 39454 53170
rect 39506 53118 39508 53170
rect 39452 53106 39508 53118
rect 39676 52386 39732 53676
rect 39788 53172 39844 55412
rect 39900 55188 39956 55198
rect 39900 55186 40292 55188
rect 39900 55134 39902 55186
rect 39954 55134 40292 55186
rect 39900 55132 40292 55134
rect 39900 55122 39956 55132
rect 40236 54738 40292 55132
rect 40236 54686 40238 54738
rect 40290 54686 40292 54738
rect 40236 54674 40292 54686
rect 40460 55076 40516 55086
rect 39788 53106 39844 53116
rect 40012 54516 40068 54526
rect 40012 52946 40068 54460
rect 40348 54402 40404 54414
rect 40348 54350 40350 54402
rect 40402 54350 40404 54402
rect 40012 52894 40014 52946
rect 40066 52894 40068 52946
rect 40012 52882 40068 52894
rect 40124 53732 40180 53742
rect 39676 52334 39678 52386
rect 39730 52334 39732 52386
rect 39676 52322 39732 52334
rect 39788 52052 39844 52062
rect 39788 52050 40068 52052
rect 39788 51998 39790 52050
rect 39842 51998 40068 52050
rect 39788 51996 40068 51998
rect 39788 51986 39844 51996
rect 38892 51772 39284 51828
rect 38780 51268 38836 51278
rect 38780 51174 38836 51212
rect 38668 51154 38724 51166
rect 38668 51102 38670 51154
rect 38722 51102 38724 51154
rect 38668 50706 38724 51102
rect 38668 50654 38670 50706
rect 38722 50654 38724 50706
rect 38668 50642 38724 50654
rect 38668 49698 38724 49710
rect 38668 49646 38670 49698
rect 38722 49646 38724 49698
rect 38668 49588 38724 49646
rect 38668 49522 38724 49532
rect 38892 49028 38948 51772
rect 39340 51716 39396 51726
rect 39228 51604 39284 51614
rect 39228 50820 39284 51548
rect 39228 50754 39284 50764
rect 39340 51602 39396 51660
rect 39340 51550 39342 51602
rect 39394 51550 39396 51602
rect 39228 50036 39284 50046
rect 39340 50036 39396 51550
rect 40012 51604 40068 51996
rect 40124 51828 40180 53676
rect 40236 53620 40292 53630
rect 40236 52050 40292 53564
rect 40236 51998 40238 52050
rect 40290 51998 40292 52050
rect 40236 51986 40292 51998
rect 40348 51938 40404 54350
rect 40348 51886 40350 51938
rect 40402 51886 40404 51938
rect 40348 51874 40404 51886
rect 40460 52162 40516 55020
rect 41132 54740 41188 56028
rect 41244 55468 41300 59200
rect 42812 57428 42868 59200
rect 44380 59108 44436 59200
rect 44716 59108 44772 59276
rect 44380 59052 44772 59108
rect 42812 57372 43428 57428
rect 42812 56194 42868 56206
rect 42812 56142 42814 56194
rect 42866 56142 42868 56194
rect 41244 55412 41412 55468
rect 41244 54740 41300 54750
rect 41132 54738 41300 54740
rect 41132 54686 41246 54738
rect 41298 54686 41300 54738
rect 41132 54684 41300 54686
rect 41244 54674 41300 54684
rect 41020 54628 41076 54638
rect 41020 54534 41076 54572
rect 40908 54514 40964 54526
rect 40908 54462 40910 54514
rect 40962 54462 40964 54514
rect 40908 53396 40964 54462
rect 41356 54180 41412 55412
rect 41468 55412 41524 55422
rect 41468 54404 41524 55356
rect 42028 55410 42084 55422
rect 42028 55358 42030 55410
rect 42082 55358 42084 55410
rect 42028 55188 42084 55358
rect 42700 55298 42756 55310
rect 42700 55246 42702 55298
rect 42754 55246 42756 55298
rect 42364 55188 42420 55198
rect 42028 55132 42364 55188
rect 42364 55122 42420 55132
rect 42476 55074 42532 55086
rect 42476 55022 42478 55074
rect 42530 55022 42532 55074
rect 42364 54852 42420 54862
rect 41468 54310 41524 54348
rect 42140 54796 42364 54852
rect 41356 54124 41524 54180
rect 41356 53844 41412 53854
rect 40908 53330 40964 53340
rect 41244 53842 41412 53844
rect 41244 53790 41358 53842
rect 41410 53790 41412 53842
rect 41244 53788 41412 53790
rect 41244 52164 41300 53788
rect 41356 53778 41412 53788
rect 41468 53508 41524 54124
rect 41692 53730 41748 53742
rect 41692 53678 41694 53730
rect 41746 53678 41748 53730
rect 41692 53620 41748 53678
rect 41692 53554 41748 53564
rect 41468 53442 41524 53452
rect 41916 53172 41972 53182
rect 41916 53078 41972 53116
rect 40460 52110 40462 52162
rect 40514 52110 40516 52162
rect 40124 51772 40292 51828
rect 40124 51604 40180 51614
rect 40012 51602 40180 51604
rect 40012 51550 40126 51602
rect 40178 51550 40180 51602
rect 40012 51548 40180 51550
rect 40124 51538 40180 51548
rect 39228 50034 39396 50036
rect 39228 49982 39230 50034
rect 39282 49982 39396 50034
rect 39228 49980 39396 49982
rect 39452 51378 39508 51390
rect 39452 51326 39454 51378
rect 39506 51326 39508 51378
rect 39228 49970 39284 49980
rect 38780 48972 38948 49028
rect 39004 49812 39060 49822
rect 39004 49140 39060 49756
rect 39116 49810 39172 49822
rect 39116 49758 39118 49810
rect 39170 49758 39172 49810
rect 39116 49588 39172 49758
rect 39452 49812 39508 51326
rect 39788 51380 39844 51390
rect 39788 51286 39844 51324
rect 39676 51268 39732 51278
rect 39676 50036 39732 51212
rect 40124 51266 40180 51278
rect 40124 51214 40126 51266
rect 40178 51214 40180 51266
rect 40124 50372 40180 51214
rect 40012 50316 40124 50372
rect 39788 50036 39844 50046
rect 39676 50034 39844 50036
rect 39676 49982 39790 50034
rect 39842 49982 39844 50034
rect 39676 49980 39844 49982
rect 39788 49970 39844 49980
rect 39452 49810 39620 49812
rect 39452 49758 39454 49810
rect 39506 49758 39620 49810
rect 39452 49756 39620 49758
rect 39452 49746 39508 49756
rect 39116 49522 39172 49532
rect 39452 49476 39508 49486
rect 39452 49140 39508 49420
rect 38780 47012 38836 48972
rect 38892 48020 38948 48030
rect 38892 47570 38948 47964
rect 38892 47518 38894 47570
rect 38946 47518 38948 47570
rect 38892 47506 38948 47518
rect 38780 46898 38836 46956
rect 38780 46846 38782 46898
rect 38834 46846 38836 46898
rect 38780 46834 38836 46846
rect 38332 46732 38612 46788
rect 37772 45780 37828 45790
rect 37772 45778 38052 45780
rect 37772 45726 37774 45778
rect 37826 45726 38052 45778
rect 37772 45724 38052 45726
rect 37772 45714 37828 45724
rect 37996 44548 38052 45724
rect 38332 45220 38388 46732
rect 38892 46676 38948 46686
rect 38668 46674 38948 46676
rect 38668 46622 38894 46674
rect 38946 46622 38948 46674
rect 38668 46620 38948 46622
rect 38556 46564 38612 46574
rect 38332 45154 38388 45164
rect 38444 46508 38556 46564
rect 38108 45108 38164 45118
rect 38108 44994 38164 45052
rect 38108 44942 38110 44994
rect 38162 44942 38164 44994
rect 38108 44930 38164 44942
rect 38220 44996 38276 45006
rect 38444 44996 38500 46508
rect 38556 46498 38612 46508
rect 38668 45332 38724 46620
rect 38892 46610 38948 46620
rect 39004 45444 39060 49084
rect 39228 49138 39508 49140
rect 39228 49086 39454 49138
rect 39506 49086 39508 49138
rect 39228 49084 39508 49086
rect 39228 48244 39284 49084
rect 39452 49074 39508 49084
rect 39564 48356 39620 49756
rect 39116 48242 39284 48244
rect 39116 48190 39230 48242
rect 39282 48190 39284 48242
rect 39116 48188 39284 48190
rect 39116 46564 39172 48188
rect 39228 48178 39284 48188
rect 39340 48300 39620 48356
rect 39788 49810 39844 49822
rect 39788 49758 39790 49810
rect 39842 49758 39844 49810
rect 39340 47684 39396 48300
rect 39676 48130 39732 48142
rect 39676 48078 39678 48130
rect 39730 48078 39732 48130
rect 39564 48020 39620 48030
rect 39564 47926 39620 47964
rect 39228 47628 39396 47684
rect 39228 46900 39284 47628
rect 39564 47460 39620 47470
rect 39228 46844 39508 46900
rect 39228 46674 39284 46844
rect 39228 46622 39230 46674
rect 39282 46622 39284 46674
rect 39228 46610 39284 46622
rect 39340 46674 39396 46686
rect 39340 46622 39342 46674
rect 39394 46622 39396 46674
rect 39116 46498 39172 46508
rect 39228 46340 39284 46350
rect 39228 45892 39284 46284
rect 39340 46004 39396 46622
rect 39452 46116 39508 46844
rect 39564 46562 39620 47404
rect 39676 46898 39732 48078
rect 39676 46846 39678 46898
rect 39730 46846 39732 46898
rect 39676 46834 39732 46846
rect 39788 47572 39844 49758
rect 40012 49810 40068 50316
rect 40124 50306 40180 50316
rect 40012 49758 40014 49810
rect 40066 49758 40068 49810
rect 40012 49746 40068 49758
rect 40124 49140 40180 49150
rect 40236 49140 40292 51772
rect 40460 51716 40516 52110
rect 40460 51650 40516 51660
rect 40572 52162 41300 52164
rect 40572 52110 41246 52162
rect 41298 52110 41300 52162
rect 40572 52108 41300 52110
rect 40460 51268 40516 51278
rect 40572 51268 40628 52108
rect 41244 52098 41300 52108
rect 41356 52946 41412 52958
rect 41356 52894 41358 52946
rect 41410 52894 41412 52946
rect 41356 51604 41412 52894
rect 41692 52276 41748 52286
rect 41692 52162 41748 52220
rect 41692 52110 41694 52162
rect 41746 52110 41748 52162
rect 41692 52098 41748 52110
rect 42140 52050 42196 54796
rect 42364 54786 42420 54796
rect 42476 54516 42532 55022
rect 42588 55076 42644 55086
rect 42588 54982 42644 55020
rect 42476 54450 42532 54460
rect 42140 51998 42142 52050
rect 42194 51998 42196 52050
rect 41468 51716 41524 51726
rect 41524 51660 41636 51716
rect 41468 51650 41524 51660
rect 41356 51538 41412 51548
rect 41244 51492 41300 51502
rect 41244 51398 41300 51436
rect 40460 51266 40628 51268
rect 40460 51214 40462 51266
rect 40514 51214 40628 51266
rect 40460 51212 40628 51214
rect 40796 51380 40852 51390
rect 41468 51380 41524 51390
rect 40460 51202 40516 51212
rect 40796 50708 40852 51324
rect 40348 50706 40852 50708
rect 40348 50654 40798 50706
rect 40850 50654 40852 50706
rect 40348 50652 40852 50654
rect 40348 49698 40404 50652
rect 40796 50642 40852 50652
rect 41356 51378 41524 51380
rect 41356 51326 41470 51378
rect 41522 51326 41524 51378
rect 41356 51324 41524 51326
rect 40348 49646 40350 49698
rect 40402 49646 40404 49698
rect 40348 49634 40404 49646
rect 40460 50484 40516 50494
rect 40124 49138 40236 49140
rect 40124 49086 40126 49138
rect 40178 49086 40236 49138
rect 40124 49084 40236 49086
rect 40124 49074 40180 49084
rect 40236 49046 40292 49084
rect 40012 48356 40068 48366
rect 40068 48300 40180 48356
rect 40012 48262 40068 48300
rect 39788 46676 39844 47516
rect 39900 46676 39956 46686
rect 39788 46674 39956 46676
rect 39788 46622 39902 46674
rect 39954 46622 39956 46674
rect 39788 46620 39956 46622
rect 39900 46610 39956 46620
rect 39564 46510 39566 46562
rect 39618 46510 39620 46562
rect 39564 46340 39620 46510
rect 39564 46274 39620 46284
rect 39788 46172 40068 46228
rect 39788 46116 39844 46172
rect 39452 46060 39844 46116
rect 39900 46004 39956 46014
rect 39340 46002 39956 46004
rect 39340 45950 39902 46002
rect 39954 45950 39956 46002
rect 39340 45948 39956 45950
rect 39228 45836 39508 45892
rect 39004 45388 39396 45444
rect 38668 45238 38724 45276
rect 38556 45220 38612 45230
rect 38556 45126 38612 45164
rect 38780 45220 38836 45230
rect 38780 45106 38836 45164
rect 39116 45108 39172 45118
rect 38780 45054 38782 45106
rect 38834 45054 38836 45106
rect 38780 45042 38836 45054
rect 38892 45052 39116 45108
rect 38444 44940 38724 44996
rect 38108 44548 38164 44558
rect 37996 44546 38164 44548
rect 37996 44494 38110 44546
rect 38162 44494 38164 44546
rect 37996 44492 38164 44494
rect 38108 44482 38164 44492
rect 38220 44434 38276 44940
rect 38220 44382 38222 44434
rect 38274 44382 38276 44434
rect 38220 44370 38276 44382
rect 38668 44434 38724 44940
rect 38668 44382 38670 44434
rect 38722 44382 38724 44434
rect 38668 44370 38724 44382
rect 37548 43764 37604 43774
rect 37324 43558 37380 43596
rect 37436 43708 37548 43764
rect 36988 42702 36990 42754
rect 37042 42702 37044 42754
rect 36988 42690 37044 42702
rect 37100 42532 37156 42542
rect 37100 42438 37156 42476
rect 37212 42530 37268 42542
rect 37212 42478 37214 42530
rect 37266 42478 37268 42530
rect 37212 42196 37268 42478
rect 37212 42130 37268 42140
rect 36764 41794 36820 41804
rect 36540 41682 36596 41692
rect 35308 41298 35588 41300
rect 35308 41246 35310 41298
rect 35362 41246 35588 41298
rect 35308 41244 35588 41246
rect 37212 41412 37268 41422
rect 34636 40674 34692 40684
rect 34972 40964 35028 40974
rect 34524 40350 34526 40402
rect 34578 40350 34580 40402
rect 34524 40338 34580 40350
rect 34748 40516 34804 40526
rect 34188 39778 34244 39788
rect 34076 39666 34132 39676
rect 33964 39116 34244 39172
rect 33740 38782 33742 38834
rect 33794 38782 33796 38834
rect 33740 38668 33796 38782
rect 33964 38948 34020 38958
rect 33740 38612 33908 38668
rect 33068 38110 33070 38162
rect 33122 38110 33124 38162
rect 33068 38098 33124 38110
rect 32172 38050 32228 38062
rect 32172 37998 32174 38050
rect 32226 37998 32228 38050
rect 32172 37268 32228 37998
rect 32396 38052 32452 38062
rect 33628 38052 33684 38062
rect 32396 37958 32452 37996
rect 33292 37996 33628 38052
rect 33068 37828 33124 37838
rect 32172 37202 32228 37212
rect 32508 37268 32564 37278
rect 32508 37174 32564 37212
rect 32956 37266 33012 37278
rect 32956 37214 32958 37266
rect 33010 37214 33012 37266
rect 32956 37044 33012 37214
rect 32956 36978 33012 36988
rect 32172 36596 32228 36606
rect 32060 36540 32172 36596
rect 32060 36482 32116 36540
rect 32172 36530 32228 36540
rect 32060 36430 32062 36482
rect 32114 36430 32116 36482
rect 32060 36418 32116 36430
rect 31948 36204 32228 36260
rect 31164 35700 31220 35710
rect 31500 35700 31556 35710
rect 30828 35644 31164 35700
rect 30828 35586 30884 35644
rect 31164 35606 31220 35644
rect 31276 35698 31556 35700
rect 31276 35646 31502 35698
rect 31554 35646 31556 35698
rect 31276 35644 31556 35646
rect 30828 35534 30830 35586
rect 30882 35534 30884 35586
rect 30828 35522 30884 35534
rect 30828 34916 30884 34926
rect 30828 34244 30884 34860
rect 31052 34802 31108 34814
rect 31052 34750 31054 34802
rect 31106 34750 31108 34802
rect 31052 34354 31108 34750
rect 31052 34302 31054 34354
rect 31106 34302 31108 34354
rect 31052 34290 31108 34302
rect 31276 34356 31332 35644
rect 31500 35634 31556 35644
rect 31724 35700 31780 35710
rect 31724 35698 31892 35700
rect 31724 35646 31726 35698
rect 31778 35646 31892 35698
rect 31724 35644 31892 35646
rect 31724 35634 31780 35644
rect 30828 34130 30884 34188
rect 31276 34242 31332 34300
rect 31612 35586 31668 35598
rect 31612 35534 31614 35586
rect 31666 35534 31668 35586
rect 31276 34190 31278 34242
rect 31330 34190 31332 34242
rect 31276 34178 31332 34190
rect 31500 34244 31556 34254
rect 31612 34244 31668 35534
rect 31500 34242 31668 34244
rect 31500 34190 31502 34242
rect 31554 34190 31668 34242
rect 31500 34188 31668 34190
rect 31836 34244 31892 35644
rect 31948 34356 32004 34366
rect 31948 34262 32004 34300
rect 31500 34178 31556 34188
rect 31836 34150 31892 34188
rect 30828 34078 30830 34130
rect 30882 34078 30884 34130
rect 30828 34066 30884 34078
rect 30828 33908 30884 33918
rect 30828 33570 30884 33852
rect 30828 33518 30830 33570
rect 30882 33518 30884 33570
rect 30828 33506 30884 33518
rect 31052 33908 31108 33918
rect 31052 33346 31108 33852
rect 31948 33908 32004 33918
rect 31948 33814 32004 33852
rect 31052 33294 31054 33346
rect 31106 33294 31108 33346
rect 31052 32562 31108 33294
rect 31052 32510 31054 32562
rect 31106 32510 31108 32562
rect 31052 32498 31108 32510
rect 31164 33460 31220 33470
rect 30940 31780 30996 31790
rect 30940 31218 30996 31724
rect 30940 31166 30942 31218
rect 30994 31166 30996 31218
rect 30940 31154 30996 31166
rect 31164 31444 31220 33404
rect 31836 33122 31892 33134
rect 31836 33070 31838 33122
rect 31890 33070 31892 33122
rect 31836 32676 31892 33070
rect 31836 32610 31892 32620
rect 31724 32452 31780 32462
rect 32060 32452 32116 32462
rect 31724 32450 32116 32452
rect 31724 32398 31726 32450
rect 31778 32398 32062 32450
rect 32114 32398 32116 32450
rect 31724 32396 32116 32398
rect 31724 32386 31780 32396
rect 32060 32386 32116 32396
rect 32172 32228 32228 36204
rect 33068 34242 33124 37772
rect 33292 37266 33348 37996
rect 33628 37958 33684 37996
rect 33292 37214 33294 37266
rect 33346 37214 33348 37266
rect 33292 37202 33348 37214
rect 33404 37828 33460 37838
rect 33180 37154 33236 37166
rect 33180 37102 33182 37154
rect 33234 37102 33236 37154
rect 33180 36596 33236 37102
rect 33404 37044 33460 37772
rect 33516 37826 33572 37838
rect 33516 37774 33518 37826
rect 33570 37774 33572 37826
rect 33516 37604 33572 37774
rect 33852 37826 33908 38612
rect 33852 37774 33854 37826
rect 33906 37774 33908 37826
rect 33516 37548 33684 37604
rect 33628 37378 33684 37548
rect 33628 37326 33630 37378
rect 33682 37326 33684 37378
rect 33628 37314 33684 37326
rect 33404 36978 33460 36988
rect 33852 37268 33908 37774
rect 33964 37828 34020 38892
rect 33964 37762 34020 37772
rect 34076 38946 34132 38958
rect 34076 38894 34078 38946
rect 34130 38894 34132 38946
rect 34076 38052 34132 38894
rect 34188 38668 34244 39116
rect 34300 38836 34356 38846
rect 34300 38834 34468 38836
rect 34300 38782 34302 38834
rect 34354 38782 34468 38834
rect 34300 38780 34468 38782
rect 34300 38770 34356 38780
rect 34188 38612 34356 38668
rect 33180 36530 33236 36540
rect 33628 36484 33684 36494
rect 33628 35588 33684 36428
rect 33180 35026 33236 35038
rect 33180 34974 33182 35026
rect 33234 34974 33236 35026
rect 33180 34356 33236 34974
rect 33180 34290 33236 34300
rect 33628 35026 33684 35532
rect 33628 34974 33630 35026
rect 33682 34974 33684 35026
rect 33068 34190 33070 34242
rect 33122 34190 33124 34242
rect 33068 34178 33124 34190
rect 33292 34132 33348 34142
rect 32508 33684 32564 33694
rect 32284 33348 32340 33358
rect 32284 33254 32340 33292
rect 32396 32564 32452 32574
rect 32396 32470 32452 32508
rect 30716 31052 30884 31108
rect 30380 29538 30436 29596
rect 30604 29540 30660 31052
rect 30380 29486 30382 29538
rect 30434 29486 30436 29538
rect 30380 29474 30436 29486
rect 30492 29538 30660 29540
rect 30492 29486 30606 29538
rect 30658 29486 30660 29538
rect 30492 29484 30660 29486
rect 30156 28914 30212 28924
rect 30380 29316 30436 29326
rect 30380 28756 30436 29260
rect 29820 28478 29822 28530
rect 29874 28478 29876 28530
rect 29820 28466 29876 28478
rect 30156 28532 30212 28542
rect 30156 28438 30212 28476
rect 30156 28084 30212 28094
rect 29708 27860 29764 27870
rect 29708 27766 29764 27804
rect 29708 27300 29764 27310
rect 29596 27298 29764 27300
rect 29596 27246 29710 27298
rect 29762 27246 29764 27298
rect 29596 27244 29764 27246
rect 29372 27234 29428 27244
rect 29708 27234 29764 27244
rect 29148 27076 29204 27086
rect 29148 26982 29204 27020
rect 29260 26292 29316 26302
rect 29260 26198 29316 26236
rect 29932 26178 29988 26190
rect 29932 26126 29934 26178
rect 29986 26126 29988 26178
rect 29932 25618 29988 26126
rect 29932 25566 29934 25618
rect 29986 25566 29988 25618
rect 29932 25554 29988 25566
rect 30044 26068 30100 26078
rect 29820 25394 29876 25406
rect 29820 25342 29822 25394
rect 29874 25342 29876 25394
rect 29708 24834 29764 24846
rect 29708 24782 29710 24834
rect 29762 24782 29764 24834
rect 29036 24610 29092 24668
rect 29596 24724 29652 24734
rect 29036 24558 29038 24610
rect 29090 24558 29092 24610
rect 29036 24546 29092 24558
rect 29260 24612 29316 24622
rect 29260 23938 29316 24556
rect 29260 23886 29262 23938
rect 29314 23886 29316 23938
rect 29260 23874 29316 23886
rect 29148 23714 29204 23726
rect 29148 23662 29150 23714
rect 29202 23662 29204 23714
rect 29148 23548 29204 23662
rect 29148 23492 29316 23548
rect 29036 23044 29092 23054
rect 29036 22950 29092 22988
rect 29260 22708 29316 23492
rect 29596 23492 29652 24668
rect 29708 24612 29764 24782
rect 29708 24546 29764 24556
rect 29708 24164 29764 24174
rect 29820 24164 29876 25342
rect 29932 25394 29988 25406
rect 29932 25342 29934 25394
rect 29986 25342 29988 25394
rect 29932 24946 29988 25342
rect 30044 25394 30100 26012
rect 30044 25342 30046 25394
rect 30098 25342 30100 25394
rect 30044 25330 30100 25342
rect 29932 24894 29934 24946
rect 29986 24894 29988 24946
rect 29932 24882 29988 24894
rect 29764 24108 29876 24164
rect 29708 24050 29764 24108
rect 29708 23998 29710 24050
rect 29762 23998 29764 24050
rect 29708 23986 29764 23998
rect 30044 23714 30100 23726
rect 30044 23662 30046 23714
rect 30098 23662 30100 23714
rect 30044 23492 30100 23662
rect 29596 23436 30100 23492
rect 29148 22652 29316 22708
rect 29484 23044 29540 23054
rect 29148 22484 29204 22652
rect 29372 22596 29428 22606
rect 29148 21810 29204 22428
rect 29148 21758 29150 21810
rect 29202 21758 29204 21810
rect 29148 21746 29204 21758
rect 29260 22540 29372 22596
rect 29260 20916 29316 22540
rect 29372 22530 29428 22540
rect 29484 22482 29540 22988
rect 29484 22430 29486 22482
rect 29538 22430 29540 22482
rect 29484 22418 29540 22430
rect 29372 22260 29428 22270
rect 29596 22260 29652 23436
rect 30156 23044 30212 28028
rect 30380 27746 30436 28700
rect 30380 27694 30382 27746
rect 30434 27694 30436 27746
rect 30380 27682 30436 27694
rect 30492 26628 30548 29484
rect 30604 29474 30660 29484
rect 30604 28644 30660 28654
rect 30604 28550 30660 28588
rect 30716 27860 30772 27870
rect 30716 27074 30772 27804
rect 30716 27022 30718 27074
rect 30770 27022 30772 27074
rect 30716 27010 30772 27022
rect 30828 26908 30884 31052
rect 31164 30324 31220 31388
rect 32060 32172 32228 32228
rect 32284 32450 32340 32462
rect 32284 32398 32286 32450
rect 32338 32398 32340 32450
rect 31388 31332 31444 31342
rect 31276 31276 31388 31332
rect 31276 31106 31332 31276
rect 31388 31266 31444 31276
rect 31612 31108 31668 31118
rect 31276 31054 31278 31106
rect 31330 31054 31332 31106
rect 31276 31042 31332 31054
rect 31388 31106 31668 31108
rect 31388 31054 31614 31106
rect 31666 31054 31668 31106
rect 31388 31052 31668 31054
rect 31164 30258 31220 30268
rect 31276 30100 31332 30110
rect 30940 29986 30996 29998
rect 30940 29934 30942 29986
rect 30994 29934 30996 29986
rect 30940 29428 30996 29934
rect 31052 29988 31108 29998
rect 31052 29894 31108 29932
rect 31164 29986 31220 29998
rect 31164 29934 31166 29986
rect 31218 29934 31220 29986
rect 30940 29362 30996 29372
rect 31052 29652 31108 29662
rect 30940 29204 30996 29214
rect 30940 28530 30996 29148
rect 30940 28478 30942 28530
rect 30994 28478 30996 28530
rect 30940 28466 30996 28478
rect 31052 27524 31108 29596
rect 31164 29540 31220 29934
rect 31164 29474 31220 29484
rect 31276 29538 31332 30044
rect 31276 29486 31278 29538
rect 31330 29486 31332 29538
rect 31276 29474 31332 29486
rect 31388 29316 31444 31052
rect 31612 31042 31668 31052
rect 31836 30994 31892 31006
rect 31836 30942 31838 30994
rect 31890 30942 31892 30994
rect 31500 30324 31556 30334
rect 31500 30210 31556 30268
rect 31500 30158 31502 30210
rect 31554 30158 31556 30210
rect 31500 30146 31556 30158
rect 31836 29652 31892 30942
rect 31836 29586 31892 29596
rect 31948 30212 32004 30222
rect 31612 29426 31668 29438
rect 31612 29374 31614 29426
rect 31666 29374 31668 29426
rect 31164 29260 31444 29316
rect 31500 29316 31556 29326
rect 31164 27748 31220 29260
rect 31500 29222 31556 29260
rect 31612 28868 31668 29374
rect 31948 29204 32004 30156
rect 31948 29138 32004 29148
rect 32060 29092 32116 32172
rect 32060 29026 32116 29036
rect 32172 32004 32228 32014
rect 31276 28812 31668 28868
rect 31276 28196 31332 28812
rect 32060 28756 32116 28766
rect 32172 28756 32228 31948
rect 32284 31890 32340 32398
rect 32284 31838 32286 31890
rect 32338 31838 32340 31890
rect 32284 31826 32340 31838
rect 32508 31668 32564 33628
rect 33180 33460 33236 33470
rect 33180 33366 33236 33404
rect 32732 33348 32788 33358
rect 32732 33254 32788 33292
rect 33292 32674 33348 34076
rect 33404 33572 33460 33582
rect 33404 32786 33460 33516
rect 33628 33348 33684 34974
rect 33852 34244 33908 37212
rect 34076 36596 34132 37996
rect 34300 37938 34356 38612
rect 34412 38052 34468 38780
rect 34748 38722 34804 40460
rect 34748 38670 34750 38722
rect 34802 38670 34804 38722
rect 34748 38658 34804 38670
rect 34860 38162 34916 38174
rect 34860 38110 34862 38162
rect 34914 38110 34916 38162
rect 34748 38052 34804 38062
rect 34412 38050 34804 38052
rect 34412 37998 34750 38050
rect 34802 37998 34804 38050
rect 34412 37996 34804 37998
rect 34300 37886 34302 37938
rect 34354 37886 34356 37938
rect 34300 37874 34356 37886
rect 34636 37378 34692 37390
rect 34636 37326 34638 37378
rect 34690 37326 34692 37378
rect 34524 37156 34580 37166
rect 34524 36706 34580 37100
rect 34524 36654 34526 36706
rect 34578 36654 34580 36706
rect 34524 36642 34580 36654
rect 34188 36596 34244 36606
rect 34076 36594 34244 36596
rect 34076 36542 34190 36594
rect 34242 36542 34244 36594
rect 34076 36540 34244 36542
rect 34188 36530 34244 36540
rect 34636 36372 34692 37326
rect 34748 37266 34804 37996
rect 34748 37214 34750 37266
rect 34802 37214 34804 37266
rect 34748 37202 34804 37214
rect 34860 36706 34916 38110
rect 34860 36654 34862 36706
rect 34914 36654 34916 36706
rect 34860 36642 34916 36654
rect 34748 36372 34804 36382
rect 34636 36316 34748 36372
rect 34748 36278 34804 36316
rect 34412 35588 34468 35598
rect 34412 35494 34468 35532
rect 33852 34178 33908 34188
rect 34860 34242 34916 34254
rect 34860 34190 34862 34242
rect 34914 34190 34916 34242
rect 33404 32734 33406 32786
rect 33458 32734 33460 32786
rect 33404 32722 33460 32734
rect 33516 33346 33684 33348
rect 33516 33294 33630 33346
rect 33682 33294 33684 33346
rect 33516 33292 33684 33294
rect 33292 32622 33294 32674
rect 33346 32622 33348 32674
rect 33292 32610 33348 32622
rect 33404 32340 33460 32350
rect 33404 32246 33460 32284
rect 33180 32004 33236 32014
rect 33404 32004 33460 32014
rect 33236 32002 33460 32004
rect 33236 31950 33406 32002
rect 33458 31950 33460 32002
rect 33236 31948 33460 31950
rect 33180 31938 33236 31948
rect 33404 31938 33460 31948
rect 33516 32004 33572 33292
rect 33628 33282 33684 33292
rect 33740 34130 33796 34142
rect 33740 34078 33742 34130
rect 33794 34078 33796 34130
rect 33740 33348 33796 34078
rect 34524 34132 34580 34142
rect 34524 34038 34580 34076
rect 34748 34130 34804 34142
rect 34748 34078 34750 34130
rect 34802 34078 34804 34130
rect 33852 34018 33908 34030
rect 33852 33966 33854 34018
rect 33906 33966 33908 34018
rect 33852 33684 33908 33966
rect 33852 33628 34020 33684
rect 33740 32788 33796 33292
rect 33740 32722 33796 32732
rect 33852 33460 33908 33470
rect 33852 32674 33908 33404
rect 33964 33348 34020 33628
rect 34748 33460 34804 34078
rect 34748 33394 34804 33404
rect 33964 33282 34020 33292
rect 34300 33236 34356 33246
rect 34300 33234 34692 33236
rect 34300 33182 34302 33234
rect 34354 33182 34692 33234
rect 34300 33180 34692 33182
rect 34300 33170 34356 33180
rect 34636 32786 34692 33180
rect 34636 32734 34638 32786
rect 34690 32734 34692 32786
rect 34636 32722 34692 32734
rect 33852 32622 33854 32674
rect 33906 32622 33908 32674
rect 33852 32610 33908 32622
rect 34076 32674 34132 32686
rect 34076 32622 34078 32674
rect 34130 32622 34132 32674
rect 33068 31780 33124 31790
rect 33516 31780 33572 31948
rect 33068 31778 33572 31780
rect 33068 31726 33070 31778
rect 33122 31726 33572 31778
rect 33068 31724 33572 31726
rect 33628 32452 33684 32462
rect 33068 31714 33124 31724
rect 32284 31612 32564 31668
rect 32284 29764 32340 31612
rect 33516 31556 33572 31566
rect 33628 31556 33684 32396
rect 34076 32452 34132 32622
rect 34748 32674 34804 32686
rect 34748 32622 34750 32674
rect 34802 32622 34804 32674
rect 34748 32564 34804 32622
rect 34076 32386 34132 32396
rect 34188 32508 34804 32564
rect 34188 32450 34244 32508
rect 34188 32398 34190 32450
rect 34242 32398 34244 32450
rect 34188 32386 34244 32398
rect 34860 32452 34916 34190
rect 34860 32386 34916 32396
rect 34524 32340 34580 32350
rect 34524 32246 34580 32284
rect 34860 32002 34916 32014
rect 34860 31950 34862 32002
rect 34914 31950 34916 32002
rect 34860 31892 34916 31950
rect 34636 31836 34916 31892
rect 33516 31554 33684 31556
rect 33516 31502 33518 31554
rect 33570 31502 33684 31554
rect 33516 31500 33684 31502
rect 33740 31666 33796 31678
rect 33740 31614 33742 31666
rect 33794 31614 33796 31666
rect 32508 31220 32564 31230
rect 32396 31108 32452 31118
rect 32396 31014 32452 31052
rect 32508 31106 32564 31164
rect 32508 31054 32510 31106
rect 32562 31054 32564 31106
rect 32508 31042 32564 31054
rect 33180 30994 33236 31006
rect 33180 30942 33182 30994
rect 33234 30942 33236 30994
rect 33180 30884 33236 30942
rect 33404 30884 33460 30894
rect 32620 30828 33404 30884
rect 32396 30772 32452 30782
rect 32396 30678 32452 30716
rect 32396 30210 32452 30222
rect 32396 30158 32398 30210
rect 32450 30158 32452 30210
rect 32396 30100 32452 30158
rect 32396 30034 32452 30044
rect 32284 29698 32340 29708
rect 32508 29428 32564 29438
rect 32508 29334 32564 29372
rect 32060 28754 32228 28756
rect 32060 28702 32062 28754
rect 32114 28702 32228 28754
rect 32060 28700 32228 28702
rect 32060 28690 32116 28700
rect 31388 28642 31444 28654
rect 31388 28590 31390 28642
rect 31442 28590 31444 28642
rect 31388 28532 31444 28590
rect 32620 28532 32676 30828
rect 33404 30818 33460 30828
rect 33516 30436 33572 31500
rect 33516 30370 33572 30380
rect 33628 30324 33684 30334
rect 33740 30324 33796 31614
rect 34300 31668 34356 31678
rect 34300 31666 34468 31668
rect 34300 31614 34302 31666
rect 34354 31614 34468 31666
rect 34300 31612 34468 31614
rect 34300 31602 34356 31612
rect 33964 31556 34020 31566
rect 33964 31462 34020 31500
rect 34188 31554 34244 31566
rect 34188 31502 34190 31554
rect 34242 31502 34244 31554
rect 34188 31332 34244 31502
rect 34188 31266 34244 31276
rect 33964 31108 34020 31118
rect 33852 30996 33908 31006
rect 33964 30996 34020 31052
rect 33852 30994 34020 30996
rect 33852 30942 33854 30994
rect 33906 30942 34020 30994
rect 33852 30940 34020 30942
rect 33852 30930 33908 30940
rect 33628 30322 33796 30324
rect 33628 30270 33630 30322
rect 33682 30270 33796 30322
rect 33628 30268 33796 30270
rect 33628 30258 33684 30268
rect 32844 30212 32900 30222
rect 32844 30118 32900 30156
rect 33964 30212 34020 30222
rect 34020 30156 34132 30212
rect 33964 30146 34020 30156
rect 33516 29986 33572 29998
rect 33516 29934 33518 29986
rect 33570 29934 33572 29986
rect 33180 29876 33236 29886
rect 33180 29650 33236 29820
rect 33180 29598 33182 29650
rect 33234 29598 33236 29650
rect 33180 29586 33236 29598
rect 33516 29764 33572 29934
rect 32956 29540 33012 29550
rect 32956 29428 33012 29484
rect 31388 28476 32676 28532
rect 31276 28130 31332 28140
rect 31836 27972 31892 27982
rect 31724 27916 31836 27972
rect 31164 27682 31220 27692
rect 31276 27746 31332 27758
rect 31276 27694 31278 27746
rect 31330 27694 31332 27746
rect 31276 27524 31332 27694
rect 31052 27468 31332 27524
rect 31276 27188 31332 27198
rect 31276 27094 31332 27132
rect 31724 27186 31780 27916
rect 31836 27878 31892 27916
rect 32172 27970 32228 27982
rect 32172 27918 32174 27970
rect 32226 27918 32228 27970
rect 32172 27412 32228 27918
rect 32508 27860 32564 27870
rect 32508 27636 32564 27804
rect 32508 27570 32564 27580
rect 32172 27346 32228 27356
rect 31724 27134 31726 27186
rect 31778 27134 31780 27186
rect 31724 27122 31780 27134
rect 32620 27074 32676 28476
rect 32620 27022 32622 27074
rect 32674 27022 32676 27074
rect 30492 26562 30548 26572
rect 30604 26852 30884 26908
rect 32172 26962 32228 26974
rect 32172 26910 32174 26962
rect 32226 26910 32228 26962
rect 30268 25282 30324 25294
rect 30268 25230 30270 25282
rect 30322 25230 30324 25282
rect 30268 24724 30324 25230
rect 30492 24724 30548 24734
rect 30268 24668 30492 24724
rect 30492 24630 30548 24668
rect 30604 24164 30660 26852
rect 32172 26628 32228 26910
rect 32172 26562 32228 26572
rect 32508 26404 32564 26414
rect 32060 26348 32508 26404
rect 30716 26292 30772 26302
rect 30716 25506 30772 26236
rect 32060 26178 32116 26348
rect 32508 26310 32564 26348
rect 32620 26292 32676 27022
rect 32620 26226 32676 26236
rect 32844 29426 33012 29428
rect 32844 29374 32958 29426
rect 33010 29374 33012 29426
rect 32844 29372 33012 29374
rect 32060 26126 32062 26178
rect 32114 26126 32116 26178
rect 32060 26114 32116 26126
rect 32396 26068 32452 26078
rect 32396 25974 32452 26012
rect 30716 25454 30718 25506
rect 30770 25454 30772 25506
rect 30716 25442 30772 25454
rect 31612 25732 31668 25742
rect 31500 25396 31556 25406
rect 30828 25394 31556 25396
rect 30828 25342 31502 25394
rect 31554 25342 31556 25394
rect 30828 25340 31556 25342
rect 30716 24948 30772 24958
rect 30828 24948 30884 25340
rect 31500 25330 31556 25340
rect 31500 24948 31556 24958
rect 30716 24946 30884 24948
rect 30716 24894 30718 24946
rect 30770 24894 30884 24946
rect 30716 24892 30884 24894
rect 31052 24946 31556 24948
rect 31052 24894 31502 24946
rect 31554 24894 31556 24946
rect 31052 24892 31556 24894
rect 30716 24882 30772 24892
rect 31052 24834 31108 24892
rect 31500 24882 31556 24892
rect 31612 24946 31668 25676
rect 31612 24894 31614 24946
rect 31666 24894 31668 24946
rect 31612 24882 31668 24894
rect 31052 24782 31054 24834
rect 31106 24782 31108 24834
rect 31052 24770 31108 24782
rect 31836 24834 31892 24846
rect 31836 24782 31838 24834
rect 31890 24782 31892 24834
rect 30828 24724 30884 24734
rect 31388 24724 31444 24734
rect 30828 24722 30996 24724
rect 30828 24670 30830 24722
rect 30882 24670 30996 24722
rect 30828 24668 30996 24670
rect 30828 24658 30884 24668
rect 30156 22978 30212 22988
rect 30268 24108 30660 24164
rect 30940 24276 30996 24668
rect 29372 22258 29652 22260
rect 29372 22206 29374 22258
rect 29426 22206 29652 22258
rect 29372 22204 29652 22206
rect 29708 22258 29764 22270
rect 29708 22206 29710 22258
rect 29762 22206 29764 22258
rect 29372 22194 29428 22204
rect 29596 21474 29652 21486
rect 29596 21422 29598 21474
rect 29650 21422 29652 21474
rect 29596 21140 29652 21422
rect 29708 21140 29764 22206
rect 29932 22258 29988 22270
rect 29932 22206 29934 22258
rect 29986 22206 29988 22258
rect 29932 22148 29988 22206
rect 29932 22082 29988 22092
rect 30268 21700 30324 24108
rect 30380 23940 30436 23950
rect 30604 23940 30660 23950
rect 30380 23938 30660 23940
rect 30380 23886 30382 23938
rect 30434 23886 30606 23938
rect 30658 23886 30660 23938
rect 30380 23884 30660 23886
rect 30380 22370 30436 23884
rect 30604 23874 30660 23884
rect 30940 23828 30996 24220
rect 31164 24722 31444 24724
rect 31164 24670 31390 24722
rect 31442 24670 31444 24722
rect 31164 24668 31444 24670
rect 31052 24164 31108 24174
rect 31164 24164 31220 24668
rect 31388 24658 31444 24668
rect 31052 24162 31220 24164
rect 31052 24110 31054 24162
rect 31106 24110 31220 24162
rect 31052 24108 31220 24110
rect 31052 24098 31108 24108
rect 30828 23716 30884 23726
rect 30828 23622 30884 23660
rect 30380 22318 30382 22370
rect 30434 22318 30436 22370
rect 30380 22306 30436 22318
rect 30604 23044 30660 23054
rect 30604 22370 30660 22988
rect 30604 22318 30606 22370
rect 30658 22318 30660 22370
rect 30604 22306 30660 22318
rect 30492 22148 30548 22158
rect 30492 22054 30548 22092
rect 30828 22146 30884 22158
rect 30828 22094 30830 22146
rect 30882 22094 30884 22146
rect 30828 21924 30884 22094
rect 30828 21858 30884 21868
rect 30268 21634 30324 21644
rect 29652 21084 29876 21140
rect 29596 21074 29652 21084
rect 29820 20916 29876 21084
rect 29260 20860 29428 20916
rect 29260 20692 29316 20702
rect 28924 19842 28980 19852
rect 29036 20580 29092 20590
rect 28588 19124 28644 19134
rect 28588 19122 28868 19124
rect 28588 19070 28590 19122
rect 28642 19070 28868 19122
rect 28588 19068 28868 19070
rect 28588 19058 28644 19068
rect 28812 18674 28868 19068
rect 29036 18788 29092 20524
rect 29260 19234 29316 20636
rect 29260 19182 29262 19234
rect 29314 19182 29316 19234
rect 29260 19170 29316 19182
rect 29036 18722 29092 18732
rect 28812 18622 28814 18674
rect 28866 18622 28868 18674
rect 28812 18610 28868 18622
rect 29148 18676 29204 18686
rect 28924 18562 28980 18574
rect 28924 18510 28926 18562
rect 28978 18510 28980 18562
rect 28476 17826 28532 17836
rect 28700 18450 28756 18462
rect 28700 18398 28702 18450
rect 28754 18398 28756 18450
rect 28588 17780 28644 17790
rect 28700 17780 28756 18398
rect 28644 17724 28756 17780
rect 28924 17780 28980 18510
rect 29148 17780 29204 18620
rect 28588 17666 28644 17724
rect 28924 17714 28980 17724
rect 29036 17724 29204 17780
rect 29260 18450 29316 18462
rect 29260 18398 29262 18450
rect 29314 18398 29316 18450
rect 28588 17614 28590 17666
rect 28642 17614 28644 17666
rect 28588 17602 28644 17614
rect 28476 17556 28532 17566
rect 28476 17462 28532 17500
rect 28364 17442 28420 17454
rect 28364 17390 28366 17442
rect 28418 17390 28420 17442
rect 28364 16996 28420 17390
rect 28364 16930 28420 16940
rect 29036 16324 29092 17724
rect 29148 17556 29204 17566
rect 29148 17462 29204 17500
rect 29260 17444 29316 18398
rect 29260 17378 29316 17388
rect 29372 18338 29428 20860
rect 29820 20914 30436 20916
rect 29820 20862 29822 20914
rect 29874 20862 30436 20914
rect 29820 20860 30436 20862
rect 29820 20850 29876 20860
rect 30156 20018 30212 20030
rect 30156 19966 30158 20018
rect 30210 19966 30212 20018
rect 29820 19906 29876 19918
rect 29820 19854 29822 19906
rect 29874 19854 29876 19906
rect 29708 19796 29764 19806
rect 29372 18286 29374 18338
rect 29426 18286 29428 18338
rect 29372 17666 29428 18286
rect 29372 17614 29374 17666
rect 29426 17614 29428 17666
rect 29372 17332 29428 17614
rect 29596 19740 29708 19796
rect 29596 17668 29652 19740
rect 29708 19730 29764 19740
rect 29708 18338 29764 18350
rect 29708 18286 29710 18338
rect 29762 18286 29764 18338
rect 29708 18226 29764 18286
rect 29708 18174 29710 18226
rect 29762 18174 29764 18226
rect 29708 18162 29764 18174
rect 29820 17780 29876 19854
rect 30156 19796 30212 19966
rect 30380 20018 30436 20860
rect 30940 20468 30996 23772
rect 31164 23268 31220 24108
rect 31276 24052 31332 24062
rect 31276 23826 31332 23996
rect 31836 24052 31892 24782
rect 32396 24612 32452 24622
rect 32396 24164 32452 24556
rect 31836 23986 31892 23996
rect 32172 24108 32452 24164
rect 31612 23940 31668 23950
rect 31612 23846 31668 23884
rect 31276 23774 31278 23826
rect 31330 23774 31332 23826
rect 31276 23762 31332 23774
rect 32060 23828 32116 23838
rect 32060 23734 32116 23772
rect 31164 23212 31332 23268
rect 31164 23044 31220 23054
rect 31164 22950 31220 22988
rect 31052 21700 31108 21710
rect 31052 21606 31108 21644
rect 31276 21474 31332 23212
rect 31612 23042 31668 23054
rect 31612 22990 31614 23042
rect 31666 22990 31668 23042
rect 31612 22596 31668 22990
rect 32172 22596 32228 24108
rect 31612 22540 32228 22596
rect 32284 23940 32340 23950
rect 31724 22370 31780 22382
rect 31724 22318 31726 22370
rect 31778 22318 31780 22370
rect 31388 22148 31444 22158
rect 31724 22148 31780 22318
rect 31388 22146 31780 22148
rect 31388 22094 31390 22146
rect 31442 22094 31780 22146
rect 31388 22092 31780 22094
rect 31388 21924 31444 22092
rect 31388 21858 31444 21868
rect 31612 21812 31668 21822
rect 31388 21698 31444 21710
rect 31388 21646 31390 21698
rect 31442 21646 31444 21698
rect 31388 21588 31444 21646
rect 31612 21698 31668 21756
rect 31612 21646 31614 21698
rect 31666 21646 31668 21698
rect 31612 21634 31668 21646
rect 31388 21522 31444 21532
rect 31276 21422 31278 21474
rect 31330 21422 31332 21474
rect 31276 21410 31332 21422
rect 31500 20802 31556 20814
rect 31500 20750 31502 20802
rect 31554 20750 31556 20802
rect 31500 20692 31556 20750
rect 31500 20626 31556 20636
rect 30940 20412 31556 20468
rect 30716 20132 31220 20188
rect 30716 20130 30772 20132
rect 30716 20078 30718 20130
rect 30770 20078 30772 20130
rect 30716 20066 30772 20078
rect 31164 20130 31220 20132
rect 31164 20078 31166 20130
rect 31218 20078 31220 20130
rect 31164 20066 31220 20078
rect 30380 19966 30382 20018
rect 30434 19966 30436 20018
rect 30380 19954 30436 19966
rect 31052 20018 31108 20030
rect 31052 19966 31054 20018
rect 31106 19966 31108 20018
rect 30156 19730 30212 19740
rect 30268 19906 30324 19918
rect 30268 19854 30270 19906
rect 30322 19854 30324 19906
rect 30268 19572 30324 19854
rect 29932 19516 30324 19572
rect 29932 19346 29988 19516
rect 29932 19294 29934 19346
rect 29986 19294 29988 19346
rect 29932 19282 29988 19294
rect 30380 19460 30436 19470
rect 30268 18788 30324 18798
rect 29820 17714 29876 17724
rect 30044 18340 30100 18350
rect 29708 17668 29764 17678
rect 29596 17666 29764 17668
rect 29596 17614 29710 17666
rect 29762 17614 29764 17666
rect 29596 17612 29764 17614
rect 29708 17556 29764 17612
rect 29932 17666 29988 17678
rect 29932 17614 29934 17666
rect 29986 17614 29988 17666
rect 29932 17556 29988 17614
rect 29708 17500 29988 17556
rect 29596 17444 29652 17454
rect 30044 17444 30100 18284
rect 29372 17266 29428 17276
rect 29484 17442 29652 17444
rect 29484 17390 29598 17442
rect 29650 17390 29652 17442
rect 29484 17388 29652 17390
rect 29372 16996 29428 17006
rect 29484 16996 29540 17388
rect 29596 17378 29652 17388
rect 29932 17388 30100 17444
rect 30156 17442 30212 17454
rect 30156 17390 30158 17442
rect 30210 17390 30212 17442
rect 29372 16994 29540 16996
rect 29372 16942 29374 16994
rect 29426 16942 29540 16994
rect 29372 16940 29540 16942
rect 29708 17332 29764 17342
rect 29372 16930 29428 16940
rect 29036 16268 29652 16324
rect 29372 16098 29428 16110
rect 29372 16046 29374 16098
rect 29426 16046 29428 16098
rect 28252 15092 28420 15148
rect 27020 13694 27022 13746
rect 27074 13694 27076 13746
rect 27020 13524 27076 13694
rect 27916 13692 28084 13748
rect 27692 13636 27748 13646
rect 27692 13542 27748 13580
rect 27020 11618 27076 13468
rect 27580 13524 27636 13534
rect 27132 13412 27188 13422
rect 27132 12290 27188 13356
rect 27132 12238 27134 12290
rect 27186 12238 27188 12290
rect 27132 12226 27188 12238
rect 27020 11566 27022 11618
rect 27074 11566 27076 11618
rect 27020 11554 27076 11566
rect 27132 11284 27188 11294
rect 27132 11170 27188 11228
rect 27132 11118 27134 11170
rect 27186 11118 27188 11170
rect 27132 10164 27188 11118
rect 27132 10098 27188 10108
rect 27468 10500 27524 10510
rect 27356 9940 27412 9950
rect 26908 9938 27412 9940
rect 26908 9886 27358 9938
rect 27410 9886 27412 9938
rect 26908 9884 27412 9886
rect 26908 9826 26964 9884
rect 27356 9874 27412 9884
rect 26908 9774 26910 9826
rect 26962 9774 26964 9826
rect 26908 9762 26964 9774
rect 26572 9716 26628 9726
rect 26572 9622 26628 9660
rect 27468 9154 27524 10444
rect 27468 9102 27470 9154
rect 27522 9102 27524 9154
rect 27468 9090 27524 9102
rect 26684 9044 26740 9054
rect 26460 9042 26740 9044
rect 26460 8990 26686 9042
rect 26738 8990 26740 9042
rect 26460 8988 26740 8990
rect 26124 6692 26180 6702
rect 26124 6598 26180 6636
rect 26012 6514 26068 6524
rect 25004 6300 25172 6356
rect 24668 6132 24724 6142
rect 24668 6038 24724 6076
rect 24556 4958 24558 5010
rect 24610 4958 24612 5010
rect 24556 4946 24612 4958
rect 24780 5684 24836 5694
rect 24780 5010 24836 5628
rect 25004 5236 25060 5246
rect 25004 5142 25060 5180
rect 24780 4958 24782 5010
rect 24834 4958 24836 5010
rect 24780 4946 24836 4958
rect 25116 5122 25172 6300
rect 25564 6290 25620 6300
rect 25116 5070 25118 5122
rect 25170 5070 25172 5122
rect 25116 4788 25172 5070
rect 24444 4732 25172 4788
rect 25340 6132 25396 6142
rect 24444 4226 24500 4732
rect 25340 4562 25396 6076
rect 26012 5908 26068 5918
rect 26012 5814 26068 5852
rect 26236 5908 26292 5918
rect 25452 5796 25508 5806
rect 25452 5572 25508 5740
rect 25788 5684 25844 5694
rect 26236 5684 26292 5852
rect 26348 5796 26404 5806
rect 26348 5702 26404 5740
rect 25788 5682 26292 5684
rect 25788 5630 25790 5682
rect 25842 5630 26292 5682
rect 25788 5628 26292 5630
rect 26460 5682 26516 5694
rect 26460 5630 26462 5682
rect 26514 5630 26516 5682
rect 25788 5618 25844 5628
rect 25452 5506 25508 5516
rect 26460 5572 26516 5630
rect 26460 5506 26516 5516
rect 25564 5122 25620 5134
rect 25564 5070 25566 5122
rect 25618 5070 25620 5122
rect 25564 5012 25620 5070
rect 25564 4946 25620 4956
rect 26236 5012 26292 5022
rect 26572 5012 26628 8988
rect 26684 8978 26740 8988
rect 26684 8372 26740 8382
rect 26684 8146 26740 8316
rect 26684 8094 26686 8146
rect 26738 8094 26740 8146
rect 26684 7364 26740 8094
rect 27020 8034 27076 8046
rect 27020 7982 27022 8034
rect 27074 7982 27076 8034
rect 27020 7700 27076 7982
rect 27020 7606 27076 7644
rect 27468 7588 27524 7598
rect 27580 7588 27636 13468
rect 27804 13522 27860 13534
rect 27804 13470 27806 13522
rect 27858 13470 27860 13522
rect 27804 13412 27860 13470
rect 27804 13346 27860 13356
rect 27692 13188 27748 13198
rect 27692 13074 27748 13132
rect 27692 13022 27694 13074
rect 27746 13022 27748 13074
rect 27692 13010 27748 13022
rect 27916 12292 27972 13692
rect 28028 13524 28084 13534
rect 28252 13524 28308 13534
rect 28028 13522 28252 13524
rect 28028 13470 28030 13522
rect 28082 13470 28252 13522
rect 28028 13468 28252 13470
rect 28028 13458 28084 13468
rect 28252 13458 28308 13468
rect 28140 12292 28196 12302
rect 27916 12178 27972 12236
rect 27916 12126 27918 12178
rect 27970 12126 27972 12178
rect 27916 12114 27972 12126
rect 28028 12290 28196 12292
rect 28028 12238 28142 12290
rect 28194 12238 28196 12290
rect 28028 12236 28196 12238
rect 27804 11620 27860 11630
rect 27804 11618 27972 11620
rect 27804 11566 27806 11618
rect 27858 11566 27972 11618
rect 27804 11564 27972 11566
rect 27804 11554 27860 11564
rect 27804 11396 27860 11406
rect 27804 11302 27860 11340
rect 27468 7586 27636 7588
rect 27468 7534 27470 7586
rect 27522 7534 27636 7586
rect 27468 7532 27636 7534
rect 27804 10164 27860 10174
rect 27468 7522 27524 7532
rect 26684 7308 27076 7364
rect 27020 6690 27076 7308
rect 27804 7140 27860 10108
rect 27916 7474 27972 11564
rect 28028 11282 28084 12236
rect 28140 12226 28196 12236
rect 28364 11396 28420 15092
rect 28588 14532 28644 14542
rect 29372 14532 29428 16046
rect 29596 15538 29652 16268
rect 29596 15486 29598 15538
rect 29650 15486 29652 15538
rect 29596 14644 29652 15486
rect 29596 14550 29652 14588
rect 28588 14530 29428 14532
rect 28588 14478 28590 14530
rect 28642 14478 29428 14530
rect 28588 14476 29428 14478
rect 28588 14466 28644 14476
rect 29372 12962 29428 14476
rect 29372 12910 29374 12962
rect 29426 12910 29428 12962
rect 29372 12852 29428 12910
rect 29372 12786 29428 12796
rect 29596 12628 29652 12638
rect 29596 12402 29652 12572
rect 29596 12350 29598 12402
rect 29650 12350 29652 12402
rect 29596 12338 29652 12350
rect 28476 12292 28532 12302
rect 28476 12198 28532 12236
rect 28812 12292 28868 12302
rect 28812 12290 29204 12292
rect 28812 12238 28814 12290
rect 28866 12238 29204 12290
rect 28812 12236 29204 12238
rect 28812 12226 28868 12236
rect 28364 11302 28420 11340
rect 29148 11844 29204 12236
rect 28028 11230 28030 11282
rect 28082 11230 28084 11282
rect 28028 10612 28084 11230
rect 28588 11284 28644 11294
rect 28588 11282 29092 11284
rect 28588 11230 28590 11282
rect 28642 11230 29092 11282
rect 28588 11228 29092 11230
rect 28588 11218 28644 11228
rect 28140 11170 28196 11182
rect 28140 11118 28142 11170
rect 28194 11118 28196 11170
rect 28140 10724 28196 11118
rect 29036 10948 29092 11228
rect 29148 11170 29204 11788
rect 29708 11732 29764 17276
rect 29932 15148 29988 17388
rect 30156 17108 30212 17390
rect 30044 17052 30212 17108
rect 30044 16212 30100 17052
rect 30156 16884 30212 16894
rect 30156 16790 30212 16828
rect 30268 16772 30324 18732
rect 30380 17666 30436 19404
rect 30380 17614 30382 17666
rect 30434 17614 30436 17666
rect 30380 17220 30436 17614
rect 30492 19348 30548 19358
rect 30492 17444 30548 19292
rect 31052 19348 31108 19966
rect 31052 19282 31108 19292
rect 31276 20018 31332 20030
rect 31276 19966 31278 20018
rect 31330 19966 31332 20018
rect 31276 19348 31332 19966
rect 31276 19282 31332 19292
rect 31052 17780 31108 17790
rect 30716 17778 31108 17780
rect 30716 17726 31054 17778
rect 31106 17726 31108 17778
rect 30716 17724 31108 17726
rect 30604 17668 30660 17678
rect 30716 17668 30772 17724
rect 31052 17714 31108 17724
rect 30604 17666 30772 17668
rect 30604 17614 30606 17666
rect 30658 17614 30772 17666
rect 30604 17612 30772 17614
rect 30604 17602 30660 17612
rect 31388 17556 31444 17566
rect 31388 17462 31444 17500
rect 30940 17444 30996 17454
rect 30492 17442 30996 17444
rect 30492 17390 30942 17442
rect 30994 17390 30996 17442
rect 30492 17388 30996 17390
rect 30940 17378 30996 17388
rect 31164 17444 31220 17454
rect 31164 17350 31220 17388
rect 30380 17164 30884 17220
rect 30492 16772 30548 16782
rect 30268 16716 30492 16772
rect 30492 16706 30548 16716
rect 30156 16212 30212 16222
rect 30044 16210 30212 16212
rect 30044 16158 30158 16210
rect 30210 16158 30212 16210
rect 30044 16156 30212 16158
rect 30156 16146 30212 16156
rect 30156 15316 30212 15326
rect 30604 15316 30660 17164
rect 30828 17106 30884 17164
rect 31500 17108 31556 20412
rect 31724 20020 31780 20030
rect 31724 19926 31780 19964
rect 31948 18676 32004 22540
rect 32284 22372 32340 23884
rect 32620 22372 32676 22382
rect 32284 22370 32676 22372
rect 32284 22318 32286 22370
rect 32338 22318 32622 22370
rect 32674 22318 32676 22370
rect 32284 22316 32676 22318
rect 32284 22306 32340 22316
rect 32620 22306 32676 22316
rect 32172 22260 32228 22270
rect 32060 21700 32116 21710
rect 32060 21586 32116 21644
rect 32060 21534 32062 21586
rect 32114 21534 32116 21586
rect 32060 21522 32116 21534
rect 32172 20130 32228 22204
rect 32284 21474 32340 21486
rect 32284 21422 32286 21474
rect 32338 21422 32340 21474
rect 32284 20914 32340 21422
rect 32284 20862 32286 20914
rect 32338 20862 32340 20914
rect 32284 20850 32340 20862
rect 32396 21362 32452 21374
rect 32396 21310 32398 21362
rect 32450 21310 32452 21362
rect 32172 20078 32174 20130
rect 32226 20078 32228 20130
rect 32172 20020 32228 20078
rect 32172 19954 32228 19964
rect 32060 19348 32116 19358
rect 32060 18788 32116 19292
rect 32396 19234 32452 21310
rect 32508 20692 32564 20702
rect 32508 20130 32564 20636
rect 32508 20078 32510 20130
rect 32562 20078 32564 20130
rect 32508 20066 32564 20078
rect 32396 19182 32398 19234
rect 32450 19182 32452 19234
rect 32396 19170 32452 19182
rect 32060 18722 32116 18732
rect 31836 18620 32004 18676
rect 31836 18228 31892 18620
rect 32844 18564 32900 29372
rect 32956 29362 33012 29372
rect 33292 29428 33348 29438
rect 33292 29334 33348 29372
rect 33404 29092 33460 29102
rect 32956 28980 33012 28990
rect 32956 28082 33012 28924
rect 32956 28030 32958 28082
rect 33010 28030 33012 28082
rect 32956 28018 33012 28030
rect 33068 28308 33124 28318
rect 33068 28082 33124 28252
rect 33068 28030 33070 28082
rect 33122 28030 33124 28082
rect 33068 28018 33124 28030
rect 33292 27860 33348 27870
rect 33180 27858 33348 27860
rect 33180 27806 33294 27858
rect 33346 27806 33348 27858
rect 33180 27804 33348 27806
rect 33180 27748 33236 27804
rect 33292 27794 33348 27804
rect 33180 27682 33236 27692
rect 33292 27636 33348 27646
rect 32956 27412 33012 27422
rect 32956 26908 33012 27356
rect 33292 27186 33348 27580
rect 33292 27134 33294 27186
rect 33346 27134 33348 27186
rect 33292 27122 33348 27134
rect 33404 26908 33460 29036
rect 33516 28868 33572 29708
rect 33628 29988 33684 29998
rect 33628 29538 33684 29932
rect 33740 29988 33796 29998
rect 33964 29988 34020 29998
rect 33740 29986 33908 29988
rect 33740 29934 33742 29986
rect 33794 29934 33908 29986
rect 33740 29932 33908 29934
rect 33740 29922 33796 29932
rect 33628 29486 33630 29538
rect 33682 29486 33684 29538
rect 33628 29474 33684 29486
rect 33740 29428 33796 29438
rect 33740 28980 33796 29372
rect 33852 29092 33908 29932
rect 33964 29894 34020 29932
rect 34076 29428 34132 30156
rect 34076 29334 34132 29372
rect 33852 29036 34244 29092
rect 33740 28924 34132 28980
rect 33516 28802 33572 28812
rect 34076 28196 34132 28924
rect 34188 28756 34244 29036
rect 34188 28662 34244 28700
rect 34076 28082 34132 28140
rect 34076 28030 34078 28082
rect 34130 28030 34132 28082
rect 34076 28018 34132 28030
rect 33628 27972 33684 27982
rect 33516 27916 33628 27972
rect 33516 27858 33572 27916
rect 33628 27906 33684 27916
rect 34412 27972 34468 31612
rect 34636 31108 34692 31836
rect 34972 31780 35028 40908
rect 35308 40404 35364 41244
rect 36988 41188 37044 41198
rect 36988 41094 37044 41132
rect 35756 41076 35812 41086
rect 35756 40516 35812 41020
rect 37100 41076 37156 41086
rect 37100 40982 37156 41020
rect 37212 40852 37268 41356
rect 37436 41076 37492 43708
rect 37548 43698 37604 43708
rect 38780 43764 38836 43774
rect 38892 43764 38948 45052
rect 39116 45014 39172 45052
rect 38780 43762 38948 43764
rect 38780 43710 38782 43762
rect 38834 43710 38948 43762
rect 38780 43708 38948 43710
rect 39228 44884 39284 44894
rect 39228 43708 39284 44828
rect 38780 43698 38836 43708
rect 37772 43652 37828 43662
rect 37772 43558 37828 43596
rect 39116 43652 39284 43708
rect 39340 43708 39396 45388
rect 39452 45106 39508 45836
rect 39452 45054 39454 45106
rect 39506 45054 39508 45106
rect 39452 44660 39508 45054
rect 39676 45106 39732 45948
rect 39900 45938 39956 45948
rect 40012 45330 40068 46172
rect 40012 45278 40014 45330
rect 40066 45278 40068 45330
rect 40012 45220 40068 45278
rect 40012 45154 40068 45164
rect 39676 45054 39678 45106
rect 39730 45054 39732 45106
rect 39676 45042 39732 45054
rect 39564 44996 39620 45006
rect 39564 44902 39620 44940
rect 39452 44604 40068 44660
rect 39676 44436 39732 44446
rect 39676 43708 39732 44380
rect 39340 43652 39508 43708
rect 39676 43652 39956 43708
rect 38556 43538 38612 43550
rect 38556 43486 38558 43538
rect 38610 43486 38612 43538
rect 38444 43428 38500 43438
rect 38108 42868 38164 42878
rect 37660 42866 38164 42868
rect 37660 42814 38110 42866
rect 38162 42814 38164 42866
rect 37660 42812 38164 42814
rect 37660 42754 37716 42812
rect 38108 42802 38164 42812
rect 37660 42702 37662 42754
rect 37714 42702 37716 42754
rect 37660 42690 37716 42702
rect 38220 42756 38276 42766
rect 38276 42700 38388 42756
rect 38220 42662 38276 42700
rect 38108 42532 38164 42542
rect 38108 41186 38164 42476
rect 38332 41860 38388 42700
rect 38444 42754 38500 43372
rect 38444 42702 38446 42754
rect 38498 42702 38500 42754
rect 38444 42690 38500 42702
rect 38556 43316 38612 43486
rect 38780 43540 38836 43550
rect 38780 43426 38836 43484
rect 39004 43540 39060 43550
rect 39004 43446 39060 43484
rect 38780 43374 38782 43426
rect 38834 43374 38836 43426
rect 38780 43362 38836 43374
rect 38556 42532 38612 43260
rect 38780 42980 38836 42990
rect 38556 42466 38612 42476
rect 38668 42642 38724 42654
rect 38668 42590 38670 42642
rect 38722 42590 38724 42642
rect 38444 41860 38500 41870
rect 38332 41858 38500 41860
rect 38332 41806 38446 41858
rect 38498 41806 38500 41858
rect 38332 41804 38500 41806
rect 38444 41794 38500 41804
rect 38108 41134 38110 41186
rect 38162 41134 38164 41186
rect 38108 41122 38164 41134
rect 36988 40796 37268 40852
rect 37324 41020 37492 41076
rect 37660 41076 37716 41086
rect 35756 40422 35812 40460
rect 36428 40628 36484 40638
rect 35308 40338 35364 40348
rect 35756 40292 35812 40302
rect 35980 40292 36036 40302
rect 35196 40012 35460 40022
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35196 39946 35460 39956
rect 35644 39844 35700 39854
rect 35644 39750 35700 39788
rect 35308 39732 35364 39742
rect 35308 39638 35364 39676
rect 35756 39396 35812 40236
rect 35868 40290 36036 40292
rect 35868 40238 35982 40290
rect 36034 40238 36036 40290
rect 35868 40236 36036 40238
rect 35868 39620 35924 40236
rect 35980 40226 36036 40236
rect 35980 39844 36036 39854
rect 36204 39844 36260 39854
rect 35980 39842 36260 39844
rect 35980 39790 35982 39842
rect 36034 39790 36206 39842
rect 36258 39790 36260 39842
rect 35980 39788 36260 39790
rect 35980 39778 36036 39788
rect 36204 39778 36260 39788
rect 36428 39620 36484 40572
rect 36540 40404 36596 40414
rect 36540 40310 36596 40348
rect 36540 39844 36596 39854
rect 36540 39842 36932 39844
rect 36540 39790 36542 39842
rect 36594 39790 36932 39842
rect 36540 39788 36932 39790
rect 36540 39778 36596 39788
rect 35868 39564 36148 39620
rect 35868 39396 35924 39406
rect 35756 39394 35924 39396
rect 35756 39342 35870 39394
rect 35922 39342 35924 39394
rect 35756 39340 35924 39342
rect 35196 38444 35460 38454
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35196 38378 35460 38388
rect 35532 38050 35588 38062
rect 35532 37998 35534 38050
rect 35586 37998 35588 38050
rect 35084 37156 35140 37166
rect 35084 36484 35140 37100
rect 35196 36876 35460 36886
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35196 36810 35460 36820
rect 35196 36484 35252 36494
rect 35084 36482 35252 36484
rect 35084 36430 35198 36482
rect 35250 36430 35252 36482
rect 35084 36428 35252 36430
rect 35196 36418 35252 36428
rect 35532 36482 35588 37998
rect 35644 37266 35700 37278
rect 35644 37214 35646 37266
rect 35698 37214 35700 37266
rect 35644 37156 35700 37214
rect 35644 37090 35700 37100
rect 35532 36430 35534 36482
rect 35586 36430 35588 36482
rect 35532 36418 35588 36430
rect 35308 36372 35364 36382
rect 35868 36372 35924 39340
rect 35980 39284 36036 39294
rect 35980 37940 36036 39228
rect 36092 38274 36148 39564
rect 36316 39564 36484 39620
rect 36316 38668 36372 39564
rect 36428 39396 36484 39406
rect 36428 39302 36484 39340
rect 36876 38946 36932 39788
rect 36988 39730 37044 40796
rect 37100 40292 37156 40302
rect 37100 40198 37156 40236
rect 36988 39678 36990 39730
rect 37042 39678 37044 39730
rect 36988 39666 37044 39678
rect 36876 38894 36878 38946
rect 36930 38894 36932 38946
rect 36876 38882 36932 38894
rect 36092 38222 36094 38274
rect 36146 38222 36148 38274
rect 36092 38210 36148 38222
rect 36204 38612 36372 38668
rect 36204 38050 36260 38612
rect 36204 37998 36206 38050
rect 36258 37998 36260 38050
rect 36204 37986 36260 37998
rect 36988 38050 37044 38062
rect 36988 37998 36990 38050
rect 37042 37998 37044 38050
rect 36092 37940 36148 37950
rect 35980 37938 36148 37940
rect 35980 37886 36094 37938
rect 36146 37886 36148 37938
rect 35980 37884 36148 37886
rect 36092 37874 36148 37884
rect 36988 37604 37044 37998
rect 36764 37548 36988 37604
rect 36092 37490 36148 37502
rect 36092 37438 36094 37490
rect 36146 37438 36148 37490
rect 36092 36706 36148 37438
rect 36092 36654 36094 36706
rect 36146 36654 36148 36706
rect 36092 36642 36148 36654
rect 35364 36316 35476 36372
rect 35308 36278 35364 36316
rect 35420 35588 35476 36316
rect 35868 36306 35924 36316
rect 36316 36372 36372 36382
rect 36316 36278 36372 36316
rect 36204 36260 36260 36270
rect 36204 36166 36260 36204
rect 36540 35700 36596 35710
rect 35644 35588 35700 35598
rect 35420 35586 35700 35588
rect 35420 35534 35646 35586
rect 35698 35534 35700 35586
rect 35420 35532 35700 35534
rect 35644 35522 35700 35532
rect 35196 35308 35460 35318
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35196 35242 35460 35252
rect 36092 34692 36148 34702
rect 36092 34354 36148 34636
rect 36092 34302 36094 34354
rect 36146 34302 36148 34354
rect 36092 34290 36148 34302
rect 35084 34132 35140 34142
rect 35084 34038 35140 34076
rect 35532 34018 35588 34030
rect 35532 33966 35534 34018
rect 35586 33966 35588 34018
rect 35196 33740 35460 33750
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35196 33674 35460 33684
rect 35532 32564 35588 33966
rect 36428 33460 36484 33470
rect 35868 33458 36484 33460
rect 35868 33406 36430 33458
rect 36482 33406 36484 33458
rect 35868 33404 36484 33406
rect 35756 32788 35812 32798
rect 35756 32694 35812 32732
rect 35868 32674 35924 33404
rect 36428 33394 36484 33404
rect 35868 32622 35870 32674
rect 35922 32622 35924 32674
rect 35868 32610 35924 32622
rect 35196 32172 35460 32182
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35196 32106 35460 32116
rect 35532 32004 35588 32508
rect 36540 32228 36596 35644
rect 36540 32162 36596 32172
rect 36652 32450 36708 32462
rect 36652 32398 36654 32450
rect 36706 32398 36708 32450
rect 35420 31948 35588 32004
rect 35756 32004 35812 32014
rect 34636 31042 34692 31052
rect 34748 31724 35028 31780
rect 35308 31780 35364 31790
rect 34524 30100 34580 30110
rect 34524 30006 34580 30044
rect 34748 29652 34804 31724
rect 35196 31666 35252 31678
rect 35196 31614 35198 31666
rect 35250 31614 35252 31666
rect 34972 31556 35028 31566
rect 34972 31462 35028 31500
rect 35196 31108 35252 31614
rect 34860 31052 35252 31108
rect 34860 30322 34916 31052
rect 35308 30772 35364 31724
rect 34860 30270 34862 30322
rect 34914 30270 34916 30322
rect 34860 30258 34916 30270
rect 35084 30716 35364 30772
rect 35420 30772 35476 31948
rect 35756 31890 35812 31948
rect 36652 32004 36708 32398
rect 36652 31938 36708 31948
rect 35756 31838 35758 31890
rect 35810 31838 35812 31890
rect 35756 31826 35812 31838
rect 36092 31780 36148 31790
rect 36764 31780 36820 37548
rect 36988 37538 37044 37548
rect 36988 36372 37044 36382
rect 36988 36260 37044 36316
rect 37100 36260 37156 36270
rect 36988 36258 37156 36260
rect 36988 36206 37102 36258
rect 37154 36206 37156 36258
rect 36988 36204 37156 36206
rect 36988 34914 37044 36204
rect 37100 36194 37156 36204
rect 36988 34862 36990 34914
rect 37042 34862 37044 34914
rect 36988 33684 37044 34862
rect 37324 34468 37380 41020
rect 37660 40982 37716 41020
rect 38444 41076 38500 41086
rect 38444 40982 38500 41020
rect 37772 40964 37828 40974
rect 38332 40964 38388 40974
rect 37772 40962 38164 40964
rect 37772 40910 37774 40962
rect 37826 40910 38164 40962
rect 37772 40908 38164 40910
rect 37772 40898 37828 40908
rect 38108 40516 38164 40908
rect 38332 40870 38388 40908
rect 38556 40962 38612 40974
rect 38556 40910 38558 40962
rect 38610 40910 38612 40962
rect 38220 40516 38276 40526
rect 38108 40514 38276 40516
rect 38108 40462 38222 40514
rect 38274 40462 38276 40514
rect 38108 40460 38276 40462
rect 38220 40450 38276 40460
rect 37436 40404 37492 40414
rect 37436 38836 37492 40348
rect 37548 39508 37604 39518
rect 37548 39414 37604 39452
rect 37996 39508 38052 39518
rect 37548 38836 37604 38846
rect 37436 38834 37604 38836
rect 37436 38782 37550 38834
rect 37602 38782 37604 38834
rect 37436 38780 37604 38782
rect 37436 37492 37492 38780
rect 37548 38770 37604 38780
rect 37996 38668 38052 39452
rect 38332 39394 38388 39406
rect 38332 39342 38334 39394
rect 38386 39342 38388 39394
rect 38332 38948 38388 39342
rect 38444 38948 38500 38958
rect 38332 38946 38500 38948
rect 38332 38894 38446 38946
rect 38498 38894 38500 38946
rect 38332 38892 38500 38894
rect 38108 38722 38164 38734
rect 38108 38670 38110 38722
rect 38162 38670 38164 38722
rect 38108 38668 38164 38670
rect 37884 38612 38164 38668
rect 38332 38668 38388 38892
rect 38444 38882 38500 38892
rect 38556 38948 38612 40910
rect 38668 40964 38724 42590
rect 38780 41524 38836 42924
rect 39004 42756 39060 42766
rect 39116 42756 39172 43652
rect 39228 43538 39284 43550
rect 39228 43486 39230 43538
rect 39282 43486 39284 43538
rect 39228 42980 39284 43486
rect 39228 42914 39284 42924
rect 39228 42756 39284 42766
rect 39116 42754 39284 42756
rect 39116 42702 39230 42754
rect 39282 42702 39284 42754
rect 39116 42700 39284 42702
rect 39004 42662 39060 42700
rect 39228 42690 39284 42700
rect 39340 42754 39396 42766
rect 39340 42702 39342 42754
rect 39394 42702 39396 42754
rect 39340 42196 39396 42702
rect 39340 42130 39396 42140
rect 38780 41458 38836 41468
rect 38892 41858 38948 41870
rect 38892 41806 38894 41858
rect 38946 41806 38948 41858
rect 38892 41746 38948 41806
rect 39116 41860 39172 41870
rect 39116 41748 39172 41804
rect 39340 41858 39396 41870
rect 39340 41806 39342 41858
rect 39394 41806 39396 41858
rect 39340 41748 39396 41806
rect 38892 41694 38894 41746
rect 38946 41694 38948 41746
rect 38780 41188 38836 41198
rect 38780 41094 38836 41132
rect 38668 40898 38724 40908
rect 38892 40404 38948 41694
rect 39004 41692 39396 41748
rect 39004 41188 39060 41692
rect 39340 41524 39396 41534
rect 39340 41298 39396 41468
rect 39340 41246 39342 41298
rect 39394 41246 39396 41298
rect 39340 41234 39396 41246
rect 39004 41132 39172 41188
rect 38892 40338 38948 40348
rect 38556 38882 38612 38892
rect 39004 39956 39060 39966
rect 39004 38836 39060 39900
rect 39116 39618 39172 41132
rect 39452 39620 39508 43652
rect 39788 43426 39844 43438
rect 39788 43374 39790 43426
rect 39842 43374 39844 43426
rect 39788 42868 39844 43374
rect 39564 42812 39844 42868
rect 39564 41746 39620 42812
rect 39564 41694 39566 41746
rect 39618 41694 39620 41746
rect 39564 41682 39620 41694
rect 39676 42644 39732 42654
rect 39900 42644 39956 43652
rect 40012 42866 40068 44604
rect 40124 43426 40180 48300
rect 40348 48244 40404 48254
rect 40348 48150 40404 48188
rect 40460 48132 40516 50428
rect 41132 50372 41188 50382
rect 41356 50372 41412 51324
rect 41468 51314 41524 51324
rect 41580 51156 41636 51660
rect 41468 51100 41636 51156
rect 42028 51492 42084 51502
rect 41468 50482 41524 51100
rect 42028 50708 42084 51436
rect 42028 50614 42084 50652
rect 41468 50430 41470 50482
rect 41522 50430 41524 50482
rect 41468 50418 41524 50430
rect 41020 50370 41412 50372
rect 41020 50318 41134 50370
rect 41186 50318 41412 50370
rect 41020 50316 41412 50318
rect 41580 50372 41636 50382
rect 42140 50372 42196 51998
rect 42252 54404 42308 54414
rect 42252 51378 42308 54348
rect 42700 53732 42756 55246
rect 42812 54628 42868 56142
rect 42924 55972 42980 55982
rect 42924 55878 42980 55916
rect 43036 55858 43092 55870
rect 43036 55806 43038 55858
rect 43090 55806 43092 55858
rect 43036 55468 43092 55806
rect 43260 55524 43316 55534
rect 43372 55524 43428 57372
rect 44604 57092 44660 57102
rect 44604 56306 44660 57036
rect 44604 56254 44606 56306
rect 44658 56254 44660 56306
rect 44604 56242 44660 56254
rect 43820 56082 43876 56094
rect 43820 56030 43822 56082
rect 43874 56030 43876 56082
rect 43596 55524 43652 55534
rect 43372 55468 43540 55524
rect 43036 55412 43204 55468
rect 42812 53844 42868 54572
rect 42812 53778 42868 53788
rect 43036 55188 43092 55198
rect 42588 53676 42756 53732
rect 42588 52948 42644 53676
rect 42700 53508 42756 53518
rect 42700 53414 42756 53452
rect 42364 52892 42644 52948
rect 42364 52276 42420 52892
rect 42364 51828 42420 52220
rect 42476 52164 42532 52174
rect 43036 52164 43092 55132
rect 43148 53284 43204 55412
rect 43260 55412 43316 55468
rect 43260 55346 43316 55356
rect 43372 55298 43428 55310
rect 43372 55246 43374 55298
rect 43426 55246 43428 55298
rect 43372 54852 43428 55246
rect 43372 54786 43428 54796
rect 43484 54740 43540 55468
rect 43596 55410 43652 55468
rect 43596 55358 43598 55410
rect 43650 55358 43652 55410
rect 43596 55346 43652 55358
rect 43708 55188 43764 55198
rect 43484 54674 43540 54684
rect 43596 55076 43652 55086
rect 43596 54626 43652 55020
rect 43708 55074 43764 55132
rect 43708 55022 43710 55074
rect 43762 55022 43764 55074
rect 43708 55010 43764 55022
rect 43596 54574 43598 54626
rect 43650 54574 43652 54626
rect 43596 54562 43652 54574
rect 43148 53218 43204 53228
rect 43820 53060 43876 56030
rect 44044 55972 44100 55982
rect 44044 55298 44100 55916
rect 44044 55246 44046 55298
rect 44098 55246 44100 55298
rect 44044 53508 44100 55246
rect 44940 55188 44996 55198
rect 44940 55094 44996 55132
rect 44268 55074 44324 55086
rect 44268 55022 44270 55074
rect 44322 55022 44324 55074
rect 44268 54852 44324 55022
rect 44828 55076 44884 55086
rect 44828 54982 44884 55020
rect 44268 54786 44324 54796
rect 44268 54514 44324 54526
rect 44268 54462 44270 54514
rect 44322 54462 44324 54514
rect 44268 53732 44324 54462
rect 44716 54516 44772 54526
rect 44716 54422 44772 54460
rect 44828 54068 44884 54078
rect 44268 53666 44324 53676
rect 44716 54012 44828 54068
rect 44044 53442 44100 53452
rect 43820 52994 43876 53004
rect 44156 53396 44212 53406
rect 42476 52162 43092 52164
rect 42476 52110 42478 52162
rect 42530 52110 43092 52162
rect 42476 52108 43092 52110
rect 43596 52836 43652 52846
rect 43820 52836 43876 52846
rect 42476 52098 42532 52108
rect 43484 52052 43540 52062
rect 43484 51958 43540 51996
rect 42924 51940 42980 51950
rect 42924 51846 42980 51884
rect 42364 51772 42532 51828
rect 42252 51326 42254 51378
rect 42306 51326 42308 51378
rect 42252 51314 42308 51326
rect 42476 51378 42532 51772
rect 42476 51326 42478 51378
rect 42530 51326 42532 51378
rect 42364 51268 42420 51278
rect 42364 50594 42420 51212
rect 42364 50542 42366 50594
rect 42418 50542 42420 50594
rect 42364 50530 42420 50542
rect 41636 50316 42196 50372
rect 41020 48914 41076 50316
rect 41132 50306 41188 50316
rect 41468 50260 41524 50270
rect 41356 49812 41412 49822
rect 41468 49812 41524 50204
rect 41580 50034 41636 50316
rect 41580 49982 41582 50034
rect 41634 49982 41636 50034
rect 41580 49970 41636 49982
rect 42140 49924 42196 49934
rect 42140 49830 42196 49868
rect 41356 49810 41524 49812
rect 41356 49758 41358 49810
rect 41410 49758 41524 49810
rect 41356 49756 41524 49758
rect 41356 49746 41412 49756
rect 41020 48862 41022 48914
rect 41074 48862 41076 48914
rect 40572 48804 40628 48814
rect 40908 48804 40964 48814
rect 40628 48802 40964 48804
rect 40628 48750 40910 48802
rect 40962 48750 40964 48802
rect 40628 48748 40964 48750
rect 40572 48710 40628 48748
rect 40908 48738 40964 48748
rect 41020 48580 41076 48862
rect 40460 48066 40516 48076
rect 40908 48524 41076 48580
rect 41244 49588 41300 49598
rect 40908 48020 40964 48524
rect 41020 48356 41076 48366
rect 41244 48356 41300 49532
rect 41356 49140 41412 49150
rect 41356 49026 41412 49084
rect 41356 48974 41358 49026
rect 41410 48974 41412 49026
rect 41356 48962 41412 48974
rect 41020 48354 41300 48356
rect 41020 48302 41022 48354
rect 41074 48302 41300 48354
rect 41020 48300 41300 48302
rect 41020 48290 41076 48300
rect 41468 48244 41524 49756
rect 41916 49810 41972 49822
rect 41916 49758 41918 49810
rect 41970 49758 41972 49810
rect 41916 48804 41972 49758
rect 42028 49698 42084 49710
rect 42028 49646 42030 49698
rect 42082 49646 42084 49698
rect 42028 49364 42084 49646
rect 42476 49476 42532 51326
rect 43036 51490 43092 51502
rect 43036 51438 43038 51490
rect 43090 51438 43092 51490
rect 42812 51268 42868 51278
rect 42812 51266 42980 51268
rect 42812 51214 42814 51266
rect 42866 51214 42980 51266
rect 42812 51212 42980 51214
rect 42812 51202 42868 51212
rect 42924 49924 42980 51212
rect 43036 50484 43092 51438
rect 43484 51380 43540 51390
rect 43036 50418 43092 50428
rect 43148 51378 43540 51380
rect 43148 51326 43486 51378
rect 43538 51326 43540 51378
rect 43148 51324 43540 51326
rect 42924 49858 42980 49868
rect 42252 49420 42532 49476
rect 42588 49810 42644 49822
rect 42588 49758 42590 49810
rect 42642 49758 42644 49810
rect 42028 49308 42196 49364
rect 41916 48738 41972 48748
rect 42028 49140 42084 49150
rect 41244 48132 41300 48142
rect 40908 47964 41188 48020
rect 41020 47572 41076 47582
rect 41020 47478 41076 47516
rect 41020 47012 41076 47022
rect 41020 46898 41076 46956
rect 41020 46846 41022 46898
rect 41074 46846 41076 46898
rect 41020 46834 41076 46846
rect 40348 46562 40404 46574
rect 40348 46510 40350 46562
rect 40402 46510 40404 46562
rect 40348 45892 40404 46510
rect 40348 45798 40404 45836
rect 40236 45332 40292 45342
rect 40236 44436 40292 45276
rect 40908 45332 40964 45342
rect 40908 45238 40964 45276
rect 40348 45108 40404 45118
rect 40348 45014 40404 45052
rect 41132 45106 41188 47964
rect 41244 47124 41300 48076
rect 41468 47348 41524 48188
rect 41692 48356 41748 48366
rect 41468 47282 41524 47292
rect 41580 47458 41636 47470
rect 41580 47406 41582 47458
rect 41634 47406 41636 47458
rect 41356 47236 41412 47246
rect 41356 47142 41412 47180
rect 41244 46564 41300 47068
rect 41356 46564 41412 46574
rect 41244 46562 41412 46564
rect 41244 46510 41358 46562
rect 41410 46510 41412 46562
rect 41244 46508 41412 46510
rect 41356 46498 41412 46508
rect 41132 45054 41134 45106
rect 41186 45054 41188 45106
rect 41132 44546 41188 45054
rect 41580 45108 41636 47406
rect 41692 47460 41748 48300
rect 41692 47394 41748 47404
rect 42028 47572 42084 49084
rect 42140 49138 42196 49308
rect 42140 49086 42142 49138
rect 42194 49086 42196 49138
rect 42140 49074 42196 49086
rect 42140 47572 42196 47582
rect 42028 47570 42196 47572
rect 42028 47518 42142 47570
rect 42194 47518 42196 47570
rect 42028 47516 42196 47518
rect 42028 47012 42084 47516
rect 42140 47506 42196 47516
rect 42252 47348 42308 49420
rect 42476 48692 42532 48702
rect 42476 48466 42532 48636
rect 42476 48414 42478 48466
rect 42530 48414 42532 48466
rect 42476 48402 42532 48414
rect 42588 48466 42644 49758
rect 42588 48414 42590 48466
rect 42642 48414 42644 48466
rect 42588 48402 42644 48414
rect 42924 49700 42980 49710
rect 43148 49700 43204 51324
rect 43484 51314 43540 51324
rect 43596 50594 43652 52780
rect 43596 50542 43598 50594
rect 43650 50542 43652 50594
rect 43596 50530 43652 50542
rect 43708 52834 43876 52836
rect 43708 52782 43822 52834
rect 43874 52782 43876 52834
rect 43708 52780 43876 52782
rect 43708 50260 43764 52780
rect 43820 52770 43876 52780
rect 44156 52834 44212 53340
rect 44716 53284 44772 54012
rect 44828 54002 44884 54012
rect 45052 53844 45108 53854
rect 44940 53732 44996 53742
rect 44940 53638 44996 53676
rect 44156 52782 44158 52834
rect 44210 52782 44212 52834
rect 44156 52276 44212 52782
rect 44156 52210 44212 52220
rect 44268 53228 44772 53284
rect 44268 52162 44324 53228
rect 44268 52110 44270 52162
rect 44322 52110 44324 52162
rect 44268 52098 44324 52110
rect 44380 53060 44436 53070
rect 43932 52052 43988 52062
rect 43820 52050 43988 52052
rect 43820 51998 43934 52050
rect 43986 51998 43988 52050
rect 43820 51996 43988 51998
rect 43820 50818 43876 51996
rect 43932 51986 43988 51996
rect 44044 51938 44100 51950
rect 44044 51886 44046 51938
rect 44098 51886 44100 51938
rect 44044 51492 44100 51886
rect 44044 51426 44100 51436
rect 44268 51940 44324 51950
rect 44156 51380 44212 51390
rect 44268 51380 44324 51884
rect 44156 51378 44324 51380
rect 44156 51326 44158 51378
rect 44210 51326 44324 51378
rect 44156 51324 44324 51326
rect 44156 51314 44212 51324
rect 43932 51268 43988 51278
rect 43932 51174 43988 51212
rect 43820 50766 43822 50818
rect 43874 50766 43876 50818
rect 43820 50754 43876 50766
rect 43708 50194 43764 50204
rect 42924 49698 43204 49700
rect 42924 49646 42926 49698
rect 42978 49646 43204 49698
rect 42924 49644 43204 49646
rect 42364 48356 42420 48366
rect 42364 48262 42420 48300
rect 42924 48354 42980 49644
rect 44380 49588 44436 53004
rect 44604 52946 44660 52958
rect 44604 52894 44606 52946
rect 44658 52894 44660 52946
rect 44604 52052 44660 52894
rect 44492 51154 44548 51166
rect 44492 51102 44494 51154
rect 44546 51102 44548 51154
rect 44492 49812 44548 51102
rect 44604 50484 44660 51996
rect 44604 50418 44660 50428
rect 44716 51828 44772 53228
rect 44828 53284 44884 53294
rect 44828 52164 44884 53228
rect 44828 52050 44884 52108
rect 44828 51998 44830 52050
rect 44882 51998 44884 52050
rect 44828 51986 44884 51998
rect 44716 51772 44996 51828
rect 44716 50148 44772 51772
rect 44940 51602 44996 51772
rect 44940 51550 44942 51602
rect 44994 51550 44996 51602
rect 44940 51538 44996 51550
rect 45052 51380 45108 53788
rect 45164 53172 45220 59276
rect 45920 59200 46032 60000
rect 45276 55412 45332 55422
rect 45276 55318 45332 55356
rect 45500 54852 45556 54862
rect 45276 53844 45332 53854
rect 45276 53750 45332 53788
rect 45500 53396 45556 54796
rect 45724 54740 45780 54750
rect 45724 54646 45780 54684
rect 45500 53340 45780 53396
rect 45612 53172 45668 53182
rect 45164 53170 45668 53172
rect 45164 53118 45614 53170
rect 45666 53118 45668 53170
rect 45164 53116 45668 53118
rect 45612 53106 45668 53116
rect 45164 52276 45220 52286
rect 45164 51938 45220 52220
rect 45612 52164 45668 52174
rect 45612 52070 45668 52108
rect 45164 51886 45166 51938
rect 45218 51886 45220 51938
rect 45164 51492 45220 51886
rect 45164 51436 45444 51492
rect 45052 51324 45220 51380
rect 45052 50484 45108 50494
rect 45052 50260 45108 50428
rect 45164 50482 45220 51324
rect 45164 50430 45166 50482
rect 45218 50430 45220 50482
rect 45164 50418 45220 50430
rect 45276 51268 45332 51278
rect 45052 50204 45220 50260
rect 44716 50082 44772 50092
rect 44492 49746 44548 49756
rect 45052 49700 45108 49710
rect 45052 49606 45108 49644
rect 44380 49522 44436 49532
rect 45052 49252 45108 49262
rect 45164 49252 45220 50204
rect 45052 49250 45220 49252
rect 45052 49198 45054 49250
rect 45106 49198 45220 49250
rect 45052 49196 45220 49198
rect 45052 49186 45108 49196
rect 44268 49138 44324 49150
rect 44268 49086 44270 49138
rect 44322 49086 44324 49138
rect 44268 48692 44324 49086
rect 44828 49028 44884 49038
rect 45276 49028 45332 51212
rect 45388 50596 45444 51436
rect 45500 50596 45556 50606
rect 45388 50594 45556 50596
rect 45388 50542 45502 50594
rect 45554 50542 45556 50594
rect 45388 50540 45556 50542
rect 45500 50530 45556 50540
rect 45388 49252 45444 49262
rect 45388 49158 45444 49196
rect 44828 49026 45332 49028
rect 44828 48974 44830 49026
rect 44882 48974 45332 49026
rect 44828 48972 45332 48974
rect 44828 48962 44884 48972
rect 44268 48626 44324 48636
rect 44940 48692 44996 48702
rect 43372 48468 43428 48478
rect 43372 48374 43428 48412
rect 44044 48468 44100 48478
rect 44492 48468 44548 48478
rect 44940 48468 44996 48636
rect 44100 48466 44996 48468
rect 44100 48414 44494 48466
rect 44546 48414 44942 48466
rect 44994 48414 44996 48466
rect 44100 48412 44996 48414
rect 44044 48374 44100 48412
rect 44492 48402 44548 48412
rect 42924 48302 42926 48354
rect 42978 48302 42980 48354
rect 42924 48290 42980 48302
rect 42700 48242 42756 48254
rect 42700 48190 42702 48242
rect 42754 48190 42756 48242
rect 42700 47572 42756 48190
rect 41916 46956 42028 47012
rect 41916 46002 41972 46956
rect 42028 46946 42084 46956
rect 42140 47292 42308 47348
rect 42364 47516 42756 47572
rect 41916 45950 41918 46002
rect 41970 45950 41972 46002
rect 41916 45938 41972 45950
rect 41580 45014 41636 45052
rect 42028 44996 42084 45006
rect 42140 44996 42196 47292
rect 42364 47236 42420 47516
rect 42812 47404 43092 47460
rect 42364 47124 42420 47180
rect 42028 44994 42196 44996
rect 42028 44942 42030 44994
rect 42082 44942 42196 44994
rect 42028 44940 42196 44942
rect 42252 47068 42420 47124
rect 42476 47346 42532 47358
rect 42476 47294 42478 47346
rect 42530 47294 42532 47346
rect 42476 47124 42532 47294
rect 42028 44884 42084 44940
rect 42028 44818 42084 44828
rect 41132 44494 41134 44546
rect 41186 44494 41188 44546
rect 41132 44482 41188 44494
rect 40236 44370 40292 44380
rect 41916 44436 41972 44446
rect 40796 44322 40852 44334
rect 40796 44270 40798 44322
rect 40850 44270 40852 44322
rect 40236 44098 40292 44110
rect 40236 44046 40238 44098
rect 40290 44046 40292 44098
rect 40236 43876 40292 44046
rect 40236 43810 40292 43820
rect 40796 43708 40852 44270
rect 41132 44324 41188 44334
rect 41132 44230 41188 44268
rect 41580 44324 41636 44334
rect 41580 44230 41636 44268
rect 41916 44322 41972 44380
rect 41916 44270 41918 44322
rect 41970 44270 41972 44322
rect 41916 44258 41972 44270
rect 41692 44098 41748 44110
rect 41692 44046 41694 44098
rect 41746 44046 41748 44098
rect 41020 43764 41076 43774
rect 40124 43374 40126 43426
rect 40178 43374 40180 43426
rect 40124 43316 40180 43374
rect 40124 43250 40180 43260
rect 40460 43652 40964 43708
rect 40012 42814 40014 42866
rect 40066 42814 40068 42866
rect 40012 42802 40068 42814
rect 40236 42980 40292 42990
rect 40236 42866 40292 42924
rect 40236 42814 40238 42866
rect 40290 42814 40292 42866
rect 40236 42802 40292 42814
rect 39676 42642 39956 42644
rect 39676 42590 39678 42642
rect 39730 42590 39956 42642
rect 39676 42588 39956 42590
rect 39564 41188 39620 41198
rect 39676 41188 39732 42588
rect 40012 42530 40068 42542
rect 40012 42478 40014 42530
rect 40066 42478 40068 42530
rect 40012 42082 40068 42478
rect 40012 42030 40014 42082
rect 40066 42030 40068 42082
rect 40012 42018 40068 42030
rect 40124 41748 40180 41758
rect 40124 41654 40180 41692
rect 39620 41132 39732 41188
rect 39564 41122 39620 41132
rect 40348 40964 40404 40974
rect 40348 40290 40404 40908
rect 40348 40238 40350 40290
rect 40402 40238 40404 40290
rect 40348 40226 40404 40238
rect 39116 39566 39118 39618
rect 39170 39566 39172 39618
rect 39116 39554 39172 39566
rect 39340 39564 39508 39620
rect 39004 38834 39172 38836
rect 39004 38782 39006 38834
rect 39058 38782 39172 38834
rect 39004 38780 39172 38782
rect 39004 38770 39060 38780
rect 38892 38724 38948 38734
rect 38332 38612 38612 38668
rect 37548 37826 37604 37838
rect 37548 37774 37550 37826
rect 37602 37774 37604 37826
rect 37548 37604 37604 37774
rect 37548 37538 37604 37548
rect 37884 37826 37940 38612
rect 37884 37774 37886 37826
rect 37938 37774 37940 37826
rect 37436 37426 37492 37436
rect 37884 37490 37940 37774
rect 38220 37828 38276 37838
rect 38220 37734 38276 37772
rect 37884 37438 37886 37490
rect 37938 37438 37940 37490
rect 37884 37426 37940 37438
rect 38220 37492 38276 37502
rect 38220 37156 38276 37436
rect 38556 37492 38612 38612
rect 38556 37398 38612 37436
rect 38780 38164 38836 38174
rect 38780 38050 38836 38108
rect 38780 37998 38782 38050
rect 38834 37998 38836 38050
rect 38780 37156 38836 37998
rect 38220 37100 38836 37156
rect 38892 37266 38948 38668
rect 38892 37214 38894 37266
rect 38946 37214 38948 37266
rect 38556 36596 38612 37100
rect 38892 36820 38948 37214
rect 39116 36820 39172 38780
rect 39228 37492 39284 37502
rect 39228 37398 39284 37436
rect 38892 36764 39060 36820
rect 39116 36764 39284 36820
rect 38556 36594 38724 36596
rect 38556 36542 38558 36594
rect 38610 36542 38724 36594
rect 38556 36540 38724 36542
rect 38556 36502 38612 36540
rect 38668 36484 38724 36540
rect 38892 36484 38948 36494
rect 38668 36482 38948 36484
rect 38668 36430 38894 36482
rect 38946 36430 38948 36482
rect 38668 36428 38948 36430
rect 38892 36418 38948 36428
rect 37772 36260 37828 36270
rect 37772 35810 37828 36204
rect 37772 35758 37774 35810
rect 37826 35758 37828 35810
rect 37772 35746 37828 35758
rect 38556 35698 38612 35710
rect 38556 35646 38558 35698
rect 38610 35646 38612 35698
rect 38556 35252 38612 35646
rect 38556 35186 38612 35196
rect 38892 35698 38948 35710
rect 38892 35646 38894 35698
rect 38946 35646 38948 35698
rect 37436 34914 37492 34926
rect 37436 34862 37438 34914
rect 37490 34862 37492 34914
rect 37436 34692 37492 34862
rect 38444 34916 38500 34926
rect 38556 34916 38612 34926
rect 38444 34914 38556 34916
rect 38444 34862 38446 34914
rect 38498 34862 38556 34914
rect 38444 34860 38556 34862
rect 38444 34850 38500 34860
rect 37436 34626 37492 34636
rect 37884 34692 37940 34702
rect 37884 34598 37940 34636
rect 37324 34412 37716 34468
rect 37324 34244 37380 34254
rect 37212 34132 37268 34142
rect 36988 33618 37044 33628
rect 37100 34130 37268 34132
rect 37100 34078 37214 34130
rect 37266 34078 37268 34130
rect 37100 34076 37268 34078
rect 37324 34132 37380 34188
rect 37324 34076 37492 34132
rect 36092 31686 36148 31724
rect 36316 31724 36820 31780
rect 36988 33458 37044 33470
rect 36988 33406 36990 33458
rect 37042 33406 37044 33458
rect 35980 30884 36036 30894
rect 35084 30324 35140 30716
rect 35420 30706 35476 30716
rect 35532 30882 36036 30884
rect 35532 30830 35982 30882
rect 36034 30830 36036 30882
rect 35532 30828 36036 30830
rect 35196 30604 35460 30614
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35196 30538 35460 30548
rect 35084 30268 35252 30324
rect 35084 30100 35140 30110
rect 34748 29596 35028 29652
rect 34524 29540 34580 29550
rect 34524 29426 34580 29484
rect 34524 29374 34526 29426
rect 34578 29374 34580 29426
rect 34524 29362 34580 29374
rect 34748 29428 34804 29438
rect 34636 28644 34692 28654
rect 34748 28644 34804 29372
rect 34636 28642 34804 28644
rect 34636 28590 34638 28642
rect 34690 28590 34804 28642
rect 34636 28588 34804 28590
rect 34972 28754 35028 29596
rect 35084 29538 35140 30044
rect 35084 29486 35086 29538
rect 35138 29486 35140 29538
rect 35084 29474 35140 29486
rect 35196 29204 35252 30268
rect 35532 30210 35588 30828
rect 35980 30818 36036 30828
rect 36092 30772 36148 30782
rect 35980 30436 36036 30446
rect 35756 30324 35812 30334
rect 35756 30230 35812 30268
rect 35532 30158 35534 30210
rect 35586 30158 35588 30210
rect 35532 30100 35588 30158
rect 35532 30034 35588 30044
rect 35420 29428 35476 29438
rect 35420 29426 35588 29428
rect 35420 29374 35422 29426
rect 35474 29374 35588 29426
rect 35420 29372 35588 29374
rect 35420 29362 35476 29372
rect 34972 28702 34974 28754
rect 35026 28702 35028 28754
rect 34636 28578 34692 28588
rect 34972 28308 35028 28702
rect 34972 28242 35028 28252
rect 35084 29148 35252 29204
rect 34412 27906 34468 27916
rect 34748 27860 34804 27870
rect 35084 27860 35140 29148
rect 35196 29036 35460 29046
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35196 28970 35460 28980
rect 35420 28756 35476 28766
rect 35420 28662 35476 28700
rect 35532 28084 35588 29372
rect 35868 29426 35924 29438
rect 35868 29374 35870 29426
rect 35922 29374 35924 29426
rect 35644 28868 35700 28878
rect 35644 28774 35700 28812
rect 35532 28018 35588 28028
rect 35644 28196 35700 28206
rect 35868 28196 35924 29374
rect 35980 28866 36036 30380
rect 36092 29650 36148 30716
rect 36092 29598 36094 29650
rect 36146 29598 36148 29650
rect 36092 29586 36148 29598
rect 35980 28814 35982 28866
rect 36034 28814 36036 28866
rect 35980 28802 36036 28814
rect 35700 28140 35924 28196
rect 35644 28082 35700 28140
rect 35644 28030 35646 28082
rect 35698 28030 35700 28082
rect 35644 28018 35700 28030
rect 33516 27806 33518 27858
rect 33570 27806 33572 27858
rect 33516 27794 33572 27806
rect 34636 27858 34804 27860
rect 34636 27806 34750 27858
rect 34802 27806 34804 27858
rect 34636 27804 34804 27806
rect 34412 27748 34468 27758
rect 34412 27654 34468 27692
rect 34636 27300 34692 27804
rect 34748 27794 34804 27804
rect 34972 27804 35140 27860
rect 34748 27636 34804 27646
rect 34748 27542 34804 27580
rect 34636 27234 34692 27244
rect 32956 26852 33124 26908
rect 33404 26852 33572 26908
rect 33068 26514 33124 26852
rect 33068 26462 33070 26514
rect 33122 26462 33124 26514
rect 33068 23940 33124 26462
rect 33180 26292 33236 26302
rect 33180 25620 33236 26236
rect 33180 24722 33236 25564
rect 33180 24670 33182 24722
rect 33234 24670 33236 24722
rect 33180 24658 33236 24670
rect 33516 26178 33572 26852
rect 34860 26516 34916 26526
rect 34972 26516 35028 27804
rect 36204 27748 36260 27758
rect 36092 27746 36260 27748
rect 36092 27694 36206 27746
rect 36258 27694 36260 27746
rect 36092 27692 36260 27694
rect 35084 27636 35140 27646
rect 35084 27542 35140 27580
rect 35868 27636 35924 27646
rect 35196 27468 35460 27478
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35196 27402 35460 27412
rect 34860 26514 35028 26516
rect 34860 26462 34862 26514
rect 34914 26462 35028 26514
rect 34860 26460 35028 26462
rect 35196 27300 35252 27310
rect 35196 27076 35252 27244
rect 35420 27188 35476 27198
rect 35420 27186 35700 27188
rect 35420 27134 35422 27186
rect 35474 27134 35700 27186
rect 35420 27132 35700 27134
rect 35420 27122 35476 27132
rect 35196 26514 35252 27020
rect 35196 26462 35198 26514
rect 35250 26462 35252 26514
rect 34860 26292 34916 26460
rect 35196 26450 35252 26462
rect 35532 26852 35588 26862
rect 34636 26236 34916 26292
rect 33516 26126 33518 26178
rect 33570 26126 33572 26178
rect 33068 23874 33124 23884
rect 33516 23716 33572 26126
rect 34076 26178 34132 26190
rect 34076 26126 34078 26178
rect 34130 26126 34132 26178
rect 33628 25732 33684 25742
rect 33628 25618 33684 25676
rect 33628 25566 33630 25618
rect 33682 25566 33684 25618
rect 33628 25554 33684 25566
rect 34076 25620 34132 26126
rect 34524 25620 34580 25630
rect 34076 25526 34132 25564
rect 34188 25618 34580 25620
rect 34188 25566 34526 25618
rect 34578 25566 34580 25618
rect 34188 25564 34580 25566
rect 34188 24948 34244 25564
rect 34524 25554 34580 25564
rect 33852 24892 34244 24948
rect 34524 25396 34580 25406
rect 33852 24834 33908 24892
rect 33852 24782 33854 24834
rect 33906 24782 33908 24834
rect 33852 24770 33908 24782
rect 33516 23650 33572 23660
rect 34188 22482 34244 22494
rect 34188 22430 34190 22482
rect 34242 22430 34244 22482
rect 33852 22370 33908 22382
rect 33852 22318 33854 22370
rect 33906 22318 33908 22370
rect 32956 22148 33012 22158
rect 33404 22148 33460 22158
rect 33852 22148 33908 22318
rect 34188 22372 34244 22430
rect 34188 22306 34244 22316
rect 32956 22146 33908 22148
rect 32956 22094 32958 22146
rect 33010 22094 33406 22146
rect 33458 22094 33908 22146
rect 32956 22092 33908 22094
rect 32956 22082 33012 22092
rect 33404 22082 33460 22092
rect 33852 20580 33908 22092
rect 33964 21588 34020 21598
rect 34020 21532 34132 21588
rect 33964 21522 34020 21532
rect 33852 20514 33908 20524
rect 33628 20356 33684 20366
rect 33180 19346 33236 19358
rect 33180 19294 33182 19346
rect 33234 19294 33236 19346
rect 33180 18674 33236 19294
rect 33292 19348 33348 19358
rect 33292 19234 33348 19292
rect 33292 19182 33294 19234
rect 33346 19182 33348 19234
rect 33292 19170 33348 19182
rect 33180 18622 33182 18674
rect 33234 18622 33236 18674
rect 33180 18610 33236 18622
rect 31948 18508 32900 18564
rect 31948 18450 32004 18508
rect 31948 18398 31950 18450
rect 32002 18398 32004 18450
rect 31948 18386 32004 18398
rect 32844 18452 32900 18508
rect 32956 18452 33012 18462
rect 32844 18450 33012 18452
rect 32844 18398 32958 18450
rect 33010 18398 33012 18450
rect 32844 18396 33012 18398
rect 32956 18386 33012 18396
rect 33292 18452 33348 18462
rect 33292 18358 33348 18396
rect 33628 18450 33684 20300
rect 33740 20132 33796 20142
rect 33740 20038 33796 20076
rect 33964 20132 34020 20142
rect 34076 20132 34132 21532
rect 34412 20914 34468 20926
rect 34412 20862 34414 20914
rect 34466 20862 34468 20914
rect 34188 20356 34244 20366
rect 34412 20356 34468 20862
rect 34244 20300 34468 20356
rect 34188 20290 34244 20300
rect 34524 20244 34580 25340
rect 34636 25394 34692 26236
rect 34636 25342 34638 25394
rect 34690 25342 34692 25394
rect 34636 25330 34692 25342
rect 34748 26068 34804 26078
rect 34636 23940 34692 23950
rect 34636 23846 34692 23884
rect 34636 22370 34692 22382
rect 34636 22318 34638 22370
rect 34690 22318 34692 22370
rect 34636 21812 34692 22318
rect 34748 22260 34804 26012
rect 35532 26066 35588 26796
rect 35644 26628 35700 27132
rect 35868 27186 35924 27580
rect 35868 27134 35870 27186
rect 35922 27134 35924 27186
rect 35868 27122 35924 27134
rect 36092 26964 36148 27692
rect 36204 27682 36260 27692
rect 36092 26898 36148 26908
rect 36316 26908 36372 31724
rect 36988 31668 37044 33406
rect 36988 31218 37044 31612
rect 36988 31166 36990 31218
rect 37042 31166 37044 31218
rect 36540 30884 36596 30894
rect 36428 29988 36484 29998
rect 36428 29894 36484 29932
rect 36428 28756 36484 28766
rect 36540 28756 36596 30828
rect 36764 29426 36820 29438
rect 36764 29374 36766 29426
rect 36818 29374 36820 29426
rect 36428 28754 36708 28756
rect 36428 28702 36430 28754
rect 36482 28702 36708 28754
rect 36428 28700 36708 28702
rect 36428 28690 36484 28700
rect 35756 26852 35812 26862
rect 35756 26758 35812 26796
rect 35980 26850 36036 26862
rect 35980 26798 35982 26850
rect 36034 26798 36036 26850
rect 35980 26628 36036 26798
rect 35644 26572 36036 26628
rect 36204 26850 36260 26862
rect 36316 26852 36596 26908
rect 36204 26798 36206 26850
rect 36258 26798 36260 26850
rect 35756 26290 35812 26572
rect 35756 26238 35758 26290
rect 35810 26238 35812 26290
rect 35756 26226 35812 26238
rect 36204 26180 36260 26798
rect 36204 26178 36372 26180
rect 36204 26126 36206 26178
rect 36258 26126 36372 26178
rect 36204 26124 36372 26126
rect 36204 26114 36260 26124
rect 35532 26014 35534 26066
rect 35586 26014 35588 26066
rect 35196 25900 35460 25910
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35196 25834 35460 25844
rect 35532 25508 35588 26014
rect 35532 25414 35588 25452
rect 35980 25620 36036 25630
rect 34860 25396 34916 25406
rect 35644 25396 35700 25406
rect 35868 25396 35924 25406
rect 34860 25394 35140 25396
rect 34860 25342 34862 25394
rect 34914 25342 35140 25394
rect 34860 25340 35140 25342
rect 34860 25330 34916 25340
rect 34860 25060 34916 25070
rect 34860 22708 34916 25004
rect 35084 24050 35140 25340
rect 35644 25394 35924 25396
rect 35644 25342 35646 25394
rect 35698 25342 35870 25394
rect 35922 25342 35924 25394
rect 35644 25340 35924 25342
rect 35644 25330 35700 25340
rect 35868 25330 35924 25340
rect 35980 25394 36036 25564
rect 35980 25342 35982 25394
rect 36034 25342 36036 25394
rect 35980 25330 36036 25342
rect 36204 25282 36260 25294
rect 36204 25230 36206 25282
rect 36258 25230 36260 25282
rect 35868 25172 35924 25182
rect 35196 24332 35460 24342
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35196 24266 35460 24276
rect 35084 23998 35086 24050
rect 35138 23998 35140 24050
rect 35084 23986 35140 23998
rect 35868 24052 35924 25116
rect 35980 24612 36036 24622
rect 36204 24612 36260 25230
rect 36316 25172 36372 26124
rect 36428 26066 36484 26078
rect 36428 26014 36430 26066
rect 36482 26014 36484 26066
rect 36428 25396 36484 26014
rect 36428 25302 36484 25340
rect 36316 25116 36484 25172
rect 35980 24610 36260 24612
rect 35980 24558 35982 24610
rect 36034 24558 36260 24610
rect 35980 24556 36260 24558
rect 36316 24612 36372 24622
rect 35980 24546 36036 24556
rect 35980 24052 36036 24062
rect 35868 24050 36036 24052
rect 35868 23998 35982 24050
rect 36034 23998 36036 24050
rect 35868 23996 36036 23998
rect 35980 23986 36036 23996
rect 34972 23938 35028 23950
rect 35756 23940 35812 23950
rect 36092 23940 36148 24556
rect 34972 23886 34974 23938
rect 35026 23886 35028 23938
rect 34972 23604 35028 23886
rect 35644 23938 35924 23940
rect 35644 23886 35758 23938
rect 35810 23886 35924 23938
rect 35644 23884 35924 23886
rect 35196 23828 35252 23838
rect 34972 23538 35028 23548
rect 35084 23772 35196 23828
rect 34860 22642 34916 22652
rect 35084 22596 35140 23772
rect 35196 23762 35252 23772
rect 35644 23826 35700 23884
rect 35756 23874 35812 23884
rect 35644 23774 35646 23826
rect 35698 23774 35700 23826
rect 35644 23762 35700 23774
rect 35532 23604 35588 23614
rect 35196 22764 35460 22774
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35196 22698 35460 22708
rect 35196 22596 35252 22606
rect 35084 22594 35252 22596
rect 35084 22542 35198 22594
rect 35250 22542 35252 22594
rect 35084 22540 35252 22542
rect 35196 22530 35252 22540
rect 34748 22194 34804 22204
rect 34860 22370 34916 22382
rect 34860 22318 34862 22370
rect 34914 22318 34916 22370
rect 34636 21746 34692 21756
rect 34860 21588 34916 22318
rect 35084 22372 35140 22382
rect 35084 22278 35140 22316
rect 35532 22260 35588 23548
rect 35868 22708 35924 23884
rect 36092 23846 36148 23884
rect 36316 23938 36372 24556
rect 36316 23886 36318 23938
rect 36370 23886 36372 23938
rect 36316 23874 36372 23886
rect 35868 22642 35924 22652
rect 36316 23492 36372 23502
rect 36316 22482 36372 23436
rect 36316 22430 36318 22482
rect 36370 22430 36372 22482
rect 35756 22372 35812 22382
rect 35532 22258 35700 22260
rect 35532 22206 35534 22258
rect 35586 22206 35700 22258
rect 35532 22204 35700 22206
rect 35532 22194 35588 22204
rect 35196 21588 35252 21598
rect 34860 21522 34916 21532
rect 35084 21586 35252 21588
rect 35084 21534 35198 21586
rect 35250 21534 35252 21586
rect 35084 21532 35252 21534
rect 34860 20692 34916 20702
rect 35084 20692 35140 21532
rect 35196 21522 35252 21532
rect 35196 21196 35460 21206
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35196 21130 35460 21140
rect 35644 20916 35700 22204
rect 35756 21028 35812 22316
rect 36316 22372 36372 22430
rect 36428 22484 36484 25116
rect 36428 22418 36484 22428
rect 36316 22306 36372 22316
rect 35868 22148 35924 22158
rect 35868 21700 35924 22092
rect 35868 21644 36372 21700
rect 35980 21476 36036 21486
rect 35980 21474 36148 21476
rect 35980 21422 35982 21474
rect 36034 21422 36148 21474
rect 35980 21420 36148 21422
rect 35980 21410 36036 21420
rect 35756 20934 35812 20972
rect 35420 20860 35700 20916
rect 36092 20914 36148 21420
rect 36092 20862 36094 20914
rect 36146 20862 36148 20914
rect 34916 20636 35140 20692
rect 35308 20690 35364 20702
rect 35308 20638 35310 20690
rect 35362 20638 35364 20690
rect 34860 20598 34916 20636
rect 33964 20130 34132 20132
rect 33964 20078 33966 20130
rect 34018 20078 34132 20130
rect 33964 20076 34132 20078
rect 34300 20188 34580 20244
rect 34972 20244 35028 20636
rect 33964 20066 34020 20076
rect 33852 19906 33908 19918
rect 33852 19854 33854 19906
rect 33906 19854 33908 19906
rect 33628 18398 33630 18450
rect 33682 18398 33684 18450
rect 32508 18338 32564 18350
rect 32508 18286 32510 18338
rect 32562 18286 32564 18338
rect 31836 18172 32004 18228
rect 31724 18004 31780 18014
rect 31724 17108 31780 17948
rect 30828 17054 30830 17106
rect 30882 17054 30884 17106
rect 30828 17042 30884 17054
rect 31052 17052 31556 17108
rect 31612 17106 31780 17108
rect 31612 17054 31726 17106
rect 31778 17054 31780 17106
rect 31612 17052 31780 17054
rect 30828 16660 30884 16670
rect 30716 16658 30884 16660
rect 30716 16606 30830 16658
rect 30882 16606 30884 16658
rect 30716 16604 30884 16606
rect 30716 15426 30772 16604
rect 30828 16594 30884 16604
rect 30716 15374 30718 15426
rect 30770 15374 30772 15426
rect 30716 15362 30772 15374
rect 30940 15428 30996 15438
rect 30156 15314 30660 15316
rect 30156 15262 30158 15314
rect 30210 15262 30660 15314
rect 30156 15260 30660 15262
rect 30156 15250 30212 15260
rect 29820 15092 29988 15148
rect 29820 12628 29876 15092
rect 30268 14754 30324 14766
rect 30268 14702 30270 14754
rect 30322 14702 30324 14754
rect 30044 14306 30100 14318
rect 30044 14254 30046 14306
rect 30098 14254 30100 14306
rect 30044 14084 30100 14254
rect 29932 13748 29988 13758
rect 30044 13748 30100 14028
rect 29932 13746 30100 13748
rect 29932 13694 29934 13746
rect 29986 13694 30100 13746
rect 29932 13692 30100 13694
rect 29932 13682 29988 13692
rect 30268 13634 30324 14702
rect 30492 14644 30548 14654
rect 30492 14550 30548 14588
rect 30268 13582 30270 13634
rect 30322 13582 30324 13634
rect 30268 13300 30324 13582
rect 30268 13234 30324 13244
rect 29820 12562 29876 12572
rect 29932 12852 29988 12862
rect 29484 11676 29764 11732
rect 29148 11118 29150 11170
rect 29202 11118 29204 11170
rect 29148 11106 29204 11118
rect 29260 11170 29316 11182
rect 29260 11118 29262 11170
rect 29314 11118 29316 11170
rect 29260 10948 29316 11118
rect 29036 10892 29316 10948
rect 29372 11170 29428 11182
rect 29372 11118 29374 11170
rect 29426 11118 29428 11170
rect 29372 10836 29428 11118
rect 28140 10658 28196 10668
rect 29036 10780 29428 10836
rect 28028 10546 28084 10556
rect 28812 10500 28868 10510
rect 29036 10500 29092 10780
rect 29484 10724 29540 11676
rect 29596 11172 29652 11182
rect 29596 11078 29652 11116
rect 29372 10722 29540 10724
rect 29372 10670 29486 10722
rect 29538 10670 29540 10722
rect 29372 10668 29540 10670
rect 29148 10612 29204 10622
rect 29148 10518 29204 10556
rect 28588 10498 29092 10500
rect 28588 10446 28814 10498
rect 28866 10446 29092 10498
rect 28588 10444 29092 10446
rect 29260 10500 29316 10510
rect 28588 10164 28644 10444
rect 28812 10434 28868 10444
rect 29260 10406 29316 10444
rect 29372 10276 29428 10668
rect 29484 10658 29540 10668
rect 29820 10836 29876 10846
rect 29708 10612 29764 10622
rect 29820 10612 29876 10780
rect 29708 10610 29876 10612
rect 29708 10558 29710 10610
rect 29762 10558 29876 10610
rect 29708 10556 29876 10558
rect 29708 10546 29764 10556
rect 28588 10098 28644 10108
rect 28700 10220 29428 10276
rect 28700 9938 28756 10220
rect 28700 9886 28702 9938
rect 28754 9886 28756 9938
rect 28700 9874 28756 9886
rect 29596 9828 29652 9838
rect 29932 9828 29988 12796
rect 30044 12852 30100 12862
rect 30044 12850 30324 12852
rect 30044 12798 30046 12850
rect 30098 12798 30324 12850
rect 30044 12796 30324 12798
rect 30044 12786 30100 12796
rect 30156 12628 30212 12638
rect 30044 12516 30100 12526
rect 30044 12068 30100 12460
rect 30156 12290 30212 12572
rect 30156 12238 30158 12290
rect 30210 12238 30212 12290
rect 30156 12226 30212 12238
rect 30268 12068 30324 12796
rect 30604 12628 30660 15260
rect 30940 15314 30996 15372
rect 30940 15262 30942 15314
rect 30994 15262 30996 15314
rect 30940 15250 30996 15262
rect 30828 15202 30884 15214
rect 30828 15150 30830 15202
rect 30882 15150 30884 15202
rect 30828 14420 30884 15150
rect 31052 14754 31108 17052
rect 31388 16884 31444 16894
rect 31388 16790 31444 16828
rect 31052 14702 31054 14754
rect 31106 14702 31108 14754
rect 31052 14690 31108 14702
rect 31164 16772 31220 16782
rect 30828 14354 30884 14364
rect 31052 14306 31108 14318
rect 31052 14254 31054 14306
rect 31106 14254 31108 14306
rect 30828 14084 30884 14094
rect 31052 14084 31108 14254
rect 30884 14028 31108 14084
rect 30828 13970 30884 14028
rect 30828 13918 30830 13970
rect 30882 13918 30884 13970
rect 30828 13906 30884 13918
rect 30604 12572 31108 12628
rect 30380 12292 30436 12302
rect 30380 12198 30436 12236
rect 30492 12234 30548 12246
rect 30492 12182 30494 12234
rect 30546 12182 30548 12234
rect 30492 12180 30548 12182
rect 30604 12180 30660 12190
rect 30492 12124 30604 12180
rect 30604 12114 30660 12124
rect 30716 12180 30772 12190
rect 30716 12178 30884 12180
rect 30716 12126 30718 12178
rect 30770 12126 30884 12178
rect 30716 12124 30884 12126
rect 30716 12114 30772 12124
rect 30380 12068 30436 12078
rect 30044 12012 30212 12068
rect 30268 12066 30436 12068
rect 30268 12014 30382 12066
rect 30434 12014 30436 12066
rect 30268 12012 30436 12014
rect 30044 11844 30100 11854
rect 30044 10610 30100 11788
rect 30156 11788 30212 12012
rect 30380 12002 30436 12012
rect 30156 11732 30548 11788
rect 30156 10836 30212 10846
rect 30156 10742 30212 10780
rect 30268 10612 30324 10622
rect 30044 10558 30046 10610
rect 30098 10558 30100 10610
rect 30044 10546 30100 10558
rect 30156 10610 30324 10612
rect 30156 10558 30270 10610
rect 30322 10558 30324 10610
rect 30156 10556 30324 10558
rect 29596 9826 29988 9828
rect 29596 9774 29598 9826
rect 29650 9774 29988 9826
rect 29596 9772 29988 9774
rect 29596 9762 29652 9772
rect 30156 9044 30212 10556
rect 30268 10546 30324 10556
rect 30268 9716 30324 9726
rect 30268 9622 30324 9660
rect 29596 8988 30212 9044
rect 29596 8930 29652 8988
rect 29596 8878 29598 8930
rect 29650 8878 29652 8930
rect 29036 7700 29092 7710
rect 28924 7588 28980 7598
rect 28924 7494 28980 7532
rect 27916 7422 27918 7474
rect 27970 7422 27972 7474
rect 27916 7410 27972 7422
rect 27580 7084 27860 7140
rect 27356 6804 27412 6814
rect 27020 6638 27022 6690
rect 27074 6638 27076 6690
rect 27020 6626 27076 6638
rect 27244 6748 27356 6804
rect 26684 6580 26740 6590
rect 26684 6018 26740 6524
rect 26684 5966 26686 6018
rect 26738 5966 26740 6018
rect 26684 5954 26740 5966
rect 27020 6244 27076 6254
rect 27020 6018 27076 6188
rect 27020 5966 27022 6018
rect 27074 5966 27076 6018
rect 27020 5684 27076 5966
rect 27244 6018 27300 6748
rect 27356 6738 27412 6748
rect 27468 6692 27524 6702
rect 27580 6692 27636 7084
rect 27468 6690 27636 6692
rect 27468 6638 27470 6690
rect 27522 6638 27636 6690
rect 27468 6636 27636 6638
rect 27692 6804 27748 6814
rect 27692 6690 27748 6748
rect 28476 6804 28532 6814
rect 27692 6638 27694 6690
rect 27746 6638 27748 6690
rect 27468 6626 27524 6636
rect 27692 6626 27748 6638
rect 28364 6692 28420 6702
rect 28364 6598 28420 6636
rect 27244 5966 27246 6018
rect 27298 5966 27300 6018
rect 27244 5954 27300 5966
rect 27356 6466 27412 6478
rect 27356 6414 27358 6466
rect 27410 6414 27412 6466
rect 27020 5618 27076 5628
rect 27132 5906 27188 5918
rect 27132 5854 27134 5906
rect 27186 5854 27188 5906
rect 27132 5124 27188 5854
rect 27356 5908 27412 6414
rect 28028 6466 28084 6478
rect 28028 6414 28030 6466
rect 28082 6414 28084 6466
rect 27916 6132 27972 6142
rect 28028 6132 28084 6414
rect 27972 6076 28084 6132
rect 28364 6468 28420 6478
rect 27916 6038 27972 6076
rect 27356 5842 27412 5852
rect 27692 5908 27748 5918
rect 27692 5814 27748 5852
rect 28364 5906 28420 6412
rect 28364 5854 28366 5906
rect 28418 5854 28420 5906
rect 28364 5842 28420 5854
rect 27804 5796 27860 5806
rect 27804 5702 27860 5740
rect 28364 5236 28420 5246
rect 28476 5236 28532 6748
rect 28588 6690 28644 6702
rect 28588 6638 28590 6690
rect 28642 6638 28644 6690
rect 28588 6580 28644 6638
rect 29036 6690 29092 7644
rect 29036 6638 29038 6690
rect 29090 6638 29092 6690
rect 29036 6626 29092 6638
rect 29260 6692 29316 6702
rect 29260 6598 29316 6636
rect 29484 6692 29540 6702
rect 29596 6692 29652 8878
rect 30268 8258 30324 8270
rect 30268 8206 30270 8258
rect 30322 8206 30324 8258
rect 30268 7700 30324 8206
rect 30492 8146 30548 11732
rect 30716 11172 30772 11182
rect 30716 10724 30772 11116
rect 30716 10610 30772 10668
rect 30716 10558 30718 10610
rect 30770 10558 30772 10610
rect 30716 10546 30772 10558
rect 30828 10612 30884 12124
rect 30940 12178 30996 12190
rect 30940 12126 30942 12178
rect 30994 12126 30996 12178
rect 30940 11956 30996 12126
rect 30940 11890 30996 11900
rect 31052 11732 31108 12572
rect 31164 12290 31220 16716
rect 31612 16658 31668 17052
rect 31724 17042 31780 17052
rect 31612 16606 31614 16658
rect 31666 16606 31668 16658
rect 31612 15538 31668 16606
rect 31948 16324 32004 18172
rect 32284 18226 32340 18238
rect 32284 18174 32286 18226
rect 32338 18174 32340 18226
rect 32284 17892 32340 18174
rect 32284 17826 32340 17836
rect 31948 16258 32004 16268
rect 32284 17444 32340 17454
rect 32284 16772 32340 17388
rect 32284 16210 32340 16716
rect 32508 16772 32564 18286
rect 33516 18340 33572 18350
rect 33404 18228 33460 18238
rect 33180 17892 33236 17902
rect 33180 17798 33236 17836
rect 32956 17780 33012 17790
rect 32956 17686 33012 17724
rect 33404 17220 33460 18172
rect 33516 17890 33572 18284
rect 33516 17838 33518 17890
rect 33570 17838 33572 17890
rect 33516 17826 33572 17838
rect 33516 17220 33572 17230
rect 33404 17164 33516 17220
rect 33292 16994 33348 17006
rect 33292 16942 33294 16994
rect 33346 16942 33348 16994
rect 32508 16716 33236 16772
rect 32508 16660 32564 16716
rect 32508 16594 32564 16604
rect 32284 16158 32286 16210
rect 32338 16158 32340 16210
rect 32284 16146 32340 16158
rect 31612 15486 31614 15538
rect 31666 15486 31668 15538
rect 31612 15474 31668 15486
rect 32172 15988 32228 15998
rect 31276 15314 31332 15326
rect 31276 15262 31278 15314
rect 31330 15262 31332 15314
rect 31276 15148 31332 15262
rect 32172 15314 32228 15932
rect 32172 15262 32174 15314
rect 32226 15262 32228 15314
rect 32172 15250 32228 15262
rect 32396 15540 32452 15550
rect 31276 15092 31444 15148
rect 31164 12238 31166 12290
rect 31218 12238 31220 12290
rect 31164 12180 31220 12238
rect 31388 14642 31444 15092
rect 31388 14590 31390 14642
rect 31442 14590 31444 14642
rect 31164 12114 31220 12124
rect 31276 12178 31332 12190
rect 31276 12126 31278 12178
rect 31330 12126 31332 12178
rect 31052 11666 31108 11676
rect 31164 11844 31220 11854
rect 31276 11844 31332 12126
rect 31388 12068 31444 14590
rect 31948 15090 32004 15102
rect 31948 15038 31950 15090
rect 32002 15038 32004 15090
rect 31948 14644 32004 15038
rect 31948 14578 32004 14588
rect 31948 14420 32004 14430
rect 31836 13972 31892 13982
rect 31836 13746 31892 13916
rect 31836 13694 31838 13746
rect 31890 13694 31892 13746
rect 31836 13682 31892 13694
rect 31948 13634 32004 14364
rect 31948 13582 31950 13634
rect 32002 13582 32004 13634
rect 31948 13570 32004 13582
rect 32172 13074 32228 13086
rect 32172 13022 32174 13074
rect 32226 13022 32228 13074
rect 31724 12516 31780 12526
rect 31612 12292 31668 12302
rect 31612 12198 31668 12236
rect 31724 12290 31780 12460
rect 32172 12516 32228 13022
rect 32172 12450 32228 12460
rect 31724 12238 31726 12290
rect 31778 12238 31780 12290
rect 31724 12226 31780 12238
rect 32172 12292 32228 12302
rect 32172 12198 32228 12236
rect 31388 12012 31668 12068
rect 31220 11788 31332 11844
rect 31164 11394 31220 11788
rect 31164 11342 31166 11394
rect 31218 11342 31220 11394
rect 31164 11330 31220 11342
rect 30940 11170 30996 11182
rect 30940 11118 30942 11170
rect 30994 11118 30996 11170
rect 30940 10724 30996 11118
rect 31052 11170 31108 11182
rect 31052 11118 31054 11170
rect 31106 11118 31108 11170
rect 31052 10836 31108 11118
rect 31052 10780 31444 10836
rect 30940 10668 31220 10724
rect 30828 10518 30884 10556
rect 31052 10498 31108 10510
rect 31052 10446 31054 10498
rect 31106 10446 31108 10498
rect 31052 9716 31108 10446
rect 31164 10052 31220 10668
rect 31276 10612 31332 10622
rect 31276 10518 31332 10556
rect 31388 10610 31444 10780
rect 31388 10558 31390 10610
rect 31442 10558 31444 10610
rect 31388 10546 31444 10558
rect 31164 9986 31220 9996
rect 31052 9650 31108 9660
rect 31500 9156 31556 9166
rect 31500 8372 31556 9100
rect 31164 8370 31556 8372
rect 31164 8318 31502 8370
rect 31554 8318 31556 8370
rect 31164 8316 31556 8318
rect 31164 8260 31220 8316
rect 31500 8306 31556 8316
rect 31612 8372 31668 12012
rect 31948 11732 32004 11742
rect 31948 10612 32004 11676
rect 32396 11508 32452 15484
rect 33068 15092 33124 15102
rect 32620 15090 33124 15092
rect 32620 15038 33070 15090
rect 33122 15038 33124 15090
rect 32620 15036 33124 15038
rect 32508 13860 32564 13870
rect 32620 13860 32676 15036
rect 33068 15026 33124 15036
rect 32508 13858 32676 13860
rect 32508 13806 32510 13858
rect 32562 13806 32676 13858
rect 32508 13804 32676 13806
rect 32732 14644 32788 14654
rect 32508 13794 32564 13804
rect 32396 11442 32452 11452
rect 32732 11618 32788 14588
rect 32732 11566 32734 11618
rect 32786 11566 32788 11618
rect 31948 10518 32004 10556
rect 32508 11394 32564 11406
rect 32508 11342 32510 11394
rect 32562 11342 32564 11394
rect 32508 10276 32564 11342
rect 32508 10210 32564 10220
rect 31612 8306 31668 8316
rect 31948 10052 32004 10062
rect 30492 8094 30494 8146
rect 30546 8094 30548 8146
rect 30492 8082 30548 8094
rect 30940 8258 31220 8260
rect 30940 8206 31166 8258
rect 31218 8206 31220 8258
rect 30940 8204 31220 8206
rect 30268 7634 30324 7644
rect 30044 7476 30100 7486
rect 30940 7476 30996 8204
rect 31164 8194 31220 8204
rect 31052 8036 31108 8046
rect 31052 8034 31332 8036
rect 31052 7982 31054 8034
rect 31106 7982 31332 8034
rect 31052 7980 31332 7982
rect 31052 7970 31108 7980
rect 31052 7476 31108 7486
rect 30940 7474 31108 7476
rect 30940 7422 31054 7474
rect 31106 7422 31108 7474
rect 30940 7420 31108 7422
rect 30044 7382 30100 7420
rect 31052 7410 31108 7420
rect 30380 7362 30436 7374
rect 30380 7310 30382 7362
rect 30434 7310 30436 7362
rect 30380 6804 30436 7310
rect 30380 6738 30436 6748
rect 30604 7250 30660 7262
rect 30604 7198 30606 7250
rect 30658 7198 30660 7250
rect 29484 6690 29652 6692
rect 29484 6638 29486 6690
rect 29538 6638 29652 6690
rect 29484 6636 29652 6638
rect 30044 6692 30100 6702
rect 29484 6626 29540 6636
rect 30044 6598 30100 6636
rect 28588 6514 28644 6524
rect 29708 6578 29764 6590
rect 29708 6526 29710 6578
rect 29762 6526 29764 6578
rect 29260 6244 29316 6254
rect 29260 6018 29316 6188
rect 29260 5966 29262 6018
rect 29314 5966 29316 6018
rect 29260 5954 29316 5966
rect 29596 6020 29652 6030
rect 29596 5926 29652 5964
rect 29036 5908 29092 5918
rect 29036 5814 29092 5852
rect 29148 5906 29204 5918
rect 29148 5854 29150 5906
rect 29202 5854 29204 5906
rect 28364 5234 28532 5236
rect 28364 5182 28366 5234
rect 28418 5182 28532 5234
rect 28364 5180 28532 5182
rect 29148 5236 29204 5854
rect 29708 5908 29764 6526
rect 30268 6580 30324 6590
rect 30268 6486 30324 6524
rect 30156 6466 30212 6478
rect 30156 6414 30158 6466
rect 30210 6414 30212 6466
rect 29708 5842 29764 5852
rect 29820 6132 29876 6142
rect 29820 5906 29876 6076
rect 29820 5854 29822 5906
rect 29874 5854 29876 5906
rect 29820 5842 29876 5854
rect 29932 5908 29988 5918
rect 30156 5908 30212 6414
rect 30492 6468 30548 6478
rect 30492 6374 30548 6412
rect 29932 5906 30212 5908
rect 29932 5854 29934 5906
rect 29986 5854 30212 5906
rect 29932 5852 30212 5854
rect 30268 5908 30324 5918
rect 30604 5908 30660 7198
rect 30324 5852 30660 5908
rect 30828 7252 30884 7262
rect 30828 5908 30884 7196
rect 31276 6804 31332 7980
rect 31612 7700 31668 7710
rect 31500 7476 31556 7486
rect 31500 7382 31556 7420
rect 31612 7474 31668 7644
rect 31612 7422 31614 7474
rect 31666 7422 31668 7474
rect 31612 7410 31668 7422
rect 31948 7474 32004 9996
rect 32396 10052 32452 10062
rect 32396 9938 32452 9996
rect 32396 9886 32398 9938
rect 32450 9886 32452 9938
rect 32396 9874 32452 9886
rect 32732 8260 32788 11566
rect 33180 11508 33236 16716
rect 33292 15988 33348 16942
rect 33516 16882 33572 17164
rect 33516 16830 33518 16882
rect 33570 16830 33572 16882
rect 33516 16818 33572 16830
rect 33628 16660 33684 18398
rect 33628 16594 33684 16604
rect 33740 19684 33796 19694
rect 33516 16100 33572 16110
rect 33292 15922 33348 15932
rect 33404 16044 33516 16100
rect 33292 15540 33348 15550
rect 33292 15446 33348 15484
rect 33404 15316 33460 16044
rect 33516 16006 33572 16044
rect 33292 15260 33460 15316
rect 33292 11620 33348 15260
rect 33740 15148 33796 19628
rect 33852 16772 33908 19854
rect 34188 19010 34244 19022
rect 34188 18958 34190 19010
rect 34242 18958 34244 19010
rect 34188 18004 34244 18958
rect 34300 18228 34356 20188
rect 34972 20178 35028 20188
rect 34748 20130 34804 20142
rect 34748 20078 34750 20130
rect 34802 20078 34804 20130
rect 34412 19908 34468 19918
rect 34412 19814 34468 19852
rect 34748 19684 34804 20078
rect 35084 20132 35140 20142
rect 35084 20038 35140 20076
rect 35308 19796 35364 20638
rect 35420 20020 35476 20860
rect 36092 20850 36148 20862
rect 35980 20802 36036 20814
rect 35980 20750 35982 20802
rect 36034 20750 36036 20802
rect 35532 20690 35588 20702
rect 35532 20638 35534 20690
rect 35586 20638 35588 20690
rect 35532 20356 35588 20638
rect 35980 20580 36036 20750
rect 36204 20692 36260 20702
rect 36204 20598 36260 20636
rect 35980 20514 36036 20524
rect 35532 20290 35588 20300
rect 35868 20356 35924 20366
rect 35924 20300 36260 20356
rect 35868 20290 35924 20300
rect 35756 20244 35812 20254
rect 35644 20132 35700 20142
rect 35756 20132 36036 20188
rect 35644 20038 35700 20076
rect 35420 19964 35588 20020
rect 35532 19908 35588 19964
rect 35868 20018 35924 20030
rect 35868 19966 35870 20018
rect 35922 19966 35924 20018
rect 35756 19908 35812 19918
rect 35868 19908 35924 19966
rect 35532 19852 35700 19908
rect 35308 19740 35588 19796
rect 34748 19618 34804 19628
rect 35196 19628 35460 19638
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35196 19562 35460 19572
rect 35532 19460 35588 19740
rect 35308 19404 35588 19460
rect 34524 19348 34580 19358
rect 34524 19254 34580 19292
rect 35308 19346 35364 19404
rect 35308 19294 35310 19346
rect 35362 19294 35364 19346
rect 35308 19282 35364 19294
rect 34748 19234 34804 19246
rect 34748 19182 34750 19234
rect 34802 19182 34804 19234
rect 34412 19122 34468 19134
rect 34412 19070 34414 19122
rect 34466 19070 34468 19122
rect 34412 18900 34468 19070
rect 34412 18834 34468 18844
rect 34636 19124 34692 19134
rect 34636 18340 34692 19068
rect 34636 18246 34692 18284
rect 34300 18162 34356 18172
rect 34748 18116 34804 19182
rect 35196 19234 35252 19246
rect 35196 19182 35198 19234
rect 35250 19182 35252 19234
rect 35084 19124 35140 19134
rect 35196 19124 35252 19182
rect 35420 19124 35476 19134
rect 35140 19068 35252 19124
rect 35308 19068 35420 19124
rect 35084 19058 35140 19068
rect 35196 18900 35252 18910
rect 35196 18676 35252 18844
rect 35084 18452 35140 18462
rect 35084 18358 35140 18396
rect 35196 18228 35252 18620
rect 35308 18452 35364 19068
rect 35420 19030 35476 19068
rect 35308 18386 35364 18396
rect 35532 18452 35588 18462
rect 35532 18358 35588 18396
rect 34636 18060 34804 18116
rect 35084 18172 35252 18228
rect 34188 17948 34468 18004
rect 33964 17892 34020 17902
rect 33964 17666 34020 17836
rect 33964 17614 33966 17666
rect 34018 17614 34020 17666
rect 33964 17602 34020 17614
rect 34188 17780 34244 17790
rect 34188 17442 34244 17724
rect 34300 17556 34356 17566
rect 34300 17462 34356 17500
rect 34188 17390 34190 17442
rect 34242 17390 34244 17442
rect 34188 17378 34244 17390
rect 34412 17332 34468 17948
rect 34636 17780 34692 18060
rect 35084 17890 35140 18172
rect 35196 18060 35460 18070
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35644 18004 35700 19852
rect 35812 19852 35924 19908
rect 35980 19908 36036 20132
rect 35756 19842 35812 19852
rect 35756 19234 35812 19246
rect 35756 19182 35758 19234
rect 35810 19182 35812 19234
rect 35756 18452 35812 19182
rect 35868 18676 35924 18714
rect 35868 18610 35924 18620
rect 35868 18452 35924 18462
rect 35756 18396 35868 18452
rect 35980 18452 36036 19852
rect 36092 20132 36148 20142
rect 36092 19460 36148 20076
rect 36092 19394 36148 19404
rect 36204 19346 36260 20300
rect 36316 20132 36372 21644
rect 36316 20066 36372 20076
rect 36204 19294 36206 19346
rect 36258 19294 36260 19346
rect 36204 19282 36260 19294
rect 36316 19796 36372 19806
rect 36092 19122 36148 19134
rect 36092 19070 36094 19122
rect 36146 19070 36148 19122
rect 36092 18676 36148 19070
rect 36316 19122 36372 19740
rect 36316 19070 36318 19122
rect 36370 19070 36372 19122
rect 36316 19058 36372 19070
rect 36092 18610 36148 18620
rect 36204 18900 36260 18910
rect 36092 18452 36148 18462
rect 35980 18450 36148 18452
rect 35980 18398 36094 18450
rect 36146 18398 36148 18450
rect 35980 18396 36148 18398
rect 35196 17994 35460 18004
rect 35532 17948 35700 18004
rect 35084 17838 35086 17890
rect 35138 17838 35140 17890
rect 35084 17826 35140 17838
rect 35308 17892 35364 17902
rect 35532 17892 35588 17948
rect 35308 17890 35588 17892
rect 35308 17838 35310 17890
rect 35362 17838 35588 17890
rect 35308 17836 35588 17838
rect 34636 17714 34692 17724
rect 34972 17780 35028 17790
rect 34860 17668 34916 17678
rect 34860 17574 34916 17612
rect 34524 17556 34580 17566
rect 34524 17462 34580 17500
rect 34412 17276 34692 17332
rect 34188 17220 34244 17230
rect 34188 17106 34244 17164
rect 34188 17054 34190 17106
rect 34242 17054 34244 17106
rect 34188 17042 34244 17054
rect 34412 17108 34468 17118
rect 34412 17014 34468 17052
rect 33852 16716 34580 16772
rect 33964 16098 34020 16110
rect 33964 16046 33966 16098
rect 34018 16046 34020 16098
rect 33964 15876 34020 16046
rect 34300 15988 34356 15998
rect 34300 15894 34356 15932
rect 33852 15540 33908 15550
rect 33852 15446 33908 15484
rect 33964 15316 34020 15820
rect 33964 15250 34020 15260
rect 34188 15316 34244 15326
rect 34188 15148 34244 15260
rect 33404 15092 33460 15102
rect 33740 15092 33908 15148
rect 34188 15092 34356 15148
rect 33404 15090 33572 15092
rect 33404 15038 33406 15090
rect 33458 15038 33572 15090
rect 33404 15036 33572 15038
rect 33404 15026 33460 15036
rect 33404 14644 33460 14654
rect 33404 13858 33460 14588
rect 33516 14642 33572 15036
rect 33516 14590 33518 14642
rect 33570 14590 33572 14642
rect 33516 14578 33572 14590
rect 33404 13806 33406 13858
rect 33458 13806 33460 13858
rect 33404 13794 33460 13806
rect 33628 13970 33684 13982
rect 33628 13918 33630 13970
rect 33682 13918 33684 13970
rect 33628 13748 33684 13918
rect 33740 13860 33796 13870
rect 33740 13766 33796 13804
rect 33628 13682 33684 13692
rect 33740 13636 33796 13646
rect 33628 12180 33684 12190
rect 33292 11564 33572 11620
rect 33180 11452 33460 11508
rect 33068 11396 33124 11406
rect 33068 11302 33124 11340
rect 33180 10722 33236 11452
rect 33404 11394 33460 11452
rect 33404 11342 33406 11394
rect 33458 11342 33460 11394
rect 33404 11330 33460 11342
rect 33516 10948 33572 11564
rect 33628 11172 33684 12124
rect 33740 11396 33796 13580
rect 33852 12404 33908 15092
rect 34188 14980 34244 14990
rect 34076 14756 34132 14766
rect 33964 13746 34020 13758
rect 33964 13694 33966 13746
rect 34018 13694 34020 13746
rect 33964 12964 34020 13694
rect 34076 13636 34132 14700
rect 34076 13570 34132 13580
rect 34188 13524 34244 14924
rect 34188 13458 34244 13468
rect 34300 14530 34356 15092
rect 34524 14980 34580 16716
rect 34636 16100 34692 17276
rect 34636 15986 34692 16044
rect 34636 15934 34638 15986
rect 34690 15934 34692 15986
rect 34636 15148 34692 15934
rect 34860 16884 34916 16894
rect 34860 15316 34916 16828
rect 34972 16882 35028 17724
rect 34972 16830 34974 16882
rect 35026 16830 35028 16882
rect 34972 16818 35028 16830
rect 35308 16660 35364 17836
rect 35420 17556 35476 17566
rect 35756 17556 35812 17566
rect 35420 17554 35812 17556
rect 35420 17502 35422 17554
rect 35474 17502 35758 17554
rect 35810 17502 35812 17554
rect 35420 17500 35812 17502
rect 35420 17490 35476 17500
rect 35756 17490 35812 17500
rect 35868 17332 35924 18396
rect 36092 18386 36148 18396
rect 36204 17778 36260 18844
rect 36204 17726 36206 17778
rect 36258 17726 36260 17778
rect 36204 17714 36260 17726
rect 36316 18004 36372 18014
rect 36092 17668 36148 17678
rect 36092 17574 36148 17612
rect 36316 17666 36372 17948
rect 36316 17614 36318 17666
rect 36370 17614 36372 17666
rect 36316 17602 36372 17614
rect 36428 17892 36484 17902
rect 36428 17332 36484 17836
rect 35756 17276 35924 17332
rect 36092 17276 36484 17332
rect 35420 17108 35476 17118
rect 35420 17014 35476 17052
rect 35084 16604 35364 16660
rect 35084 15988 35140 16604
rect 35196 16492 35460 16502
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35196 16426 35460 16436
rect 35196 16268 35364 16324
rect 35196 16210 35252 16268
rect 35196 16158 35198 16210
rect 35250 16158 35252 16210
rect 35196 16146 35252 16158
rect 35308 16212 35364 16268
rect 35420 16212 35476 16222
rect 35308 16156 35420 16212
rect 35420 16146 35476 16156
rect 35532 16100 35588 16110
rect 35756 16100 35812 17276
rect 36092 16994 36148 17276
rect 36316 17108 36372 17118
rect 36092 16942 36094 16994
rect 36146 16942 36148 16994
rect 36092 16930 36148 16942
rect 36204 17052 36316 17108
rect 35980 16884 36036 16894
rect 35532 16098 35812 16100
rect 35532 16046 35534 16098
rect 35586 16046 35812 16098
rect 35532 16044 35812 16046
rect 35868 16324 35924 16334
rect 35868 16098 35924 16268
rect 35868 16046 35870 16098
rect 35922 16046 35924 16098
rect 35532 16034 35588 16044
rect 35868 16034 35924 16046
rect 35980 16100 36036 16828
rect 36092 16324 36148 16334
rect 36204 16324 36260 17052
rect 36316 17014 36372 17052
rect 36428 16996 36484 17006
rect 36428 16902 36484 16940
rect 36092 16322 36260 16324
rect 36092 16270 36094 16322
rect 36146 16270 36260 16322
rect 36092 16268 36260 16270
rect 36428 16660 36484 16670
rect 36540 16660 36596 26852
rect 36652 26178 36708 28700
rect 36652 26126 36654 26178
rect 36706 26126 36708 26178
rect 36652 25284 36708 26126
rect 36764 25732 36820 29374
rect 36988 29428 37044 31166
rect 37100 30882 37156 34076
rect 37212 34066 37268 34076
rect 37324 33906 37380 33918
rect 37324 33854 37326 33906
rect 37378 33854 37380 33906
rect 37324 32676 37380 33854
rect 37436 33572 37492 34076
rect 37436 33506 37492 33516
rect 37548 33236 37604 33246
rect 37548 32786 37604 33180
rect 37548 32734 37550 32786
rect 37602 32734 37604 32786
rect 37548 32722 37604 32734
rect 37436 32676 37492 32686
rect 37324 32674 37492 32676
rect 37324 32622 37438 32674
rect 37490 32622 37492 32674
rect 37324 32620 37492 32622
rect 37436 32610 37492 32620
rect 37660 32004 37716 34412
rect 37772 32564 37828 32574
rect 37772 32562 38276 32564
rect 37772 32510 37774 32562
rect 37826 32510 38276 32562
rect 37772 32508 38276 32510
rect 37772 32498 37828 32508
rect 37660 31948 38052 32004
rect 37548 31668 37604 31678
rect 37772 31668 37828 31678
rect 37604 31666 37828 31668
rect 37604 31614 37774 31666
rect 37826 31614 37828 31666
rect 37604 31612 37828 31614
rect 37548 31602 37604 31612
rect 37772 31602 37828 31612
rect 37436 31554 37492 31566
rect 37436 31502 37438 31554
rect 37490 31502 37492 31554
rect 37436 31444 37492 31502
rect 37492 31388 37716 31444
rect 37436 31378 37492 31388
rect 37212 31220 37268 31230
rect 37212 31126 37268 31164
rect 37100 30830 37102 30882
rect 37154 30830 37156 30882
rect 37100 30324 37156 30830
rect 37100 30258 37156 30268
rect 37436 30994 37492 31006
rect 37436 30942 37438 30994
rect 37490 30942 37492 30994
rect 37100 29428 37156 29438
rect 36988 29426 37156 29428
rect 36988 29374 37102 29426
rect 37154 29374 37156 29426
rect 36988 29372 37156 29374
rect 37100 29362 37156 29372
rect 37436 28868 37492 30942
rect 37660 30994 37716 31388
rect 37660 30942 37662 30994
rect 37714 30942 37716 30994
rect 37660 30930 37716 30942
rect 37548 30436 37604 30446
rect 37548 30322 37604 30380
rect 37548 30270 37550 30322
rect 37602 30270 37604 30322
rect 37548 30258 37604 30270
rect 37548 28868 37604 28878
rect 37436 28866 37940 28868
rect 37436 28814 37550 28866
rect 37602 28814 37940 28866
rect 37436 28812 37940 28814
rect 37548 28802 37604 28812
rect 36988 28642 37044 28654
rect 36988 28590 36990 28642
rect 37042 28590 37044 28642
rect 36988 27748 37044 28590
rect 36876 27692 37044 27748
rect 37212 28642 37268 28654
rect 37212 28590 37214 28642
rect 37266 28590 37268 28642
rect 36876 26964 36932 27692
rect 37212 27412 37268 28590
rect 37884 28642 37940 28812
rect 37884 28590 37886 28642
rect 37938 28590 37940 28642
rect 37884 28578 37940 28590
rect 37996 27748 38052 31948
rect 38220 31890 38276 32508
rect 38220 31838 38222 31890
rect 38274 31838 38276 31890
rect 38220 31826 38276 31838
rect 38108 31778 38164 31790
rect 38108 31726 38110 31778
rect 38162 31726 38164 31778
rect 38108 31220 38164 31726
rect 38108 31126 38164 31164
rect 38332 31666 38388 31678
rect 38332 31614 38334 31666
rect 38386 31614 38388 31666
rect 38332 31108 38388 31614
rect 38220 30996 38276 31006
rect 38220 30902 38276 30940
rect 38332 30994 38388 31052
rect 38332 30942 38334 30994
rect 38386 30942 38388 30994
rect 38108 30436 38164 30446
rect 38108 29426 38164 30380
rect 38108 29374 38110 29426
rect 38162 29374 38164 29426
rect 38108 29362 38164 29374
rect 38220 28420 38276 28430
rect 38332 28420 38388 30942
rect 37996 27682 38052 27692
rect 38108 28418 38388 28420
rect 38108 28366 38222 28418
rect 38274 28366 38388 28418
rect 38108 28364 38388 28366
rect 36988 27356 37268 27412
rect 36988 27076 37044 27356
rect 36988 26982 37044 27020
rect 37100 27076 37156 27086
rect 37884 27076 37940 27086
rect 37100 27074 37940 27076
rect 37100 27022 37102 27074
rect 37154 27022 37886 27074
rect 37938 27022 37940 27074
rect 37100 27020 37940 27022
rect 37100 27010 37156 27020
rect 37884 27010 37940 27020
rect 37996 26964 38052 26974
rect 36876 26898 36932 26908
rect 36988 26852 37044 26862
rect 37212 26852 37268 26862
rect 37436 26852 37492 26862
rect 37044 26796 37156 26852
rect 36988 26786 37044 26796
rect 36764 25666 36820 25676
rect 37100 26628 37156 26796
rect 37212 26758 37268 26796
rect 37324 26850 37492 26852
rect 37324 26798 37438 26850
rect 37490 26798 37492 26850
rect 37324 26796 37492 26798
rect 37324 26628 37380 26796
rect 37436 26786 37492 26796
rect 37548 26852 38052 26908
rect 38108 26962 38164 28364
rect 38220 28354 38276 28364
rect 38332 27746 38388 27758
rect 38332 27694 38334 27746
rect 38386 27694 38388 27746
rect 38220 27300 38276 27310
rect 38332 27300 38388 27694
rect 38220 27298 38388 27300
rect 38220 27246 38222 27298
rect 38274 27246 38388 27298
rect 38220 27244 38388 27246
rect 38220 27234 38276 27244
rect 38108 26910 38110 26962
rect 38162 26910 38164 26962
rect 38108 26898 38164 26910
rect 37100 26572 37380 26628
rect 37100 26514 37156 26572
rect 37100 26462 37102 26514
rect 37154 26462 37156 26514
rect 36988 25508 37044 25518
rect 36988 25414 37044 25452
rect 36652 25228 37044 25284
rect 36988 23716 37044 25228
rect 37100 25060 37156 26462
rect 37436 26516 37492 26526
rect 37436 25730 37492 26460
rect 37548 26178 37604 26852
rect 38220 26628 38276 26638
rect 37996 26516 38052 26526
rect 37996 26422 38052 26460
rect 37548 26126 37550 26178
rect 37602 26126 37604 26178
rect 37548 26066 37604 26126
rect 37548 26014 37550 26066
rect 37602 26014 37604 26066
rect 37548 26002 37604 26014
rect 37436 25678 37438 25730
rect 37490 25678 37492 25730
rect 37212 25506 37268 25518
rect 37212 25454 37214 25506
rect 37266 25454 37268 25506
rect 37212 25284 37268 25454
rect 37212 25218 37268 25228
rect 37100 25004 37268 25060
rect 37100 23716 37156 23726
rect 36988 23714 37156 23716
rect 36988 23662 37102 23714
rect 37154 23662 37156 23714
rect 36988 23660 37156 23662
rect 36764 23042 36820 23054
rect 36764 22990 36766 23042
rect 36818 22990 36820 23042
rect 36652 20580 36708 20590
rect 36764 20580 36820 22990
rect 37100 22372 37156 23660
rect 37212 23268 37268 25004
rect 37436 23492 37492 25678
rect 38220 25618 38276 26572
rect 38220 25566 38222 25618
rect 38274 25566 38276 25618
rect 38220 25554 38276 25566
rect 37548 25394 37604 25406
rect 37548 25342 37550 25394
rect 37602 25342 37604 25394
rect 37548 24836 37604 25342
rect 38444 24836 38500 24846
rect 37548 24834 38500 24836
rect 37548 24782 38446 24834
rect 38498 24782 38500 24834
rect 37548 24780 38500 24782
rect 38444 24770 38500 24780
rect 38556 24052 38612 34860
rect 38780 34804 38836 34814
rect 38892 34804 38948 35646
rect 38836 34748 38948 34804
rect 39004 34804 39060 36764
rect 39116 34804 39172 34814
rect 39004 34802 39172 34804
rect 39004 34750 39118 34802
rect 39170 34750 39172 34802
rect 39004 34748 39172 34750
rect 38780 34710 38836 34748
rect 39116 33572 39172 34748
rect 39116 33506 39172 33516
rect 39116 33236 39172 33246
rect 39116 33142 39172 33180
rect 39228 32788 39284 36764
rect 39340 35586 39396 39564
rect 39676 38946 39732 38958
rect 39676 38894 39678 38946
rect 39730 38894 39732 38946
rect 39564 38610 39620 38622
rect 39564 38558 39566 38610
rect 39618 38558 39620 38610
rect 39452 38164 39508 38174
rect 39564 38164 39620 38558
rect 39452 38162 39620 38164
rect 39452 38110 39454 38162
rect 39506 38110 39620 38162
rect 39452 38108 39620 38110
rect 39452 38098 39508 38108
rect 39676 37828 39732 38894
rect 40348 38724 40404 38734
rect 40236 38722 40404 38724
rect 40236 38670 40350 38722
rect 40402 38670 40404 38722
rect 40236 38668 40404 38670
rect 39900 38610 39956 38622
rect 39900 38558 39902 38610
rect 39954 38558 39956 38610
rect 39900 38276 39956 38558
rect 39900 38210 39956 38220
rect 40124 38612 40292 38668
rect 40348 38658 40404 38668
rect 40460 38724 40516 43652
rect 40908 43650 40964 43652
rect 40908 43598 40910 43650
rect 40962 43598 40964 43650
rect 40908 43586 40964 43598
rect 41020 43650 41076 43708
rect 41468 43764 41524 43802
rect 41692 43764 41748 44046
rect 41524 43708 41748 43764
rect 42252 43708 42308 47068
rect 42476 47058 42532 47068
rect 42588 47348 42644 47358
rect 42476 45892 42532 45902
rect 42364 44996 42420 45006
rect 42364 44436 42420 44940
rect 42364 44322 42420 44380
rect 42364 44270 42366 44322
rect 42418 44270 42420 44322
rect 42364 44258 42420 44270
rect 41468 43698 41524 43708
rect 41020 43598 41022 43650
rect 41074 43598 41076 43650
rect 41020 43586 41076 43598
rect 42028 43652 42308 43708
rect 42028 43540 42084 43652
rect 40684 43316 40740 43326
rect 40684 42868 40740 43260
rect 40684 42866 41076 42868
rect 40684 42814 40686 42866
rect 40738 42814 41076 42866
rect 40684 42812 41076 42814
rect 40684 42802 40740 42812
rect 41020 42194 41076 42812
rect 42028 42866 42084 43484
rect 42028 42814 42030 42866
rect 42082 42814 42084 42866
rect 42028 42802 42084 42814
rect 41020 42142 41022 42194
rect 41074 42142 41076 42194
rect 41020 42130 41076 42142
rect 41244 42754 41300 42766
rect 41244 42702 41246 42754
rect 41298 42702 41300 42754
rect 40908 40404 40964 40414
rect 40908 40310 40964 40348
rect 41132 40404 41188 40414
rect 41244 40404 41300 42702
rect 41188 40348 41300 40404
rect 41356 42084 41412 42094
rect 41356 40404 41412 42028
rect 41468 41748 41524 41758
rect 41468 41298 41524 41692
rect 41468 41246 41470 41298
rect 41522 41246 41524 41298
rect 41468 41234 41524 41246
rect 42252 41186 42308 41198
rect 42252 41134 42254 41186
rect 42306 41134 42308 41186
rect 41916 40516 41972 40526
rect 41916 40422 41972 40460
rect 41468 40404 41524 40414
rect 41356 40402 41524 40404
rect 41356 40350 41470 40402
rect 41522 40350 41524 40402
rect 41356 40348 41524 40350
rect 41132 39730 41188 40348
rect 41132 39678 41134 39730
rect 41186 39678 41188 39730
rect 41132 38834 41188 39678
rect 41132 38782 41134 38834
rect 41186 38782 41188 38834
rect 41132 38770 41188 38782
rect 40460 38658 40516 38668
rect 40124 38164 40180 38612
rect 40124 38098 40180 38108
rect 39676 37762 39732 37772
rect 40236 37828 40292 37838
rect 39788 37380 39844 37390
rect 39788 37266 39844 37324
rect 39788 37214 39790 37266
rect 39842 37214 39844 37266
rect 39788 37202 39844 37214
rect 40236 37154 40292 37772
rect 40236 37102 40238 37154
rect 40290 37102 40292 37154
rect 40236 36596 40292 37102
rect 40012 36540 40292 36596
rect 40348 37380 40404 37390
rect 41468 37380 41524 40348
rect 42252 40404 42308 41134
rect 42252 40338 42308 40348
rect 42476 39956 42532 45836
rect 42588 45668 42644 47292
rect 42700 47346 42756 47358
rect 42700 47294 42702 47346
rect 42754 47294 42756 47346
rect 42700 47236 42756 47294
rect 42700 47170 42756 47180
rect 42812 46004 42868 47404
rect 43036 47346 43092 47404
rect 43036 47294 43038 47346
rect 43090 47294 43092 47346
rect 43036 47282 43092 47294
rect 42924 47234 42980 47246
rect 42924 47182 42926 47234
rect 42978 47182 42980 47234
rect 42924 46788 42980 47182
rect 43484 47234 43540 47246
rect 43484 47182 43486 47234
rect 43538 47182 43540 47234
rect 43484 47124 43540 47182
rect 43484 47058 43540 47068
rect 43596 47236 43652 47246
rect 43596 47012 43652 47180
rect 44268 47234 44324 47246
rect 44268 47182 44270 47234
rect 44322 47182 44324 47234
rect 43596 46956 43708 47012
rect 43652 46900 43708 46956
rect 44268 46900 44324 47182
rect 44716 46900 44772 48412
rect 44940 48402 44996 48412
rect 45276 48130 45332 48142
rect 45276 48078 45278 48130
rect 45330 48078 45332 48130
rect 45276 47684 45332 48078
rect 44940 47628 45332 47684
rect 44828 47460 44884 47470
rect 44940 47460 44996 47628
rect 44828 47458 44996 47460
rect 44828 47406 44830 47458
rect 44882 47406 44996 47458
rect 44828 47404 44996 47406
rect 44828 47348 44884 47404
rect 44828 47282 44884 47292
rect 43652 46844 43876 46900
rect 43820 46788 43876 46844
rect 44268 46898 44772 46900
rect 44268 46846 44718 46898
rect 44770 46846 44772 46898
rect 44268 46844 44772 46846
rect 42924 46732 43652 46788
rect 43820 46732 43988 46788
rect 43484 46564 43540 46574
rect 43148 46562 43540 46564
rect 43148 46510 43486 46562
rect 43538 46510 43540 46562
rect 43148 46508 43540 46510
rect 43148 46114 43204 46508
rect 43484 46498 43540 46508
rect 43148 46062 43150 46114
rect 43202 46062 43204 46114
rect 43148 46050 43204 46062
rect 43484 46116 43540 46126
rect 43596 46116 43652 46732
rect 43484 46114 43652 46116
rect 43484 46062 43486 46114
rect 43538 46062 43652 46114
rect 43484 46060 43652 46062
rect 43708 46676 43764 46686
rect 43484 46050 43540 46060
rect 42812 45938 42868 45948
rect 43260 45892 43316 45902
rect 43260 45798 43316 45836
rect 43596 45892 43652 45902
rect 43596 45798 43652 45836
rect 42588 45612 43540 45668
rect 43372 45220 43428 45230
rect 42812 45108 42868 45118
rect 42812 45014 42868 45052
rect 43036 45108 43092 45118
rect 43036 45106 43204 45108
rect 43036 45054 43038 45106
rect 43090 45054 43204 45106
rect 43036 45052 43204 45054
rect 43036 45042 43092 45052
rect 42700 44884 42756 44894
rect 42588 44828 42700 44884
rect 42588 44210 42644 44828
rect 42700 44790 42756 44828
rect 42924 44548 42980 44558
rect 42924 44454 42980 44492
rect 43036 44436 43092 44446
rect 43148 44436 43204 45052
rect 43372 44436 43428 45164
rect 43484 44882 43540 45612
rect 43596 44996 43652 45006
rect 43596 44902 43652 44940
rect 43484 44830 43486 44882
rect 43538 44830 43540 44882
rect 43484 44818 43540 44830
rect 43708 44436 43764 46620
rect 43932 45106 43988 46732
rect 44268 46676 44324 46844
rect 44716 46834 44772 46844
rect 44268 46582 44324 46620
rect 43932 45054 43934 45106
rect 43986 45054 43988 45106
rect 43932 44548 43988 45054
rect 43932 44482 43988 44492
rect 44044 46004 44100 46014
rect 43036 44434 43428 44436
rect 43036 44382 43038 44434
rect 43090 44382 43428 44434
rect 43036 44380 43428 44382
rect 43036 44370 43092 44380
rect 42588 44158 42590 44210
rect 42642 44158 42644 44210
rect 42588 44146 42644 44158
rect 43372 43876 43428 44380
rect 43372 43810 43428 43820
rect 43596 44380 43764 44436
rect 43260 43652 43316 43662
rect 43596 43652 43652 44380
rect 44044 44324 44100 45948
rect 44828 46004 44884 46014
rect 44828 45910 44884 45948
rect 44940 45780 44996 47404
rect 45052 47460 45108 47470
rect 45108 47404 45332 47460
rect 45052 47366 45108 47404
rect 45276 46562 45332 47404
rect 45388 47236 45444 47246
rect 45388 47142 45444 47180
rect 45276 46510 45278 46562
rect 45330 46510 45332 46562
rect 45276 45890 45332 46510
rect 45276 45838 45278 45890
rect 45330 45838 45332 45890
rect 45276 45826 45332 45838
rect 45164 45780 45220 45790
rect 44940 45778 45220 45780
rect 44940 45726 45166 45778
rect 45218 45726 45220 45778
rect 44940 45724 45220 45726
rect 45164 45714 45220 45724
rect 44156 45668 44212 45678
rect 44156 45574 44212 45612
rect 45052 45556 45108 45566
rect 44828 45332 44884 45342
rect 44604 45330 44884 45332
rect 44604 45278 44830 45330
rect 44882 45278 44884 45330
rect 44604 45276 44884 45278
rect 44492 45108 44548 45118
rect 44156 45106 44548 45108
rect 44156 45054 44494 45106
rect 44546 45054 44548 45106
rect 44156 45052 44548 45054
rect 44156 44434 44212 45052
rect 44492 45042 44548 45052
rect 44156 44382 44158 44434
rect 44210 44382 44212 44434
rect 44156 44370 44212 44382
rect 43932 44268 44044 44324
rect 43260 43650 43652 43652
rect 43260 43598 43262 43650
rect 43314 43598 43652 43650
rect 43260 43596 43652 43598
rect 43260 43586 43316 43596
rect 43596 43540 43652 43596
rect 43596 43446 43652 43484
rect 43820 44212 43876 44222
rect 43484 41748 43540 41758
rect 42812 41412 42868 41422
rect 42812 41300 42868 41356
rect 43484 41410 43540 41692
rect 43484 41358 43486 41410
rect 43538 41358 43540 41410
rect 43484 41346 43540 41358
rect 42812 41298 43204 41300
rect 42812 41246 42814 41298
rect 42866 41246 43204 41298
rect 42812 41244 43204 41246
rect 42812 41234 42868 41244
rect 43148 41186 43204 41244
rect 43148 41134 43150 41186
rect 43202 41134 43204 41186
rect 43148 41122 43204 41134
rect 43372 40962 43428 40974
rect 43372 40910 43374 40962
rect 43426 40910 43428 40962
rect 43372 40514 43428 40910
rect 43372 40462 43374 40514
rect 43426 40462 43428 40514
rect 43372 40450 43428 40462
rect 43820 40516 43876 44156
rect 43932 44210 43988 44268
rect 44044 44258 44100 44268
rect 44268 44324 44324 44334
rect 44268 44230 44324 44268
rect 43932 44158 43934 44210
rect 43986 44158 43988 44210
rect 43932 44146 43988 44158
rect 44044 44100 44100 44138
rect 44044 44034 44100 44044
rect 44044 43876 44100 43886
rect 44044 42868 44100 43820
rect 44604 43708 44660 45276
rect 44828 45266 44884 45276
rect 44940 45332 44996 45342
rect 44828 45108 44884 45118
rect 44940 45108 44996 45276
rect 44828 45106 44996 45108
rect 44828 45054 44830 45106
rect 44882 45054 44996 45106
rect 44828 45052 44996 45054
rect 44828 45042 44884 45052
rect 44940 44212 44996 44222
rect 44940 44118 44996 44156
rect 44380 43652 44660 43708
rect 45052 43708 45108 45500
rect 45388 45332 45444 45342
rect 45388 45238 45444 45276
rect 45612 45220 45668 45230
rect 45164 45108 45220 45118
rect 45164 44324 45220 45052
rect 45612 45106 45668 45164
rect 45612 45054 45614 45106
rect 45666 45054 45668 45106
rect 45612 45042 45668 45054
rect 45276 44436 45332 44446
rect 45276 44342 45332 44380
rect 45164 44258 45220 44268
rect 45052 43652 45220 43708
rect 44380 43650 44436 43652
rect 44380 43598 44382 43650
rect 44434 43598 44436 43650
rect 44380 43586 44436 43598
rect 45052 43540 45108 43550
rect 44156 42868 44212 42878
rect 44044 42866 44212 42868
rect 44044 42814 44158 42866
rect 44210 42814 44212 42866
rect 44044 42812 44212 42814
rect 44156 42802 44212 42812
rect 45052 42866 45108 43484
rect 45052 42814 45054 42866
rect 45106 42814 45108 42866
rect 45052 42802 45108 42814
rect 43820 40450 43876 40460
rect 42700 40404 42756 40414
rect 42756 40348 42868 40404
rect 42700 40310 42756 40348
rect 42476 39890 42532 39900
rect 42476 39732 42532 39742
rect 42028 39730 42532 39732
rect 42028 39678 42478 39730
rect 42530 39678 42532 39730
rect 42028 39676 42532 39678
rect 42028 39618 42084 39676
rect 42476 39666 42532 39676
rect 42028 39566 42030 39618
rect 42082 39566 42084 39618
rect 42028 39554 42084 39566
rect 41692 39506 41748 39518
rect 41692 39454 41694 39506
rect 41746 39454 41748 39506
rect 41580 38162 41636 38174
rect 41580 38110 41582 38162
rect 41634 38110 41636 38162
rect 41580 38052 41636 38110
rect 41580 37986 41636 37996
rect 39676 36372 39732 36382
rect 39676 36370 39844 36372
rect 39676 36318 39678 36370
rect 39730 36318 39844 36370
rect 39676 36316 39844 36318
rect 39676 36306 39732 36316
rect 39340 35534 39342 35586
rect 39394 35534 39396 35586
rect 39340 35522 39396 35534
rect 39788 35586 39844 36316
rect 39788 35534 39790 35586
rect 39842 35534 39844 35586
rect 39788 35522 39844 35534
rect 39900 35812 39956 35822
rect 40012 35812 40068 36540
rect 40348 36484 40404 37324
rect 41356 37378 41524 37380
rect 41356 37326 41470 37378
rect 41522 37326 41524 37378
rect 41356 37324 41524 37326
rect 40236 36428 40404 36484
rect 40460 37044 40516 37054
rect 39900 35810 40068 35812
rect 39900 35758 39902 35810
rect 39954 35758 40068 35810
rect 39900 35756 40068 35758
rect 40124 36372 40180 36382
rect 40124 35810 40180 36316
rect 40124 35758 40126 35810
rect 40178 35758 40180 35810
rect 38892 32732 39284 32788
rect 39564 34692 39620 34702
rect 39900 34692 39956 35756
rect 40124 35746 40180 35758
rect 39564 34690 39956 34692
rect 39564 34638 39566 34690
rect 39618 34638 39956 34690
rect 39564 34636 39956 34638
rect 38668 31668 38724 31678
rect 38668 31666 38836 31668
rect 38668 31614 38670 31666
rect 38722 31614 38836 31666
rect 38668 31612 38836 31614
rect 38668 31602 38724 31612
rect 38668 30996 38724 31006
rect 38668 30902 38724 30940
rect 38780 30436 38836 31612
rect 38780 30370 38836 30380
rect 38892 26516 38948 32732
rect 39564 31780 39620 34636
rect 39900 33348 39956 33358
rect 39900 33254 39956 33292
rect 40012 33236 40068 33246
rect 40012 32786 40068 33180
rect 40012 32734 40014 32786
rect 40066 32734 40068 32786
rect 40012 32722 40068 32734
rect 40236 32676 40292 36428
rect 40348 33348 40404 33358
rect 40348 33254 40404 33292
rect 40124 32620 40292 32676
rect 39676 32564 39732 32574
rect 40124 32564 40180 32620
rect 39676 32562 40180 32564
rect 39676 32510 39678 32562
rect 39730 32510 40180 32562
rect 39676 32508 40180 32510
rect 40236 32562 40292 32620
rect 40236 32510 40238 32562
rect 40290 32510 40292 32562
rect 39676 32498 39732 32508
rect 40236 32498 40292 32510
rect 39900 32338 39956 32350
rect 39900 32286 39902 32338
rect 39954 32286 39956 32338
rect 39900 31892 39956 32286
rect 39564 31714 39620 31724
rect 39676 31836 39900 31892
rect 39004 31554 39060 31566
rect 39004 31502 39006 31554
rect 39058 31502 39060 31554
rect 39004 31220 39060 31502
rect 39004 30994 39060 31164
rect 39676 31218 39732 31836
rect 39900 31826 39956 31836
rect 40012 32340 40068 32350
rect 39676 31166 39678 31218
rect 39730 31166 39732 31218
rect 39676 31154 39732 31166
rect 39228 31108 39284 31118
rect 39228 31014 39284 31052
rect 39004 30942 39006 30994
rect 39058 30942 39060 30994
rect 39004 30930 39060 30942
rect 39116 30882 39172 30894
rect 39116 30830 39118 30882
rect 39170 30830 39172 30882
rect 39116 30548 39172 30830
rect 39564 30884 39620 30894
rect 39564 30790 39620 30828
rect 39116 30492 39732 30548
rect 39676 30322 39732 30492
rect 39676 30270 39678 30322
rect 39730 30270 39732 30322
rect 39676 30258 39732 30270
rect 39228 29428 39284 29438
rect 39004 28642 39060 28654
rect 39004 28590 39006 28642
rect 39058 28590 39060 28642
rect 39004 26908 39060 28590
rect 39228 28642 39284 29372
rect 39228 28590 39230 28642
rect 39282 28590 39284 28642
rect 39228 28578 39284 28590
rect 39900 28532 39956 28542
rect 39900 28438 39956 28476
rect 39116 27858 39172 27870
rect 39116 27806 39118 27858
rect 39170 27806 39172 27858
rect 39116 27748 39172 27806
rect 39564 27748 39620 27758
rect 39116 27692 39564 27748
rect 39564 27074 39620 27692
rect 39564 27022 39566 27074
rect 39618 27022 39620 27074
rect 39564 27010 39620 27022
rect 39004 26852 39172 26908
rect 38892 26450 38948 26460
rect 39116 26514 39172 26852
rect 39116 26462 39118 26514
rect 39170 26462 39172 26514
rect 39116 26450 39172 26462
rect 39340 26404 39396 26414
rect 39340 26310 39396 26348
rect 39452 26290 39508 26302
rect 39452 26238 39454 26290
rect 39506 26238 39508 26290
rect 39452 25508 39508 26238
rect 39452 25442 39508 25452
rect 39228 24722 39284 24734
rect 39228 24670 39230 24722
rect 39282 24670 39284 24722
rect 39228 24612 39284 24670
rect 39228 24546 39284 24556
rect 39676 24612 39732 24622
rect 39676 24518 39732 24556
rect 37996 23996 38612 24052
rect 37436 23426 37492 23436
rect 37884 23938 37940 23950
rect 37884 23886 37886 23938
rect 37938 23886 37940 23938
rect 37212 23212 37716 23268
rect 37548 22372 37604 22382
rect 37100 22370 37604 22372
rect 37100 22318 37550 22370
rect 37602 22318 37604 22370
rect 37100 22316 37604 22318
rect 37100 22148 37156 22158
rect 37100 22054 37156 22092
rect 37548 21812 37604 22316
rect 37660 22260 37716 23212
rect 37660 22204 37828 22260
rect 36988 20692 37044 20702
rect 36988 20598 37044 20636
rect 37100 20690 37156 20702
rect 37100 20638 37102 20690
rect 37154 20638 37156 20690
rect 36708 20524 36820 20580
rect 36652 20514 36708 20524
rect 36988 20468 37044 20478
rect 36988 19684 37044 20412
rect 37100 20132 37156 20638
rect 37100 20066 37156 20076
rect 37100 19908 37156 19918
rect 37548 19908 37604 21756
rect 37660 21028 37716 21038
rect 37660 20914 37716 20972
rect 37660 20862 37662 20914
rect 37714 20862 37716 20914
rect 37660 20850 37716 20862
rect 37772 20692 37828 22204
rect 37884 21812 37940 23886
rect 37884 21746 37940 21756
rect 37156 19852 37604 19908
rect 37100 19814 37156 19852
rect 36988 19628 37380 19684
rect 36876 19234 36932 19246
rect 36876 19182 36878 19234
rect 36930 19182 36932 19234
rect 36876 18900 36932 19182
rect 37212 19236 37268 19246
rect 37212 19142 37268 19180
rect 36876 18834 36932 18844
rect 37100 19010 37156 19022
rect 37100 18958 37102 19010
rect 37154 18958 37156 19010
rect 36876 18452 36932 18462
rect 37100 18452 37156 18958
rect 36876 18450 37156 18452
rect 36876 18398 36878 18450
rect 36930 18398 37156 18450
rect 36876 18396 37156 18398
rect 37212 18452 37268 18462
rect 36876 18386 36932 18396
rect 36876 18004 36932 18014
rect 36652 17220 36708 17230
rect 36708 17164 36820 17220
rect 36652 17154 36708 17164
rect 36652 16884 36708 16894
rect 36652 16790 36708 16828
rect 36540 16604 36708 16660
rect 36428 16322 36484 16604
rect 36428 16270 36430 16322
rect 36482 16270 36484 16322
rect 36092 16258 36148 16268
rect 36428 16258 36484 16270
rect 36316 16212 36372 16222
rect 35980 16044 36148 16100
rect 35084 15932 35476 15988
rect 35084 15316 35140 15326
rect 34860 15260 35084 15316
rect 34636 15092 35028 15148
rect 34524 14924 34804 14980
rect 34300 14478 34302 14530
rect 34354 14478 34356 14530
rect 34188 13076 34244 13086
rect 34188 12982 34244 13020
rect 33964 12898 34020 12908
rect 33852 12178 33908 12348
rect 34076 12852 34132 12862
rect 34076 12292 34132 12796
rect 34300 12740 34356 14478
rect 34524 14530 34580 14542
rect 34524 14478 34526 14530
rect 34578 14478 34580 14530
rect 34412 13748 34468 13758
rect 34524 13748 34580 14478
rect 34748 14196 34804 14924
rect 34972 14420 35028 15092
rect 35084 14756 35140 15260
rect 35420 15092 35476 15932
rect 35644 15874 35700 15886
rect 35644 15822 35646 15874
rect 35698 15822 35700 15874
rect 35644 15764 35700 15822
rect 35644 15698 35700 15708
rect 35980 15764 36036 15774
rect 35868 15652 35924 15662
rect 35756 15596 35868 15652
rect 35756 15148 35812 15596
rect 35868 15586 35924 15596
rect 35420 15026 35476 15036
rect 35644 15092 35812 15148
rect 35868 15204 35924 15242
rect 35868 15138 35924 15148
rect 35196 14924 35460 14934
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35196 14858 35460 14868
rect 35084 14700 35588 14756
rect 35532 14642 35588 14700
rect 35532 14590 35534 14642
rect 35586 14590 35588 14642
rect 35532 14578 35588 14590
rect 35084 14420 35140 14430
rect 34972 14418 35140 14420
rect 34972 14366 35086 14418
rect 35138 14366 35140 14418
rect 34972 14364 35140 14366
rect 35084 14354 35140 14364
rect 34748 14130 34804 14140
rect 34860 14306 34916 14318
rect 34860 14254 34862 14306
rect 34914 14254 34916 14306
rect 34860 13748 34916 14254
rect 35196 14306 35252 14318
rect 35196 14254 35198 14306
rect 35250 14254 35252 14306
rect 35196 13972 35252 14254
rect 35196 13906 35252 13916
rect 35420 13970 35476 13982
rect 35420 13918 35422 13970
rect 35474 13918 35476 13970
rect 34468 13692 34580 13748
rect 34636 13692 34916 13748
rect 35084 13746 35140 13758
rect 35084 13694 35086 13746
rect 35138 13694 35140 13746
rect 34412 13654 34468 13692
rect 34524 13524 34580 13534
rect 34636 13524 34692 13692
rect 34524 13522 34692 13524
rect 34524 13470 34526 13522
rect 34578 13470 34692 13522
rect 34524 13468 34692 13470
rect 34748 13524 34804 13534
rect 34412 12964 34468 12974
rect 34412 12870 34468 12908
rect 34300 12674 34356 12684
rect 34524 12516 34580 13468
rect 34748 13430 34804 13468
rect 34860 13522 34916 13534
rect 34860 13470 34862 13522
rect 34914 13470 34916 13522
rect 34636 12964 34692 12974
rect 34860 12964 34916 13470
rect 35084 13076 35140 13694
rect 35420 13524 35476 13918
rect 35532 13972 35588 13982
rect 35532 13858 35588 13916
rect 35532 13806 35534 13858
rect 35586 13806 35588 13858
rect 35532 13794 35588 13806
rect 35420 13468 35588 13524
rect 35196 13356 35460 13366
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35196 13290 35460 13300
rect 35084 13010 35140 13020
rect 34636 12962 34916 12964
rect 34636 12910 34638 12962
rect 34690 12910 34916 12962
rect 34636 12908 34916 12910
rect 34636 12898 34692 12908
rect 35084 12852 35140 12862
rect 35532 12852 35588 13468
rect 35084 12758 35140 12796
rect 35308 12796 35588 12852
rect 35644 12852 35700 15092
rect 35756 13860 35812 13870
rect 35756 13766 35812 13804
rect 33852 12126 33854 12178
rect 33906 12126 33908 12178
rect 33852 12114 33908 12126
rect 33964 12236 34132 12292
rect 34188 12460 34580 12516
rect 34636 12740 34692 12750
rect 33740 11340 33908 11396
rect 33740 11172 33796 11182
rect 33628 11170 33796 11172
rect 33628 11118 33742 11170
rect 33794 11118 33796 11170
rect 33628 11116 33796 11118
rect 33180 10670 33182 10722
rect 33234 10670 33236 10722
rect 33180 10658 33236 10670
rect 33292 10892 33572 10948
rect 33180 10052 33236 10062
rect 33180 9042 33236 9996
rect 33180 8990 33182 9042
rect 33234 8990 33236 9042
rect 33180 8978 33236 8990
rect 32732 8194 32788 8204
rect 33180 7588 33236 7598
rect 33180 7494 33236 7532
rect 31948 7422 31950 7474
rect 32002 7422 32004 7474
rect 31948 7410 32004 7422
rect 32172 7474 32228 7486
rect 32172 7422 32174 7474
rect 32226 7422 32228 7474
rect 31836 7362 31892 7374
rect 31836 7310 31838 7362
rect 31890 7310 31892 7362
rect 31388 6916 31444 6926
rect 31836 6916 31892 7310
rect 32172 7252 32228 7422
rect 32172 7186 32228 7196
rect 33068 7474 33124 7486
rect 33068 7422 33070 7474
rect 33122 7422 33124 7474
rect 31388 6914 31892 6916
rect 31388 6862 31390 6914
rect 31442 6862 31892 6914
rect 31388 6860 31892 6862
rect 31388 6850 31444 6860
rect 31276 6692 31332 6748
rect 31612 6692 31668 6702
rect 31276 6690 31668 6692
rect 31276 6638 31614 6690
rect 31666 6638 31668 6690
rect 31276 6636 31668 6638
rect 31836 6692 31892 6860
rect 32172 6804 32228 6814
rect 31948 6692 32004 6702
rect 31836 6690 32004 6692
rect 31836 6638 31950 6690
rect 32002 6638 32004 6690
rect 31836 6636 32004 6638
rect 31612 6626 31668 6636
rect 31948 6626 32004 6636
rect 32172 6690 32228 6748
rect 33068 6804 33124 7422
rect 33068 6738 33124 6748
rect 32172 6638 32174 6690
rect 32226 6638 32228 6690
rect 32172 6626 32228 6638
rect 33180 6692 33236 6702
rect 33292 6692 33348 10892
rect 33516 10722 33572 10734
rect 33516 10670 33518 10722
rect 33570 10670 33572 10722
rect 33516 9380 33572 10670
rect 33740 9492 33796 11116
rect 33852 10052 33908 11340
rect 33852 9986 33908 9996
rect 33964 9604 34020 12236
rect 34076 12068 34132 12078
rect 34076 11974 34132 12012
rect 34188 11954 34244 12460
rect 34636 12292 34692 12684
rect 34524 12236 34692 12292
rect 35308 12290 35364 12796
rect 35644 12786 35700 12796
rect 35308 12238 35310 12290
rect 35362 12238 35364 12290
rect 34524 12180 34580 12236
rect 35308 12226 35364 12238
rect 34188 11902 34190 11954
rect 34242 11902 34244 11954
rect 34188 11618 34244 11902
rect 34188 11566 34190 11618
rect 34242 11566 34244 11618
rect 34188 11554 34244 11566
rect 34412 12178 34580 12180
rect 34412 12126 34526 12178
rect 34578 12126 34580 12178
rect 34412 12124 34580 12126
rect 34300 11506 34356 11518
rect 34300 11454 34302 11506
rect 34354 11454 34356 11506
rect 34300 11396 34356 11454
rect 34300 11330 34356 11340
rect 34412 10610 34468 12124
rect 34524 12114 34580 12124
rect 34636 12068 34692 12078
rect 34692 12012 34916 12068
rect 34636 12002 34692 12012
rect 34636 11394 34692 11406
rect 34636 11342 34638 11394
rect 34690 11342 34692 11394
rect 34636 11060 34692 11342
rect 34636 10994 34692 11004
rect 34748 11284 34804 11294
rect 34412 10558 34414 10610
rect 34466 10558 34468 10610
rect 33964 9548 34244 9604
rect 33740 9436 34020 9492
rect 33516 9314 33572 9324
rect 33404 9044 33460 9054
rect 33404 8950 33460 8988
rect 33740 9042 33796 9054
rect 33740 8990 33742 9042
rect 33794 8990 33796 9042
rect 33516 8930 33572 8942
rect 33516 8878 33518 8930
rect 33570 8878 33572 8930
rect 33516 8372 33572 8878
rect 33628 8372 33684 8382
rect 33516 8370 33684 8372
rect 33516 8318 33630 8370
rect 33682 8318 33684 8370
rect 33516 8316 33684 8318
rect 33628 8306 33684 8316
rect 33740 8148 33796 8990
rect 33852 9044 33908 9054
rect 33852 8950 33908 8988
rect 33404 8092 33796 8148
rect 33404 7698 33460 8092
rect 33404 7646 33406 7698
rect 33458 7646 33460 7698
rect 33404 7634 33460 7646
rect 33740 7588 33796 7598
rect 33740 7494 33796 7532
rect 33964 6692 34020 9436
rect 34188 9268 34244 9548
rect 34076 9156 34132 9166
rect 34076 9062 34132 9100
rect 34188 9154 34244 9212
rect 34188 9102 34190 9154
rect 34242 9102 34244 9154
rect 34188 9090 34244 9102
rect 34412 8258 34468 10558
rect 34636 10388 34692 10398
rect 34524 10052 34580 10062
rect 34524 9156 34580 9996
rect 34636 9826 34692 10332
rect 34636 9774 34638 9826
rect 34690 9774 34692 9826
rect 34636 9762 34692 9774
rect 34748 9268 34804 11228
rect 34860 9826 34916 12012
rect 35196 11788 35460 11798
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35196 11722 35460 11732
rect 34972 11394 35028 11406
rect 34972 11342 34974 11394
rect 35026 11342 35028 11394
rect 34972 11284 35028 11342
rect 35644 11396 35700 11406
rect 35644 11302 35700 11340
rect 34972 11218 35028 11228
rect 35532 11172 35588 11182
rect 35196 10498 35252 10510
rect 35196 10446 35198 10498
rect 35250 10446 35252 10498
rect 35196 10388 35252 10446
rect 34860 9774 34862 9826
rect 34914 9774 34916 9826
rect 34860 9762 34916 9774
rect 34972 10332 35252 10388
rect 34972 9602 35028 10332
rect 35196 10220 35460 10230
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35196 10154 35460 10164
rect 35420 10052 35476 10062
rect 35308 9996 35420 10052
rect 35308 9938 35364 9996
rect 35420 9986 35476 9996
rect 35308 9886 35310 9938
rect 35362 9886 35364 9938
rect 35308 9874 35364 9886
rect 35084 9828 35140 9838
rect 35084 9734 35140 9772
rect 35532 9826 35588 11116
rect 35756 11170 35812 11182
rect 35756 11118 35758 11170
rect 35810 11118 35812 11170
rect 35756 10388 35812 11118
rect 35868 11170 35924 11182
rect 35868 11118 35870 11170
rect 35922 11118 35924 11170
rect 35868 11060 35924 11118
rect 35868 10500 35924 11004
rect 35868 10434 35924 10444
rect 35756 10322 35812 10332
rect 35532 9774 35534 9826
rect 35586 9774 35588 9826
rect 35532 9762 35588 9774
rect 35980 9604 36036 15708
rect 36092 11508 36148 16044
rect 36316 15986 36372 16156
rect 36540 16100 36596 16110
rect 36316 15934 36318 15986
rect 36370 15934 36372 15986
rect 36316 15922 36372 15934
rect 36428 16044 36540 16100
rect 36204 15092 36260 15102
rect 36204 14756 36260 15036
rect 36204 13970 36260 14700
rect 36428 14642 36484 16044
rect 36540 16034 36596 16044
rect 36428 14590 36430 14642
rect 36482 14590 36484 14642
rect 36428 14578 36484 14590
rect 36204 13918 36206 13970
rect 36258 13918 36260 13970
rect 36204 13860 36260 13918
rect 36204 13794 36260 13804
rect 36092 11452 36260 11508
rect 36092 11284 36148 11294
rect 36092 11190 36148 11228
rect 36092 10948 36148 10958
rect 36204 10948 36260 11452
rect 36148 10892 36260 10948
rect 36092 10164 36148 10892
rect 36092 9938 36148 10108
rect 36092 9886 36094 9938
rect 36146 9886 36148 9938
rect 36092 9874 36148 9886
rect 36316 10388 36372 10398
rect 34972 9550 34974 9602
rect 35026 9550 35028 9602
rect 34972 9538 35028 9550
rect 35644 9548 36036 9604
rect 35084 9268 35140 9278
rect 34748 9212 35028 9268
rect 34524 9100 34804 9156
rect 34748 9042 34804 9100
rect 34748 8990 34750 9042
rect 34802 8990 34804 9042
rect 34748 8978 34804 8990
rect 34412 8206 34414 8258
rect 34466 8206 34468 8258
rect 34412 8036 34468 8206
rect 34636 8260 34692 8270
rect 34636 8166 34692 8204
rect 34412 7970 34468 7980
rect 34860 8034 34916 8046
rect 34860 7982 34862 8034
rect 34914 7982 34916 8034
rect 34860 7812 34916 7982
rect 34076 7756 34356 7812
rect 34076 7586 34132 7756
rect 34300 7700 34356 7756
rect 34636 7756 34916 7812
rect 34636 7700 34692 7756
rect 34300 7644 34692 7700
rect 34076 7534 34078 7586
rect 34130 7534 34132 7586
rect 34076 7522 34132 7534
rect 34188 7588 34244 7598
rect 34188 7586 34356 7588
rect 34188 7534 34190 7586
rect 34242 7534 34356 7586
rect 34188 7532 34356 7534
rect 34188 7522 34244 7532
rect 33180 6690 33348 6692
rect 33180 6638 33182 6690
rect 33234 6638 33348 6690
rect 33180 6636 33348 6638
rect 33404 6636 34020 6692
rect 34300 6692 34356 7532
rect 34412 7476 34468 7486
rect 34412 7382 34468 7420
rect 34524 7474 34580 7486
rect 34524 7422 34526 7474
rect 34578 7422 34580 7474
rect 34412 6804 34468 6814
rect 34412 6710 34468 6748
rect 33180 6626 33236 6636
rect 31052 6580 31108 6590
rect 31052 6486 31108 6524
rect 31724 6580 31780 6590
rect 31276 6132 31332 6142
rect 31276 6018 31332 6076
rect 31276 5966 31278 6018
rect 31330 5966 31332 6018
rect 31276 5954 31332 5966
rect 31500 6020 31556 6030
rect 31500 5926 31556 5964
rect 31052 5908 31108 5918
rect 30828 5906 31108 5908
rect 30828 5854 31054 5906
rect 31106 5854 31108 5906
rect 30828 5852 31108 5854
rect 29932 5842 29988 5852
rect 29260 5236 29316 5246
rect 29148 5234 29316 5236
rect 29148 5182 29262 5234
rect 29314 5182 29316 5234
rect 29148 5180 29316 5182
rect 28364 5170 28420 5180
rect 29260 5170 29316 5180
rect 26236 5010 26516 5012
rect 26236 4958 26238 5010
rect 26290 4958 26516 5010
rect 26236 4956 26516 4958
rect 26236 4946 26292 4956
rect 25340 4510 25342 4562
rect 25394 4510 25396 4562
rect 25340 4498 25396 4510
rect 26460 4564 26516 4956
rect 26572 4946 26628 4956
rect 26684 5068 27188 5124
rect 28140 5124 28196 5134
rect 26572 4564 26628 4574
rect 26460 4562 26628 4564
rect 26460 4510 26574 4562
rect 26626 4510 26628 4562
rect 26460 4508 26628 4510
rect 26572 4498 26628 4508
rect 26684 4450 26740 5068
rect 26684 4398 26686 4450
rect 26738 4398 26740 4450
rect 26684 4386 26740 4398
rect 27356 5012 27412 5022
rect 27356 4338 27412 4956
rect 28140 4450 28196 5068
rect 29036 5124 29092 5134
rect 29932 5124 29988 5134
rect 29092 5068 29204 5124
rect 29036 5058 29092 5068
rect 29148 5010 29204 5068
rect 29932 5030 29988 5068
rect 29148 4958 29150 5010
rect 29202 4958 29204 5010
rect 29148 4946 29204 4958
rect 28140 4398 28142 4450
rect 28194 4398 28196 4450
rect 28140 4386 28196 4398
rect 27356 4286 27358 4338
rect 27410 4286 27412 4338
rect 27356 4274 27412 4286
rect 24444 4174 24446 4226
rect 24498 4174 24500 4226
rect 24444 4162 24500 4174
rect 30268 4226 30324 5852
rect 31052 5236 31108 5852
rect 31052 5170 31108 5180
rect 31164 5906 31220 5918
rect 31164 5854 31166 5906
rect 31218 5854 31220 5906
rect 30604 5012 30660 5022
rect 30604 5010 31108 5012
rect 30604 4958 30606 5010
rect 30658 4958 31108 5010
rect 30604 4956 31108 4958
rect 30604 4946 30660 4956
rect 31052 4562 31108 4956
rect 31052 4510 31054 4562
rect 31106 4510 31108 4562
rect 31052 4498 31108 4510
rect 31164 4450 31220 5854
rect 31724 5908 31780 6524
rect 32060 6466 32116 6478
rect 32060 6414 32062 6466
rect 32114 6414 32116 6466
rect 31836 5908 31892 5918
rect 31724 5906 31892 5908
rect 31724 5854 31838 5906
rect 31890 5854 31892 5906
rect 31724 5852 31892 5854
rect 31836 5842 31892 5852
rect 31948 5908 32004 5918
rect 32060 5908 32116 6414
rect 31948 5906 32116 5908
rect 31948 5854 31950 5906
rect 32002 5854 32116 5906
rect 31948 5852 32116 5854
rect 32396 6466 32452 6478
rect 32396 6414 32398 6466
rect 32450 6414 32452 6466
rect 31948 5842 32004 5852
rect 32396 5348 32452 6414
rect 32844 6468 32900 6478
rect 32844 6374 32900 6412
rect 32620 6244 32676 6254
rect 32620 6130 32676 6188
rect 32620 6078 32622 6130
rect 32674 6078 32676 6130
rect 32620 6066 32676 6078
rect 33068 6132 33124 6142
rect 33068 6038 33124 6076
rect 32396 5282 32452 5292
rect 33404 5906 33460 6636
rect 34300 6626 34356 6636
rect 34076 6244 34132 6254
rect 33740 6020 33796 6030
rect 33740 5926 33796 5964
rect 34076 6018 34132 6188
rect 34076 5966 34078 6018
rect 34130 5966 34132 6018
rect 34076 5954 34132 5966
rect 33404 5854 33406 5906
rect 33458 5854 33460 5906
rect 32732 5236 32788 5246
rect 32732 5142 32788 5180
rect 31164 4398 31166 4450
rect 31218 4398 31220 4450
rect 31164 4386 31220 4398
rect 33180 5124 33236 5134
rect 33180 4338 33236 5068
rect 33404 5012 33460 5854
rect 33516 5908 33572 5918
rect 34524 5908 34580 7422
rect 34636 6914 34692 7644
rect 34636 6862 34638 6914
rect 34690 6862 34692 6914
rect 34636 6850 34692 6862
rect 34748 7588 34804 7598
rect 34748 6804 34804 7532
rect 34860 7588 34916 7598
rect 34972 7588 35028 9212
rect 35084 9174 35140 9212
rect 35644 9266 35700 9548
rect 35644 9214 35646 9266
rect 35698 9214 35700 9266
rect 35644 9202 35700 9214
rect 35196 8652 35460 8662
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35196 8586 35460 8596
rect 35644 8260 35700 8270
rect 35084 8146 35140 8158
rect 35084 8094 35086 8146
rect 35138 8094 35140 8146
rect 35084 7812 35140 8094
rect 35084 7746 35140 7756
rect 35308 8146 35364 8158
rect 35308 8094 35310 8146
rect 35362 8094 35364 8146
rect 35308 7812 35364 8094
rect 35644 8146 35700 8204
rect 35644 8094 35646 8146
rect 35698 8094 35700 8146
rect 35644 8082 35700 8094
rect 35364 7756 35588 7812
rect 35308 7746 35364 7756
rect 34860 7586 35028 7588
rect 34860 7534 34862 7586
rect 34914 7534 35028 7586
rect 34860 7532 35028 7534
rect 35420 7588 35476 7598
rect 34860 7476 34916 7532
rect 35420 7494 35476 7532
rect 34860 7410 34916 7420
rect 35196 7084 35460 7094
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35196 7018 35460 7028
rect 34748 6738 34804 6748
rect 34860 6692 34916 6702
rect 34860 6578 34916 6636
rect 35308 6692 35364 6702
rect 35308 6598 35364 6636
rect 34860 6526 34862 6578
rect 34914 6526 34916 6578
rect 34860 6514 34916 6526
rect 34748 6466 34804 6478
rect 34748 6414 34750 6466
rect 34802 6414 34804 6466
rect 34636 5908 34692 5918
rect 34524 5906 34692 5908
rect 34524 5854 34638 5906
rect 34690 5854 34692 5906
rect 34524 5852 34692 5854
rect 33516 5234 33572 5852
rect 34636 5842 34692 5852
rect 34748 5906 34804 6414
rect 34972 6020 35028 6030
rect 34972 5926 35028 5964
rect 35532 6018 35588 7756
rect 35532 5966 35534 6018
rect 35586 5966 35588 6018
rect 34748 5854 34750 5906
rect 34802 5854 34804 5906
rect 34748 5842 34804 5854
rect 35308 5906 35364 5918
rect 35308 5854 35310 5906
rect 35362 5854 35364 5906
rect 35308 5796 35364 5854
rect 35420 5908 35476 5918
rect 35420 5814 35476 5852
rect 35308 5730 35364 5740
rect 35532 5684 35588 5966
rect 35532 5618 35588 5628
rect 35644 7698 35700 7710
rect 35644 7646 35646 7698
rect 35698 7646 35700 7698
rect 35644 6802 35700 7646
rect 35756 7700 35812 9548
rect 35868 9380 35924 9390
rect 35868 9042 35924 9324
rect 35868 8990 35870 9042
rect 35922 8990 35924 9042
rect 35868 8978 35924 8990
rect 35980 8036 36036 8046
rect 36204 8036 36260 8046
rect 35980 8034 36148 8036
rect 35980 7982 35982 8034
rect 36034 7982 36148 8034
rect 35980 7980 36148 7982
rect 35980 7970 36036 7980
rect 35756 7634 35812 7644
rect 36092 7588 36148 7980
rect 36092 7522 36148 7532
rect 35756 7476 35812 7486
rect 35756 7382 35812 7420
rect 35980 7474 36036 7486
rect 35980 7422 35982 7474
rect 36034 7422 36036 7474
rect 35644 6750 35646 6802
rect 35698 6750 35700 6802
rect 35196 5516 35460 5526
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35196 5450 35460 5460
rect 33516 5182 33518 5234
rect 33570 5182 33572 5234
rect 33516 5170 33572 5182
rect 35308 5348 35364 5358
rect 35644 5348 35700 6750
rect 35868 6690 35924 6702
rect 35868 6638 35870 6690
rect 35922 6638 35924 6690
rect 35868 6132 35924 6638
rect 35980 6692 36036 7422
rect 35980 6626 36036 6636
rect 35868 6066 35924 6076
rect 36092 6580 36148 6590
rect 36092 5906 36148 6524
rect 36092 5854 36094 5906
rect 36146 5854 36148 5906
rect 36092 5842 36148 5854
rect 35980 5682 36036 5694
rect 35980 5630 35982 5682
rect 36034 5630 36036 5682
rect 35980 5572 36036 5630
rect 33516 5012 33572 5022
rect 33404 4956 33516 5012
rect 33516 4946 33572 4956
rect 33628 4900 33684 4910
rect 33628 4898 33908 4900
rect 33628 4846 33630 4898
rect 33682 4846 33908 4898
rect 33628 4844 33908 4846
rect 33628 4834 33684 4844
rect 33852 4450 33908 4844
rect 35308 4788 35364 5292
rect 35420 5292 35700 5348
rect 35756 5516 36036 5572
rect 36092 5684 36148 5694
rect 35420 5122 35476 5292
rect 35756 5236 35812 5516
rect 36092 5460 36148 5628
rect 35980 5404 36148 5460
rect 35420 5070 35422 5122
rect 35474 5070 35476 5122
rect 35420 5058 35476 5070
rect 35532 5180 35812 5236
rect 35868 5236 35924 5246
rect 35532 5122 35588 5180
rect 35868 5124 35924 5180
rect 35532 5070 35534 5122
rect 35586 5070 35588 5122
rect 35532 5058 35588 5070
rect 35644 5068 35924 5124
rect 35644 5010 35700 5068
rect 35644 4958 35646 5010
rect 35698 4958 35700 5010
rect 35644 4946 35700 4958
rect 35868 4898 35924 4910
rect 35868 4846 35870 4898
rect 35922 4846 35924 4898
rect 35868 4788 35924 4846
rect 35308 4732 35924 4788
rect 33852 4398 33854 4450
rect 33906 4398 33908 4450
rect 33852 4386 33908 4398
rect 33180 4286 33182 4338
rect 33234 4286 33236 4338
rect 33180 4274 33236 4286
rect 30268 4174 30270 4226
rect 30322 4174 30324 4226
rect 30268 4162 30324 4174
rect 35980 4226 36036 5404
rect 36092 5124 36148 5134
rect 36204 5124 36260 7980
rect 36316 7588 36372 10332
rect 36540 9940 36596 9950
rect 36652 9940 36708 16604
rect 36764 13524 36820 17164
rect 36876 15652 36932 17948
rect 37212 17890 37268 18396
rect 37212 17838 37214 17890
rect 37266 17838 37268 17890
rect 37212 17826 37268 17838
rect 37100 17554 37156 17566
rect 37100 17502 37102 17554
rect 37154 17502 37156 17554
rect 37100 17108 37156 17502
rect 37100 17042 37156 17052
rect 37212 17442 37268 17454
rect 37212 17390 37214 17442
rect 37266 17390 37268 17442
rect 36988 16658 37044 16670
rect 36988 16606 36990 16658
rect 37042 16606 37044 16658
rect 36988 16324 37044 16606
rect 37100 16660 37156 16670
rect 37100 16566 37156 16604
rect 36988 16258 37044 16268
rect 37212 16212 37268 17390
rect 37212 16146 37268 16156
rect 36876 15586 36932 15596
rect 37324 14532 37380 19628
rect 37548 19572 37604 19852
rect 37548 19506 37604 19516
rect 37660 20636 37828 20692
rect 37548 19122 37604 19134
rect 37548 19070 37550 19122
rect 37602 19070 37604 19122
rect 37548 19012 37604 19070
rect 37548 18946 37604 18956
rect 37660 17780 37716 20636
rect 37660 17714 37716 17724
rect 37772 20132 37828 20142
rect 37772 19124 37828 20076
rect 37772 17778 37828 19068
rect 37884 19010 37940 19022
rect 37884 18958 37886 19010
rect 37938 18958 37940 19010
rect 37884 17892 37940 18958
rect 37996 19012 38052 23996
rect 38556 23828 38612 23838
rect 38556 23734 38612 23772
rect 39564 23380 39620 23390
rect 39564 23286 39620 23324
rect 38556 23268 38612 23278
rect 38332 22258 38388 22270
rect 38332 22206 38334 22258
rect 38386 22206 38388 22258
rect 38332 21588 38388 22206
rect 38332 21522 38388 21532
rect 38556 21586 38612 23212
rect 39116 23042 39172 23054
rect 39116 22990 39118 23042
rect 39170 22990 39172 23042
rect 39116 21812 39172 22990
rect 40012 22932 40068 32284
rect 40012 22866 40068 22876
rect 40124 32228 40180 32238
rect 39116 21756 39620 21812
rect 38556 21534 38558 21586
rect 38610 21534 38612 21586
rect 38108 21474 38164 21486
rect 38108 21422 38110 21474
rect 38162 21422 38164 21474
rect 38108 20132 38164 21422
rect 38220 21364 38276 21374
rect 38220 20804 38276 21308
rect 38556 21364 38612 21534
rect 38556 21298 38612 21308
rect 38668 21588 38724 21598
rect 38668 21252 38724 21532
rect 38668 21186 38724 21196
rect 38892 21476 38948 21486
rect 39116 21476 39172 21756
rect 39564 21698 39620 21756
rect 39564 21646 39566 21698
rect 39618 21646 39620 21698
rect 39564 21634 39620 21646
rect 40012 21700 40068 21710
rect 38892 21474 39172 21476
rect 38892 21422 38894 21474
rect 38946 21422 39172 21474
rect 38892 21420 39172 21422
rect 39228 21588 39284 21598
rect 38220 20802 38500 20804
rect 38220 20750 38222 20802
rect 38274 20750 38500 20802
rect 38220 20748 38500 20750
rect 38220 20738 38276 20748
rect 38444 20188 38500 20748
rect 38556 20692 38612 20702
rect 38556 20598 38612 20636
rect 38892 20244 38948 21420
rect 39228 21252 39284 21532
rect 39228 21186 39284 21196
rect 39340 21586 39396 21598
rect 39340 21534 39342 21586
rect 39394 21534 39396 21586
rect 39340 20914 39396 21534
rect 39788 21588 39844 21598
rect 39788 21494 39844 21532
rect 40012 21586 40068 21644
rect 40012 21534 40014 21586
rect 40066 21534 40068 21586
rect 40012 21522 40068 21534
rect 40124 21140 40180 32172
rect 40460 30436 40516 36988
rect 41356 36708 41412 37324
rect 41468 37314 41524 37324
rect 41580 37268 41636 37278
rect 41580 37174 41636 37212
rect 41468 37044 41524 37054
rect 41692 37044 41748 39454
rect 42364 39506 42420 39518
rect 42700 39508 42756 39518
rect 42364 39454 42366 39506
rect 42418 39454 42420 39506
rect 41804 39394 41860 39406
rect 41804 39342 41806 39394
rect 41858 39342 41860 39394
rect 41804 38946 41860 39342
rect 41804 38894 41806 38946
rect 41858 38894 41860 38946
rect 41804 38882 41860 38894
rect 42028 38276 42084 38286
rect 42028 38182 42084 38220
rect 42364 38276 42420 39454
rect 42364 38162 42420 38220
rect 42364 38110 42366 38162
rect 42418 38110 42420 38162
rect 41916 37492 41972 37502
rect 41916 37398 41972 37436
rect 42364 37378 42420 38110
rect 42476 39506 42756 39508
rect 42476 39454 42702 39506
rect 42754 39454 42756 39506
rect 42476 39452 42756 39454
rect 42476 38052 42532 39452
rect 42700 39442 42756 39452
rect 42812 38836 42868 40348
rect 44156 40180 44212 40190
rect 44044 40124 44156 40180
rect 43372 39732 43428 39742
rect 43260 39620 43316 39630
rect 42476 37986 42532 37996
rect 42588 38780 42868 38836
rect 42924 39506 42980 39518
rect 42924 39454 42926 39506
rect 42978 39454 42980 39506
rect 42364 37326 42366 37378
rect 42418 37326 42420 37378
rect 42364 37314 42420 37326
rect 42140 37266 42196 37278
rect 42140 37214 42142 37266
rect 42194 37214 42196 37266
rect 42140 37156 42196 37214
rect 42140 37090 42196 37100
rect 42252 37268 42308 37278
rect 41468 37042 41748 37044
rect 41468 36990 41470 37042
rect 41522 36990 41748 37042
rect 41468 36988 41748 36990
rect 42252 37042 42308 37212
rect 42252 36990 42254 37042
rect 42306 36990 42308 37042
rect 41468 36978 41524 36988
rect 41356 36652 41524 36708
rect 41356 35252 41412 35262
rect 41020 34132 41076 34142
rect 41356 34132 41412 35196
rect 41468 34244 41524 36652
rect 41804 36596 41860 36606
rect 41804 36502 41860 36540
rect 42252 36482 42308 36990
rect 42588 36708 42644 38780
rect 42924 38724 42980 39454
rect 42700 38668 42924 38724
rect 42700 37492 42756 38668
rect 42924 38658 42980 38668
rect 42812 38052 42868 38062
rect 42868 37996 42980 38052
rect 42812 37958 42868 37996
rect 42700 37266 42756 37436
rect 42700 37214 42702 37266
rect 42754 37214 42756 37266
rect 42700 37202 42756 37214
rect 42924 37156 42980 37996
rect 42924 37062 42980 37100
rect 43148 37044 43204 37054
rect 43036 37042 43204 37044
rect 43036 36990 43150 37042
rect 43202 36990 43204 37042
rect 43036 36988 43204 36990
rect 42588 36652 42756 36708
rect 42252 36430 42254 36482
rect 42306 36430 42308 36482
rect 42252 36418 42308 36430
rect 42140 36372 42196 36382
rect 42140 36278 42196 36316
rect 42700 35698 42756 36652
rect 42812 36596 42868 36606
rect 42812 36484 42868 36540
rect 43036 36484 43092 36988
rect 43148 36978 43204 36988
rect 42812 36482 43092 36484
rect 42812 36430 42814 36482
rect 42866 36430 43092 36482
rect 42812 36428 43092 36430
rect 42812 36418 42868 36428
rect 43260 35700 43316 39564
rect 43372 37380 43428 39676
rect 43932 38724 43988 38734
rect 43932 38630 43988 38668
rect 43820 38276 43876 38286
rect 43820 38182 43876 38220
rect 43932 38276 43988 38286
rect 44044 38276 44100 40124
rect 44156 40114 44212 40124
rect 43932 38274 44100 38276
rect 43932 38222 43934 38274
rect 43986 38222 44100 38274
rect 43932 38220 44100 38222
rect 44156 39732 44212 39742
rect 44156 38274 44212 39676
rect 45164 38668 45220 43652
rect 45724 41972 45780 53340
rect 45948 52388 46004 59200
rect 47404 56308 47460 56318
rect 47404 56306 47572 56308
rect 47404 56254 47406 56306
rect 47458 56254 47572 56306
rect 47404 56252 47572 56254
rect 47404 56242 47460 56252
rect 46844 56084 46900 56094
rect 46732 56082 46900 56084
rect 46732 56030 46846 56082
rect 46898 56030 46900 56082
rect 46732 56028 46900 56030
rect 46508 55858 46564 55870
rect 46508 55806 46510 55858
rect 46562 55806 46564 55858
rect 46508 54068 46564 55806
rect 46732 55468 46788 56028
rect 46844 56018 46900 56028
rect 46844 55860 46900 55870
rect 46844 55858 47348 55860
rect 46844 55806 46846 55858
rect 46898 55806 47348 55858
rect 46844 55804 47348 55806
rect 46844 55794 46900 55804
rect 46732 55412 47124 55468
rect 46508 54002 46564 54012
rect 46620 52388 46676 52398
rect 45948 52386 46676 52388
rect 45948 52334 46622 52386
rect 46674 52334 46676 52386
rect 45948 52332 46676 52334
rect 46620 52322 46676 52332
rect 47068 50706 47124 55412
rect 47292 53732 47348 55804
rect 47516 55468 47572 56252
rect 47628 56252 48468 56308
rect 47628 56082 47684 56252
rect 47628 56030 47630 56082
rect 47682 56030 47684 56082
rect 47628 56018 47684 56030
rect 47852 56084 47908 56094
rect 47852 55990 47908 56028
rect 48188 56082 48244 56094
rect 48188 56030 48190 56082
rect 48242 56030 48244 56082
rect 47628 55860 47684 55870
rect 47628 55766 47684 55804
rect 47404 55412 47572 55468
rect 47404 55410 47460 55412
rect 47404 55358 47406 55410
rect 47458 55358 47460 55410
rect 47404 55346 47460 55358
rect 48076 55298 48132 55310
rect 48076 55246 48078 55298
rect 48130 55246 48132 55298
rect 47852 54514 47908 54526
rect 47852 54462 47854 54514
rect 47906 54462 47908 54514
rect 47404 53732 47460 53742
rect 47292 53730 47460 53732
rect 47292 53678 47406 53730
rect 47458 53678 47460 53730
rect 47292 53676 47460 53678
rect 47404 53666 47460 53676
rect 47516 52836 47572 52846
rect 47516 52742 47572 52780
rect 47740 52612 47796 52622
rect 47404 51492 47460 51502
rect 47404 51398 47460 51436
rect 47068 50654 47070 50706
rect 47122 50654 47124 50706
rect 47068 50642 47124 50654
rect 47516 50818 47572 50830
rect 47516 50766 47518 50818
rect 47570 50766 47572 50818
rect 47516 50706 47572 50766
rect 47516 50654 47518 50706
rect 47570 50654 47572 50706
rect 47516 50642 47572 50654
rect 46844 50484 46900 50494
rect 46844 50390 46900 50428
rect 46396 49924 46452 49934
rect 46396 49830 46452 49868
rect 45836 49810 45892 49822
rect 45836 49758 45838 49810
rect 45890 49758 45892 49810
rect 45836 48804 45892 49758
rect 46732 49812 46788 49822
rect 46732 49718 46788 49756
rect 47740 49810 47796 52556
rect 47852 50484 47908 54462
rect 48076 53732 48132 55246
rect 48188 54738 48244 56030
rect 48188 54686 48190 54738
rect 48242 54686 48244 54738
rect 48188 54674 48244 54686
rect 48076 53730 48244 53732
rect 48076 53678 48078 53730
rect 48130 53678 48244 53730
rect 48076 53676 48244 53678
rect 48076 53666 48132 53676
rect 48076 53508 48132 53518
rect 47964 52946 48020 52958
rect 47964 52894 47966 52946
rect 48018 52894 48020 52946
rect 47964 52612 48020 52894
rect 47964 52546 48020 52556
rect 48076 50706 48132 53452
rect 48076 50654 48078 50706
rect 48130 50654 48132 50706
rect 48076 50642 48132 50654
rect 48188 51378 48244 53676
rect 48188 51326 48190 51378
rect 48242 51326 48244 51378
rect 48188 50818 48244 51326
rect 48188 50766 48190 50818
rect 48242 50766 48244 50818
rect 47852 49922 47908 50428
rect 47852 49870 47854 49922
rect 47906 49870 47908 49922
rect 47852 49858 47908 49870
rect 47740 49758 47742 49810
rect 47794 49758 47796 49810
rect 47740 49746 47796 49758
rect 46284 49700 46340 49710
rect 46284 49606 46340 49644
rect 47404 49698 47460 49710
rect 47404 49646 47406 49698
rect 47458 49646 47460 49698
rect 47404 49252 47460 49646
rect 47404 49186 47460 49196
rect 45836 48710 45892 48748
rect 46396 49028 46452 49038
rect 45948 48580 46004 48590
rect 45948 46114 46004 48524
rect 46060 47236 46116 47246
rect 46116 47180 46340 47236
rect 46060 47170 46116 47180
rect 45948 46062 45950 46114
rect 46002 46062 46004 46114
rect 45948 46050 46004 46062
rect 46284 46114 46340 47180
rect 46284 46062 46286 46114
rect 46338 46062 46340 46114
rect 46284 46050 46340 46062
rect 45836 45892 45892 45902
rect 45836 45798 45892 45836
rect 46172 45890 46228 45902
rect 46172 45838 46174 45890
rect 46226 45838 46228 45890
rect 46172 45332 46228 45838
rect 46172 44100 46228 45276
rect 46284 45220 46340 45230
rect 46284 45106 46340 45164
rect 46284 45054 46286 45106
rect 46338 45054 46340 45106
rect 46284 45042 46340 45054
rect 46172 44034 46228 44044
rect 46396 43708 46452 48972
rect 47628 49028 47684 49038
rect 48188 49028 48244 50766
rect 47628 48934 47684 48972
rect 48076 48972 48244 49028
rect 48300 50260 48356 50270
rect 46732 48914 46788 48926
rect 46732 48862 46734 48914
rect 46786 48862 46788 48914
rect 46508 48802 46564 48814
rect 46508 48750 46510 48802
rect 46562 48750 46564 48802
rect 46508 45892 46564 48750
rect 46620 48802 46676 48814
rect 46620 48750 46622 48802
rect 46674 48750 46676 48802
rect 46620 48356 46676 48750
rect 46620 48290 46676 48300
rect 46732 47682 46788 48862
rect 47404 48804 47460 48814
rect 47404 48710 47460 48748
rect 48076 48692 48132 48972
rect 48188 48804 48244 48814
rect 48300 48804 48356 50204
rect 48244 48748 48356 48804
rect 48188 48710 48244 48748
rect 47404 48356 47460 48366
rect 47404 48262 47460 48300
rect 46732 47630 46734 47682
rect 46786 47630 46788 47682
rect 46732 47618 46788 47630
rect 48076 48242 48132 48636
rect 48076 48190 48078 48242
rect 48130 48190 48132 48242
rect 46844 47572 46900 47582
rect 46844 47478 46900 47516
rect 47964 47572 48020 47582
rect 46620 47458 46676 47470
rect 46620 47406 46622 47458
rect 46674 47406 46676 47458
rect 46620 47348 46676 47406
rect 47404 47460 47460 47470
rect 47404 47366 47460 47404
rect 47964 47458 48020 47516
rect 47964 47406 47966 47458
rect 48018 47406 48020 47458
rect 46620 47282 46676 47292
rect 47628 47348 47684 47358
rect 47628 47254 47684 47292
rect 47740 47234 47796 47246
rect 47740 47182 47742 47234
rect 47794 47182 47796 47234
rect 47404 46564 47460 46574
rect 46956 46562 47460 46564
rect 46956 46510 47406 46562
rect 47458 46510 47460 46562
rect 46956 46508 47460 46510
rect 46956 46002 47012 46508
rect 47404 46498 47460 46508
rect 47740 46340 47796 47182
rect 47068 46284 47796 46340
rect 47068 46114 47124 46284
rect 47068 46062 47070 46114
rect 47122 46062 47124 46114
rect 47068 46050 47124 46062
rect 46956 45950 46958 46002
rect 47010 45950 47012 46002
rect 46956 45938 47012 45950
rect 46732 45892 46788 45902
rect 46508 45890 46788 45892
rect 46508 45838 46734 45890
rect 46786 45838 46788 45890
rect 46508 45836 46788 45838
rect 46284 43652 46452 43708
rect 46508 45108 46564 45118
rect 45724 41906 45780 41916
rect 46060 42084 46116 42094
rect 45724 41748 45780 41758
rect 45724 41654 45780 41692
rect 46060 41298 46116 42028
rect 46060 41246 46062 41298
rect 46114 41246 46116 41298
rect 46060 41234 46116 41246
rect 45388 41186 45444 41198
rect 45388 41134 45390 41186
rect 45442 41134 45444 41186
rect 45388 40404 45444 41134
rect 45388 40338 45444 40348
rect 45612 40516 45668 40526
rect 45500 40292 45556 40302
rect 45500 40198 45556 40236
rect 45612 39842 45668 40460
rect 45948 40514 46004 40526
rect 45948 40462 45950 40514
rect 46002 40462 46004 40514
rect 45836 40180 45892 40190
rect 45836 40086 45892 40124
rect 45612 39790 45614 39842
rect 45666 39790 45668 39842
rect 45612 39778 45668 39790
rect 45836 39620 45892 39630
rect 45948 39620 46004 40462
rect 46172 40516 46228 40526
rect 46172 40290 46228 40460
rect 46172 40238 46174 40290
rect 46226 40238 46228 40290
rect 46172 40226 46228 40238
rect 46284 39620 46340 43652
rect 46508 43540 46564 45052
rect 46620 45106 46676 45118
rect 46620 45054 46622 45106
rect 46674 45054 46676 45106
rect 46620 44436 46676 45054
rect 46732 44996 46788 45836
rect 47628 45890 47684 45902
rect 47628 45838 47630 45890
rect 47682 45838 47684 45890
rect 47628 45556 47684 45838
rect 47628 45490 47684 45500
rect 47068 45332 47124 45342
rect 47964 45332 48020 47406
rect 47068 45330 48020 45332
rect 47068 45278 47070 45330
rect 47122 45278 48020 45330
rect 47068 45276 48020 45278
rect 47068 45266 47124 45276
rect 47964 45106 48020 45276
rect 47964 45054 47966 45106
rect 48018 45054 48020 45106
rect 47964 45042 48020 45054
rect 48076 46674 48132 48190
rect 48076 46622 48078 46674
rect 48130 46622 48132 46674
rect 46732 44930 46788 44940
rect 47516 44996 47572 45006
rect 47516 44902 47572 44940
rect 46620 44370 46676 44380
rect 47180 44884 47236 44894
rect 47180 44324 47236 44828
rect 47404 44882 47460 44894
rect 47404 44830 47406 44882
rect 47458 44830 47460 44882
rect 47068 44268 47236 44324
rect 47292 44436 47348 44446
rect 47068 43762 47124 44268
rect 47068 43710 47070 43762
rect 47122 43710 47124 43762
rect 47068 43698 47124 43710
rect 47180 44100 47236 44110
rect 47180 43650 47236 44044
rect 47180 43598 47182 43650
rect 47234 43598 47236 43650
rect 47180 43586 47236 43598
rect 46732 43540 46788 43550
rect 46508 43538 46788 43540
rect 46508 43486 46734 43538
rect 46786 43486 46788 43538
rect 46508 43484 46788 43486
rect 46508 43426 46564 43484
rect 46732 43474 46788 43484
rect 47292 43538 47348 44380
rect 47404 44434 47460 44830
rect 47740 44884 47796 44894
rect 47740 44790 47796 44828
rect 47404 44382 47406 44434
rect 47458 44382 47460 44434
rect 47404 44370 47460 44382
rect 48076 44322 48132 46622
rect 48076 44270 48078 44322
rect 48130 44270 48132 44322
rect 48076 44258 48132 44270
rect 48188 45666 48244 45678
rect 48188 45614 48190 45666
rect 48242 45614 48244 45666
rect 48188 44436 48244 45614
rect 48188 43652 48244 44380
rect 48300 43652 48356 43662
rect 48188 43650 48356 43652
rect 48188 43598 48302 43650
rect 48354 43598 48356 43650
rect 48188 43596 48356 43598
rect 48300 43586 48356 43596
rect 47292 43486 47294 43538
rect 47346 43486 47348 43538
rect 47292 43474 47348 43486
rect 46508 43374 46510 43426
rect 46562 43374 46564 43426
rect 46508 43362 46564 43374
rect 46732 42532 46788 42542
rect 47180 42532 47236 42542
rect 46732 42530 47180 42532
rect 46732 42478 46734 42530
rect 46786 42478 47180 42530
rect 46732 42476 47180 42478
rect 46732 42466 46788 42476
rect 47068 42084 47124 42094
rect 47068 41990 47124 42028
rect 46508 41972 46564 41982
rect 46508 41970 46788 41972
rect 46508 41918 46510 41970
rect 46562 41918 46788 41970
rect 46508 41916 46788 41918
rect 46508 41906 46564 41916
rect 46396 41858 46452 41870
rect 46396 41806 46398 41858
rect 46450 41806 46452 41858
rect 46396 40292 46452 41806
rect 46396 40226 46452 40236
rect 46732 40402 46788 41916
rect 47180 41746 47236 42476
rect 48300 42530 48356 42542
rect 48300 42478 48302 42530
rect 48354 42478 48356 42530
rect 48076 41972 48132 41982
rect 47964 41916 48076 41972
rect 47404 41748 47460 41758
rect 47180 41694 47182 41746
rect 47234 41694 47236 41746
rect 46732 40350 46734 40402
rect 46786 40350 46788 40402
rect 46732 39732 46788 40350
rect 46956 40402 47012 40414
rect 46956 40350 46958 40402
rect 47010 40350 47012 40402
rect 46956 40180 47012 40350
rect 46956 40114 47012 40124
rect 47068 40402 47124 40414
rect 47068 40350 47070 40402
rect 47122 40350 47124 40402
rect 47068 40068 47124 40350
rect 47068 39956 47124 40012
rect 45836 39618 46004 39620
rect 45836 39566 45838 39618
rect 45890 39566 46004 39618
rect 45836 39564 46004 39566
rect 45836 39554 45892 39564
rect 45500 39508 45556 39518
rect 44156 38222 44158 38274
rect 44210 38222 44212 38274
rect 43932 38210 43988 38220
rect 44156 38210 44212 38222
rect 45052 38612 45220 38668
rect 45276 39394 45332 39406
rect 45276 39342 45278 39394
rect 45330 39342 45332 39394
rect 44268 37940 44324 37950
rect 44268 37938 44660 37940
rect 44268 37886 44270 37938
rect 44322 37886 44660 37938
rect 44268 37884 44660 37886
rect 44268 37874 44324 37884
rect 43372 37314 43428 37324
rect 43596 37380 43652 37390
rect 43596 37286 43652 37324
rect 44604 37378 44660 37884
rect 44604 37326 44606 37378
rect 44658 37326 44660 37378
rect 44604 37314 44660 37326
rect 42700 35646 42702 35698
rect 42754 35646 42756 35698
rect 42700 35364 42756 35646
rect 42700 35298 42756 35308
rect 42924 35644 43316 35700
rect 43820 37266 43876 37278
rect 43820 37214 43822 37266
rect 43874 37214 43876 37266
rect 41468 34178 41524 34188
rect 41020 34130 41412 34132
rect 41020 34078 41022 34130
rect 41074 34078 41412 34130
rect 41020 34076 41412 34078
rect 41020 34066 41076 34076
rect 40348 30380 40516 30436
rect 40796 33572 40852 33582
rect 40236 27188 40292 27198
rect 40236 27094 40292 27132
rect 40348 26964 40404 30380
rect 40796 30322 40852 33516
rect 41244 33460 41300 33470
rect 41020 33236 41076 33246
rect 41020 33142 41076 33180
rect 41244 32674 41300 33404
rect 41244 32622 41246 32674
rect 41298 32622 41300 32674
rect 41244 32610 41300 32622
rect 41356 33348 41412 34076
rect 41692 34020 41748 34030
rect 41692 33926 41748 33964
rect 41356 31778 41412 33292
rect 41692 33460 41748 33470
rect 41356 31726 41358 31778
rect 41410 31726 41412 31778
rect 41356 31714 41412 31726
rect 41468 32338 41524 32350
rect 41468 32286 41470 32338
rect 41522 32286 41524 32338
rect 41468 31892 41524 32286
rect 41356 31108 41412 31118
rect 41468 31108 41524 31836
rect 41356 31106 41524 31108
rect 41356 31054 41358 31106
rect 41410 31054 41524 31106
rect 41356 31052 41524 31054
rect 41580 31780 41636 31790
rect 41356 31042 41412 31052
rect 41580 30882 41636 31724
rect 41692 30994 41748 33404
rect 41804 32338 41860 32350
rect 41804 32286 41806 32338
rect 41858 32286 41860 32338
rect 41804 31220 41860 32286
rect 42028 31668 42084 31678
rect 42028 31574 42084 31612
rect 41804 31154 41860 31164
rect 42476 31220 42532 31230
rect 42532 31164 42756 31220
rect 42476 31126 42532 31164
rect 41692 30942 41694 30994
rect 41746 30942 41748 30994
rect 41692 30930 41748 30942
rect 41580 30830 41582 30882
rect 41634 30830 41636 30882
rect 41580 30818 41636 30830
rect 40796 30270 40798 30322
rect 40850 30270 40852 30322
rect 40796 30258 40852 30270
rect 40460 30210 40516 30222
rect 41020 30212 41076 30222
rect 40460 30158 40462 30210
rect 40514 30158 40516 30210
rect 40460 29204 40516 30158
rect 40908 30210 41076 30212
rect 40908 30158 41022 30210
rect 41074 30158 41076 30210
rect 40908 30156 41076 30158
rect 40796 29204 40852 29214
rect 40460 29202 40852 29204
rect 40460 29150 40798 29202
rect 40850 29150 40852 29202
rect 40460 29148 40852 29150
rect 40796 29138 40852 29148
rect 40908 28756 40964 30156
rect 41020 30146 41076 30156
rect 42252 30210 42308 30222
rect 42252 30158 42254 30210
rect 42306 30158 42308 30210
rect 41356 29988 41412 29998
rect 41356 29894 41412 29932
rect 42028 29986 42084 29998
rect 42028 29934 42030 29986
rect 42082 29934 42084 29986
rect 40348 26898 40404 26908
rect 40796 28700 40964 28756
rect 41020 29314 41076 29326
rect 41020 29262 41022 29314
rect 41074 29262 41076 29314
rect 41020 29202 41076 29262
rect 41020 29150 41022 29202
rect 41074 29150 41076 29202
rect 40348 25956 40404 25966
rect 40348 25618 40404 25900
rect 40348 25566 40350 25618
rect 40402 25566 40404 25618
rect 40348 25554 40404 25566
rect 40684 24052 40740 24062
rect 40796 24052 40852 28700
rect 41020 28644 41076 29150
rect 41356 28644 41412 28654
rect 41020 28642 41412 28644
rect 41020 28590 41358 28642
rect 41410 28590 41412 28642
rect 41020 28588 41412 28590
rect 40908 28532 40964 28542
rect 40908 28082 40964 28476
rect 40908 28030 40910 28082
rect 40962 28030 40964 28082
rect 40908 28018 40964 28030
rect 41132 27858 41188 27870
rect 41132 27806 41134 27858
rect 41186 27806 41188 27858
rect 41020 27746 41076 27758
rect 41020 27694 41022 27746
rect 41074 27694 41076 27746
rect 41020 27188 41076 27694
rect 41020 27122 41076 27132
rect 41132 27524 41188 27806
rect 41356 27748 41412 28588
rect 41916 28084 41972 28094
rect 41580 28082 41972 28084
rect 41580 28030 41918 28082
rect 41970 28030 41972 28082
rect 41580 28028 41972 28030
rect 41580 27858 41636 28028
rect 41916 28018 41972 28028
rect 41580 27806 41582 27858
rect 41634 27806 41636 27858
rect 41580 27794 41636 27806
rect 41692 27858 41748 27870
rect 41692 27806 41694 27858
rect 41746 27806 41748 27858
rect 41356 27682 41412 27692
rect 41692 27524 41748 27806
rect 41132 27468 41748 27524
rect 42028 27748 42084 29934
rect 42252 29988 42308 30158
rect 42700 30210 42756 31164
rect 42812 31108 42868 31118
rect 42812 31014 42868 31052
rect 42700 30158 42702 30210
rect 42754 30158 42756 30210
rect 42700 30146 42756 30158
rect 42252 29922 42308 29932
rect 42924 29764 42980 35644
rect 43372 35588 43428 35598
rect 43372 35586 43652 35588
rect 43372 35534 43374 35586
rect 43426 35534 43652 35586
rect 43372 35532 43652 35534
rect 43372 35522 43428 35532
rect 43260 35476 43316 35486
rect 43260 35140 43316 35420
rect 43596 35140 43652 35532
rect 43820 35252 43876 37214
rect 43820 35186 43876 35196
rect 43596 35084 43764 35140
rect 43260 35074 43316 35084
rect 43708 35028 43764 35084
rect 44156 35084 44996 35140
rect 43820 35028 43876 35038
rect 43708 35026 43876 35028
rect 43708 34974 43822 35026
rect 43874 34974 43876 35026
rect 43708 34972 43876 34974
rect 43820 34962 43876 34972
rect 44044 34916 44100 34926
rect 44156 34916 44212 35084
rect 44044 34914 44212 34916
rect 44044 34862 44046 34914
rect 44098 34862 44212 34914
rect 44044 34860 44212 34862
rect 44268 34916 44324 34926
rect 44268 34914 44660 34916
rect 44268 34862 44270 34914
rect 44322 34862 44660 34914
rect 44268 34860 44660 34862
rect 44044 34850 44100 34860
rect 44268 34850 44324 34860
rect 43148 34802 43204 34814
rect 43148 34750 43150 34802
rect 43202 34750 43204 34802
rect 43148 33684 43204 34750
rect 43708 34802 43764 34814
rect 43708 34750 43710 34802
rect 43762 34750 43764 34802
rect 43260 34690 43316 34702
rect 43260 34638 43262 34690
rect 43314 34638 43316 34690
rect 43260 34132 43316 34638
rect 43484 34692 43540 34702
rect 43484 34598 43540 34636
rect 43316 34076 43428 34132
rect 43260 34066 43316 34076
rect 43148 33628 43316 33684
rect 43148 33460 43204 33470
rect 43148 33366 43204 33404
rect 43260 33348 43316 33628
rect 43260 31108 43316 33292
rect 43372 32452 43428 34076
rect 43708 33572 43764 34750
rect 44380 34692 44436 34702
rect 43820 34132 43876 34142
rect 43820 34018 43876 34076
rect 43820 33966 43822 34018
rect 43874 33966 43876 34018
rect 43820 33954 43876 33966
rect 44044 34130 44100 34142
rect 44044 34078 44046 34130
rect 44098 34078 44100 34130
rect 43708 33516 43876 33572
rect 43596 33234 43652 33246
rect 43596 33182 43598 33234
rect 43650 33182 43652 33234
rect 43596 32900 43652 33182
rect 43484 32844 43652 32900
rect 43708 33122 43764 33134
rect 43708 33070 43710 33122
rect 43762 33070 43764 33122
rect 43484 32676 43540 32844
rect 43484 32582 43540 32620
rect 43596 32674 43652 32686
rect 43596 32622 43598 32674
rect 43650 32622 43652 32674
rect 43596 32452 43652 32622
rect 43372 32396 43652 32452
rect 43596 32228 43652 32238
rect 43372 31780 43428 31790
rect 43428 31724 43540 31780
rect 43372 31714 43428 31724
rect 43260 31042 43316 31052
rect 43484 30212 43540 31724
rect 43596 31668 43652 32172
rect 43708 32004 43764 33070
rect 43820 32786 43876 33516
rect 43932 33348 43988 33358
rect 44044 33348 44100 34078
rect 44380 34130 44436 34636
rect 44380 34078 44382 34130
rect 44434 34078 44436 34130
rect 44380 34066 44436 34078
rect 44604 34130 44660 34860
rect 44604 34078 44606 34130
rect 44658 34078 44660 34130
rect 44268 34020 44324 34030
rect 44268 33926 44324 33964
rect 43932 33346 44100 33348
rect 43932 33294 43934 33346
rect 43986 33294 44100 33346
rect 43932 33292 44100 33294
rect 43932 33282 43988 33292
rect 44604 33124 44660 34078
rect 44940 33570 44996 35084
rect 44940 33518 44942 33570
rect 44994 33518 44996 33570
rect 44940 33506 44996 33518
rect 44716 33348 44772 33358
rect 44772 33292 44884 33348
rect 44716 33282 44772 33292
rect 44828 33234 44884 33292
rect 44828 33182 44830 33234
rect 44882 33182 44884 33234
rect 44828 33170 44884 33182
rect 44940 33236 44996 33246
rect 44940 33142 44996 33180
rect 44604 33058 44660 33068
rect 43820 32734 43822 32786
rect 43874 32734 43876 32786
rect 43820 32722 43876 32734
rect 44044 32676 44100 32686
rect 44044 32582 44100 32620
rect 44828 32674 44884 32686
rect 44828 32622 44830 32674
rect 44882 32622 44884 32674
rect 44268 32562 44324 32574
rect 44268 32510 44270 32562
rect 44322 32510 44324 32562
rect 44268 32116 44324 32510
rect 44604 32562 44660 32574
rect 44604 32510 44606 32562
rect 44658 32510 44660 32562
rect 44604 32228 44660 32510
rect 44604 32162 44660 32172
rect 44268 32050 44324 32060
rect 43708 31948 44212 32004
rect 44156 31892 44212 31948
rect 44156 31890 44436 31892
rect 44156 31838 44158 31890
rect 44210 31838 44436 31890
rect 44156 31836 44436 31838
rect 44156 31826 44212 31836
rect 43820 31668 43876 31678
rect 43596 31612 43764 31668
rect 43596 31108 43652 31118
rect 43596 30772 43652 31052
rect 43708 31106 43764 31612
rect 43820 31218 43876 31612
rect 44380 31556 44436 31836
rect 44828 31556 44884 32622
rect 44940 32676 44996 32686
rect 44940 32582 44996 32620
rect 44380 31500 44772 31556
rect 44828 31500 44996 31556
rect 44492 31220 44548 31230
rect 43820 31166 43822 31218
rect 43874 31166 43876 31218
rect 43820 31154 43876 31166
rect 44156 31218 44548 31220
rect 44156 31166 44494 31218
rect 44546 31166 44548 31218
rect 44156 31164 44548 31166
rect 43708 31054 43710 31106
rect 43762 31054 43764 31106
rect 43708 31042 43764 31054
rect 44044 31108 44100 31118
rect 44156 31108 44212 31164
rect 44492 31154 44548 31164
rect 44604 31220 44660 31230
rect 44044 31106 44212 31108
rect 44044 31054 44046 31106
rect 44098 31054 44212 31106
rect 44044 31052 44212 31054
rect 44044 31042 44100 31052
rect 44268 30996 44324 31006
rect 44604 30996 44660 31164
rect 44716 31218 44772 31500
rect 44716 31166 44718 31218
rect 44770 31166 44772 31218
rect 44716 31154 44772 31166
rect 44828 31108 44884 31118
rect 44828 31014 44884 31052
rect 44268 30994 44660 30996
rect 44268 30942 44270 30994
rect 44322 30942 44660 30994
rect 44268 30940 44660 30942
rect 44268 30930 44324 30940
rect 43596 30716 43876 30772
rect 43484 30156 43652 30212
rect 43148 30044 43540 30100
rect 42476 29708 42980 29764
rect 43036 29986 43092 29998
rect 43036 29934 43038 29986
rect 43090 29934 43092 29986
rect 43036 29764 43092 29934
rect 42364 29316 42420 29326
rect 42140 29260 42364 29316
rect 42140 28754 42196 29260
rect 42364 29250 42420 29260
rect 42140 28702 42142 28754
rect 42194 28702 42196 28754
rect 42140 28690 42196 28702
rect 42476 28196 42532 29708
rect 43036 29698 43092 29708
rect 42812 29540 42868 29550
rect 42812 29538 43092 29540
rect 42812 29486 42814 29538
rect 42866 29486 43092 29538
rect 42812 29484 43092 29486
rect 42812 29474 42868 29484
rect 42924 29316 42980 29326
rect 42924 29222 42980 29260
rect 42364 28140 42532 28196
rect 42588 28644 42644 28654
rect 42140 27972 42196 27982
rect 42140 27878 42196 27916
rect 42252 27858 42308 27870
rect 42252 27806 42254 27858
rect 42306 27806 42308 27858
rect 42252 27748 42308 27806
rect 42028 27692 42308 27748
rect 41132 26516 41188 27468
rect 42028 26908 42084 27692
rect 42364 27636 42420 28140
rect 41916 26852 42084 26908
rect 42140 27580 42420 27636
rect 42476 27972 42532 27982
rect 41804 26796 41916 26852
rect 41020 26460 41132 26516
rect 41020 26402 41076 26460
rect 41132 26450 41188 26460
rect 41244 26740 41300 26750
rect 41020 26350 41022 26402
rect 41074 26350 41076 26402
rect 41020 26338 41076 26350
rect 41244 26402 41300 26684
rect 41244 26350 41246 26402
rect 41298 26350 41300 26402
rect 41244 26338 41300 26350
rect 41804 26290 41860 26796
rect 41916 26786 41972 26796
rect 41804 26238 41806 26290
rect 41858 26238 41860 26290
rect 41804 26226 41860 26238
rect 41132 26178 41188 26190
rect 41132 26126 41134 26178
rect 41186 26126 41188 26178
rect 41132 25956 41188 26126
rect 41580 26068 41636 26078
rect 41580 26066 41972 26068
rect 41580 26014 41582 26066
rect 41634 26014 41972 26066
rect 41580 26012 41972 26014
rect 41580 26002 41636 26012
rect 41132 25890 41188 25900
rect 41132 25676 41636 25732
rect 41132 25506 41188 25676
rect 41132 25454 41134 25506
rect 41186 25454 41188 25506
rect 41132 25442 41188 25454
rect 41356 25508 41412 25518
rect 41356 24610 41412 25452
rect 41356 24558 41358 24610
rect 41410 24558 41412 24610
rect 41356 24546 41412 24558
rect 41580 25282 41636 25676
rect 41916 25730 41972 26012
rect 41916 25678 41918 25730
rect 41970 25678 41972 25730
rect 41916 25666 41972 25678
rect 41916 25508 41972 25518
rect 41916 25414 41972 25452
rect 41580 25230 41582 25282
rect 41634 25230 41636 25282
rect 41580 24612 41636 25230
rect 40684 24050 40852 24052
rect 40684 23998 40686 24050
rect 40738 23998 40852 24050
rect 40684 23996 40852 23998
rect 40684 23986 40740 23996
rect 41132 23716 41188 23726
rect 41020 23714 41188 23716
rect 41020 23662 41134 23714
rect 41186 23662 41188 23714
rect 41020 23660 41188 23662
rect 40908 23154 40964 23166
rect 40908 23102 40910 23154
rect 40962 23102 40964 23154
rect 40460 23042 40516 23054
rect 40460 22990 40462 23042
rect 40514 22990 40516 23042
rect 40460 22708 40516 22990
rect 40908 23044 40964 23102
rect 40908 22978 40964 22988
rect 40460 22642 40516 22652
rect 40460 22482 40516 22494
rect 40908 22484 40964 22494
rect 41020 22484 41076 23660
rect 41132 23650 41188 23660
rect 41580 23044 41636 24556
rect 41580 22978 41636 22988
rect 41692 23042 41748 23054
rect 41692 22990 41694 23042
rect 41746 22990 41748 23042
rect 40460 22430 40462 22482
rect 40514 22430 40516 22482
rect 40460 22372 40516 22430
rect 39340 20862 39342 20914
rect 39394 20862 39396 20914
rect 39340 20850 39396 20862
rect 39564 21084 40180 21140
rect 40236 22316 40516 22372
rect 40572 22482 41076 22484
rect 40572 22430 40910 22482
rect 40962 22430 41076 22482
rect 40572 22428 41076 22430
rect 39004 20804 39060 20814
rect 39004 20690 39060 20748
rect 39004 20638 39006 20690
rect 39058 20638 39060 20690
rect 39004 20626 39060 20638
rect 39564 20804 39620 21084
rect 39228 20580 39284 20590
rect 39228 20486 39284 20524
rect 39452 20578 39508 20590
rect 39452 20526 39454 20578
rect 39506 20526 39508 20578
rect 39452 20356 39508 20526
rect 39228 20300 39508 20356
rect 38444 20132 38836 20188
rect 38892 20178 38948 20188
rect 39116 20244 39172 20254
rect 39228 20244 39284 20300
rect 39116 20242 39284 20244
rect 39116 20190 39118 20242
rect 39170 20190 39284 20242
rect 39116 20188 39284 20190
rect 39116 20178 39172 20188
rect 38108 20066 38164 20076
rect 38780 20130 38836 20132
rect 38780 20078 38782 20130
rect 38834 20078 38836 20130
rect 38780 20066 38836 20078
rect 38892 19908 38948 19918
rect 37996 18946 38052 18956
rect 38220 19122 38276 19134
rect 38220 19070 38222 19122
rect 38274 19070 38276 19122
rect 38220 18452 38276 19070
rect 38220 18386 38276 18396
rect 38668 19012 38724 19022
rect 37884 17826 37940 17836
rect 37772 17726 37774 17778
rect 37826 17726 37828 17778
rect 37772 17714 37828 17726
rect 37996 17668 38052 17678
rect 37884 17666 38052 17668
rect 37884 17614 37998 17666
rect 38050 17614 38052 17666
rect 37884 17612 38052 17614
rect 37436 16994 37492 17006
rect 37436 16942 37438 16994
rect 37490 16942 37492 16994
rect 37436 15540 37492 16942
rect 37660 16882 37716 16894
rect 37660 16830 37662 16882
rect 37714 16830 37716 16882
rect 37548 16100 37604 16110
rect 37548 16006 37604 16044
rect 37660 15764 37716 16830
rect 37660 15698 37716 15708
rect 37884 16884 37940 17612
rect 37996 17602 38052 17612
rect 38220 17666 38276 17678
rect 38220 17614 38222 17666
rect 38274 17614 38276 17666
rect 38220 16996 38276 17614
rect 38444 17666 38500 17678
rect 38444 17614 38446 17666
rect 38498 17614 38500 17666
rect 38444 17220 38500 17614
rect 38444 17154 38500 17164
rect 38332 16996 38388 17006
rect 38220 16994 38388 16996
rect 38220 16942 38334 16994
rect 38386 16942 38388 16994
rect 38220 16940 38388 16942
rect 37436 15148 37492 15484
rect 37884 15204 37940 16828
rect 37996 16772 38052 16782
rect 37996 16770 38276 16772
rect 37996 16718 37998 16770
rect 38050 16718 38276 16770
rect 37996 16716 38276 16718
rect 37996 16706 38052 16716
rect 38220 15652 38276 16716
rect 38332 16436 38388 16940
rect 38556 16882 38612 16894
rect 38556 16830 38558 16882
rect 38610 16830 38612 16882
rect 38556 16772 38612 16830
rect 38556 16706 38612 16716
rect 38668 16660 38724 18956
rect 38780 18452 38836 18462
rect 38780 17332 38836 18396
rect 38892 18116 38948 19852
rect 39228 19684 39284 20188
rect 39564 20242 39620 20748
rect 39564 20190 39566 20242
rect 39618 20190 39620 20242
rect 39564 20178 39620 20190
rect 40012 20802 40068 20814
rect 40012 20750 40014 20802
rect 40066 20750 40068 20802
rect 39228 19618 39284 19628
rect 39676 20132 39732 20142
rect 39116 19572 39172 19582
rect 39116 19346 39172 19516
rect 39116 19294 39118 19346
rect 39170 19294 39172 19346
rect 39116 19282 39172 19294
rect 39564 19236 39620 19246
rect 39676 19236 39732 20076
rect 40012 19908 40068 20750
rect 40236 20580 40292 22316
rect 40572 22260 40628 22428
rect 40908 22418 40964 22428
rect 41692 22372 41748 22990
rect 41132 22316 41748 22372
rect 40348 22204 40628 22260
rect 41020 22260 41076 22270
rect 40348 21812 40404 22204
rect 40348 21718 40404 21756
rect 40236 20514 40292 20524
rect 40796 21700 40852 21710
rect 40796 21586 40852 21644
rect 40796 21534 40798 21586
rect 40850 21534 40852 21586
rect 40796 20692 40852 21534
rect 41020 21588 41076 22204
rect 41132 21810 41188 22316
rect 41916 22260 41972 22270
rect 41580 22148 41636 22158
rect 41580 22054 41636 22092
rect 41692 22146 41748 22158
rect 41692 22094 41694 22146
rect 41746 22094 41748 22146
rect 41132 21758 41134 21810
rect 41186 21758 41188 21810
rect 41132 21746 41188 21758
rect 41468 21700 41524 21710
rect 41692 21700 41748 22094
rect 41804 22148 41860 22158
rect 41804 22054 41860 22092
rect 41916 21812 41972 22204
rect 42140 22036 42196 27580
rect 42364 27188 42420 27198
rect 42476 27188 42532 27916
rect 42364 27186 42532 27188
rect 42364 27134 42366 27186
rect 42418 27134 42532 27186
rect 42364 27132 42532 27134
rect 42364 27122 42420 27132
rect 42364 26516 42420 26526
rect 42364 26422 42420 26460
rect 42588 26290 42644 28588
rect 42924 28532 42980 28542
rect 42812 27972 42868 27982
rect 42812 27878 42868 27916
rect 42924 27970 42980 28476
rect 42924 27918 42926 27970
rect 42978 27918 42980 27970
rect 42924 27906 42980 27918
rect 42812 27636 42868 27646
rect 43036 27636 43092 29484
rect 43148 29538 43204 30044
rect 43484 29986 43540 30044
rect 43484 29934 43486 29986
rect 43538 29934 43540 29986
rect 43484 29922 43540 29934
rect 43148 29486 43150 29538
rect 43202 29486 43204 29538
rect 43148 29474 43204 29486
rect 43484 29764 43540 29774
rect 43260 29426 43316 29438
rect 43260 29374 43262 29426
rect 43314 29374 43316 29426
rect 43260 28196 43316 29374
rect 43484 28644 43540 29708
rect 43484 28578 43540 28588
rect 43596 28532 43652 30156
rect 43820 30210 43876 30716
rect 44940 30324 44996 31500
rect 43820 30158 43822 30210
rect 43874 30158 43876 30210
rect 43820 30146 43876 30158
rect 43932 30268 44996 30324
rect 43708 29988 43764 29998
rect 43932 29988 43988 30268
rect 43708 29986 43988 29988
rect 43708 29934 43710 29986
rect 43762 29934 43988 29986
rect 43708 29932 43988 29934
rect 44044 30100 44100 30110
rect 43708 29922 43764 29932
rect 43596 28466 43652 28476
rect 42812 27634 43092 27636
rect 42812 27582 42814 27634
rect 42866 27582 43092 27634
rect 42812 27580 43092 27582
rect 43148 28140 43316 28196
rect 42812 27570 42868 27580
rect 42924 26962 42980 26974
rect 42924 26910 42926 26962
rect 42978 26910 42980 26962
rect 42924 26516 42980 26910
rect 42924 26450 42980 26460
rect 43036 26850 43092 26862
rect 43036 26798 43038 26850
rect 43090 26798 43092 26850
rect 42588 26238 42590 26290
rect 42642 26238 42644 26290
rect 42252 25732 42308 25742
rect 42588 25732 42644 26238
rect 42252 25730 42644 25732
rect 42252 25678 42254 25730
rect 42306 25678 42644 25730
rect 42252 25676 42644 25678
rect 42252 25666 42308 25676
rect 43036 25508 43092 26798
rect 43148 26852 43204 28140
rect 43596 27748 43652 27758
rect 43596 27186 43652 27692
rect 43596 27134 43598 27186
rect 43650 27134 43652 27186
rect 43596 27122 43652 27134
rect 43148 26404 43204 26796
rect 43260 26852 43316 26862
rect 43260 26850 43540 26852
rect 43260 26798 43262 26850
rect 43314 26798 43540 26850
rect 43260 26796 43540 26798
rect 43260 26786 43316 26796
rect 43372 26404 43428 26414
rect 43148 26402 43428 26404
rect 43148 26350 43374 26402
rect 43426 26350 43428 26402
rect 43148 26348 43428 26350
rect 43372 26338 43428 26348
rect 43036 25442 43092 25452
rect 43372 25508 43428 25518
rect 43372 25414 43428 25452
rect 43484 25506 43540 26796
rect 43484 25454 43486 25506
rect 43538 25454 43540 25506
rect 43484 25442 43540 25454
rect 43708 26402 43764 26414
rect 43708 26350 43710 26402
rect 43762 26350 43764 26402
rect 43708 25508 43764 26350
rect 43596 25282 43652 25294
rect 43596 25230 43598 25282
rect 43650 25230 43652 25282
rect 43484 24836 43540 24846
rect 43596 24836 43652 25230
rect 43484 24834 43652 24836
rect 43484 24782 43486 24834
rect 43538 24782 43652 24834
rect 43484 24780 43652 24782
rect 43484 24770 43540 24780
rect 43708 23380 43764 25452
rect 43932 25506 43988 25518
rect 43932 25454 43934 25506
rect 43986 25454 43988 25506
rect 43932 24948 43988 25454
rect 43932 24882 43988 24892
rect 43708 23314 43764 23324
rect 43148 23044 43204 23054
rect 43820 23044 43876 23054
rect 43148 22482 43204 22988
rect 43148 22430 43150 22482
rect 43202 22430 43204 22482
rect 43148 22418 43204 22430
rect 43708 23042 43876 23044
rect 43708 22990 43822 23042
rect 43874 22990 43876 23042
rect 43708 22988 43876 22990
rect 42140 21970 42196 21980
rect 42252 22370 42308 22382
rect 42252 22318 42254 22370
rect 42306 22318 42308 22370
rect 41468 21698 41748 21700
rect 41468 21646 41470 21698
rect 41522 21646 41748 21698
rect 41468 21644 41748 21646
rect 41804 21756 41972 21812
rect 41468 21634 41524 21644
rect 41132 21588 41188 21598
rect 41020 21586 41188 21588
rect 41020 21534 41134 21586
rect 41186 21534 41188 21586
rect 41020 21532 41188 21534
rect 40796 20018 40852 20636
rect 41132 20580 41188 21532
rect 40796 19966 40798 20018
rect 40850 19966 40852 20018
rect 40796 19954 40852 19966
rect 40908 20524 41188 20580
rect 41244 20580 41300 20590
rect 40012 19814 40068 19852
rect 40236 19908 40292 19918
rect 40236 19346 40292 19852
rect 40908 19796 40964 20524
rect 41132 20018 41188 20030
rect 41132 19966 41134 20018
rect 41186 19966 41188 20018
rect 41020 19908 41076 19918
rect 41020 19814 41076 19852
rect 40684 19740 40964 19796
rect 41132 19796 41188 19966
rect 40236 19294 40238 19346
rect 40290 19294 40292 19346
rect 40236 19282 40292 19294
rect 40460 19572 40516 19582
rect 39564 19234 39732 19236
rect 39564 19182 39566 19234
rect 39618 19182 39732 19234
rect 39564 19180 39732 19182
rect 39564 19170 39620 19180
rect 40012 18562 40068 18574
rect 40012 18510 40014 18562
rect 40066 18510 40068 18562
rect 40012 18452 40068 18510
rect 40012 18386 40068 18396
rect 40348 18450 40404 18462
rect 40348 18398 40350 18450
rect 40402 18398 40404 18450
rect 39004 18340 39060 18350
rect 39004 18338 39172 18340
rect 39004 18286 39006 18338
rect 39058 18286 39172 18338
rect 39004 18284 39172 18286
rect 39004 18274 39060 18284
rect 38892 18060 39060 18116
rect 38892 17556 38948 17566
rect 38892 17462 38948 17500
rect 38780 17276 38948 17332
rect 38892 16994 38948 17276
rect 38892 16942 38894 16994
rect 38946 16942 38948 16994
rect 38892 16930 38948 16942
rect 38780 16884 38836 16894
rect 38780 16790 38836 16828
rect 38668 16604 38836 16660
rect 38332 16380 38724 16436
rect 38556 15764 38612 15774
rect 38220 15596 38500 15652
rect 38108 15428 38164 15438
rect 37996 15204 38052 15214
rect 37884 15202 38052 15204
rect 37884 15150 37998 15202
rect 38050 15150 38052 15202
rect 37884 15148 38052 15150
rect 37436 15092 37716 15148
rect 37996 15138 38052 15148
rect 36764 13458 36820 13468
rect 36988 14530 37380 14532
rect 36988 14478 37326 14530
rect 37378 14478 37380 14530
rect 36988 14476 37380 14478
rect 36988 13970 37044 14476
rect 37324 14466 37380 14476
rect 37660 14418 37716 15092
rect 38108 14642 38164 15372
rect 38444 15426 38500 15596
rect 38444 15374 38446 15426
rect 38498 15374 38500 15426
rect 38444 15362 38500 15374
rect 38332 15204 38388 15242
rect 38556 15204 38612 15708
rect 38668 15428 38724 16380
rect 38668 15362 38724 15372
rect 38332 15138 38388 15148
rect 38108 14590 38110 14642
rect 38162 14590 38164 14642
rect 38108 14578 38164 14590
rect 38444 15092 38612 15148
rect 37660 14366 37662 14418
rect 37714 14366 37716 14418
rect 37660 14354 37716 14366
rect 36988 13918 36990 13970
rect 37042 13918 37044 13970
rect 36988 11396 37044 13918
rect 37772 13076 37828 13086
rect 36876 11340 37044 11396
rect 37436 12964 37492 12974
rect 37436 12066 37492 12908
rect 37772 12180 37828 13020
rect 38444 12964 38500 15092
rect 38780 13636 38836 16604
rect 39004 16100 39060 18060
rect 39116 17668 39172 18284
rect 39452 18338 39508 18350
rect 39452 18286 39454 18338
rect 39506 18286 39508 18338
rect 39452 18116 39508 18286
rect 39452 18050 39508 18060
rect 40348 18340 40404 18398
rect 40348 17778 40404 18284
rect 40348 17726 40350 17778
rect 40402 17726 40404 17778
rect 40348 17714 40404 17726
rect 39116 17574 39172 17612
rect 39228 17554 39284 17566
rect 39228 17502 39230 17554
rect 39282 17502 39284 17554
rect 39228 16884 39284 17502
rect 39788 16996 39844 17006
rect 39116 16828 39284 16884
rect 39564 16884 39620 16894
rect 39116 16548 39172 16828
rect 39564 16790 39620 16828
rect 39788 16882 39844 16940
rect 39788 16830 39790 16882
rect 39842 16830 39844 16882
rect 39788 16818 39844 16830
rect 40236 16770 40292 16782
rect 40236 16718 40238 16770
rect 40290 16718 40292 16770
rect 39116 16482 39172 16492
rect 39228 16658 39284 16670
rect 39228 16606 39230 16658
rect 39282 16606 39284 16658
rect 39228 16436 39284 16606
rect 39228 16380 39620 16436
rect 39004 16034 39060 16044
rect 39228 16210 39284 16222
rect 39228 16158 39230 16210
rect 39282 16158 39284 16210
rect 39228 15540 39284 16158
rect 39564 16212 39620 16380
rect 39228 15474 39284 15484
rect 39452 15876 39508 15886
rect 38892 15428 38948 15438
rect 38892 15334 38948 15372
rect 39452 15426 39508 15820
rect 39452 15374 39454 15426
rect 39506 15374 39508 15426
rect 39452 15362 39508 15374
rect 39004 15314 39060 15326
rect 39004 15262 39006 15314
rect 39058 15262 39060 15314
rect 38780 13570 38836 13580
rect 38892 14980 38948 14990
rect 37772 12086 37828 12124
rect 38108 12908 38500 12964
rect 38556 13524 38612 13534
rect 38108 12402 38164 12908
rect 38108 12350 38110 12402
rect 38162 12350 38164 12402
rect 37436 12014 37438 12066
rect 37490 12014 37492 12066
rect 36876 10948 36932 11340
rect 37100 11282 37156 11294
rect 37100 11230 37102 11282
rect 37154 11230 37156 11282
rect 36988 11172 37044 11182
rect 36988 11078 37044 11116
rect 36876 10892 37044 10948
rect 36540 9938 36708 9940
rect 36540 9886 36542 9938
rect 36594 9886 36708 9938
rect 36540 9884 36708 9886
rect 36540 9828 36596 9884
rect 36540 9762 36596 9772
rect 36428 8036 36484 8046
rect 36428 7942 36484 7980
rect 36540 7812 36596 7822
rect 36596 7756 36708 7812
rect 36540 7746 36596 7756
rect 36428 7588 36484 7598
rect 36316 7586 36484 7588
rect 36316 7534 36430 7586
rect 36482 7534 36484 7586
rect 36316 7532 36484 7534
rect 36428 7522 36484 7532
rect 36652 7474 36708 7756
rect 36652 7422 36654 7474
rect 36706 7422 36708 7474
rect 36652 7410 36708 7422
rect 36876 7250 36932 7262
rect 36876 7198 36878 7250
rect 36930 7198 36932 7250
rect 36876 6692 36932 7198
rect 36540 6580 36596 6590
rect 36540 6466 36596 6524
rect 36540 6414 36542 6466
rect 36594 6414 36596 6466
rect 36540 6356 36596 6414
rect 36540 6290 36596 6300
rect 36316 6020 36372 6030
rect 36316 5926 36372 5964
rect 36652 5906 36708 5918
rect 36652 5854 36654 5906
rect 36706 5854 36708 5906
rect 36652 5796 36708 5854
rect 36652 5730 36708 5740
rect 36764 5906 36820 5918
rect 36764 5854 36766 5906
rect 36818 5854 36820 5906
rect 36764 5348 36820 5854
rect 36316 5292 36820 5348
rect 36876 5908 36932 6636
rect 36988 6244 37044 10892
rect 37100 10500 37156 11230
rect 37324 10500 37380 10510
rect 37100 10498 37380 10500
rect 37100 10446 37326 10498
rect 37378 10446 37380 10498
rect 37100 10444 37380 10446
rect 37324 10388 37380 10444
rect 37324 10322 37380 10332
rect 37212 10164 37268 10174
rect 37212 9828 37268 10108
rect 37100 9826 37268 9828
rect 37100 9774 37214 9826
rect 37266 9774 37268 9826
rect 37100 9772 37268 9774
rect 37100 8036 37156 9772
rect 37212 9762 37268 9772
rect 37324 9380 37380 9390
rect 37324 9266 37380 9324
rect 37324 9214 37326 9266
rect 37378 9214 37380 9266
rect 37324 9202 37380 9214
rect 37436 8260 37492 12014
rect 38108 11620 38164 12350
rect 38556 12180 38612 13468
rect 38108 11554 38164 11564
rect 38220 12178 38612 12180
rect 38220 12126 38558 12178
rect 38610 12126 38612 12178
rect 38220 12124 38612 12126
rect 37660 11508 37716 11518
rect 37660 11172 37716 11452
rect 37548 11170 37716 11172
rect 37548 11118 37662 11170
rect 37714 11118 37716 11170
rect 37548 11116 37716 11118
rect 37548 10164 37604 11116
rect 37660 11106 37716 11116
rect 38108 11396 38164 11406
rect 38220 11396 38276 12124
rect 38556 12114 38612 12124
rect 38780 12290 38836 12302
rect 38780 12238 38782 12290
rect 38834 12238 38836 12290
rect 38780 11732 38836 12238
rect 38780 11666 38836 11676
rect 38108 11394 38276 11396
rect 38108 11342 38110 11394
rect 38162 11342 38276 11394
rect 38108 11340 38276 11342
rect 38780 11508 38836 11518
rect 37996 10836 38052 10846
rect 38108 10836 38164 11340
rect 38556 11284 38612 11294
rect 38556 11190 38612 11228
rect 38668 11170 38724 11182
rect 38668 11118 38670 11170
rect 38722 11118 38724 11170
rect 38444 10836 38500 10846
rect 37996 10834 38500 10836
rect 37996 10782 37998 10834
rect 38050 10782 38446 10834
rect 38498 10782 38500 10834
rect 37996 10780 38500 10782
rect 37996 10770 38052 10780
rect 38444 10770 38500 10780
rect 37660 10724 37716 10734
rect 37660 10630 37716 10668
rect 38668 10276 38724 11118
rect 38780 10836 38836 11452
rect 38892 11396 38948 14924
rect 39004 13860 39060 15262
rect 39116 15314 39172 15326
rect 39116 15262 39118 15314
rect 39170 15262 39172 15314
rect 39116 15204 39172 15262
rect 39564 15316 39620 16156
rect 39900 16100 39956 16110
rect 40236 16100 40292 16718
rect 39956 16044 40292 16100
rect 39900 16006 39956 16044
rect 39788 15652 39844 15662
rect 39676 15316 39732 15326
rect 39564 15314 39732 15316
rect 39564 15262 39678 15314
rect 39730 15262 39732 15314
rect 39564 15260 39732 15262
rect 39676 15250 39732 15260
rect 39788 15314 39844 15596
rect 40236 15540 40292 15550
rect 40236 15446 40292 15484
rect 39788 15262 39790 15314
rect 39842 15262 39844 15314
rect 39788 15250 39844 15262
rect 40460 15148 40516 19516
rect 39116 15138 39172 15148
rect 40348 15092 40516 15148
rect 40684 15148 40740 19740
rect 41132 19730 41188 19740
rect 41244 18562 41300 20524
rect 41804 20130 41860 21756
rect 41916 21586 41972 21598
rect 41916 21534 41918 21586
rect 41970 21534 41972 21586
rect 41916 20914 41972 21534
rect 41916 20862 41918 20914
rect 41970 20862 41972 20914
rect 41916 20188 41972 20862
rect 41916 20132 42196 20188
rect 41804 20078 41806 20130
rect 41858 20078 41860 20130
rect 41356 20020 41412 20030
rect 41356 19926 41412 19964
rect 41804 19684 41860 20078
rect 42140 20066 42196 20076
rect 42252 20130 42308 22318
rect 42476 22260 42532 22270
rect 42476 22166 42532 22204
rect 43596 22258 43652 22270
rect 43596 22206 43598 22258
rect 43650 22206 43652 22258
rect 42588 22146 42644 22158
rect 42588 22094 42590 22146
rect 42642 22094 42644 22146
rect 42588 22036 42644 22094
rect 42812 22148 42868 22158
rect 43484 22148 43540 22158
rect 42812 22146 43092 22148
rect 42812 22094 42814 22146
rect 42866 22094 43092 22146
rect 42812 22092 43092 22094
rect 42812 22082 42868 22092
rect 42588 21700 42644 21980
rect 42252 20078 42254 20130
rect 42306 20078 42308 20130
rect 41916 20020 41972 20030
rect 41916 19926 41972 19964
rect 42028 20018 42084 20030
rect 42028 19966 42030 20018
rect 42082 19966 42084 20018
rect 41804 19618 41860 19628
rect 42028 19348 42084 19966
rect 42252 19572 42308 20078
rect 42476 21644 42644 21700
rect 42252 19506 42308 19516
rect 42364 19906 42420 19918
rect 42364 19854 42366 19906
rect 42418 19854 42420 19906
rect 42364 19348 42420 19854
rect 42028 19346 42420 19348
rect 42028 19294 42366 19346
rect 42418 19294 42420 19346
rect 42028 19292 42420 19294
rect 42364 19282 42420 19292
rect 42476 19124 42532 21644
rect 42588 21474 42644 21486
rect 42588 21422 42590 21474
rect 42642 21422 42644 21474
rect 42588 20916 42644 21422
rect 42812 20916 42868 20926
rect 42588 20914 42868 20916
rect 42588 20862 42814 20914
rect 42866 20862 42868 20914
rect 42588 20860 42868 20862
rect 42812 20850 42868 20860
rect 42700 20692 42756 20702
rect 42700 20598 42756 20636
rect 43036 20690 43092 22092
rect 43260 22146 43540 22148
rect 43260 22094 43486 22146
rect 43538 22094 43540 22146
rect 43260 22092 43540 22094
rect 43036 20638 43038 20690
rect 43090 20638 43092 20690
rect 43036 20626 43092 20638
rect 43148 20692 43204 20702
rect 43148 20598 43204 20636
rect 42924 20578 42980 20590
rect 42924 20526 42926 20578
rect 42978 20526 42980 20578
rect 42924 20468 42980 20526
rect 43260 20468 43316 22092
rect 43484 22082 43540 22092
rect 43596 21476 43652 22206
rect 43596 21410 43652 21420
rect 43708 22148 43764 22988
rect 43820 22978 43876 22988
rect 43708 21252 43764 22092
rect 42924 20412 43316 20468
rect 43596 21196 43764 21252
rect 43260 20132 43316 20142
rect 43260 20038 43316 20076
rect 42812 19906 42868 19918
rect 42812 19854 42814 19906
rect 42866 19854 42868 19906
rect 42812 19796 42868 19854
rect 42812 19730 42868 19740
rect 43260 19794 43316 19806
rect 43260 19742 43262 19794
rect 43314 19742 43316 19794
rect 42364 19068 42532 19124
rect 42140 19012 42196 19022
rect 41804 18788 41860 18798
rect 41860 18732 41972 18788
rect 41804 18722 41860 18732
rect 41244 18510 41246 18562
rect 41298 18510 41300 18562
rect 41244 18498 41300 18510
rect 40908 18452 40964 18462
rect 40908 18358 40964 18396
rect 41468 18450 41524 18462
rect 41468 18398 41470 18450
rect 41522 18398 41524 18450
rect 41020 18338 41076 18350
rect 41020 18286 41022 18338
rect 41074 18286 41076 18338
rect 41020 17332 41076 18286
rect 41020 17266 41076 17276
rect 41356 17220 41412 17230
rect 41132 16996 41188 17006
rect 41132 16902 41188 16940
rect 40908 16884 40964 16894
rect 40908 16790 40964 16828
rect 41020 16770 41076 16782
rect 41020 16718 41022 16770
rect 41074 16718 41076 16770
rect 41020 15652 41076 16718
rect 41020 15586 41076 15596
rect 41356 15540 41412 17164
rect 41468 16660 41524 18398
rect 41692 18452 41748 18462
rect 41468 16594 41524 16604
rect 41580 16882 41636 16894
rect 41580 16830 41582 16882
rect 41634 16830 41636 16882
rect 41580 16436 41636 16830
rect 41692 16882 41748 18396
rect 41916 17780 41972 18732
rect 42140 18450 42196 18956
rect 42140 18398 42142 18450
rect 42194 18398 42196 18450
rect 41916 17724 42084 17780
rect 41804 17556 41860 17566
rect 41804 17462 41860 17500
rect 41692 16830 41694 16882
rect 41746 16830 41748 16882
rect 41692 16818 41748 16830
rect 42028 16882 42084 17724
rect 42028 16830 42030 16882
rect 42082 16830 42084 16882
rect 42028 16818 42084 16830
rect 41916 16770 41972 16782
rect 41916 16718 41918 16770
rect 41970 16718 41972 16770
rect 41580 16370 41636 16380
rect 41692 16548 41748 16558
rect 41580 15540 41636 15578
rect 41356 15484 41524 15540
rect 41468 15426 41524 15484
rect 41580 15474 41636 15484
rect 41468 15374 41470 15426
rect 41522 15374 41524 15426
rect 41468 15316 41524 15374
rect 41356 15260 41524 15316
rect 41692 15426 41748 16492
rect 41692 15374 41694 15426
rect 41746 15374 41748 15426
rect 41020 15204 41076 15214
rect 40684 15092 40964 15148
rect 40236 14420 40292 14430
rect 39228 14418 40292 14420
rect 39228 14366 40238 14418
rect 40290 14366 40292 14418
rect 39228 14364 40292 14366
rect 39228 13970 39284 14364
rect 40236 14354 40292 14364
rect 39228 13918 39230 13970
rect 39282 13918 39284 13970
rect 39228 13906 39284 13918
rect 39340 14196 39396 14206
rect 40348 14196 40404 15092
rect 39116 13860 39172 13870
rect 39004 13858 39172 13860
rect 39004 13806 39118 13858
rect 39170 13806 39172 13858
rect 39004 13804 39172 13806
rect 39116 13794 39172 13804
rect 39340 12404 39396 14140
rect 40236 14140 40404 14196
rect 39788 12404 39844 12414
rect 39340 12402 39844 12404
rect 39340 12350 39790 12402
rect 39842 12350 39844 12402
rect 39340 12348 39844 12350
rect 39116 12290 39172 12302
rect 39116 12238 39118 12290
rect 39170 12238 39172 12290
rect 39116 11620 39172 12238
rect 39340 12178 39396 12348
rect 39788 12338 39844 12348
rect 40124 12292 40180 12302
rect 39340 12126 39342 12178
rect 39394 12126 39396 12178
rect 39340 12114 39396 12126
rect 40012 12290 40180 12292
rect 40012 12238 40126 12290
rect 40178 12238 40180 12290
rect 40012 12236 40180 12238
rect 39116 11554 39172 11564
rect 39116 11396 39172 11406
rect 39900 11396 39956 11406
rect 38948 11340 39060 11396
rect 38892 11302 38948 11340
rect 39004 11172 39060 11340
rect 39116 11394 39956 11396
rect 39116 11342 39118 11394
rect 39170 11342 39902 11394
rect 39954 11342 39956 11394
rect 39116 11340 39956 11342
rect 39116 11330 39172 11340
rect 39900 11330 39956 11340
rect 40012 11396 40068 12236
rect 40124 12226 40180 12236
rect 40012 11302 40068 11340
rect 40236 11732 40292 14140
rect 40908 12404 40964 15092
rect 41020 14530 41076 15148
rect 41356 14642 41412 15260
rect 41356 14590 41358 14642
rect 41410 14590 41412 14642
rect 41356 14578 41412 14590
rect 41020 14478 41022 14530
rect 41074 14478 41076 14530
rect 41020 14466 41076 14478
rect 41468 13972 41524 13982
rect 41692 13972 41748 15374
rect 41468 13970 41748 13972
rect 41468 13918 41470 13970
rect 41522 13918 41748 13970
rect 41468 13916 41748 13918
rect 41804 16210 41860 16222
rect 41804 16158 41806 16210
rect 41858 16158 41860 16210
rect 41804 15204 41860 16158
rect 41916 15428 41972 16718
rect 42140 16100 42196 18398
rect 42364 18340 42420 19068
rect 42700 19012 42756 19022
rect 42924 19012 42980 19022
rect 42756 19010 42980 19012
rect 42756 18958 42926 19010
rect 42978 18958 42980 19010
rect 42756 18956 42980 18958
rect 42700 18946 42756 18956
rect 42924 18946 42980 18956
rect 42476 18564 42532 18574
rect 42476 18470 42532 18508
rect 42700 18452 42756 18462
rect 42924 18452 42980 18462
rect 42700 18450 42868 18452
rect 42700 18398 42702 18450
rect 42754 18398 42868 18450
rect 42700 18396 42868 18398
rect 42700 18386 42756 18396
rect 42588 18340 42644 18350
rect 42364 18284 42532 18340
rect 42252 17220 42308 17230
rect 42308 17164 42420 17220
rect 42252 17154 42308 17164
rect 42140 16034 42196 16044
rect 42252 16996 42308 17006
rect 41916 15362 41972 15372
rect 42028 15876 42084 15886
rect 42028 15426 42084 15820
rect 42028 15374 42030 15426
rect 42082 15374 42084 15426
rect 42028 15362 42084 15374
rect 42252 15316 42308 16940
rect 42364 16994 42420 17164
rect 42364 16942 42366 16994
rect 42418 16942 42420 16994
rect 42364 16930 42420 16942
rect 42252 15222 42308 15260
rect 42364 15988 42420 15998
rect 42364 15314 42420 15932
rect 42364 15262 42366 15314
rect 42418 15262 42420 15314
rect 42364 15250 42420 15262
rect 41916 15204 41972 15214
rect 41804 15148 41916 15204
rect 42476 15148 42532 18284
rect 42588 18246 42644 18284
rect 42812 18228 42868 18396
rect 42924 18358 42980 18396
rect 43260 18450 43316 19742
rect 43596 19234 43652 21196
rect 43932 20692 43988 20702
rect 43932 20598 43988 20636
rect 44044 20356 44100 30044
rect 44268 28754 44324 30268
rect 44828 29426 44884 29438
rect 44828 29374 44830 29426
rect 44882 29374 44884 29426
rect 44268 28702 44270 28754
rect 44322 28702 44324 28754
rect 44268 28690 44324 28702
rect 44492 29316 44548 29326
rect 44828 29316 44884 29374
rect 44492 29314 44996 29316
rect 44492 29262 44494 29314
rect 44546 29262 44996 29314
rect 44492 29260 44996 29262
rect 44268 27748 44324 27758
rect 44492 27748 44548 29260
rect 44940 28754 44996 29260
rect 44940 28702 44942 28754
rect 44994 28702 44996 28754
rect 44940 28690 44996 28702
rect 44604 28532 44660 28542
rect 44604 28084 44660 28476
rect 44604 28082 44884 28084
rect 44604 28030 44606 28082
rect 44658 28030 44884 28082
rect 44604 28028 44884 28030
rect 44604 28018 44660 28028
rect 44324 27692 44548 27748
rect 44268 24722 44324 27692
rect 44828 27074 44884 28028
rect 44828 27022 44830 27074
rect 44882 27022 44884 27074
rect 44828 27010 44884 27022
rect 44940 27970 44996 27982
rect 44940 27918 44942 27970
rect 44994 27918 44996 27970
rect 44940 27076 44996 27918
rect 44940 27010 44996 27020
rect 45052 26180 45108 38612
rect 45276 38276 45332 39342
rect 45276 38210 45332 38220
rect 45388 39058 45444 39070
rect 45388 39006 45390 39058
rect 45442 39006 45444 39058
rect 45388 37940 45444 39006
rect 45500 38946 45556 39452
rect 45500 38894 45502 38946
rect 45554 38894 45556 38946
rect 45500 38882 45556 38894
rect 45948 38836 46004 39564
rect 46172 39564 46340 39620
rect 46620 39676 46732 39732
rect 45948 38742 46004 38780
rect 46060 39394 46116 39406
rect 46060 39342 46062 39394
rect 46114 39342 46116 39394
rect 46060 38050 46116 39342
rect 46060 37998 46062 38050
rect 46114 37998 46116 38050
rect 46060 37986 46116 37998
rect 46172 38052 46228 39564
rect 46396 39508 46452 39518
rect 46396 39506 46564 39508
rect 46396 39454 46398 39506
rect 46450 39454 46564 39506
rect 46396 39452 46564 39454
rect 46396 39442 46452 39452
rect 46172 37986 46228 37996
rect 46284 39394 46340 39406
rect 46284 39342 46286 39394
rect 46338 39342 46340 39394
rect 45388 37846 45444 37884
rect 46060 37828 46116 37838
rect 45836 37826 46116 37828
rect 45836 37774 46062 37826
rect 46114 37774 46116 37826
rect 45836 37772 46116 37774
rect 45724 36258 45780 36270
rect 45724 36206 45726 36258
rect 45778 36206 45780 36258
rect 45500 35588 45556 35598
rect 45500 35586 45668 35588
rect 45500 35534 45502 35586
rect 45554 35534 45668 35586
rect 45500 35532 45668 35534
rect 45500 35522 45556 35532
rect 45388 35252 45444 35262
rect 45388 34914 45444 35196
rect 45388 34862 45390 34914
rect 45442 34862 45444 34914
rect 45388 34132 45444 34862
rect 45388 34130 45556 34132
rect 45388 34078 45390 34130
rect 45442 34078 45556 34130
rect 45388 34076 45556 34078
rect 45388 34066 45444 34076
rect 45388 33236 45444 33246
rect 45276 33124 45332 33134
rect 45164 33068 45276 33124
rect 45164 31220 45220 33068
rect 45276 33058 45332 33068
rect 45388 32786 45444 33180
rect 45388 32734 45390 32786
rect 45442 32734 45444 32786
rect 45388 32722 45444 32734
rect 45276 32676 45332 32686
rect 45276 32582 45332 32620
rect 45388 31780 45444 31790
rect 45500 31780 45556 34076
rect 45612 33236 45668 35532
rect 45724 35476 45780 36206
rect 45724 35410 45780 35420
rect 45612 33170 45668 33180
rect 45724 33346 45780 33358
rect 45724 33294 45726 33346
rect 45778 33294 45780 33346
rect 45612 32788 45668 32798
rect 45724 32788 45780 33294
rect 45612 32786 45780 32788
rect 45612 32734 45614 32786
rect 45666 32734 45780 32786
rect 45612 32732 45780 32734
rect 45612 32722 45668 32732
rect 45388 31778 45556 31780
rect 45388 31726 45390 31778
rect 45442 31726 45556 31778
rect 45388 31724 45556 31726
rect 45388 31714 45444 31724
rect 45276 31220 45332 31230
rect 45220 31218 45332 31220
rect 45220 31166 45278 31218
rect 45330 31166 45332 31218
rect 45220 31164 45332 31166
rect 45164 31126 45220 31164
rect 45276 31154 45332 31164
rect 45500 30996 45556 31006
rect 45388 30994 45556 30996
rect 45388 30942 45502 30994
rect 45554 30942 45556 30994
rect 45388 30940 45556 30942
rect 45388 30212 45444 30940
rect 45500 30930 45556 30940
rect 45388 29988 45444 30156
rect 45388 29922 45444 29932
rect 45612 29988 45668 29998
rect 45612 29538 45668 29932
rect 45612 29486 45614 29538
rect 45666 29486 45668 29538
rect 45612 29474 45668 29486
rect 45724 29764 45780 29774
rect 45724 28642 45780 29708
rect 45724 28590 45726 28642
rect 45778 28590 45780 28642
rect 45276 27748 45332 27758
rect 45276 27654 45332 27692
rect 45724 26908 45780 28590
rect 45052 26114 45108 26124
rect 45164 26850 45220 26862
rect 45164 26798 45166 26850
rect 45218 26798 45220 26850
rect 44940 25282 44996 25294
rect 44940 25230 44942 25282
rect 44994 25230 44996 25282
rect 44940 25172 44996 25230
rect 45052 25172 45108 25182
rect 44940 25116 45052 25172
rect 45052 25106 45108 25116
rect 44828 24948 44884 24958
rect 44828 24854 44884 24892
rect 45164 24948 45220 26798
rect 45612 26852 45780 26908
rect 45612 26514 45668 26852
rect 45612 26462 45614 26514
rect 45666 26462 45668 26514
rect 45612 26450 45668 26462
rect 45052 24836 45108 24846
rect 44268 24670 44270 24722
rect 44322 24670 44324 24722
rect 44268 23714 44324 24670
rect 44268 23662 44270 23714
rect 44322 23662 44324 23714
rect 44268 23044 44324 23662
rect 44604 24724 44660 24734
rect 44604 23266 44660 24668
rect 44828 24052 44884 24062
rect 45052 24052 45108 24780
rect 45164 24834 45220 24892
rect 45164 24782 45166 24834
rect 45218 24782 45220 24834
rect 45164 24770 45220 24782
rect 45276 26402 45332 26414
rect 45276 26350 45278 26402
rect 45330 26350 45332 26402
rect 45276 24724 45332 26350
rect 45276 24658 45332 24668
rect 45388 25506 45444 25518
rect 45388 25454 45390 25506
rect 45442 25454 45444 25506
rect 45388 25172 45444 25454
rect 45388 24612 45444 25116
rect 45612 24836 45668 24846
rect 45612 24742 45668 24780
rect 45724 24724 45780 24734
rect 45724 24630 45780 24668
rect 45388 24546 45444 24556
rect 45612 24500 45668 24510
rect 45836 24500 45892 37772
rect 46060 37762 46116 37772
rect 46284 37380 46340 39342
rect 46284 37314 46340 37324
rect 46508 37268 46564 39452
rect 46508 37202 46564 37212
rect 46620 36372 46676 39676
rect 46732 39666 46788 39676
rect 46844 39900 47124 39956
rect 47180 39956 47236 41694
rect 46732 39508 46788 39518
rect 46844 39508 46900 39900
rect 47180 39890 47236 39900
rect 47292 41746 47460 41748
rect 47292 41694 47406 41746
rect 47458 41694 47460 41746
rect 47292 41692 47460 41694
rect 47068 39732 47124 39742
rect 47068 39618 47124 39676
rect 47180 39732 47236 39742
rect 47292 39732 47348 41692
rect 47404 41682 47460 41692
rect 47516 41746 47572 41758
rect 47516 41694 47518 41746
rect 47570 41694 47572 41746
rect 47516 40626 47572 41694
rect 47516 40574 47518 40626
rect 47570 40574 47572 40626
rect 47516 40516 47572 40574
rect 47516 40450 47572 40460
rect 47964 40516 48020 41916
rect 48076 41878 48132 41916
rect 48188 41300 48244 41310
rect 47964 40450 48020 40460
rect 48076 41298 48244 41300
rect 48076 41246 48190 41298
rect 48242 41246 48244 41298
rect 48076 41244 48244 41246
rect 47852 40290 47908 40302
rect 47852 40238 47854 40290
rect 47906 40238 47908 40290
rect 47180 39730 47348 39732
rect 47180 39678 47182 39730
rect 47234 39678 47348 39730
rect 47180 39676 47348 39678
rect 47404 40180 47460 40190
rect 47180 39666 47236 39676
rect 47068 39566 47070 39618
rect 47122 39566 47124 39618
rect 47068 39554 47124 39566
rect 47404 39618 47460 40124
rect 47404 39566 47406 39618
rect 47458 39566 47460 39618
rect 46788 39452 46900 39508
rect 46732 39414 46788 39452
rect 46732 38836 46788 38846
rect 46732 37154 46788 38780
rect 47404 38836 47460 39566
rect 47628 39620 47684 39630
rect 47628 39526 47684 39564
rect 47404 38770 47460 38780
rect 47516 38946 47572 38958
rect 47516 38894 47518 38946
rect 47570 38894 47572 38946
rect 46732 37102 46734 37154
rect 46786 37102 46788 37154
rect 46732 37090 46788 37102
rect 46844 38052 46900 38062
rect 46844 37044 46900 37996
rect 47292 37940 47348 37950
rect 47180 37380 47236 37390
rect 47180 37286 47236 37324
rect 46844 36978 46900 36988
rect 47068 37268 47124 37278
rect 46284 36370 46676 36372
rect 46284 36318 46622 36370
rect 46674 36318 46676 36370
rect 46284 36316 46676 36318
rect 46284 35698 46340 36316
rect 46620 36306 46676 36316
rect 46956 36260 47012 36270
rect 46956 36166 47012 36204
rect 46284 35646 46286 35698
rect 46338 35646 46340 35698
rect 46284 35634 46340 35646
rect 46060 35586 46116 35598
rect 46060 35534 46062 35586
rect 46114 35534 46116 35586
rect 45948 35476 46004 35486
rect 45948 35382 46004 35420
rect 46060 35026 46116 35534
rect 47068 35588 47124 37212
rect 47180 37156 47236 37166
rect 47180 37062 47236 37100
rect 47292 36482 47348 37884
rect 47292 36430 47294 36482
rect 47346 36430 47348 36482
rect 47292 36418 47348 36430
rect 47516 36260 47572 38894
rect 47852 38668 47908 40238
rect 47964 40068 48020 40078
rect 48076 40068 48132 41244
rect 48188 41234 48244 41244
rect 48188 40516 48244 40526
rect 48188 40422 48244 40460
rect 48020 40012 48132 40068
rect 47964 40002 48020 40012
rect 48188 39396 48244 39406
rect 48300 39396 48356 42478
rect 48412 42532 48468 56252
rect 48412 42466 48468 42476
rect 48188 39394 48356 39396
rect 48188 39342 48190 39394
rect 48242 39342 48356 39394
rect 48188 39340 48356 39342
rect 48076 38836 48132 38846
rect 48076 38742 48132 38780
rect 47516 36194 47572 36204
rect 47628 38612 47908 38668
rect 48188 38724 48244 39340
rect 48188 38658 48244 38668
rect 47628 38050 47684 38612
rect 47628 37998 47630 38050
rect 47682 37998 47684 38050
rect 47628 36482 47684 37998
rect 47964 37268 48020 37278
rect 47740 37266 48020 37268
rect 47740 37214 47966 37266
rect 48018 37214 48020 37266
rect 47740 37212 48020 37214
rect 47740 36594 47796 37212
rect 47964 37202 48020 37212
rect 47740 36542 47742 36594
rect 47794 36542 47796 36594
rect 47740 36530 47796 36542
rect 47852 37044 47908 37054
rect 47628 36430 47630 36482
rect 47682 36430 47684 36482
rect 47628 36036 47684 36430
rect 47404 35980 47684 36036
rect 47852 36482 47908 36988
rect 47852 36430 47854 36482
rect 47906 36430 47908 36482
rect 47404 35922 47460 35980
rect 47404 35870 47406 35922
rect 47458 35870 47460 35922
rect 47404 35858 47460 35870
rect 47628 35812 47684 35822
rect 47852 35812 47908 36430
rect 47628 35810 47908 35812
rect 47628 35758 47630 35810
rect 47682 35758 47908 35810
rect 47628 35756 47908 35758
rect 48188 36260 48244 36270
rect 47628 35746 47684 35756
rect 47292 35588 47348 35598
rect 47068 35586 47348 35588
rect 47068 35534 47294 35586
rect 47346 35534 47348 35586
rect 47068 35532 47348 35534
rect 47292 35522 47348 35532
rect 46060 34974 46062 35026
rect 46114 34974 46116 35026
rect 46060 34962 46116 34974
rect 48188 35026 48244 36204
rect 48188 34974 48190 35026
rect 48242 34974 48244 35026
rect 48188 34962 48244 34974
rect 46060 34018 46116 34030
rect 46060 33966 46062 34018
rect 46114 33966 46116 34018
rect 46060 33122 46116 33966
rect 46844 34020 46900 34030
rect 46172 33404 46564 33460
rect 46172 33346 46228 33404
rect 46172 33294 46174 33346
rect 46226 33294 46228 33346
rect 46172 33282 46228 33294
rect 46508 33348 46564 33404
rect 46620 33348 46676 33358
rect 46508 33346 46676 33348
rect 46508 33294 46622 33346
rect 46674 33294 46676 33346
rect 46508 33292 46676 33294
rect 46620 33282 46676 33292
rect 46396 33234 46452 33246
rect 46396 33182 46398 33234
rect 46450 33182 46452 33234
rect 46060 33070 46062 33122
rect 46114 33070 46116 33122
rect 46060 33058 46116 33070
rect 46284 33124 46340 33134
rect 46396 33124 46452 33182
rect 46340 33068 46452 33124
rect 46844 33234 46900 33964
rect 48188 34020 48244 34030
rect 48188 33926 48244 33964
rect 46844 33182 46846 33234
rect 46898 33182 46900 33234
rect 46284 33058 46340 33068
rect 46844 32788 46900 33182
rect 46956 33236 47012 33246
rect 46956 33234 47460 33236
rect 46956 33182 46958 33234
rect 47010 33182 47460 33234
rect 46956 33180 47460 33182
rect 46956 33170 47012 33180
rect 46956 32788 47012 32798
rect 46844 32786 47012 32788
rect 46844 32734 46958 32786
rect 47010 32734 47012 32786
rect 46844 32732 47012 32734
rect 46956 32722 47012 32732
rect 46396 32676 46452 32686
rect 46284 32620 46396 32676
rect 46060 31668 46116 31678
rect 46060 31574 46116 31612
rect 46060 30994 46116 31006
rect 46060 30942 46062 30994
rect 46114 30942 46116 30994
rect 46060 30212 46116 30942
rect 46060 30146 46116 30156
rect 46284 28644 46340 32620
rect 46396 32610 46452 32620
rect 47404 32676 47460 33180
rect 47628 33122 47684 33134
rect 47628 33070 47630 33122
rect 47682 33070 47684 33122
rect 47628 32788 47684 33070
rect 47852 33122 47908 33134
rect 47852 33070 47854 33122
rect 47906 33070 47908 33122
rect 47852 32900 47908 33070
rect 47852 32834 47908 32844
rect 48188 33122 48244 33134
rect 48188 33070 48190 33122
rect 48242 33070 48244 33122
rect 47628 32722 47684 32732
rect 48188 32788 48244 33070
rect 48188 32722 48244 32732
rect 47404 32582 47460 32620
rect 47516 32674 47572 32686
rect 47516 32622 47518 32674
rect 47570 32622 47572 32674
rect 46732 32562 46788 32574
rect 46732 32510 46734 32562
rect 46786 32510 46788 32562
rect 46396 31106 46452 31118
rect 46396 31054 46398 31106
rect 46450 31054 46452 31106
rect 46396 30884 46452 31054
rect 46732 30994 46788 32510
rect 47068 32562 47124 32574
rect 47068 32510 47070 32562
rect 47122 32510 47124 32562
rect 46844 31668 46900 31678
rect 46900 31612 47012 31668
rect 46844 31602 46900 31612
rect 46956 31218 47012 31612
rect 46956 31166 46958 31218
rect 47010 31166 47012 31218
rect 46956 31154 47012 31166
rect 46732 30942 46734 30994
rect 46786 30942 46788 30994
rect 46732 30930 46788 30942
rect 47068 30996 47124 32510
rect 47516 32564 47572 32622
rect 47516 32508 48244 32564
rect 47516 32340 47572 32350
rect 47516 32338 47684 32340
rect 47516 32286 47518 32338
rect 47570 32286 47684 32338
rect 47516 32284 47684 32286
rect 47516 32274 47572 32284
rect 47180 31108 47236 31118
rect 47180 31014 47236 31052
rect 47628 31108 47684 32284
rect 47852 31218 47908 32508
rect 48188 31890 48244 32508
rect 48188 31838 48190 31890
rect 48242 31838 48244 31890
rect 48188 31826 48244 31838
rect 47852 31166 47854 31218
rect 47906 31166 47908 31218
rect 47852 31154 47908 31166
rect 47628 31042 47684 31052
rect 47068 30930 47124 30940
rect 47292 30994 47348 31006
rect 47292 30942 47294 30994
rect 47346 30942 47348 30994
rect 46396 30100 46452 30828
rect 47292 30884 47348 30942
rect 47740 30996 47796 31006
rect 47796 30940 48020 30996
rect 47740 30902 47796 30940
rect 47292 30818 47348 30828
rect 47852 30772 47908 30782
rect 47404 30770 47908 30772
rect 47404 30718 47854 30770
rect 47906 30718 47908 30770
rect 47404 30716 47908 30718
rect 47068 30210 47124 30222
rect 47068 30158 47070 30210
rect 47122 30158 47124 30210
rect 46732 30100 46788 30110
rect 46396 30098 46788 30100
rect 46396 30046 46734 30098
rect 46786 30046 46788 30098
rect 46396 30044 46788 30046
rect 46396 28644 46452 28654
rect 45948 28642 46452 28644
rect 45948 28590 46398 28642
rect 46450 28590 46452 28642
rect 45948 28588 46452 28590
rect 45948 28530 46004 28588
rect 45948 28478 45950 28530
rect 46002 28478 46004 28530
rect 45948 28466 46004 28478
rect 46396 28420 46452 28588
rect 46396 28354 46452 28364
rect 46508 28418 46564 28430
rect 46508 28366 46510 28418
rect 46562 28366 46564 28418
rect 46508 27748 46564 28366
rect 46620 28196 46676 30044
rect 46732 30034 46788 30044
rect 47068 28866 47124 30158
rect 47404 30210 47460 30716
rect 47852 30706 47908 30716
rect 47404 30158 47406 30210
rect 47458 30158 47460 30210
rect 47404 30146 47460 30158
rect 47180 29988 47236 29998
rect 47180 29894 47236 29932
rect 47740 29316 47796 29326
rect 47068 28814 47070 28866
rect 47122 28814 47124 28866
rect 47068 28802 47124 28814
rect 47628 29314 47796 29316
rect 47628 29262 47742 29314
rect 47794 29262 47796 29314
rect 47628 29260 47796 29262
rect 47628 28756 47684 29260
rect 47740 29250 47796 29260
rect 47180 28700 47684 28756
rect 47180 28644 47236 28700
rect 47068 28588 47236 28644
rect 47068 28530 47124 28588
rect 47068 28478 47070 28530
rect 47122 28478 47124 28530
rect 47628 28530 47684 28700
rect 47068 28466 47124 28478
rect 47180 28474 47236 28486
rect 46732 28420 46788 28430
rect 47180 28422 47182 28474
rect 47234 28422 47236 28474
rect 47628 28478 47630 28530
rect 47682 28478 47684 28530
rect 47628 28466 47684 28478
rect 47740 28532 47796 28542
rect 47964 28532 48020 30940
rect 47740 28530 48020 28532
rect 47740 28478 47742 28530
rect 47794 28478 48020 28530
rect 47740 28476 48020 28478
rect 47180 28420 47236 28422
rect 46732 28418 47012 28420
rect 46732 28366 46734 28418
rect 46786 28366 47012 28418
rect 46732 28364 47012 28366
rect 46732 28354 46788 28364
rect 46620 28140 46788 28196
rect 46284 27076 46340 27086
rect 46284 26982 46340 27020
rect 44828 24050 45108 24052
rect 44828 23998 44830 24050
rect 44882 23998 45108 24050
rect 44828 23996 45108 23998
rect 45500 24498 45668 24500
rect 45500 24446 45614 24498
rect 45666 24446 45668 24498
rect 45500 24444 45668 24446
rect 44828 23986 44884 23996
rect 44940 23492 44996 23502
rect 44940 23378 44996 23436
rect 44940 23326 44942 23378
rect 44994 23326 44996 23378
rect 44940 23314 44996 23326
rect 45164 23380 45220 23390
rect 44604 23214 44606 23266
rect 44658 23214 44660 23266
rect 44604 23202 44660 23214
rect 44716 23268 44772 23278
rect 44268 22950 44324 22988
rect 44716 22594 44772 23212
rect 45164 23266 45220 23324
rect 45164 23214 45166 23266
rect 45218 23214 45220 23266
rect 45164 23202 45220 23214
rect 45500 23154 45556 24444
rect 45612 24434 45668 24444
rect 45724 24444 45892 24500
rect 45948 26964 46004 26974
rect 45612 23828 45668 23838
rect 45612 23378 45668 23772
rect 45612 23326 45614 23378
rect 45666 23326 45668 23378
rect 45612 23314 45668 23326
rect 45500 23102 45502 23154
rect 45554 23102 45556 23154
rect 45500 23090 45556 23102
rect 44716 22542 44718 22594
rect 44770 22542 44772 22594
rect 44716 22530 44772 22542
rect 44940 23044 44996 23054
rect 44156 22146 44212 22158
rect 44156 22094 44158 22146
rect 44210 22094 44212 22146
rect 44156 22036 44212 22094
rect 44156 21970 44212 21980
rect 44940 22146 44996 22988
rect 44940 22094 44942 22146
rect 44994 22094 44996 22146
rect 44716 21476 44772 21486
rect 44380 20916 44436 20926
rect 44268 20356 44324 20366
rect 44044 20300 44268 20356
rect 44268 20290 44324 20300
rect 44380 20132 44436 20860
rect 44716 20692 44772 21420
rect 44940 20916 44996 22094
rect 45052 22594 45108 22606
rect 45052 22542 45054 22594
rect 45106 22542 45108 22594
rect 45052 20916 45108 22542
rect 45276 22482 45332 22494
rect 45276 22430 45278 22482
rect 45330 22430 45332 22482
rect 45276 21812 45332 22430
rect 45276 21746 45332 21756
rect 45500 21364 45556 21374
rect 45276 20916 45332 20926
rect 45052 20914 45332 20916
rect 45052 20862 45278 20914
rect 45330 20862 45332 20914
rect 45052 20860 45332 20862
rect 44940 20822 44996 20860
rect 45276 20850 45332 20860
rect 45388 20916 45444 20926
rect 44716 20636 44996 20692
rect 44380 20066 44436 20076
rect 43708 20020 43764 20030
rect 43708 19460 43764 19964
rect 43708 19394 43764 19404
rect 44268 19908 44324 19918
rect 44604 19908 44660 19918
rect 43820 19236 43876 19246
rect 43596 19182 43598 19234
rect 43650 19182 43652 19234
rect 43596 19170 43652 19182
rect 43708 19234 43876 19236
rect 43708 19182 43822 19234
rect 43874 19182 43876 19234
rect 43708 19180 43876 19182
rect 43260 18398 43262 18450
rect 43314 18398 43316 18450
rect 43260 18386 43316 18398
rect 43372 19124 43428 19134
rect 43372 18452 43428 19068
rect 43372 18386 43428 18396
rect 43484 19010 43540 19022
rect 43484 18958 43486 19010
rect 43538 18958 43540 19010
rect 43148 18338 43204 18350
rect 43148 18286 43150 18338
rect 43202 18286 43204 18338
rect 43148 18228 43204 18286
rect 42812 18172 43204 18228
rect 42924 17668 42980 17678
rect 42924 17666 43092 17668
rect 42924 17614 42926 17666
rect 42978 17614 43092 17666
rect 42924 17612 43092 17614
rect 42924 17602 42980 17612
rect 42924 17332 42980 17342
rect 42700 17108 42756 17118
rect 42700 16882 42756 17052
rect 42700 16830 42702 16882
rect 42754 16830 42756 16882
rect 42700 16818 42756 16830
rect 42924 16882 42980 17276
rect 43036 16996 43092 17612
rect 43036 16930 43092 16940
rect 42924 16830 42926 16882
rect 42978 16830 42980 16882
rect 42924 16818 42980 16830
rect 43148 16772 43204 18172
rect 43260 17666 43316 17678
rect 43260 17614 43262 17666
rect 43314 17614 43316 17666
rect 43260 16884 43316 17614
rect 43372 17666 43428 17678
rect 43372 17614 43374 17666
rect 43426 17614 43428 17666
rect 43372 17108 43428 17614
rect 43484 17444 43540 18958
rect 43596 18452 43652 18462
rect 43596 18358 43652 18396
rect 43708 18004 43764 19180
rect 43820 19170 43876 19180
rect 44268 19236 44324 19852
rect 44268 19170 44324 19180
rect 44380 19906 44660 19908
rect 44380 19854 44606 19906
rect 44658 19854 44660 19906
rect 44380 19852 44660 19854
rect 44268 18564 44324 18574
rect 43596 17948 43764 18004
rect 43820 18562 44324 18564
rect 43820 18510 44270 18562
rect 44322 18510 44324 18562
rect 43820 18508 44324 18510
rect 43596 17668 43652 17948
rect 43596 17602 43652 17612
rect 43708 17780 43764 17790
rect 43820 17780 43876 18508
rect 44268 18498 44324 18508
rect 43932 18340 43988 18350
rect 43932 18246 43988 18284
rect 44380 18340 44436 19852
rect 44604 19842 44660 19852
rect 44828 19234 44884 19246
rect 44828 19182 44830 19234
rect 44882 19182 44884 19234
rect 44828 19124 44884 19182
rect 44828 19058 44884 19068
rect 44940 19122 44996 20636
rect 45276 20356 45332 20366
rect 45052 20020 45108 20030
rect 45052 19926 45108 19964
rect 44940 19070 44942 19122
rect 44994 19070 44996 19122
rect 44940 19058 44996 19070
rect 45164 19346 45220 19358
rect 45164 19294 45166 19346
rect 45218 19294 45220 19346
rect 44940 18676 44996 18686
rect 44380 18274 44436 18284
rect 44604 18450 44660 18462
rect 44604 18398 44606 18450
rect 44658 18398 44660 18450
rect 44044 18228 44100 18238
rect 44044 18134 44100 18172
rect 44604 18004 44660 18398
rect 44828 18452 44884 18462
rect 44828 18358 44884 18396
rect 44940 18338 44996 18620
rect 44940 18286 44942 18338
rect 44994 18286 44996 18338
rect 44940 18274 44996 18286
rect 45164 18564 45220 19294
rect 43764 17724 43876 17780
rect 43932 17948 44660 18004
rect 45052 18228 45108 18238
rect 43708 17554 43764 17724
rect 43708 17502 43710 17554
rect 43762 17502 43764 17554
rect 43708 17490 43764 17502
rect 43932 17666 43988 17948
rect 44268 17836 44884 17892
rect 43932 17614 43934 17666
rect 43986 17614 43988 17666
rect 43484 17378 43540 17388
rect 43372 17042 43428 17052
rect 43596 17332 43652 17342
rect 43596 17106 43652 17276
rect 43596 17054 43598 17106
rect 43650 17054 43652 17106
rect 43596 17042 43652 17054
rect 43820 17108 43876 17118
rect 43820 17014 43876 17052
rect 43260 16818 43316 16828
rect 43148 16706 43204 16716
rect 43708 16770 43764 16782
rect 43708 16718 43710 16770
rect 43762 16718 43764 16770
rect 42924 16660 42980 16670
rect 42924 16098 42980 16604
rect 43260 16660 43316 16670
rect 43260 16658 43652 16660
rect 43260 16606 43262 16658
rect 43314 16606 43652 16658
rect 43260 16604 43652 16606
rect 42924 16046 42926 16098
rect 42978 16046 42980 16098
rect 42924 16034 42980 16046
rect 43148 16548 43204 16558
rect 43148 16098 43204 16492
rect 43148 16046 43150 16098
rect 43202 16046 43204 16098
rect 43148 16034 43204 16046
rect 43036 15874 43092 15886
rect 43036 15822 43038 15874
rect 43090 15822 43092 15874
rect 43036 15652 43092 15822
rect 43036 15586 43092 15596
rect 41804 13972 41860 15148
rect 41916 15138 41972 15148
rect 42252 15092 42532 15148
rect 42588 15540 42644 15550
rect 41916 13972 41972 13982
rect 41804 13970 41972 13972
rect 41804 13918 41918 13970
rect 41970 13918 41972 13970
rect 41804 13916 41972 13918
rect 41468 13906 41524 13916
rect 41132 13746 41188 13758
rect 41132 13694 41134 13746
rect 41186 13694 41188 13746
rect 41132 13076 41188 13694
rect 41132 13010 41188 13020
rect 41916 12964 41972 13916
rect 41916 12908 42196 12964
rect 41916 12738 41972 12750
rect 41916 12686 41918 12738
rect 41970 12686 41972 12738
rect 41916 12628 41972 12686
rect 41916 12562 41972 12572
rect 42028 12740 42084 12750
rect 40908 12348 41076 12404
rect 39004 11116 39508 11172
rect 38892 10836 38948 10846
rect 38780 10780 38892 10836
rect 38892 10742 38948 10780
rect 39452 10834 39508 11116
rect 39564 11170 39620 11182
rect 39564 11118 39566 11170
rect 39618 11118 39620 11170
rect 39564 11060 39620 11118
rect 39564 10994 39620 11004
rect 39676 11172 39732 11182
rect 39452 10782 39454 10834
rect 39506 10782 39508 10834
rect 39452 10770 39508 10782
rect 39676 10722 39732 11116
rect 39788 11172 39844 11182
rect 39788 11170 39956 11172
rect 39788 11118 39790 11170
rect 39842 11118 39956 11170
rect 39788 11116 39956 11118
rect 39788 11106 39844 11116
rect 39676 10670 39678 10722
rect 39730 10670 39732 10722
rect 39676 10658 39732 10670
rect 37548 10098 37604 10108
rect 37996 10220 38724 10276
rect 39564 10612 39620 10622
rect 37996 9938 38052 10220
rect 37996 9886 37998 9938
rect 38050 9886 38052 9938
rect 37996 9874 38052 9886
rect 38108 9380 38164 9390
rect 37772 8932 37828 8942
rect 37772 8838 37828 8876
rect 37660 8372 37716 8382
rect 37548 8260 37604 8270
rect 37436 8258 37604 8260
rect 37436 8206 37550 8258
rect 37602 8206 37604 8258
rect 37436 8204 37604 8206
rect 37548 8194 37604 8204
rect 37660 8146 37716 8316
rect 37660 8094 37662 8146
rect 37714 8094 37716 8146
rect 37660 8082 37716 8094
rect 37100 7970 37156 7980
rect 37548 8036 37604 8046
rect 37548 7698 37604 7980
rect 37548 7646 37550 7698
rect 37602 7646 37604 7698
rect 37548 7634 37604 7646
rect 38108 7700 38164 9324
rect 39564 9266 39620 10556
rect 39564 9214 39566 9266
rect 39618 9214 39620 9266
rect 39564 9202 39620 9214
rect 39788 10498 39844 10510
rect 39788 10446 39790 10498
rect 39842 10446 39844 10498
rect 38668 9154 38724 9166
rect 38668 9102 38670 9154
rect 38722 9102 38724 9154
rect 38556 7700 38612 7710
rect 38108 7698 38612 7700
rect 38108 7646 38558 7698
rect 38610 7646 38612 7698
rect 38108 7644 38612 7646
rect 37884 7586 37940 7598
rect 37884 7534 37886 7586
rect 37938 7534 37940 7586
rect 37100 7252 37156 7262
rect 37100 7250 37380 7252
rect 37100 7198 37102 7250
rect 37154 7198 37380 7250
rect 37100 7196 37380 7198
rect 37100 7186 37156 7196
rect 37324 6692 37380 7196
rect 37324 6690 37492 6692
rect 37324 6638 37326 6690
rect 37378 6638 37492 6690
rect 37324 6636 37492 6638
rect 37324 6626 37380 6636
rect 37436 6356 37492 6636
rect 37548 6580 37604 6590
rect 37548 6486 37604 6524
rect 37772 6580 37828 6590
rect 37772 6486 37828 6524
rect 37884 6468 37940 7534
rect 37996 7588 38052 7598
rect 37996 6690 38052 7532
rect 38108 7474 38164 7644
rect 38556 7634 38612 7644
rect 38668 7588 38724 9102
rect 39788 9156 39844 10446
rect 39900 9940 39956 11116
rect 40236 11060 40292 11676
rect 40908 12178 40964 12190
rect 40908 12126 40910 12178
rect 40962 12126 40964 12178
rect 40236 10994 40292 11004
rect 40572 11172 40628 11182
rect 40908 11172 40964 12126
rect 40572 11170 40964 11172
rect 40572 11118 40574 11170
rect 40626 11118 40964 11170
rect 40572 11116 40964 11118
rect 40572 10836 40628 11116
rect 40572 10770 40628 10780
rect 41020 11060 41076 12348
rect 42028 12292 42084 12684
rect 41692 12068 41748 12078
rect 41244 12066 41748 12068
rect 41244 12014 41694 12066
rect 41746 12014 41748 12066
rect 41244 12012 41748 12014
rect 41132 11508 41188 11518
rect 41132 11394 41188 11452
rect 41244 11506 41300 12012
rect 41692 12002 41748 12012
rect 41244 11454 41246 11506
rect 41298 11454 41300 11506
rect 41244 11442 41300 11454
rect 41132 11342 41134 11394
rect 41186 11342 41188 11394
rect 41132 11284 41188 11342
rect 41132 11218 41188 11228
rect 41356 11394 41412 11406
rect 41356 11342 41358 11394
rect 41410 11342 41412 11394
rect 41356 11060 41412 11342
rect 41020 11004 41412 11060
rect 41468 11396 41524 11406
rect 40796 10724 40852 10734
rect 40012 10612 40068 10622
rect 40012 10518 40068 10556
rect 40236 10612 40292 10622
rect 40236 10518 40292 10556
rect 40796 10610 40852 10668
rect 40796 10558 40798 10610
rect 40850 10558 40852 10610
rect 40796 10546 40852 10558
rect 40124 9940 40180 9950
rect 39900 9938 40180 9940
rect 39900 9886 40126 9938
rect 40178 9886 40180 9938
rect 39900 9884 40180 9886
rect 39788 9090 39844 9100
rect 39004 9042 39060 9054
rect 39004 8990 39006 9042
rect 39058 8990 39060 9042
rect 39004 8036 39060 8990
rect 39676 8260 39732 8270
rect 39676 8166 39732 8204
rect 39004 7970 39060 7980
rect 38892 7700 38948 7710
rect 38892 7606 38948 7644
rect 39900 7698 39956 7710
rect 39900 7646 39902 7698
rect 39954 7646 39956 7698
rect 38668 7522 38724 7532
rect 39564 7588 39620 7598
rect 38108 7422 38110 7474
rect 38162 7422 38164 7474
rect 38108 7410 38164 7422
rect 39564 7474 39620 7532
rect 39564 7422 39566 7474
rect 39618 7422 39620 7474
rect 39564 7410 39620 7422
rect 37996 6638 37998 6690
rect 38050 6638 38052 6690
rect 37996 6626 38052 6638
rect 39900 6692 39956 7646
rect 40012 7586 40068 9884
rect 40124 9874 40180 9884
rect 40908 9716 40964 9726
rect 41020 9716 41076 11004
rect 41132 10836 41188 10846
rect 41132 9940 41188 10780
rect 41468 10836 41524 11340
rect 41692 11284 41748 11294
rect 41692 11190 41748 11228
rect 41468 10834 41972 10836
rect 41468 10782 41470 10834
rect 41522 10782 41972 10834
rect 41468 10780 41972 10782
rect 41468 10770 41524 10780
rect 41916 10722 41972 10780
rect 41916 10670 41918 10722
rect 41970 10670 41972 10722
rect 41916 10658 41972 10670
rect 42028 10724 42084 12236
rect 42028 10630 42084 10668
rect 41244 10610 41300 10622
rect 41244 10558 41246 10610
rect 41298 10558 41300 10610
rect 41244 10164 41300 10558
rect 41356 10612 41412 10622
rect 41356 10518 41412 10556
rect 42140 10612 42196 12908
rect 42252 12740 42308 15092
rect 42588 14420 42644 15484
rect 43036 15428 43092 15438
rect 42700 15316 42756 15326
rect 42700 15222 42756 15260
rect 43036 15314 43092 15372
rect 43036 15262 43038 15314
rect 43090 15262 43092 15314
rect 43036 15250 43092 15262
rect 43260 15314 43316 16604
rect 43372 16100 43428 16110
rect 43596 16100 43652 16604
rect 43708 16324 43764 16718
rect 43932 16548 43988 17614
rect 44044 17780 44100 17790
rect 44044 17108 44100 17724
rect 44268 17778 44324 17836
rect 44268 17726 44270 17778
rect 44322 17726 44324 17778
rect 44268 17714 44324 17726
rect 44828 17778 44884 17836
rect 44828 17726 44830 17778
rect 44882 17726 44884 17778
rect 44828 17714 44884 17726
rect 44156 17668 44212 17678
rect 44156 17574 44212 17612
rect 44380 17556 44436 17566
rect 44044 17052 44324 17108
rect 44156 16884 44212 16894
rect 43932 16482 43988 16492
rect 44044 16882 44212 16884
rect 44044 16830 44158 16882
rect 44210 16830 44212 16882
rect 44044 16828 44212 16830
rect 44044 16548 44100 16828
rect 44156 16818 44212 16828
rect 44156 16548 44212 16558
rect 44044 16492 44156 16548
rect 43820 16324 43876 16334
rect 43708 16322 43876 16324
rect 43708 16270 43822 16322
rect 43874 16270 43876 16322
rect 43708 16268 43876 16270
rect 43820 16258 43876 16268
rect 44044 16212 44100 16492
rect 44156 16482 44212 16492
rect 44044 16146 44100 16156
rect 44268 16210 44324 17052
rect 44268 16158 44270 16210
rect 44322 16158 44324 16210
rect 43708 16100 43764 16110
rect 43428 16044 43540 16100
rect 43596 16044 43708 16100
rect 43372 16034 43428 16044
rect 43372 15876 43428 15886
rect 43372 15782 43428 15820
rect 43260 15262 43262 15314
rect 43314 15262 43316 15314
rect 43260 15250 43316 15262
rect 43484 15148 43540 16044
rect 43708 16006 43764 16044
rect 43596 15652 43652 15662
rect 43596 15426 43652 15596
rect 43596 15374 43598 15426
rect 43650 15374 43652 15426
rect 43596 15362 43652 15374
rect 43708 15316 43764 15326
rect 43708 15222 43764 15260
rect 44156 15314 44212 15326
rect 44156 15262 44158 15314
rect 44210 15262 44212 15314
rect 43372 15092 43540 15148
rect 44156 15204 44212 15262
rect 42364 14364 42644 14420
rect 42924 14868 42980 14878
rect 42364 13858 42420 14364
rect 42364 13806 42366 13858
rect 42418 13806 42420 13858
rect 42364 13794 42420 13806
rect 42476 13524 42532 13534
rect 42700 13524 42756 13534
rect 42476 13522 42756 13524
rect 42476 13470 42478 13522
rect 42530 13470 42702 13522
rect 42754 13470 42756 13522
rect 42476 13468 42756 13470
rect 42476 13458 42532 13468
rect 42700 13458 42756 13468
rect 42364 12740 42420 12750
rect 42252 12684 42364 12740
rect 42364 12646 42420 12684
rect 42700 12628 42756 12638
rect 42252 11508 42308 11518
rect 42252 11394 42308 11452
rect 42252 11342 42254 11394
rect 42306 11342 42308 11394
rect 42252 11330 42308 11342
rect 42588 11282 42644 11294
rect 42588 11230 42590 11282
rect 42642 11230 42644 11282
rect 42476 11172 42532 11182
rect 42476 11078 42532 11116
rect 42588 10948 42644 11230
rect 42700 11282 42756 12572
rect 42700 11230 42702 11282
rect 42754 11230 42756 11282
rect 42700 11218 42756 11230
rect 42924 11060 42980 14812
rect 43036 14420 43092 14430
rect 43036 13970 43092 14364
rect 43036 13918 43038 13970
rect 43090 13918 43092 13970
rect 43036 13906 43092 13918
rect 43372 13970 43428 15092
rect 44156 14530 44212 15148
rect 44156 14478 44158 14530
rect 44210 14478 44212 14530
rect 43372 13918 43374 13970
rect 43426 13918 43428 13970
rect 43372 13906 43428 13918
rect 43484 14418 43540 14430
rect 43484 14366 43486 14418
rect 43538 14366 43540 14418
rect 43484 13522 43540 14366
rect 43820 13972 43876 13982
rect 44156 13972 44212 14478
rect 44268 14420 44324 16158
rect 44380 15876 44436 17500
rect 44940 17556 44996 17566
rect 44940 17462 44996 17500
rect 44716 17332 44772 17342
rect 44380 15810 44436 15820
rect 44492 17276 44716 17332
rect 44492 16882 44548 17276
rect 44716 17266 44772 17276
rect 45052 17220 45108 18172
rect 45164 17332 45220 18508
rect 45164 17266 45220 17276
rect 45052 17106 45108 17164
rect 45052 17054 45054 17106
rect 45106 17054 45108 17106
rect 45052 17042 45108 17054
rect 44492 16830 44494 16882
rect 44546 16830 44548 16882
rect 44492 15148 44548 16830
rect 44716 16772 44772 16782
rect 44716 16678 44772 16716
rect 45164 16324 45220 16334
rect 45052 16100 45108 16110
rect 45052 16006 45108 16044
rect 44940 15988 44996 15998
rect 44940 15894 44996 15932
rect 44828 15874 44884 15886
rect 44828 15822 44830 15874
rect 44882 15822 44884 15874
rect 44828 15764 44884 15822
rect 44828 15698 44884 15708
rect 45164 15652 45220 16268
rect 44940 15596 45220 15652
rect 44604 15316 44660 15326
rect 44828 15316 44884 15326
rect 44660 15314 44884 15316
rect 44660 15262 44830 15314
rect 44882 15262 44884 15314
rect 44660 15260 44884 15262
rect 44604 15250 44660 15260
rect 44828 15250 44884 15260
rect 44268 14354 44324 14364
rect 44380 15092 44548 15148
rect 44940 15204 44996 15596
rect 43820 13970 44212 13972
rect 43820 13918 43822 13970
rect 43874 13918 44212 13970
rect 43820 13916 44212 13918
rect 43820 13906 43876 13916
rect 44380 13860 44436 15092
rect 44940 14644 44996 15148
rect 45164 15428 45220 15438
rect 45164 14980 45220 15372
rect 45276 15148 45332 20300
rect 45388 18450 45444 20860
rect 45500 20132 45556 21308
rect 45500 20066 45556 20076
rect 45724 20020 45780 24444
rect 45948 23604 46004 26908
rect 46396 26964 46452 26974
rect 46508 26964 46564 27692
rect 46396 26962 46564 26964
rect 46396 26910 46398 26962
rect 46450 26910 46564 26962
rect 46396 26908 46564 26910
rect 46732 26964 46788 28140
rect 46956 27076 47012 28364
rect 47180 28354 47236 28364
rect 47404 28420 47460 28430
rect 47404 28418 47572 28420
rect 47404 28366 47406 28418
rect 47458 28366 47572 28418
rect 47404 28364 47572 28366
rect 47404 28354 47460 28364
rect 47404 27746 47460 27758
rect 47404 27694 47406 27746
rect 47458 27694 47460 27746
rect 47292 27188 47348 27198
rect 47404 27188 47460 27694
rect 47292 27186 47460 27188
rect 47292 27134 47294 27186
rect 47346 27134 47460 27186
rect 47292 27132 47460 27134
rect 47292 27122 47348 27132
rect 47068 27076 47124 27086
rect 46956 27074 47124 27076
rect 46956 27022 47070 27074
rect 47122 27022 47124 27074
rect 46956 27020 47124 27022
rect 47068 27010 47124 27020
rect 47516 27074 47572 28364
rect 47516 27022 47518 27074
rect 47570 27022 47572 27074
rect 47516 27010 47572 27022
rect 47740 27076 47796 28476
rect 47740 27010 47796 27020
rect 48076 27858 48132 27870
rect 48076 27806 48078 27858
rect 48130 27806 48132 27858
rect 46844 26964 46900 26974
rect 46732 26962 46900 26964
rect 46732 26910 46846 26962
rect 46898 26910 46900 26962
rect 46732 26908 46900 26910
rect 47852 26964 47908 27002
rect 46396 26898 46452 26908
rect 46620 26850 46676 26862
rect 46844 26852 47236 26908
rect 47852 26898 47908 26908
rect 46620 26798 46622 26850
rect 46674 26798 46676 26850
rect 46620 26290 46676 26798
rect 46620 26238 46622 26290
rect 46674 26238 46676 26290
rect 46620 26226 46676 26238
rect 46956 26290 47012 26302
rect 46956 26238 46958 26290
rect 47010 26238 47012 26290
rect 46844 26180 46900 26190
rect 46732 26178 46900 26180
rect 46732 26126 46846 26178
rect 46898 26126 46900 26178
rect 46732 26124 46900 26126
rect 46732 25732 46788 26124
rect 46844 26114 46900 26124
rect 46060 25676 46788 25732
rect 46060 25618 46116 25676
rect 46060 25566 46062 25618
rect 46114 25566 46116 25618
rect 46060 25554 46116 25566
rect 46956 25172 47012 26238
rect 47180 26290 47236 26852
rect 47180 26238 47182 26290
rect 47234 26238 47236 26290
rect 47180 26226 47236 26238
rect 48076 25844 48132 27806
rect 48188 26964 48244 26974
rect 48300 26964 48356 26974
rect 48188 26962 48300 26964
rect 48188 26910 48190 26962
rect 48242 26910 48300 26962
rect 48188 26908 48300 26910
rect 48188 26898 48244 26908
rect 48300 26514 48356 26908
rect 48300 26462 48302 26514
rect 48354 26462 48356 26514
rect 48300 26450 48356 26462
rect 48076 25788 48356 25844
rect 48188 25620 48244 25630
rect 47628 25618 48244 25620
rect 47628 25566 48190 25618
rect 48242 25566 48244 25618
rect 47628 25564 48244 25566
rect 46956 25116 47348 25172
rect 46284 24948 46340 24958
rect 46172 24612 46228 24622
rect 46172 24518 46228 24556
rect 45948 23548 46116 23604
rect 45948 23266 46004 23278
rect 45948 23214 45950 23266
rect 46002 23214 46004 23266
rect 45836 23156 45892 23166
rect 45948 23156 46004 23214
rect 45836 23154 46004 23156
rect 45836 23102 45838 23154
rect 45890 23102 46004 23154
rect 45836 23100 46004 23102
rect 45836 23090 45892 23100
rect 46060 21700 46116 23548
rect 46172 23268 46228 23278
rect 46172 23174 46228 23212
rect 46284 23268 46340 24892
rect 47292 24946 47348 25116
rect 47628 24948 47684 25564
rect 48188 25554 48244 25564
rect 47292 24894 47294 24946
rect 47346 24894 47348 24946
rect 47292 24882 47348 24894
rect 47404 24946 47684 24948
rect 47404 24894 47630 24946
rect 47682 24894 47684 24946
rect 47404 24892 47684 24894
rect 47068 24834 47124 24846
rect 47068 24782 47070 24834
rect 47122 24782 47124 24834
rect 46732 24724 46788 24734
rect 46956 24724 47012 24734
rect 46788 24722 47012 24724
rect 46788 24670 46958 24722
rect 47010 24670 47012 24722
rect 46788 24668 47012 24670
rect 47068 24724 47124 24782
rect 47404 24724 47460 24892
rect 47628 24882 47684 24892
rect 47068 24668 47460 24724
rect 47516 24724 47572 24734
rect 46620 23380 46676 23390
rect 46284 23266 46564 23268
rect 46284 23214 46286 23266
rect 46338 23214 46564 23266
rect 46284 23212 46564 23214
rect 46284 23202 46340 23212
rect 46060 21634 46116 21644
rect 46508 21698 46564 23212
rect 46620 23266 46676 23324
rect 46620 23214 46622 23266
rect 46674 23214 46676 23266
rect 46620 23202 46676 23214
rect 46620 21812 46676 21822
rect 46620 21718 46676 21756
rect 46508 21646 46510 21698
rect 46562 21646 46564 21698
rect 46508 21634 46564 21646
rect 46732 21700 46788 24668
rect 46956 24658 47012 24668
rect 47516 24630 47572 24668
rect 48300 24612 48356 25788
rect 47628 24500 47684 24510
rect 47292 24498 47684 24500
rect 47292 24446 47630 24498
rect 47682 24446 47684 24498
rect 47292 24444 47684 24446
rect 46956 23828 47012 23838
rect 46956 23734 47012 23772
rect 46844 23156 46900 23166
rect 46844 21810 46900 23100
rect 46844 21758 46846 21810
rect 46898 21758 46900 21810
rect 46844 21746 46900 21758
rect 46956 23154 47012 23166
rect 46956 23102 46958 23154
rect 47010 23102 47012 23154
rect 46732 21634 46788 21644
rect 46284 21474 46340 21486
rect 46284 21422 46286 21474
rect 46338 21422 46340 21474
rect 46284 21140 46340 21422
rect 46956 21364 47012 23102
rect 47292 23154 47348 24444
rect 47628 24434 47684 24444
rect 48300 24052 48356 24556
rect 47740 23996 48356 24052
rect 47740 23938 47796 23996
rect 47740 23886 47742 23938
rect 47794 23886 47796 23938
rect 47740 23874 47796 23886
rect 47740 23492 47796 23502
rect 47292 23102 47294 23154
rect 47346 23102 47348 23154
rect 47292 23090 47348 23102
rect 47404 23156 47460 23166
rect 47404 23062 47460 23100
rect 47740 23154 47796 23436
rect 48076 23380 48132 23390
rect 48076 23266 48132 23324
rect 48076 23214 48078 23266
rect 48130 23214 48132 23266
rect 48076 23202 48132 23214
rect 47740 23102 47742 23154
rect 47794 23102 47796 23154
rect 47740 23090 47796 23102
rect 47068 23042 47124 23054
rect 47068 22990 47070 23042
rect 47122 22990 47124 23042
rect 47068 22708 47124 22990
rect 47628 23042 47684 23054
rect 47628 22990 47630 23042
rect 47682 22990 47684 23042
rect 47068 22652 47460 22708
rect 47404 22482 47460 22652
rect 47404 22430 47406 22482
rect 47458 22430 47460 22482
rect 47404 22418 47460 22430
rect 47628 21924 47684 22990
rect 48188 22372 48244 23996
rect 47404 21868 47684 21924
rect 48076 22370 48244 22372
rect 48076 22318 48190 22370
rect 48242 22318 48244 22370
rect 48076 22316 48244 22318
rect 47180 21812 47236 21822
rect 47180 21718 47236 21756
rect 47068 21700 47124 21710
rect 47068 21606 47124 21644
rect 47180 21364 47236 21374
rect 46956 21362 47236 21364
rect 46956 21310 47182 21362
rect 47234 21310 47236 21362
rect 46956 21308 47236 21310
rect 47180 21298 47236 21308
rect 46284 21074 46340 21084
rect 46844 20916 46900 20926
rect 45724 19926 45780 19964
rect 46172 20020 46228 20030
rect 46172 19926 46228 19964
rect 46620 19908 46676 19918
rect 46284 19292 46564 19348
rect 45948 19236 46004 19246
rect 46284 19236 46340 19292
rect 45388 18398 45390 18450
rect 45442 18398 45444 18450
rect 45388 18386 45444 18398
rect 45836 19234 46340 19236
rect 45836 19182 45950 19234
rect 46002 19182 46340 19234
rect 45836 19180 46340 19182
rect 45388 17668 45444 17678
rect 45388 17666 45780 17668
rect 45388 17614 45390 17666
rect 45442 17614 45780 17666
rect 45388 17612 45780 17614
rect 45388 17602 45444 17612
rect 45388 17444 45444 17454
rect 45388 16882 45444 17388
rect 45612 17220 45668 17230
rect 45612 17106 45668 17164
rect 45612 17054 45614 17106
rect 45666 17054 45668 17106
rect 45388 16830 45390 16882
rect 45442 16830 45444 16882
rect 45388 16660 45444 16830
rect 45500 16884 45556 16894
rect 45500 16770 45556 16828
rect 45500 16718 45502 16770
rect 45554 16718 45556 16770
rect 45500 16706 45556 16718
rect 45388 16594 45444 16604
rect 45388 16436 45444 16446
rect 45388 16098 45444 16380
rect 45388 16046 45390 16098
rect 45442 16046 45444 16098
rect 45388 16034 45444 16046
rect 45612 16100 45668 17054
rect 45724 16324 45780 17612
rect 45724 16258 45780 16268
rect 45724 16100 45780 16110
rect 45612 16098 45780 16100
rect 45612 16046 45726 16098
rect 45778 16046 45780 16098
rect 45612 16044 45780 16046
rect 45724 16034 45780 16044
rect 45836 15148 45892 19180
rect 45948 19170 46004 19180
rect 46396 19122 46452 19134
rect 46396 19070 46398 19122
rect 46450 19070 46452 19122
rect 46284 19012 46340 19022
rect 46060 19010 46340 19012
rect 46060 18958 46286 19010
rect 46338 18958 46340 19010
rect 46060 18956 46340 18958
rect 46060 18562 46116 18956
rect 46284 18946 46340 18956
rect 46396 18676 46452 19070
rect 46508 19122 46564 19292
rect 46508 19070 46510 19122
rect 46562 19070 46564 19122
rect 46508 19058 46564 19070
rect 46396 18610 46452 18620
rect 46060 18510 46062 18562
rect 46114 18510 46116 18562
rect 46060 18498 46116 18510
rect 46060 17556 46116 17566
rect 46060 17462 46116 17500
rect 46060 17220 46116 17230
rect 46060 16882 46116 17164
rect 46060 16830 46062 16882
rect 46114 16830 46116 16882
rect 45948 16660 46004 16670
rect 45948 16322 46004 16604
rect 46060 16548 46116 16830
rect 46284 16884 46340 16894
rect 46284 16790 46340 16828
rect 46508 16884 46564 16894
rect 46060 16482 46116 16492
rect 45948 16270 45950 16322
rect 46002 16270 46004 16322
rect 45948 16258 46004 16270
rect 46284 16324 46340 16334
rect 46508 16324 46564 16828
rect 46284 16322 46564 16324
rect 46284 16270 46286 16322
rect 46338 16270 46564 16322
rect 46284 16268 46564 16270
rect 46284 16258 46340 16268
rect 46620 15148 46676 19852
rect 46844 19346 46900 20860
rect 47404 20914 47460 21868
rect 47404 20862 47406 20914
rect 47458 20862 47460 20914
rect 47404 20850 47460 20862
rect 47852 21698 47908 21710
rect 47852 21646 47854 21698
rect 47906 21646 47908 21698
rect 47516 20132 47572 20142
rect 47516 20038 47572 20076
rect 47852 20130 47908 21646
rect 48076 20916 48132 22316
rect 48188 22306 48244 22316
rect 48188 21586 48244 21598
rect 48188 21534 48190 21586
rect 48242 21534 48244 21586
rect 48188 21140 48244 21534
rect 48188 21074 48244 21084
rect 48076 20802 48132 20860
rect 48076 20750 48078 20802
rect 48130 20750 48132 20802
rect 48076 20738 48132 20750
rect 47852 20078 47854 20130
rect 47906 20078 47908 20130
rect 47852 20066 47908 20078
rect 46844 19294 46846 19346
rect 46898 19294 46900 19346
rect 46844 19282 46900 19294
rect 46732 19122 46788 19134
rect 46732 19070 46734 19122
rect 46786 19070 46788 19122
rect 46732 16770 46788 19070
rect 46956 18452 47012 18462
rect 46732 16718 46734 16770
rect 46786 16718 46788 16770
rect 46732 16706 46788 16718
rect 46844 16772 46900 16782
rect 46732 16324 46788 16334
rect 46732 16210 46788 16268
rect 46732 16158 46734 16210
rect 46786 16158 46788 16210
rect 46732 16146 46788 16158
rect 46844 15204 46900 16716
rect 46956 16770 47012 18396
rect 48188 18452 48244 18462
rect 48188 18338 48244 18396
rect 48188 18286 48190 18338
rect 48242 18286 48244 18338
rect 48188 18274 48244 18286
rect 48188 17778 48244 17790
rect 48188 17726 48190 17778
rect 48242 17726 48244 17778
rect 47180 17668 47236 17678
rect 47180 16882 47236 17612
rect 48188 17668 48244 17726
rect 48188 17602 48244 17612
rect 47852 17220 47908 17230
rect 47852 17106 47908 17164
rect 47852 17054 47854 17106
rect 47906 17054 47908 17106
rect 47852 17042 47908 17054
rect 47180 16830 47182 16882
rect 47234 16830 47236 16882
rect 47180 16818 47236 16830
rect 47404 16882 47460 16894
rect 47404 16830 47406 16882
rect 47458 16830 47460 16882
rect 46956 16718 46958 16770
rect 47010 16718 47012 16770
rect 46956 16706 47012 16718
rect 47404 16772 47460 16830
rect 47404 16706 47460 16716
rect 47852 16212 47908 16222
rect 47852 15986 47908 16156
rect 47852 15934 47854 15986
rect 47906 15934 47908 15986
rect 47852 15922 47908 15934
rect 48188 15986 48244 15998
rect 48188 15934 48190 15986
rect 48242 15934 48244 15986
rect 47628 15876 47684 15886
rect 47628 15782 47684 15820
rect 48188 15876 48244 15934
rect 48188 15316 48244 15820
rect 48188 15250 48244 15260
rect 46956 15204 47012 15214
rect 46844 15202 47012 15204
rect 46844 15150 46958 15202
rect 47010 15150 47012 15202
rect 46844 15148 47012 15150
rect 45276 15082 45332 15092
rect 45612 15092 45892 15148
rect 46172 15092 46676 15148
rect 46956 15138 47012 15148
rect 45164 14924 45556 14980
rect 43484 13470 43486 13522
rect 43538 13470 43540 13522
rect 43484 13458 43540 13470
rect 43932 13804 44436 13860
rect 44828 14642 44996 14644
rect 44828 14590 44942 14642
rect 44994 14590 44996 14642
rect 44828 14588 44996 14590
rect 43932 12962 43988 13804
rect 44492 13748 44548 13758
rect 44380 13746 44548 13748
rect 44380 13694 44494 13746
rect 44546 13694 44548 13746
rect 44380 13692 44548 13694
rect 44268 13636 44324 13646
rect 44268 13542 44324 13580
rect 43932 12910 43934 12962
rect 43986 12910 43988 12962
rect 43932 12898 43988 12910
rect 44268 12964 44324 12974
rect 44380 12964 44436 13692
rect 44492 13682 44548 13692
rect 44716 13634 44772 13646
rect 44716 13582 44718 13634
rect 44770 13582 44772 13634
rect 44716 13188 44772 13582
rect 44716 13122 44772 13132
rect 44828 12964 44884 14588
rect 44940 14578 44996 14588
rect 44940 13748 44996 13758
rect 44940 13654 44996 13692
rect 45052 13746 45108 13758
rect 45052 13694 45054 13746
rect 45106 13694 45108 13746
rect 44268 12962 44436 12964
rect 44268 12910 44270 12962
rect 44322 12910 44436 12962
rect 44268 12908 44436 12910
rect 44492 12962 44884 12964
rect 44492 12910 44830 12962
rect 44882 12910 44884 12962
rect 44492 12908 44884 12910
rect 44268 12898 44324 12908
rect 43708 12740 43764 12750
rect 44044 12740 44100 12750
rect 43708 12738 44100 12740
rect 43708 12686 43710 12738
rect 43762 12686 44046 12738
rect 44098 12686 44100 12738
rect 43708 12684 44100 12686
rect 43708 12674 43764 12684
rect 43820 12068 43876 12078
rect 43708 12066 43876 12068
rect 43708 12014 43822 12066
rect 43874 12014 43876 12066
rect 43708 12012 43876 12014
rect 43036 11508 43092 11518
rect 43036 11506 43316 11508
rect 43036 11454 43038 11506
rect 43090 11454 43316 11506
rect 43036 11452 43316 11454
rect 43036 11442 43092 11452
rect 42252 10892 42644 10948
rect 42700 11004 42980 11060
rect 42252 10834 42308 10892
rect 42252 10782 42254 10834
rect 42306 10782 42308 10834
rect 42252 10770 42308 10782
rect 42476 10612 42532 10622
rect 42140 10610 42532 10612
rect 42140 10558 42478 10610
rect 42530 10558 42532 10610
rect 42140 10556 42532 10558
rect 42140 10164 42196 10556
rect 42476 10546 42532 10556
rect 41244 10098 41300 10108
rect 41804 10108 42196 10164
rect 41244 9940 41300 9950
rect 41804 9940 41860 10108
rect 42364 10052 42420 10062
rect 42420 9996 42532 10052
rect 42364 9986 42420 9996
rect 41132 9938 41300 9940
rect 41132 9886 41246 9938
rect 41298 9886 41300 9938
rect 41132 9884 41300 9886
rect 41244 9874 41300 9884
rect 41356 9938 41860 9940
rect 41356 9886 41806 9938
rect 41858 9886 41860 9938
rect 41356 9884 41860 9886
rect 40908 9714 41076 9716
rect 40908 9662 40910 9714
rect 40962 9662 41076 9714
rect 40908 9660 41076 9662
rect 40908 9650 40964 9660
rect 41020 9044 41076 9054
rect 41356 9044 41412 9884
rect 41804 9874 41860 9884
rect 41580 9716 41636 9726
rect 41020 9042 41412 9044
rect 41020 8990 41022 9042
rect 41074 8990 41412 9042
rect 41020 8988 41412 8990
rect 41020 8978 41076 8988
rect 40236 8148 40292 8158
rect 40236 8054 40292 8092
rect 41244 8148 41300 8158
rect 41244 8034 41300 8092
rect 41244 7982 41246 8034
rect 41298 7982 41300 8034
rect 41244 7970 41300 7982
rect 40012 7534 40014 7586
rect 40066 7534 40068 7586
rect 40012 7522 40068 7534
rect 40236 7474 40292 7486
rect 40236 7422 40238 7474
rect 40290 7422 40292 7474
rect 40124 6804 40180 6814
rect 40124 6692 40180 6748
rect 39900 6690 40180 6692
rect 39900 6638 40126 6690
rect 40178 6638 40180 6690
rect 39900 6636 40180 6638
rect 40124 6626 40180 6636
rect 38780 6580 38836 6590
rect 38780 6486 38836 6524
rect 39788 6580 39844 6590
rect 38332 6468 38388 6478
rect 37884 6466 38388 6468
rect 37884 6414 38334 6466
rect 38386 6414 38388 6466
rect 37884 6412 38388 6414
rect 38332 6356 38388 6412
rect 37436 6300 38276 6356
rect 37044 6188 37492 6244
rect 36988 6150 37044 6188
rect 36988 5908 37044 5918
rect 36876 5906 37044 5908
rect 36876 5854 36990 5906
rect 37042 5854 37044 5906
rect 36876 5852 37044 5854
rect 36316 5234 36372 5292
rect 36316 5182 36318 5234
rect 36370 5182 36372 5234
rect 36316 5170 36372 5182
rect 36148 5068 36260 5124
rect 36092 5058 36148 5068
rect 35980 4174 35982 4226
rect 36034 4174 36036 4226
rect 35980 4162 36036 4174
rect 35196 3948 35460 3958
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35196 3882 35460 3892
rect 22876 3614 22878 3666
rect 22930 3614 22932 3666
rect 22876 3602 22932 3614
rect 36204 3668 36260 5068
rect 36428 4900 36484 4910
rect 36428 4806 36484 4844
rect 36316 4228 36372 4238
rect 36876 4228 36932 5852
rect 36988 5842 37044 5852
rect 37212 5234 37268 6188
rect 37436 6018 37492 6188
rect 37436 5966 37438 6018
rect 37490 5966 37492 6018
rect 37436 5954 37492 5966
rect 37772 6020 37828 6030
rect 37772 5926 37828 5964
rect 38220 6018 38276 6300
rect 38220 5966 38222 6018
rect 38274 5966 38276 6018
rect 38108 5796 38164 5806
rect 37548 5794 38164 5796
rect 37548 5742 38110 5794
rect 38162 5742 38164 5794
rect 37548 5740 38164 5742
rect 37548 5348 37604 5740
rect 38108 5730 38164 5740
rect 38220 5572 38276 5966
rect 37212 5182 37214 5234
rect 37266 5182 37268 5234
rect 37212 5170 37268 5182
rect 37436 5292 37604 5348
rect 37884 5516 38276 5572
rect 37436 5234 37492 5292
rect 37436 5182 37438 5234
rect 37490 5182 37492 5234
rect 37436 5170 37492 5182
rect 37884 5234 37940 5516
rect 38332 5348 38388 6300
rect 38556 6466 38612 6478
rect 38556 6414 38558 6466
rect 38610 6414 38612 6466
rect 38556 6132 38612 6414
rect 38668 6466 38724 6478
rect 38668 6414 38670 6466
rect 38722 6414 38724 6466
rect 38668 6244 38724 6414
rect 39676 6468 39732 6478
rect 39676 6374 39732 6412
rect 38668 6188 39172 6244
rect 38556 6066 38612 6076
rect 38444 6020 38500 6030
rect 38444 5906 38500 5964
rect 38444 5854 38446 5906
rect 38498 5854 38500 5906
rect 38444 5684 38500 5854
rect 38668 6018 38724 6030
rect 38668 5966 38670 6018
rect 38722 5966 38724 6018
rect 38668 5796 38724 5966
rect 39004 5908 39060 5918
rect 39004 5814 39060 5852
rect 39116 5906 39172 6188
rect 39116 5854 39118 5906
rect 39170 5854 39172 5906
rect 39116 5842 39172 5854
rect 39452 5908 39508 5918
rect 39452 5814 39508 5852
rect 39788 5906 39844 6524
rect 39900 6466 39956 6478
rect 39900 6414 39902 6466
rect 39954 6414 39956 6466
rect 39900 6356 39956 6414
rect 40012 6468 40068 6478
rect 40012 6374 40068 6412
rect 39900 6290 39956 6300
rect 40236 6244 40292 7422
rect 41244 7252 41300 7262
rect 41244 7158 41300 7196
rect 40684 6804 40740 6814
rect 40684 6710 40740 6748
rect 40460 6690 40516 6702
rect 40460 6638 40462 6690
rect 40514 6638 40516 6690
rect 40460 6580 40516 6638
rect 41356 6692 41412 8988
rect 41356 6626 41412 6636
rect 41468 9660 41580 9716
rect 41468 7700 41524 9660
rect 41580 9650 41636 9660
rect 42140 9604 42196 9614
rect 42028 9602 42196 9604
rect 42028 9550 42142 9602
rect 42194 9550 42196 9602
rect 42028 9548 42196 9550
rect 41692 9156 41748 9166
rect 41692 9062 41748 9100
rect 41804 8372 41860 8382
rect 41468 6690 41524 7644
rect 41580 8036 41636 8046
rect 41580 7474 41636 7980
rect 41580 7422 41582 7474
rect 41634 7422 41636 7474
rect 41580 7410 41636 7422
rect 41804 7474 41860 8316
rect 42028 8036 42084 9548
rect 42140 9538 42196 9548
rect 42252 9602 42308 9614
rect 42252 9550 42254 9602
rect 42306 9550 42308 9602
rect 42252 8260 42308 9550
rect 42364 9602 42420 9614
rect 42364 9550 42366 9602
rect 42418 9550 42420 9602
rect 42364 8484 42420 9550
rect 42364 8418 42420 8428
rect 42476 8820 42532 9996
rect 42700 9826 42756 11004
rect 42700 9774 42702 9826
rect 42754 9774 42756 9826
rect 42700 9716 42756 9774
rect 42700 9650 42756 9660
rect 42812 10836 42868 10846
rect 42252 8204 42420 8260
rect 42028 7970 42084 7980
rect 42140 8148 42196 8158
rect 42140 7588 42196 8092
rect 42252 8036 42308 8046
rect 42252 7942 42308 7980
rect 42140 7522 42196 7532
rect 41804 7422 41806 7474
rect 41858 7422 41860 7474
rect 41804 7410 41860 7422
rect 41692 7252 41748 7262
rect 42140 7252 42196 7262
rect 41692 6916 41748 7196
rect 41916 7250 42196 7252
rect 41916 7198 42142 7250
rect 42194 7198 42196 7250
rect 41916 7196 42196 7198
rect 41804 6916 41860 6926
rect 41692 6860 41804 6916
rect 41468 6638 41470 6690
rect 41522 6638 41524 6690
rect 41468 6626 41524 6638
rect 41692 6692 41748 6702
rect 40460 6356 40516 6524
rect 40460 6290 40516 6300
rect 40908 6468 40964 6478
rect 40236 6178 40292 6188
rect 40012 6132 40068 6142
rect 39788 5854 39790 5906
rect 39842 5854 39844 5906
rect 39788 5842 39844 5854
rect 39900 6020 39956 6030
rect 38668 5730 38724 5740
rect 38444 5618 38500 5628
rect 38332 5282 38388 5292
rect 37884 5182 37886 5234
rect 37938 5182 37940 5234
rect 37884 5170 37940 5182
rect 37548 5124 37604 5134
rect 37548 5030 37604 5068
rect 38444 4900 38500 4910
rect 38444 4450 38500 4844
rect 39900 4562 39956 5964
rect 40012 5906 40068 6076
rect 40012 5854 40014 5906
rect 40066 5854 40068 5906
rect 40012 5842 40068 5854
rect 40908 5906 40964 6412
rect 40908 5854 40910 5906
rect 40962 5854 40964 5906
rect 40908 5842 40964 5854
rect 41020 6466 41076 6478
rect 41020 6414 41022 6466
rect 41074 6414 41076 6466
rect 41020 6132 41076 6414
rect 41020 5906 41076 6076
rect 41020 5854 41022 5906
rect 41074 5854 41076 5906
rect 41020 5842 41076 5854
rect 41244 6468 41300 6478
rect 41244 6018 41300 6412
rect 41244 5966 41246 6018
rect 41298 5966 41300 6018
rect 41244 5796 41300 5966
rect 41580 6020 41636 6030
rect 41580 5926 41636 5964
rect 41244 5730 41300 5740
rect 41468 5348 41524 5358
rect 41132 5346 41524 5348
rect 41132 5294 41470 5346
rect 41522 5294 41524 5346
rect 41132 5292 41524 5294
rect 40796 5236 40852 5246
rect 40012 5124 40068 5134
rect 40012 5030 40068 5068
rect 40796 5122 40852 5180
rect 41132 5234 41188 5292
rect 41468 5282 41524 5292
rect 41132 5182 41134 5234
rect 41186 5182 41188 5234
rect 41132 5170 41188 5182
rect 41692 5236 41748 6636
rect 41804 6690 41860 6860
rect 41916 6802 41972 7196
rect 42140 7186 42196 7196
rect 42252 7250 42308 7262
rect 42252 7198 42254 7250
rect 42306 7198 42308 7250
rect 42140 6804 42196 6814
rect 41916 6750 41918 6802
rect 41970 6750 41972 6802
rect 41916 6738 41972 6750
rect 42028 6748 42140 6804
rect 41804 6638 41806 6690
rect 41858 6638 41860 6690
rect 41804 6626 41860 6638
rect 42028 6690 42084 6748
rect 42140 6738 42196 6748
rect 42028 6638 42030 6690
rect 42082 6638 42084 6690
rect 42028 6626 42084 6638
rect 42252 6580 42308 7198
rect 42364 6914 42420 8204
rect 42476 8258 42532 8764
rect 42476 8206 42478 8258
rect 42530 8206 42532 8258
rect 42476 8194 42532 8206
rect 42700 8148 42756 8158
rect 42700 8054 42756 8092
rect 42812 7700 42868 10780
rect 43260 10722 43316 11452
rect 43372 11396 43428 11406
rect 43372 11302 43428 11340
rect 43484 11284 43540 11294
rect 43484 11190 43540 11228
rect 43260 10670 43262 10722
rect 43314 10670 43316 10722
rect 43260 10658 43316 10670
rect 43596 11172 43652 11182
rect 43708 11172 43764 12012
rect 43820 12002 43876 12012
rect 43596 11170 43764 11172
rect 43596 11118 43598 11170
rect 43650 11118 43764 11170
rect 43596 11116 43764 11118
rect 43820 11170 43876 11182
rect 43820 11118 43822 11170
rect 43874 11118 43876 11170
rect 43372 9828 43428 9838
rect 43372 9826 43540 9828
rect 43372 9774 43374 9826
rect 43426 9774 43540 9826
rect 43372 9772 43540 9774
rect 43372 9762 43428 9772
rect 43260 9602 43316 9614
rect 43260 9550 43262 9602
rect 43314 9550 43316 9602
rect 43260 8372 43316 9550
rect 43484 8932 43540 9772
rect 43596 9604 43652 11116
rect 43820 11060 43876 11118
rect 43820 10994 43876 11004
rect 43932 9826 43988 9838
rect 43932 9774 43934 9826
rect 43986 9774 43988 9826
rect 43596 9548 43764 9604
rect 43484 8484 43540 8876
rect 43596 8484 43652 8494
rect 43484 8482 43652 8484
rect 43484 8430 43598 8482
rect 43650 8430 43652 8482
rect 43484 8428 43652 8430
rect 43596 8418 43652 8428
rect 43260 8306 43316 8316
rect 43148 8260 43204 8270
rect 43148 8166 43204 8204
rect 43372 8148 43428 8158
rect 43260 8092 43372 8148
rect 42812 7644 43092 7700
rect 42588 7586 42644 7598
rect 42588 7534 42590 7586
rect 42642 7534 42644 7586
rect 42588 7140 42644 7534
rect 42812 7586 42868 7644
rect 42812 7534 42814 7586
rect 42866 7534 42868 7586
rect 42812 7522 42868 7534
rect 42924 7474 42980 7486
rect 42924 7422 42926 7474
rect 42978 7422 42980 7474
rect 42588 7084 42868 7140
rect 42364 6862 42366 6914
rect 42418 6862 42420 6914
rect 42364 6850 42420 6862
rect 42476 6972 42756 7028
rect 42476 6916 42532 6972
rect 42476 6822 42532 6860
rect 41804 6244 41860 6254
rect 41804 6020 41860 6188
rect 42252 6130 42308 6524
rect 42252 6078 42254 6130
rect 42306 6078 42308 6130
rect 42252 6066 42308 6078
rect 42588 6804 42644 6814
rect 41916 6020 41972 6030
rect 41804 5964 41916 6020
rect 41804 5906 41860 5964
rect 41916 5954 41972 5964
rect 41804 5854 41806 5906
rect 41858 5854 41860 5906
rect 41804 5842 41860 5854
rect 42588 5906 42644 6748
rect 42588 5854 42590 5906
rect 42642 5854 42644 5906
rect 42588 5842 42644 5854
rect 42700 5908 42756 6972
rect 42812 6468 42868 7084
rect 42812 6374 42868 6412
rect 42812 5908 42868 5918
rect 42700 5906 42868 5908
rect 42700 5854 42814 5906
rect 42866 5854 42868 5906
rect 42700 5852 42868 5854
rect 42812 5842 42868 5852
rect 41916 5794 41972 5806
rect 41916 5742 41918 5794
rect 41970 5742 41972 5794
rect 41804 5348 41860 5358
rect 41916 5348 41972 5742
rect 41804 5346 41972 5348
rect 41804 5294 41806 5346
rect 41858 5294 41972 5346
rect 41804 5292 41972 5294
rect 41804 5282 41860 5292
rect 41692 5142 41748 5180
rect 42812 5236 42868 5246
rect 42924 5236 42980 7422
rect 43036 6690 43092 7644
rect 43148 7476 43204 7486
rect 43148 7382 43204 7420
rect 43036 6638 43038 6690
rect 43090 6638 43092 6690
rect 43036 6626 43092 6638
rect 43260 6916 43316 8092
rect 43372 8082 43428 8092
rect 43484 7588 43540 7598
rect 43484 7494 43540 7532
rect 43708 7474 43764 9548
rect 43820 8930 43876 8942
rect 43820 8878 43822 8930
rect 43874 8878 43876 8930
rect 43820 8820 43876 8878
rect 43820 8754 43876 8764
rect 43820 8258 43876 8270
rect 43820 8206 43822 8258
rect 43874 8206 43876 8258
rect 43820 8148 43876 8206
rect 43820 8082 43876 8092
rect 43932 7588 43988 9774
rect 44044 8708 44100 12684
rect 44492 12402 44548 12908
rect 44828 12898 44884 12908
rect 45052 13636 45108 13694
rect 45388 13748 45444 13758
rect 45388 13654 45444 13692
rect 44492 12350 44494 12402
rect 44546 12350 44548 12402
rect 44492 12338 44548 12350
rect 44940 11282 44996 11294
rect 44940 11230 44942 11282
rect 44994 11230 44996 11282
rect 44828 11172 44884 11182
rect 44828 11078 44884 11116
rect 44268 10388 44324 10398
rect 44268 9714 44324 10332
rect 44940 10388 44996 11230
rect 44940 10322 44996 10332
rect 45052 10164 45108 13580
rect 45388 10498 45444 10510
rect 45388 10446 45390 10498
rect 45442 10446 45444 10498
rect 45388 10388 45444 10446
rect 45388 10322 45444 10332
rect 44828 10108 45108 10164
rect 45500 10164 45556 14924
rect 45612 13858 45668 15092
rect 46172 13972 46228 15092
rect 45612 13806 45614 13858
rect 45666 13806 45668 13858
rect 45612 13636 45668 13806
rect 45724 13970 46228 13972
rect 45724 13918 46174 13970
rect 46226 13918 46228 13970
rect 45724 13916 46228 13918
rect 45724 13858 45780 13916
rect 46172 13906 46228 13916
rect 46956 13972 47012 13982
rect 45724 13806 45726 13858
rect 45778 13806 45780 13858
rect 45724 13794 45780 13806
rect 45612 13580 45780 13636
rect 45612 13188 45668 13198
rect 45612 13074 45668 13132
rect 45612 13022 45614 13074
rect 45666 13022 45668 13074
rect 45612 13010 45668 13022
rect 45724 13076 45780 13580
rect 45724 13010 45780 13020
rect 46956 11732 47012 13916
rect 47740 13076 47796 13086
rect 47740 12982 47796 13020
rect 46956 11676 47572 11732
rect 47516 10834 47572 11676
rect 47516 10782 47518 10834
rect 47570 10782 47572 10834
rect 47516 10770 47572 10782
rect 45948 10724 46004 10734
rect 45500 10108 45668 10164
rect 44828 9940 44884 10108
rect 44828 9826 44884 9884
rect 44828 9774 44830 9826
rect 44882 9774 44884 9826
rect 44828 9762 44884 9774
rect 45164 9826 45220 9838
rect 45164 9774 45166 9826
rect 45218 9774 45220 9826
rect 44268 9662 44270 9714
rect 44322 9662 44324 9714
rect 44268 9650 44324 9662
rect 44940 9716 44996 9726
rect 44492 8932 44548 8942
rect 44492 8838 44548 8876
rect 44044 8642 44100 8652
rect 44940 8482 44996 9660
rect 45164 8820 45220 9774
rect 45388 9716 45444 9726
rect 45388 9622 45444 9660
rect 45276 9604 45332 9614
rect 45276 9510 45332 9548
rect 45164 8764 45556 8820
rect 44940 8430 44942 8482
rect 44994 8430 44996 8482
rect 44940 8418 44996 8430
rect 45052 8708 45108 8718
rect 44828 8372 44884 8382
rect 43932 7522 43988 7532
rect 44044 8258 44100 8270
rect 44044 8206 44046 8258
rect 44098 8206 44100 8258
rect 43708 7422 43710 7474
rect 43762 7422 43764 7474
rect 43708 7410 43764 7422
rect 44044 7476 44100 8206
rect 44828 8258 44884 8316
rect 44828 8206 44830 8258
rect 44882 8206 44884 8258
rect 44828 8194 44884 8206
rect 45052 8372 45108 8652
rect 45500 8482 45556 8764
rect 45500 8430 45502 8482
rect 45554 8430 45556 8482
rect 45500 8418 45556 8430
rect 44268 8148 44324 8158
rect 44044 7382 44100 7420
rect 44156 8146 44324 8148
rect 44156 8094 44270 8146
rect 44322 8094 44324 8146
rect 44156 8092 44324 8094
rect 43260 6690 43316 6860
rect 43596 7362 43652 7374
rect 43596 7310 43598 7362
rect 43650 7310 43652 7362
rect 43260 6638 43262 6690
rect 43314 6638 43316 6690
rect 43260 6626 43316 6638
rect 43372 6802 43428 6814
rect 43372 6750 43374 6802
rect 43426 6750 43428 6802
rect 43372 6468 43428 6750
rect 43596 6804 43652 7310
rect 44156 7028 44212 8092
rect 44268 8082 44324 8092
rect 44940 8148 44996 8158
rect 45052 8148 45108 8316
rect 45612 8260 45668 10108
rect 45836 9940 45892 9950
rect 45836 9846 45892 9884
rect 44940 8146 45108 8148
rect 44940 8094 44942 8146
rect 44994 8094 45108 8146
rect 44940 8092 45108 8094
rect 45388 8258 45668 8260
rect 45388 8206 45614 8258
rect 45666 8206 45668 8258
rect 45388 8204 45668 8206
rect 44940 8082 44996 8092
rect 45388 7698 45444 8204
rect 45612 8194 45668 8204
rect 45724 8932 45780 8942
rect 45500 8036 45556 8046
rect 45724 8036 45780 8876
rect 45500 8034 45780 8036
rect 45500 7982 45502 8034
rect 45554 7982 45780 8034
rect 45500 7980 45780 7982
rect 45500 7970 45556 7980
rect 45388 7646 45390 7698
rect 45442 7646 45444 7698
rect 45388 7634 45444 7646
rect 43596 6738 43652 6748
rect 43708 6972 44212 7028
rect 44380 7476 44436 7486
rect 43372 6402 43428 6412
rect 42812 5234 42980 5236
rect 42812 5182 42814 5234
rect 42866 5182 42980 5234
rect 42812 5180 42980 5182
rect 43708 6020 43764 6972
rect 43820 6692 43876 6702
rect 43876 6636 44100 6692
rect 43820 6598 43876 6636
rect 42812 5170 42868 5180
rect 40796 5070 40798 5122
rect 40850 5070 40852 5122
rect 39900 4510 39902 4562
rect 39954 4510 39956 4562
rect 39900 4498 39956 4510
rect 40124 5012 40180 5022
rect 38444 4398 38446 4450
rect 38498 4398 38500 4450
rect 38444 4386 38500 4398
rect 39228 4340 39284 4350
rect 39228 4246 39284 4284
rect 40012 4340 40068 4350
rect 36316 4226 36932 4228
rect 36316 4174 36318 4226
rect 36370 4174 36932 4226
rect 36316 4172 36932 4174
rect 36316 4162 36372 4172
rect 36316 3668 36372 3678
rect 36204 3666 36372 3668
rect 36204 3614 36318 3666
rect 36370 3614 36372 3666
rect 36204 3612 36372 3614
rect 36316 3602 36372 3612
rect 40012 3666 40068 4284
rect 40124 4338 40180 4956
rect 40124 4286 40126 4338
rect 40178 4286 40180 4338
rect 40124 4274 40180 4286
rect 40796 4340 40852 5070
rect 41244 4900 41300 4910
rect 42924 4900 42980 4910
rect 41244 4898 41748 4900
rect 41244 4846 41246 4898
rect 41298 4846 41748 4898
rect 41244 4844 41748 4846
rect 41244 4834 41300 4844
rect 41692 4450 41748 4844
rect 42924 4806 42980 4844
rect 41692 4398 41694 4450
rect 41746 4398 41748 4450
rect 41692 4386 41748 4398
rect 40908 4340 40964 4350
rect 40852 4338 40964 4340
rect 40852 4286 40910 4338
rect 40962 4286 40964 4338
rect 40852 4284 40964 4286
rect 40796 4246 40852 4284
rect 40908 4274 40964 4284
rect 43708 4228 43764 5964
rect 44044 5234 44100 6636
rect 44156 6578 44212 6590
rect 44156 6526 44158 6578
rect 44210 6526 44212 6578
rect 44156 6468 44212 6526
rect 44268 6580 44324 6590
rect 44268 6486 44324 6524
rect 44156 6402 44212 6412
rect 44044 5182 44046 5234
rect 44098 5182 44100 5234
rect 44044 5124 44100 5182
rect 43820 4228 43876 4238
rect 43708 4226 43876 4228
rect 43708 4174 43822 4226
rect 43874 4174 43876 4226
rect 43708 4172 43876 4174
rect 43820 4162 43876 4172
rect 40012 3614 40014 3666
rect 40066 3614 40068 3666
rect 40012 3602 40068 3614
rect 43932 3668 43988 3678
rect 44044 3668 44100 5068
rect 44156 4228 44212 4238
rect 44380 4228 44436 7420
rect 44492 7364 44548 7374
rect 44940 7364 44996 7374
rect 44492 7362 44996 7364
rect 44492 7310 44494 7362
rect 44546 7310 44942 7362
rect 44994 7310 44996 7362
rect 44492 7308 44996 7310
rect 44492 6692 44548 7308
rect 44940 7298 44996 7308
rect 44828 6916 44884 6926
rect 44828 6802 44884 6860
rect 44828 6750 44830 6802
rect 44882 6750 44884 6802
rect 44828 6738 44884 6750
rect 44492 6626 44548 6636
rect 45948 4340 46004 10668
rect 47628 10500 47684 10510
rect 47628 10498 47908 10500
rect 47628 10446 47630 10498
rect 47682 10446 47908 10498
rect 47628 10444 47908 10446
rect 47628 10434 47684 10444
rect 47852 9714 47908 10444
rect 47852 9662 47854 9714
rect 47906 9662 47908 9714
rect 47852 9650 47908 9662
rect 48188 9714 48244 9726
rect 48188 9662 48190 9714
rect 48242 9662 48244 9714
rect 46620 9604 46676 9614
rect 46620 9154 46676 9548
rect 47628 9602 47684 9614
rect 47628 9550 47630 9602
rect 47682 9550 47684 9602
rect 47628 9492 47684 9550
rect 47628 9426 47684 9436
rect 48188 9492 48244 9662
rect 48188 9426 48244 9436
rect 46620 9102 46622 9154
rect 46674 9102 46676 9154
rect 46620 9090 46676 9102
rect 47292 9042 47348 9054
rect 47292 8990 47294 9042
rect 47346 8990 47348 9042
rect 46060 8372 46116 8382
rect 46060 8278 46116 8316
rect 47292 6692 47348 8990
rect 47628 6692 47684 6702
rect 47292 6690 47684 6692
rect 47292 6638 47630 6690
rect 47682 6638 47684 6690
rect 47292 6636 47684 6638
rect 46956 6580 47012 6590
rect 46956 6486 47012 6524
rect 47068 5124 47124 5134
rect 47292 5124 47348 6636
rect 47628 6626 47684 6636
rect 47124 5068 47348 5124
rect 46284 4900 46340 4910
rect 46284 4450 46340 4844
rect 46284 4398 46286 4450
rect 46338 4398 46340 4450
rect 46284 4386 46340 4398
rect 45948 4274 46004 4284
rect 47068 4338 47124 5068
rect 47068 4286 47070 4338
rect 47122 4286 47124 4338
rect 47068 4274 47124 4286
rect 47628 4340 47684 4350
rect 47628 4246 47684 4284
rect 48188 4338 48244 4350
rect 48188 4286 48190 4338
rect 48242 4286 48244 4338
rect 44156 4226 44436 4228
rect 44156 4174 44158 4226
rect 44210 4174 44436 4226
rect 44156 4172 44436 4174
rect 44156 4162 44212 4172
rect 43932 3666 44100 3668
rect 43932 3614 43934 3666
rect 43986 3614 44100 3666
rect 43932 3612 44100 3614
rect 48188 3668 48244 4286
rect 48300 3668 48356 3678
rect 48188 3612 48300 3668
rect 43932 3602 43988 3612
rect 48300 3574 48356 3612
rect 19836 3164 20100 3174
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 19836 3098 20100 3108
<< via2 >>
rect 15372 56306 15428 56308
rect 15372 56254 15374 56306
rect 15374 56254 15426 56306
rect 15426 56254 15428 56306
rect 15372 56252 15428 56254
rect 16156 56252 16212 56308
rect 4476 55690 4532 55692
rect 4476 55638 4478 55690
rect 4478 55638 4530 55690
rect 4530 55638 4532 55690
rect 4476 55636 4532 55638
rect 4580 55690 4636 55692
rect 4580 55638 4582 55690
rect 4582 55638 4634 55690
rect 4634 55638 4636 55690
rect 4580 55636 4636 55638
rect 4684 55690 4740 55692
rect 4684 55638 4686 55690
rect 4686 55638 4738 55690
rect 4738 55638 4740 55690
rect 4684 55636 4740 55638
rect 6860 55020 6916 55076
rect 9324 54796 9380 54852
rect 4476 54122 4532 54124
rect 4476 54070 4478 54122
rect 4478 54070 4530 54122
rect 4530 54070 4532 54122
rect 4476 54068 4532 54070
rect 4580 54122 4636 54124
rect 4580 54070 4582 54122
rect 4582 54070 4634 54122
rect 4634 54070 4636 54122
rect 4580 54068 4636 54070
rect 4684 54122 4740 54124
rect 4684 54070 4686 54122
rect 4686 54070 4738 54122
rect 4738 54070 4740 54122
rect 4684 54068 4740 54070
rect 4172 52946 4228 52948
rect 4172 52894 4174 52946
rect 4174 52894 4226 52946
rect 4226 52894 4228 52946
rect 4172 52892 4228 52894
rect 1596 52332 1652 52388
rect 1484 48748 1540 48804
rect 1484 21756 1540 21812
rect 3724 51212 3780 51268
rect 1708 49756 1764 49812
rect 1820 50428 1876 50484
rect 1820 47516 1876 47572
rect 2156 49980 2212 50036
rect 2492 49196 2548 49252
rect 2268 48748 2324 48804
rect 10892 55132 10948 55188
rect 10332 54796 10388 54852
rect 10108 53564 10164 53620
rect 6188 52892 6244 52948
rect 4476 52554 4532 52556
rect 4476 52502 4478 52554
rect 4478 52502 4530 52554
rect 4530 52502 4532 52554
rect 4476 52500 4532 52502
rect 4580 52554 4636 52556
rect 4580 52502 4582 52554
rect 4582 52502 4634 52554
rect 4634 52502 4636 52554
rect 4580 52500 4636 52502
rect 4684 52554 4740 52556
rect 4684 52502 4686 52554
rect 4686 52502 4738 52554
rect 4738 52502 4740 52554
rect 4684 52500 4740 52502
rect 6972 52668 7028 52724
rect 4844 52220 4900 52276
rect 6076 52274 6132 52276
rect 6076 52222 6078 52274
rect 6078 52222 6130 52274
rect 6130 52222 6132 52274
rect 6076 52220 6132 52222
rect 5740 51602 5796 51604
rect 5740 51550 5742 51602
rect 5742 51550 5794 51602
rect 5794 51550 5796 51602
rect 5740 51548 5796 51550
rect 5516 51378 5572 51380
rect 5516 51326 5518 51378
rect 5518 51326 5570 51378
rect 5570 51326 5572 51378
rect 5516 51324 5572 51326
rect 6188 51548 6244 51604
rect 5964 51324 6020 51380
rect 4844 51266 4900 51268
rect 4844 51214 4846 51266
rect 4846 51214 4898 51266
rect 4898 51214 4900 51266
rect 4844 51212 4900 51214
rect 4476 50986 4532 50988
rect 4476 50934 4478 50986
rect 4478 50934 4530 50986
rect 4530 50934 4532 50986
rect 4476 50932 4532 50934
rect 4580 50986 4636 50988
rect 4580 50934 4582 50986
rect 4582 50934 4634 50986
rect 4634 50934 4636 50986
rect 4580 50932 4636 50934
rect 4684 50986 4740 50988
rect 4684 50934 4686 50986
rect 4686 50934 4738 50986
rect 4738 50934 4740 50986
rect 4684 50932 4740 50934
rect 4172 50428 4228 50484
rect 4844 50482 4900 50484
rect 4844 50430 4846 50482
rect 4846 50430 4898 50482
rect 4898 50430 4900 50482
rect 4844 50428 4900 50430
rect 4620 49698 4676 49700
rect 4620 49646 4622 49698
rect 4622 49646 4674 49698
rect 4674 49646 4676 49698
rect 4620 49644 4676 49646
rect 4956 49644 5012 49700
rect 4476 49418 4532 49420
rect 4476 49366 4478 49418
rect 4478 49366 4530 49418
rect 4530 49366 4532 49418
rect 4476 49364 4532 49366
rect 4580 49418 4636 49420
rect 4580 49366 4582 49418
rect 4582 49366 4634 49418
rect 4634 49366 4636 49418
rect 4580 49364 4636 49366
rect 4684 49418 4740 49420
rect 4684 49366 4686 49418
rect 4686 49366 4738 49418
rect 4738 49366 4740 49418
rect 4684 49364 4740 49366
rect 4732 49026 4788 49028
rect 4732 48974 4734 49026
rect 4734 48974 4786 49026
rect 4786 48974 4788 49026
rect 4732 48972 4788 48974
rect 5628 49644 5684 49700
rect 5516 49026 5572 49028
rect 5516 48974 5518 49026
rect 5518 48974 5570 49026
rect 5570 48974 5572 49026
rect 5516 48972 5572 48974
rect 5068 48914 5124 48916
rect 5068 48862 5070 48914
rect 5070 48862 5122 48914
rect 5122 48862 5124 48914
rect 5068 48860 5124 48862
rect 6860 51884 6916 51940
rect 7644 52332 7700 52388
rect 7532 51938 7588 51940
rect 7532 51886 7534 51938
rect 7534 51886 7586 51938
rect 7586 51886 7588 51938
rect 7532 51884 7588 51886
rect 7980 52946 8036 52948
rect 7980 52894 7982 52946
rect 7982 52894 8034 52946
rect 8034 52894 8036 52946
rect 7980 52892 8036 52894
rect 8988 52892 9044 52948
rect 8092 52668 8148 52724
rect 6412 51324 6468 51380
rect 6076 50428 6132 50484
rect 8092 51938 8148 51940
rect 8092 51886 8094 51938
rect 8094 51886 8146 51938
rect 8146 51886 8148 51938
rect 8092 51884 8148 51886
rect 8316 51324 8372 51380
rect 9324 51324 9380 51380
rect 8988 51266 9044 51268
rect 8988 51214 8990 51266
rect 8990 51214 9042 51266
rect 9042 51214 9044 51266
rect 8988 51212 9044 51214
rect 8876 50540 8932 50596
rect 6748 50316 6804 50372
rect 7980 50316 8036 50372
rect 5740 48860 5796 48916
rect 7420 49138 7476 49140
rect 7420 49086 7422 49138
rect 7422 49086 7474 49138
rect 7474 49086 7476 49138
rect 7420 49084 7476 49086
rect 5068 48636 5124 48692
rect 2380 48242 2436 48244
rect 2380 48190 2382 48242
rect 2382 48190 2434 48242
rect 2434 48190 2436 48242
rect 2380 48188 2436 48190
rect 3164 48242 3220 48244
rect 3164 48190 3166 48242
rect 3166 48190 3218 48242
rect 3218 48190 3220 48242
rect 3164 48188 3220 48190
rect 3276 47404 3332 47460
rect 2380 45218 2436 45220
rect 2380 45166 2382 45218
rect 2382 45166 2434 45218
rect 2434 45166 2436 45218
rect 2380 45164 2436 45166
rect 2828 45276 2884 45332
rect 2604 45052 2660 45108
rect 3276 45052 3332 45108
rect 3052 44940 3108 44996
rect 3276 44828 3332 44884
rect 3948 48188 4004 48244
rect 4172 48242 4228 48244
rect 4172 48190 4174 48242
rect 4174 48190 4226 48242
rect 4226 48190 4228 48242
rect 4172 48188 4228 48190
rect 4844 48188 4900 48244
rect 4172 47404 4228 47460
rect 3724 46674 3780 46676
rect 3724 46622 3726 46674
rect 3726 46622 3778 46674
rect 3778 46622 3780 46674
rect 3724 46620 3780 46622
rect 4476 47850 4532 47852
rect 4476 47798 4478 47850
rect 4478 47798 4530 47850
rect 4530 47798 4532 47850
rect 4476 47796 4532 47798
rect 4580 47850 4636 47852
rect 4580 47798 4582 47850
rect 4582 47798 4634 47850
rect 4634 47798 4636 47850
rect 4580 47796 4636 47798
rect 4684 47850 4740 47852
rect 4684 47798 4686 47850
rect 4686 47798 4738 47850
rect 4738 47798 4740 47850
rect 4684 47796 4740 47798
rect 4620 47404 4676 47460
rect 5852 48636 5908 48692
rect 5068 47570 5124 47572
rect 5068 47518 5070 47570
rect 5070 47518 5122 47570
rect 5122 47518 5124 47570
rect 5068 47516 5124 47518
rect 9772 51212 9828 51268
rect 9884 50594 9940 50596
rect 9884 50542 9886 50594
rect 9886 50542 9938 50594
rect 9938 50542 9940 50594
rect 9884 50540 9940 50542
rect 10332 52108 10388 52164
rect 10444 52220 10500 52276
rect 11564 55074 11620 55076
rect 11564 55022 11566 55074
rect 11566 55022 11618 55074
rect 11618 55022 11620 55074
rect 11564 55020 11620 55022
rect 11452 54908 11508 54964
rect 13468 55186 13524 55188
rect 13468 55134 13470 55186
rect 13470 55134 13522 55186
rect 13522 55134 13524 55186
rect 13468 55132 13524 55134
rect 12236 54908 12292 54964
rect 11004 54236 11060 54292
rect 12460 54290 12516 54292
rect 12460 54238 12462 54290
rect 12462 54238 12514 54290
rect 12514 54238 12516 54290
rect 12460 54236 12516 54238
rect 11116 53564 11172 53620
rect 11228 53676 11284 53732
rect 12460 53618 12516 53620
rect 12460 53566 12462 53618
rect 12462 53566 12514 53618
rect 12514 53566 12516 53618
rect 12460 53564 12516 53566
rect 12236 53340 12292 53396
rect 13804 54348 13860 54404
rect 13132 53788 13188 53844
rect 13692 53788 13748 53844
rect 12796 53452 12852 53508
rect 13580 53506 13636 53508
rect 13580 53454 13582 53506
rect 13582 53454 13634 53506
rect 13634 53454 13636 53506
rect 13580 53452 13636 53454
rect 11228 52946 11284 52948
rect 11228 52894 11230 52946
rect 11230 52894 11282 52946
rect 11282 52894 11284 52946
rect 11228 52892 11284 52894
rect 11116 52274 11172 52276
rect 11116 52222 11118 52274
rect 11118 52222 11170 52274
rect 11170 52222 11172 52274
rect 11116 52220 11172 52222
rect 13580 52220 13636 52276
rect 13580 51548 13636 51604
rect 14588 54348 14644 54404
rect 16492 54402 16548 54404
rect 16492 54350 16494 54402
rect 16494 54350 16546 54402
rect 16546 54350 16548 54402
rect 16492 54348 16548 54350
rect 17724 55970 17780 55972
rect 17724 55918 17726 55970
rect 17726 55918 17778 55970
rect 17778 55918 17780 55970
rect 17724 55916 17780 55918
rect 16940 54348 16996 54404
rect 18060 54460 18116 54516
rect 17724 54402 17780 54404
rect 17724 54350 17726 54402
rect 17726 54350 17778 54402
rect 17778 54350 17780 54402
rect 17724 54348 17780 54350
rect 14140 53618 14196 53620
rect 14140 53566 14142 53618
rect 14142 53566 14194 53618
rect 14194 53566 14196 53618
rect 14140 53564 14196 53566
rect 13804 52780 13860 52836
rect 11004 51436 11060 51492
rect 10332 51378 10388 51380
rect 10332 51326 10334 51378
rect 10334 51326 10386 51378
rect 10386 51326 10388 51378
rect 10332 51324 10388 51326
rect 7084 47458 7140 47460
rect 7084 47406 7086 47458
rect 7086 47406 7138 47458
rect 7138 47406 7140 47458
rect 7084 47404 7140 47406
rect 7308 47346 7364 47348
rect 7308 47294 7310 47346
rect 7310 47294 7362 47346
rect 7362 47294 7364 47346
rect 7308 47292 7364 47294
rect 6524 46956 6580 47012
rect 4844 46620 4900 46676
rect 4476 46282 4532 46284
rect 4476 46230 4478 46282
rect 4478 46230 4530 46282
rect 4530 46230 4532 46282
rect 4476 46228 4532 46230
rect 4580 46282 4636 46284
rect 4580 46230 4582 46282
rect 4582 46230 4634 46282
rect 4634 46230 4636 46282
rect 4580 46228 4636 46230
rect 4684 46282 4740 46284
rect 4684 46230 4686 46282
rect 4686 46230 4738 46282
rect 4738 46230 4740 46282
rect 4684 46228 4740 46230
rect 3612 45778 3668 45780
rect 3612 45726 3614 45778
rect 3614 45726 3666 45778
rect 3666 45726 3668 45778
rect 3612 45724 3668 45726
rect 3836 45330 3892 45332
rect 3836 45278 3838 45330
rect 3838 45278 3890 45330
rect 3890 45278 3892 45330
rect 3836 45276 3892 45278
rect 3724 45218 3780 45220
rect 3724 45166 3726 45218
rect 3726 45166 3778 45218
rect 3778 45166 3780 45218
rect 3724 45164 3780 45166
rect 3500 44940 3556 44996
rect 3836 45052 3892 45108
rect 3388 44716 3444 44772
rect 1820 41970 1876 41972
rect 1820 41918 1822 41970
rect 1822 41918 1874 41970
rect 1874 41918 1876 41970
rect 1820 41916 1876 41918
rect 1708 40460 1764 40516
rect 1820 36652 1876 36708
rect 1708 33628 1764 33684
rect 1820 30940 1876 30996
rect 1708 29820 1764 29876
rect 4060 44828 4116 44884
rect 4844 45778 4900 45780
rect 4844 45726 4846 45778
rect 4846 45726 4898 45778
rect 4898 45726 4900 45778
rect 4844 45724 4900 45726
rect 6300 45778 6356 45780
rect 6300 45726 6302 45778
rect 6302 45726 6354 45778
rect 6354 45726 6356 45778
rect 6300 45724 6356 45726
rect 7084 45724 7140 45780
rect 5964 45612 6020 45668
rect 6412 45612 6468 45668
rect 6860 45666 6916 45668
rect 6860 45614 6862 45666
rect 6862 45614 6914 45666
rect 6914 45614 6916 45666
rect 6860 45612 6916 45614
rect 7084 45164 7140 45220
rect 4844 45106 4900 45108
rect 4844 45054 4846 45106
rect 4846 45054 4898 45106
rect 4898 45054 4900 45106
rect 4844 45052 4900 45054
rect 4172 44940 4228 44996
rect 4396 44940 4452 44996
rect 5740 44940 5796 44996
rect 4284 44716 4340 44772
rect 4476 44714 4532 44716
rect 4476 44662 4478 44714
rect 4478 44662 4530 44714
rect 4530 44662 4532 44714
rect 4476 44660 4532 44662
rect 4580 44714 4636 44716
rect 4580 44662 4582 44714
rect 4582 44662 4634 44714
rect 4634 44662 4636 44714
rect 4580 44660 4636 44662
rect 4684 44714 4740 44716
rect 4684 44662 4686 44714
rect 4686 44662 4738 44714
rect 4738 44662 4740 44714
rect 4684 44660 4740 44662
rect 4284 43596 4340 43652
rect 3500 43372 3556 43428
rect 3164 42642 3220 42644
rect 3164 42590 3166 42642
rect 3166 42590 3218 42642
rect 3218 42590 3220 42642
rect 3164 42588 3220 42590
rect 2828 42476 2884 42532
rect 2604 42364 2660 42420
rect 3052 42476 3108 42532
rect 4172 42812 4228 42868
rect 3724 42530 3780 42532
rect 3724 42478 3726 42530
rect 3726 42478 3778 42530
rect 3778 42478 3780 42530
rect 3724 42476 3780 42478
rect 3948 42530 4004 42532
rect 3948 42478 3950 42530
rect 3950 42478 4002 42530
rect 4002 42478 4004 42530
rect 3948 42476 4004 42478
rect 3500 42028 3556 42084
rect 3164 40460 3220 40516
rect 2828 40348 2884 40404
rect 4060 42364 4116 42420
rect 3836 38722 3892 38724
rect 3836 38670 3838 38722
rect 3838 38670 3890 38722
rect 3890 38670 3892 38722
rect 3836 38668 3892 38670
rect 4396 43426 4452 43428
rect 4396 43374 4398 43426
rect 4398 43374 4450 43426
rect 4450 43374 4452 43426
rect 4396 43372 4452 43374
rect 4476 43146 4532 43148
rect 4476 43094 4478 43146
rect 4478 43094 4530 43146
rect 4530 43094 4532 43146
rect 4476 43092 4532 43094
rect 4580 43146 4636 43148
rect 4580 43094 4582 43146
rect 4582 43094 4634 43146
rect 4634 43094 4636 43146
rect 4580 43092 4636 43094
rect 4684 43146 4740 43148
rect 4684 43094 4686 43146
rect 4686 43094 4738 43146
rect 4738 43094 4740 43146
rect 4684 43092 4740 43094
rect 4844 42754 4900 42756
rect 4844 42702 4846 42754
rect 4846 42702 4898 42754
rect 4898 42702 4900 42754
rect 4844 42700 4900 42702
rect 4732 42530 4788 42532
rect 4732 42478 4734 42530
rect 4734 42478 4786 42530
rect 4786 42478 4788 42530
rect 4732 42476 4788 42478
rect 4284 42028 4340 42084
rect 6860 44322 6916 44324
rect 6860 44270 6862 44322
rect 6862 44270 6914 44322
rect 6914 44270 6916 44322
rect 6860 44268 6916 44270
rect 5404 43650 5460 43652
rect 5404 43598 5406 43650
rect 5406 43598 5458 43650
rect 5458 43598 5460 43650
rect 5404 43596 5460 43598
rect 5516 43372 5572 43428
rect 5516 42924 5572 42980
rect 5180 42700 5236 42756
rect 5740 42588 5796 42644
rect 5404 41970 5460 41972
rect 5404 41918 5406 41970
rect 5406 41918 5458 41970
rect 5458 41918 5460 41970
rect 5404 41916 5460 41918
rect 4476 41578 4532 41580
rect 4476 41526 4478 41578
rect 4478 41526 4530 41578
rect 4530 41526 4532 41578
rect 4476 41524 4532 41526
rect 4580 41578 4636 41580
rect 4580 41526 4582 41578
rect 4582 41526 4634 41578
rect 4634 41526 4636 41578
rect 4580 41524 4636 41526
rect 4684 41578 4740 41580
rect 4684 41526 4686 41578
rect 4686 41526 4738 41578
rect 4738 41526 4740 41578
rect 4684 41524 4740 41526
rect 4172 40572 4228 40628
rect 4508 40514 4564 40516
rect 4508 40462 4510 40514
rect 4510 40462 4562 40514
rect 4562 40462 4564 40514
rect 4508 40460 4564 40462
rect 4732 40460 4788 40516
rect 4476 40010 4532 40012
rect 4476 39958 4478 40010
rect 4478 39958 4530 40010
rect 4530 39958 4532 40010
rect 4476 39956 4532 39958
rect 4580 40010 4636 40012
rect 4580 39958 4582 40010
rect 4582 39958 4634 40010
rect 4634 39958 4636 40010
rect 4580 39956 4636 39958
rect 4684 40010 4740 40012
rect 4684 39958 4686 40010
rect 4686 39958 4738 40010
rect 4738 39958 4740 40010
rect 4684 39956 4740 39958
rect 2940 37378 2996 37380
rect 2940 37326 2942 37378
rect 2942 37326 2994 37378
rect 2994 37326 2996 37378
rect 2940 37324 2996 37326
rect 2828 37212 2884 37268
rect 4172 38556 4228 38612
rect 3724 37266 3780 37268
rect 3724 37214 3726 37266
rect 3726 37214 3778 37266
rect 3778 37214 3780 37266
rect 3724 37212 3780 37214
rect 2380 34524 2436 34580
rect 2492 34636 2548 34692
rect 2940 34524 2996 34580
rect 2492 33628 2548 33684
rect 2716 34076 2772 34132
rect 2604 33458 2660 33460
rect 2604 33406 2606 33458
rect 2606 33406 2658 33458
rect 2658 33406 2660 33458
rect 2604 33404 2660 33406
rect 3612 34802 3668 34804
rect 3612 34750 3614 34802
rect 3614 34750 3666 34802
rect 3666 34750 3668 34802
rect 3612 34748 3668 34750
rect 3500 34690 3556 34692
rect 3500 34638 3502 34690
rect 3502 34638 3554 34690
rect 3554 34638 3556 34690
rect 3500 34636 3556 34638
rect 2604 33068 2660 33124
rect 3612 34130 3668 34132
rect 3612 34078 3614 34130
rect 3614 34078 3666 34130
rect 3666 34078 3668 34130
rect 3612 34076 3668 34078
rect 3612 33458 3668 33460
rect 3612 33406 3614 33458
rect 3614 33406 3666 33458
rect 3666 33406 3668 33458
rect 3612 33404 3668 33406
rect 3388 33068 3444 33124
rect 3612 33180 3668 33236
rect 4844 39564 4900 39620
rect 4476 38442 4532 38444
rect 4476 38390 4478 38442
rect 4478 38390 4530 38442
rect 4530 38390 4532 38442
rect 4476 38388 4532 38390
rect 4580 38442 4636 38444
rect 4580 38390 4582 38442
rect 4582 38390 4634 38442
rect 4634 38390 4636 38442
rect 4580 38388 4636 38390
rect 4684 38442 4740 38444
rect 4684 38390 4686 38442
rect 4686 38390 4738 38442
rect 4738 38390 4740 38442
rect 4684 38388 4740 38390
rect 3948 36652 4004 36708
rect 4172 37324 4228 37380
rect 4172 36988 4228 37044
rect 5180 39116 5236 39172
rect 5068 38722 5124 38724
rect 5068 38670 5070 38722
rect 5070 38670 5122 38722
rect 5122 38670 5124 38722
rect 5068 38668 5124 38670
rect 4956 38610 5012 38612
rect 4956 38558 4958 38610
rect 4958 38558 5010 38610
rect 5010 38558 5012 38610
rect 4956 38556 5012 38558
rect 5740 40236 5796 40292
rect 5740 39618 5796 39620
rect 5740 39566 5742 39618
rect 5742 39566 5794 39618
rect 5794 39566 5796 39618
rect 5740 39564 5796 39566
rect 5292 38556 5348 38612
rect 5740 38556 5796 38612
rect 5180 37266 5236 37268
rect 5180 37214 5182 37266
rect 5182 37214 5234 37266
rect 5234 37214 5236 37266
rect 5180 37212 5236 37214
rect 4476 36874 4532 36876
rect 4476 36822 4478 36874
rect 4478 36822 4530 36874
rect 4530 36822 4532 36874
rect 4476 36820 4532 36822
rect 4580 36874 4636 36876
rect 4580 36822 4582 36874
rect 4582 36822 4634 36874
rect 4634 36822 4636 36874
rect 4580 36820 4636 36822
rect 4684 36874 4740 36876
rect 4684 36822 4686 36874
rect 4686 36822 4738 36874
rect 4738 36822 4740 36874
rect 4684 36820 4740 36822
rect 5068 36988 5124 37044
rect 4172 35868 4228 35924
rect 5404 36652 5460 36708
rect 6748 44044 6804 44100
rect 5964 42028 6020 42084
rect 6636 42642 6692 42644
rect 6636 42590 6638 42642
rect 6638 42590 6690 42642
rect 6690 42590 6692 42642
rect 6636 42588 6692 42590
rect 6748 42028 6804 42084
rect 6300 39116 6356 39172
rect 6524 39340 6580 39396
rect 6972 39116 7028 39172
rect 7308 41298 7364 41300
rect 7308 41246 7310 41298
rect 7310 41246 7362 41298
rect 7362 41246 7364 41298
rect 7308 41244 7364 41246
rect 8428 48636 8484 48692
rect 8652 48300 8708 48356
rect 7532 47404 7588 47460
rect 9100 48300 9156 48356
rect 8540 47570 8596 47572
rect 8540 47518 8542 47570
rect 8542 47518 8594 47570
rect 8594 47518 8596 47570
rect 8540 47516 8596 47518
rect 8876 47458 8932 47460
rect 8876 47406 8878 47458
rect 8878 47406 8930 47458
rect 8930 47406 8932 47458
rect 8876 47404 8932 47406
rect 9884 48748 9940 48804
rect 9660 48354 9716 48356
rect 9660 48302 9662 48354
rect 9662 48302 9714 48354
rect 9714 48302 9716 48354
rect 9660 48300 9716 48302
rect 9548 47516 9604 47572
rect 7644 47346 7700 47348
rect 7644 47294 7646 47346
rect 7646 47294 7698 47346
rect 7698 47294 7700 47346
rect 7644 47292 7700 47294
rect 7756 46956 7812 47012
rect 9772 47068 9828 47124
rect 9996 48860 10052 48916
rect 12124 51490 12180 51492
rect 12124 51438 12126 51490
rect 12126 51438 12178 51490
rect 12178 51438 12180 51490
rect 12124 51436 12180 51438
rect 11116 50540 11172 50596
rect 12908 51324 12964 51380
rect 10892 50316 10948 50372
rect 11564 50316 11620 50372
rect 11788 50092 11844 50148
rect 11116 48860 11172 48916
rect 11564 48914 11620 48916
rect 11564 48862 11566 48914
rect 11566 48862 11618 48914
rect 11618 48862 11620 48914
rect 11564 48860 11620 48862
rect 10444 48802 10500 48804
rect 10444 48750 10446 48802
rect 10446 48750 10498 48802
rect 10498 48750 10500 48802
rect 10444 48748 10500 48750
rect 11676 48802 11732 48804
rect 11676 48750 11678 48802
rect 11678 48750 11730 48802
rect 11730 48750 11732 48802
rect 11676 48748 11732 48750
rect 10668 48300 10724 48356
rect 11228 48300 11284 48356
rect 9884 46508 9940 46564
rect 8316 45164 8372 45220
rect 7644 44268 7700 44324
rect 7644 44044 7700 44100
rect 7980 44044 8036 44100
rect 8204 43538 8260 43540
rect 8204 43486 8206 43538
rect 8206 43486 8258 43538
rect 8258 43486 8260 43538
rect 8204 43484 8260 43486
rect 8988 45106 9044 45108
rect 8988 45054 8990 45106
rect 8990 45054 9042 45106
rect 9042 45054 9044 45106
rect 8988 45052 9044 45054
rect 8764 44828 8820 44884
rect 8988 43484 9044 43540
rect 8540 42924 8596 42980
rect 8204 42028 8260 42084
rect 8204 41858 8260 41860
rect 8204 41806 8206 41858
rect 8206 41806 8258 41858
rect 8258 41806 8260 41858
rect 8204 41804 8260 41806
rect 8092 41692 8148 41748
rect 8204 41356 8260 41412
rect 8652 42754 8708 42756
rect 8652 42702 8654 42754
rect 8654 42702 8706 42754
rect 8706 42702 8708 42754
rect 8652 42700 8708 42702
rect 9772 44882 9828 44884
rect 9772 44830 9774 44882
rect 9774 44830 9826 44882
rect 9826 44830 9828 44882
rect 9772 44828 9828 44830
rect 12236 48914 12292 48916
rect 12236 48862 12238 48914
rect 12238 48862 12290 48914
rect 12290 48862 12292 48914
rect 12236 48860 12292 48862
rect 13916 53340 13972 53396
rect 14924 53618 14980 53620
rect 14924 53566 14926 53618
rect 14926 53566 14978 53618
rect 14978 53566 14980 53618
rect 14924 53564 14980 53566
rect 14364 53506 14420 53508
rect 14364 53454 14366 53506
rect 14366 53454 14418 53506
rect 14418 53454 14420 53506
rect 14364 53452 14420 53454
rect 15596 53506 15652 53508
rect 15596 53454 15598 53506
rect 15598 53454 15650 53506
rect 15650 53454 15652 53506
rect 15596 53452 15652 53454
rect 15036 53340 15092 53396
rect 14588 52834 14644 52836
rect 14588 52782 14590 52834
rect 14590 52782 14642 52834
rect 14642 52782 14644 52834
rect 14588 52780 14644 52782
rect 15372 52444 15428 52500
rect 15708 52946 15764 52948
rect 15708 52894 15710 52946
rect 15710 52894 15762 52946
rect 15762 52894 15764 52946
rect 15708 52892 15764 52894
rect 16044 52444 16100 52500
rect 14364 51938 14420 51940
rect 14364 51886 14366 51938
rect 14366 51886 14418 51938
rect 14418 51886 14420 51938
rect 14364 51884 14420 51886
rect 14140 51772 14196 51828
rect 13020 50034 13076 50036
rect 13020 49982 13022 50034
rect 13022 49982 13074 50034
rect 13074 49982 13076 50034
rect 13020 49980 13076 49982
rect 13244 48860 13300 48916
rect 13580 49586 13636 49588
rect 13580 49534 13582 49586
rect 13582 49534 13634 49586
rect 13634 49534 13636 49586
rect 13580 49532 13636 49534
rect 13020 48748 13076 48804
rect 12796 48636 12852 48692
rect 11788 48354 11844 48356
rect 11788 48302 11790 48354
rect 11790 48302 11842 48354
rect 11842 48302 11844 48354
rect 11788 48300 11844 48302
rect 11900 48188 11956 48244
rect 11676 47740 11732 47796
rect 11564 47458 11620 47460
rect 11564 47406 11566 47458
rect 11566 47406 11618 47458
rect 11618 47406 11620 47458
rect 11564 47404 11620 47406
rect 10332 47068 10388 47124
rect 10220 46508 10276 46564
rect 10780 46786 10836 46788
rect 10780 46734 10782 46786
rect 10782 46734 10834 46786
rect 10834 46734 10836 46786
rect 10780 46732 10836 46734
rect 11004 46786 11060 46788
rect 11004 46734 11006 46786
rect 11006 46734 11058 46786
rect 11058 46734 11060 46786
rect 11004 46732 11060 46734
rect 11452 46786 11508 46788
rect 11452 46734 11454 46786
rect 11454 46734 11506 46786
rect 11506 46734 11508 46786
rect 11452 46732 11508 46734
rect 12684 48242 12740 48244
rect 12684 48190 12686 48242
rect 12686 48190 12738 48242
rect 12738 48190 12740 48242
rect 12684 48188 12740 48190
rect 12124 47740 12180 47796
rect 12908 48354 12964 48356
rect 12908 48302 12910 48354
rect 12910 48302 12962 48354
rect 12962 48302 12964 48354
rect 12908 48300 12964 48302
rect 12124 47404 12180 47460
rect 12236 46786 12292 46788
rect 12236 46734 12238 46786
rect 12238 46734 12290 46786
rect 12290 46734 12292 46786
rect 12236 46732 12292 46734
rect 10668 46674 10724 46676
rect 10668 46622 10670 46674
rect 10670 46622 10722 46674
rect 10722 46622 10724 46674
rect 10668 46620 10724 46622
rect 10108 45164 10164 45220
rect 10668 45836 10724 45892
rect 9548 44098 9604 44100
rect 9548 44046 9550 44098
rect 9550 44046 9602 44098
rect 9602 44046 9604 44098
rect 9548 44044 9604 44046
rect 9324 43484 9380 43540
rect 9324 42754 9380 42756
rect 9324 42702 9326 42754
rect 9326 42702 9378 42754
rect 9378 42702 9380 42754
rect 9324 42700 9380 42702
rect 8988 42140 9044 42196
rect 9100 42252 9156 42308
rect 8652 41970 8708 41972
rect 8652 41918 8654 41970
rect 8654 41918 8706 41970
rect 8706 41918 8708 41970
rect 8652 41916 8708 41918
rect 9660 41804 9716 41860
rect 9212 41692 9268 41748
rect 8988 40962 9044 40964
rect 8988 40910 8990 40962
rect 8990 40910 9042 40962
rect 9042 40910 9044 40962
rect 8988 40908 9044 40910
rect 7980 40460 8036 40516
rect 7868 40402 7924 40404
rect 7868 40350 7870 40402
rect 7870 40350 7922 40402
rect 7922 40350 7924 40402
rect 7868 40348 7924 40350
rect 7308 39116 7364 39172
rect 7420 39452 7476 39508
rect 7644 39228 7700 39284
rect 8428 40236 8484 40292
rect 8316 40178 8372 40180
rect 8316 40126 8318 40178
rect 8318 40126 8370 40178
rect 8370 40126 8372 40178
rect 8316 40124 8372 40126
rect 8988 40514 9044 40516
rect 8988 40462 8990 40514
rect 8990 40462 9042 40514
rect 9042 40462 9044 40514
rect 8988 40460 9044 40462
rect 8204 39228 8260 39284
rect 8652 40236 8708 40292
rect 8316 39058 8372 39060
rect 8316 39006 8318 39058
rect 8318 39006 8370 39058
rect 8370 39006 8372 39058
rect 8316 39004 8372 39006
rect 8092 38780 8148 38836
rect 7532 38722 7588 38724
rect 7532 38670 7534 38722
rect 7534 38670 7586 38722
rect 7586 38670 7588 38722
rect 7532 38668 7588 38670
rect 5516 36540 5572 36596
rect 4732 35922 4788 35924
rect 4732 35870 4734 35922
rect 4734 35870 4786 35922
rect 4786 35870 4788 35922
rect 4732 35868 4788 35870
rect 4396 35532 4452 35588
rect 5516 35586 5572 35588
rect 5516 35534 5518 35586
rect 5518 35534 5570 35586
rect 5570 35534 5572 35586
rect 5516 35532 5572 35534
rect 4476 35306 4532 35308
rect 4476 35254 4478 35306
rect 4478 35254 4530 35306
rect 4530 35254 4532 35306
rect 4476 35252 4532 35254
rect 4580 35306 4636 35308
rect 4580 35254 4582 35306
rect 4582 35254 4634 35306
rect 4634 35254 4636 35306
rect 4580 35252 4636 35254
rect 4684 35306 4740 35308
rect 4684 35254 4686 35306
rect 4686 35254 4738 35306
rect 4738 35254 4740 35306
rect 4684 35252 4740 35254
rect 4956 34914 5012 34916
rect 4956 34862 4958 34914
rect 4958 34862 5010 34914
rect 5010 34862 5012 34914
rect 4956 34860 5012 34862
rect 4844 34690 4900 34692
rect 4844 34638 4846 34690
rect 4846 34638 4898 34690
rect 4898 34638 4900 34690
rect 4844 34636 4900 34638
rect 5068 34524 5124 34580
rect 4476 33738 4532 33740
rect 4476 33686 4478 33738
rect 4478 33686 4530 33738
rect 4530 33686 4532 33738
rect 4476 33684 4532 33686
rect 4580 33738 4636 33740
rect 4580 33686 4582 33738
rect 4582 33686 4634 33738
rect 4634 33686 4636 33738
rect 4580 33684 4636 33686
rect 4684 33738 4740 33740
rect 4684 33686 4686 33738
rect 4686 33686 4738 33738
rect 4738 33686 4740 33738
rect 4684 33684 4740 33686
rect 5068 33628 5124 33684
rect 6188 37772 6244 37828
rect 5740 36652 5796 36708
rect 5852 36540 5908 36596
rect 6524 37884 6580 37940
rect 5628 33404 5684 33460
rect 4732 33234 4788 33236
rect 4732 33182 4734 33234
rect 4734 33182 4786 33234
rect 4786 33182 4788 33234
rect 4732 33180 4788 33182
rect 3836 32562 3892 32564
rect 3836 32510 3838 32562
rect 3838 32510 3890 32562
rect 3890 32510 3892 32562
rect 3836 32508 3892 32510
rect 4060 32732 4116 32788
rect 4620 32732 4676 32788
rect 5068 32786 5124 32788
rect 5068 32734 5070 32786
rect 5070 32734 5122 32786
rect 5122 32734 5124 32786
rect 5068 32732 5124 32734
rect 4732 32508 4788 32564
rect 4956 32396 5012 32452
rect 4476 32170 4532 32172
rect 4476 32118 4478 32170
rect 4478 32118 4530 32170
rect 4530 32118 4532 32170
rect 4476 32116 4532 32118
rect 4580 32170 4636 32172
rect 4580 32118 4582 32170
rect 4582 32118 4634 32170
rect 4634 32118 4636 32170
rect 4580 32116 4636 32118
rect 4684 32170 4740 32172
rect 4684 32118 4686 32170
rect 4686 32118 4738 32170
rect 4738 32118 4740 32170
rect 4684 32116 4740 32118
rect 4284 31836 4340 31892
rect 2716 31106 2772 31108
rect 2716 31054 2718 31106
rect 2718 31054 2770 31106
rect 2770 31054 2772 31106
rect 2716 31052 2772 31054
rect 3500 31052 3556 31108
rect 2380 30828 2436 30884
rect 3276 30828 3332 30884
rect 4284 31164 4340 31220
rect 3500 30828 3556 30884
rect 4396 30828 4452 30884
rect 4508 31276 4564 31332
rect 4956 31890 5012 31892
rect 4956 31838 4958 31890
rect 4958 31838 5010 31890
rect 5010 31838 5012 31890
rect 4956 31836 5012 31838
rect 5852 34914 5908 34916
rect 5852 34862 5854 34914
rect 5854 34862 5906 34914
rect 5906 34862 5908 34914
rect 5852 34860 5908 34862
rect 7420 37938 7476 37940
rect 7420 37886 7422 37938
rect 7422 37886 7474 37938
rect 7474 37886 7476 37938
rect 7420 37884 7476 37886
rect 7196 37826 7252 37828
rect 7196 37774 7198 37826
rect 7198 37774 7250 37826
rect 7250 37774 7252 37826
rect 7196 37772 7252 37774
rect 8540 39452 8596 39508
rect 8652 39228 8708 39284
rect 7084 37660 7140 37716
rect 6636 36988 6692 37044
rect 8204 37884 8260 37940
rect 8988 39394 9044 39396
rect 8988 39342 8990 39394
rect 8990 39342 9042 39394
rect 9042 39342 9044 39394
rect 8988 39340 9044 39342
rect 9212 39004 9268 39060
rect 8988 38946 9044 38948
rect 8988 38894 8990 38946
rect 8990 38894 9042 38946
rect 9042 38894 9044 38946
rect 8988 38892 9044 38894
rect 8652 37660 8708 37716
rect 8988 37660 9044 37716
rect 7980 36988 8036 37044
rect 8652 36988 8708 37044
rect 8988 36764 9044 36820
rect 8204 36652 8260 36708
rect 5740 34412 5796 34468
rect 5740 33628 5796 33684
rect 6972 34636 7028 34692
rect 6972 34300 7028 34356
rect 6412 33516 6468 33572
rect 7196 33516 7252 33572
rect 6636 33458 6692 33460
rect 6636 33406 6638 33458
rect 6638 33406 6690 33458
rect 6690 33406 6692 33458
rect 6636 33404 6692 33406
rect 6300 33122 6356 33124
rect 6300 33070 6302 33122
rect 6302 33070 6354 33122
rect 6354 33070 6356 33122
rect 6300 33068 6356 33070
rect 7084 33122 7140 33124
rect 7084 33070 7086 33122
rect 7086 33070 7138 33122
rect 7138 33070 7140 33122
rect 7084 33068 7140 33070
rect 6412 32450 6468 32452
rect 6412 32398 6414 32450
rect 6414 32398 6466 32450
rect 6466 32398 6468 32450
rect 6412 32396 6468 32398
rect 6188 31778 6244 31780
rect 6188 31726 6190 31778
rect 6190 31726 6242 31778
rect 6242 31726 6244 31778
rect 6188 31724 6244 31726
rect 6412 31948 6468 32004
rect 7084 31724 7140 31780
rect 5180 31164 5236 31220
rect 4508 30716 4564 30772
rect 4476 30602 4532 30604
rect 4476 30550 4478 30602
rect 4478 30550 4530 30602
rect 4530 30550 4532 30602
rect 4476 30548 4532 30550
rect 4580 30602 4636 30604
rect 4580 30550 4582 30602
rect 4582 30550 4634 30602
rect 4634 30550 4636 30602
rect 4580 30548 4636 30550
rect 4684 30602 4740 30604
rect 4684 30550 4686 30602
rect 4686 30550 4738 30602
rect 4738 30550 4740 30602
rect 4684 30548 4740 30550
rect 4956 30268 5012 30324
rect 4844 29932 4900 29988
rect 4476 29034 4532 29036
rect 4476 28982 4478 29034
rect 4478 28982 4530 29034
rect 4530 28982 4532 29034
rect 4476 28980 4532 28982
rect 4580 29034 4636 29036
rect 4580 28982 4582 29034
rect 4582 28982 4634 29034
rect 4634 28982 4636 29034
rect 4580 28980 4636 28982
rect 4684 29034 4740 29036
rect 4684 28982 4686 29034
rect 4686 28982 4738 29034
rect 4738 28982 4740 29034
rect 4684 28980 4740 28982
rect 4508 28812 4564 28868
rect 4284 27916 4340 27972
rect 4620 28642 4676 28644
rect 4620 28590 4622 28642
rect 4622 28590 4674 28642
rect 4674 28590 4676 28642
rect 4620 28588 4676 28590
rect 5740 31052 5796 31108
rect 5180 29148 5236 29204
rect 2268 27580 2324 27636
rect 4476 27466 4532 27468
rect 4476 27414 4478 27466
rect 4478 27414 4530 27466
rect 4530 27414 4532 27466
rect 4476 27412 4532 27414
rect 4580 27466 4636 27468
rect 4580 27414 4582 27466
rect 4582 27414 4634 27466
rect 4634 27414 4636 27466
rect 4580 27412 4636 27414
rect 4684 27466 4740 27468
rect 4684 27414 4686 27466
rect 4686 27414 4738 27466
rect 4738 27414 4740 27466
rect 4684 27412 4740 27414
rect 5180 27804 5236 27860
rect 4844 26124 4900 26180
rect 4476 25898 4532 25900
rect 4476 25846 4478 25898
rect 4478 25846 4530 25898
rect 4530 25846 4532 25898
rect 4476 25844 4532 25846
rect 4580 25898 4636 25900
rect 4580 25846 4582 25898
rect 4582 25846 4634 25898
rect 4634 25846 4636 25898
rect 4580 25844 4636 25846
rect 4684 25898 4740 25900
rect 4684 25846 4686 25898
rect 4686 25846 4738 25898
rect 4738 25846 4740 25898
rect 4684 25844 4740 25846
rect 4732 25564 4788 25620
rect 3164 24610 3220 24612
rect 3164 24558 3166 24610
rect 3166 24558 3218 24610
rect 3218 24558 3220 24610
rect 3164 24556 3220 24558
rect 4956 25564 5012 25620
rect 5068 25394 5124 25396
rect 5068 25342 5070 25394
rect 5070 25342 5122 25394
rect 5122 25342 5124 25394
rect 5068 25340 5124 25342
rect 4508 24444 4564 24500
rect 4476 24330 4532 24332
rect 4476 24278 4478 24330
rect 4478 24278 4530 24330
rect 4530 24278 4532 24330
rect 4476 24276 4532 24278
rect 4580 24330 4636 24332
rect 4580 24278 4582 24330
rect 4582 24278 4634 24330
rect 4634 24278 4636 24330
rect 4580 24276 4636 24278
rect 4684 24330 4740 24332
rect 4684 24278 4686 24330
rect 4686 24278 4738 24330
rect 4738 24278 4740 24330
rect 4684 24276 4740 24278
rect 5516 26796 5572 26852
rect 5404 25228 5460 25284
rect 4284 23884 4340 23940
rect 3500 23042 3556 23044
rect 3500 22990 3502 23042
rect 3502 22990 3554 23042
rect 3554 22990 3556 23042
rect 3500 22988 3556 22990
rect 4476 22762 4532 22764
rect 4476 22710 4478 22762
rect 4478 22710 4530 22762
rect 4530 22710 4532 22762
rect 4476 22708 4532 22710
rect 4580 22762 4636 22764
rect 4580 22710 4582 22762
rect 4582 22710 4634 22762
rect 4634 22710 4636 22762
rect 4580 22708 4636 22710
rect 4684 22762 4740 22764
rect 4684 22710 4686 22762
rect 4686 22710 4738 22762
rect 4738 22710 4740 22762
rect 4684 22708 4740 22710
rect 2156 22092 2212 22148
rect 4956 22988 5012 23044
rect 4844 21586 4900 21588
rect 4844 21534 4846 21586
rect 4846 21534 4898 21586
rect 4898 21534 4900 21586
rect 4844 21532 4900 21534
rect 4476 21194 4532 21196
rect 4476 21142 4478 21194
rect 4478 21142 4530 21194
rect 4530 21142 4532 21194
rect 4476 21140 4532 21142
rect 4580 21194 4636 21196
rect 4580 21142 4582 21194
rect 4582 21142 4634 21194
rect 4634 21142 4636 21194
rect 4580 21140 4636 21142
rect 4684 21194 4740 21196
rect 4684 21142 4686 21194
rect 4686 21142 4738 21194
rect 4738 21142 4740 21194
rect 4684 21140 4740 21142
rect 4732 20972 4788 21028
rect 5292 23548 5348 23604
rect 5180 21532 5236 21588
rect 4844 20914 4900 20916
rect 4844 20862 4846 20914
rect 4846 20862 4898 20914
rect 4898 20862 4900 20914
rect 4844 20860 4900 20862
rect 5628 21980 5684 22036
rect 7756 34914 7812 34916
rect 7756 34862 7758 34914
rect 7758 34862 7810 34914
rect 7810 34862 7812 34914
rect 7756 34860 7812 34862
rect 7420 34802 7476 34804
rect 7420 34750 7422 34802
rect 7422 34750 7474 34802
rect 7474 34750 7476 34802
rect 7420 34748 7476 34750
rect 8316 34748 8372 34804
rect 8204 34636 8260 34692
rect 7532 34524 7588 34580
rect 7420 34354 7476 34356
rect 7420 34302 7422 34354
rect 7422 34302 7474 34354
rect 7474 34302 7476 34354
rect 7420 34300 7476 34302
rect 7644 34188 7700 34244
rect 8764 35698 8820 35700
rect 8764 35646 8766 35698
rect 8766 35646 8818 35698
rect 8818 35646 8820 35698
rect 8764 35644 8820 35646
rect 8764 34914 8820 34916
rect 8764 34862 8766 34914
rect 8766 34862 8818 34914
rect 8818 34862 8820 34914
rect 8764 34860 8820 34862
rect 8540 34524 8596 34580
rect 7756 33122 7812 33124
rect 7756 33070 7758 33122
rect 7758 33070 7810 33122
rect 7810 33070 7812 33122
rect 7756 33068 7812 33070
rect 7756 32450 7812 32452
rect 7756 32398 7758 32450
rect 7758 32398 7810 32450
rect 7810 32398 7812 32450
rect 7756 32396 7812 32398
rect 7644 31948 7700 32004
rect 7308 31890 7364 31892
rect 7308 31838 7310 31890
rect 7310 31838 7362 31890
rect 7362 31838 7364 31890
rect 7308 31836 7364 31838
rect 7532 31724 7588 31780
rect 8876 34636 8932 34692
rect 8652 33516 8708 33572
rect 8540 33404 8596 33460
rect 8988 33628 9044 33684
rect 9100 33516 9156 33572
rect 9660 40908 9716 40964
rect 9436 40124 9492 40180
rect 9548 38780 9604 38836
rect 9324 37884 9380 37940
rect 9324 35644 9380 35700
rect 9436 35196 9492 35252
rect 9660 37938 9716 37940
rect 9660 37886 9662 37938
rect 9662 37886 9714 37938
rect 9714 37886 9716 37938
rect 9660 37884 9716 37886
rect 9660 37266 9716 37268
rect 9660 37214 9662 37266
rect 9662 37214 9714 37266
rect 9714 37214 9716 37266
rect 9660 37212 9716 37214
rect 9660 35474 9716 35476
rect 9660 35422 9662 35474
rect 9662 35422 9714 35474
rect 9714 35422 9716 35474
rect 9660 35420 9716 35422
rect 11452 45836 11508 45892
rect 12684 45890 12740 45892
rect 12684 45838 12686 45890
rect 12686 45838 12738 45890
rect 12738 45838 12740 45890
rect 12684 45836 12740 45838
rect 12908 45778 12964 45780
rect 12908 45726 12910 45778
rect 12910 45726 12962 45778
rect 12962 45726 12964 45778
rect 12908 45724 12964 45726
rect 12908 45106 12964 45108
rect 12908 45054 12910 45106
rect 12910 45054 12962 45106
rect 12962 45054 12964 45106
rect 12908 45052 12964 45054
rect 11452 44044 11508 44100
rect 9996 43596 10052 43652
rect 9884 42700 9940 42756
rect 10444 43538 10500 43540
rect 10444 43486 10446 43538
rect 10446 43486 10498 43538
rect 10498 43486 10500 43538
rect 10444 43484 10500 43486
rect 10332 42924 10388 42980
rect 9996 42252 10052 42308
rect 10332 42588 10388 42644
rect 10444 42252 10500 42308
rect 9884 41244 9940 41300
rect 11228 43650 11284 43652
rect 11228 43598 11230 43650
rect 11230 43598 11282 43650
rect 11282 43598 11284 43650
rect 11228 43596 11284 43598
rect 12236 44098 12292 44100
rect 12236 44046 12238 44098
rect 12238 44046 12290 44098
rect 12290 44046 12292 44098
rect 12236 44044 12292 44046
rect 11116 42866 11172 42868
rect 11116 42814 11118 42866
rect 11118 42814 11170 42866
rect 11170 42814 11172 42866
rect 11116 42812 11172 42814
rect 10892 42140 10948 42196
rect 11116 42028 11172 42084
rect 10780 41468 10836 41524
rect 10444 41132 10500 41188
rect 9996 40908 10052 40964
rect 10780 40908 10836 40964
rect 9884 40572 9940 40628
rect 10780 40514 10836 40516
rect 10780 40462 10782 40514
rect 10782 40462 10834 40514
rect 10834 40462 10836 40514
rect 10780 40460 10836 40462
rect 10444 39506 10500 39508
rect 10444 39454 10446 39506
rect 10446 39454 10498 39506
rect 10498 39454 10500 39506
rect 10444 39452 10500 39454
rect 10220 38834 10276 38836
rect 10220 38782 10222 38834
rect 10222 38782 10274 38834
rect 10274 38782 10276 38834
rect 10220 38780 10276 38782
rect 10108 38722 10164 38724
rect 10108 38670 10110 38722
rect 10110 38670 10162 38722
rect 10162 38670 10164 38722
rect 10108 38668 10164 38670
rect 9996 37996 10052 38052
rect 10220 37772 10276 37828
rect 9884 36988 9940 37044
rect 11004 41356 11060 41412
rect 11676 42924 11732 42980
rect 11788 42588 11844 42644
rect 12684 43596 12740 43652
rect 12236 42978 12292 42980
rect 12236 42926 12238 42978
rect 12238 42926 12290 42978
rect 12290 42926 12292 42978
rect 12236 42924 12292 42926
rect 10892 39228 10948 39284
rect 11228 41186 11284 41188
rect 11228 41134 11230 41186
rect 11230 41134 11282 41186
rect 11282 41134 11284 41186
rect 11228 41132 11284 41134
rect 11116 40626 11172 40628
rect 11116 40574 11118 40626
rect 11118 40574 11170 40626
rect 11170 40574 11172 40626
rect 11116 40572 11172 40574
rect 11564 41132 11620 41188
rect 10780 38050 10836 38052
rect 10780 37998 10782 38050
rect 10782 37998 10834 38050
rect 10834 37998 10836 38050
rect 10780 37996 10836 37998
rect 10668 36988 10724 37044
rect 10556 36652 10612 36708
rect 9884 36092 9940 36148
rect 9996 36428 10052 36484
rect 9772 34972 9828 35028
rect 8764 33292 8820 33348
rect 8428 32284 8484 32340
rect 8876 32002 8932 32004
rect 8876 31950 8878 32002
rect 8878 31950 8930 32002
rect 8930 31950 8932 32002
rect 8876 31948 8932 31950
rect 7980 31836 8036 31892
rect 8316 31778 8372 31780
rect 8316 31726 8318 31778
rect 8318 31726 8370 31778
rect 8370 31726 8372 31778
rect 8316 31724 8372 31726
rect 8988 31612 9044 31668
rect 7980 31276 8036 31332
rect 8988 31218 9044 31220
rect 8988 31166 8990 31218
rect 8990 31166 9042 31218
rect 9042 31166 9044 31218
rect 8988 31164 9044 31166
rect 6972 30716 7028 30772
rect 6860 29484 6916 29540
rect 5964 29314 6020 29316
rect 5964 29262 5966 29314
rect 5966 29262 6018 29314
rect 6018 29262 6020 29314
rect 5964 29260 6020 29262
rect 8316 30770 8372 30772
rect 8316 30718 8318 30770
rect 8318 30718 8370 30770
rect 8370 30718 8372 30770
rect 8316 30716 8372 30718
rect 9212 30716 9268 30772
rect 9212 30322 9268 30324
rect 9212 30270 9214 30322
rect 9214 30270 9266 30322
rect 9266 30270 9268 30322
rect 9212 30268 9268 30270
rect 8540 30156 8596 30212
rect 7084 29484 7140 29540
rect 6748 28642 6804 28644
rect 6748 28590 6750 28642
rect 6750 28590 6802 28642
rect 6802 28590 6804 28642
rect 6748 28588 6804 28590
rect 6972 28588 7028 28644
rect 6300 26796 6356 26852
rect 5964 26236 6020 26292
rect 6412 26178 6468 26180
rect 6412 26126 6414 26178
rect 6414 26126 6466 26178
rect 6466 26126 6468 26178
rect 6412 26124 6468 26126
rect 5964 25228 6020 25284
rect 6860 26796 6916 26852
rect 5852 24444 5908 24500
rect 5964 23324 6020 23380
rect 6524 23826 6580 23828
rect 6524 23774 6526 23826
rect 6526 23774 6578 23826
rect 6578 23774 6580 23826
rect 6524 23772 6580 23774
rect 6748 25452 6804 25508
rect 6300 21532 6356 21588
rect 5516 20188 5572 20244
rect 5068 19852 5124 19908
rect 5740 19906 5796 19908
rect 5740 19854 5742 19906
rect 5742 19854 5794 19906
rect 5794 19854 5796 19906
rect 5740 19852 5796 19854
rect 4956 19740 5012 19796
rect 4476 19626 4532 19628
rect 4476 19574 4478 19626
rect 4478 19574 4530 19626
rect 4530 19574 4532 19626
rect 4476 19572 4532 19574
rect 4580 19626 4636 19628
rect 4580 19574 4582 19626
rect 4582 19574 4634 19626
rect 4634 19574 4636 19626
rect 4580 19572 4636 19574
rect 4684 19626 4740 19628
rect 4684 19574 4686 19626
rect 4686 19574 4738 19626
rect 4738 19574 4740 19626
rect 4684 19572 4740 19574
rect 1596 19404 1652 19460
rect 5740 19068 5796 19124
rect 4476 18058 4532 18060
rect 4476 18006 4478 18058
rect 4478 18006 4530 18058
rect 4530 18006 4532 18058
rect 4476 18004 4532 18006
rect 4580 18058 4636 18060
rect 4580 18006 4582 18058
rect 4582 18006 4634 18058
rect 4634 18006 4636 18058
rect 4580 18004 4636 18006
rect 4684 18058 4740 18060
rect 4684 18006 4686 18058
rect 4686 18006 4738 18058
rect 4738 18006 4740 18058
rect 4684 18004 4740 18006
rect 4476 16490 4532 16492
rect 4476 16438 4478 16490
rect 4478 16438 4530 16490
rect 4530 16438 4532 16490
rect 4476 16436 4532 16438
rect 4580 16490 4636 16492
rect 4580 16438 4582 16490
rect 4582 16438 4634 16490
rect 4634 16438 4636 16490
rect 4580 16436 4636 16438
rect 4684 16490 4740 16492
rect 4684 16438 4686 16490
rect 4686 16438 4738 16490
rect 4738 16438 4740 16490
rect 4684 16436 4740 16438
rect 6860 25340 6916 25396
rect 7756 29986 7812 29988
rect 7756 29934 7758 29986
rect 7758 29934 7810 29986
rect 7810 29934 7812 29986
rect 7756 29932 7812 29934
rect 7756 29036 7812 29092
rect 7308 28588 7364 28644
rect 8428 29314 8484 29316
rect 8428 29262 8430 29314
rect 8430 29262 8482 29314
rect 8482 29262 8484 29314
rect 8428 29260 8484 29262
rect 8988 30098 9044 30100
rect 8988 30046 8990 30098
rect 8990 30046 9042 30098
rect 9042 30046 9044 30098
rect 8988 30044 9044 30046
rect 8764 29650 8820 29652
rect 8764 29598 8766 29650
rect 8766 29598 8818 29650
rect 8818 29598 8820 29650
rect 8764 29596 8820 29598
rect 8428 28812 8484 28868
rect 7868 28476 7924 28532
rect 9660 33122 9716 33124
rect 9660 33070 9662 33122
rect 9662 33070 9714 33122
rect 9714 33070 9716 33122
rect 9660 33068 9716 33070
rect 10444 36370 10500 36372
rect 10444 36318 10446 36370
rect 10446 36318 10498 36370
rect 10498 36318 10500 36370
rect 10444 36316 10500 36318
rect 10108 35810 10164 35812
rect 10108 35758 10110 35810
rect 10110 35758 10162 35810
rect 10162 35758 10164 35810
rect 10108 35756 10164 35758
rect 10444 35474 10500 35476
rect 10444 35422 10446 35474
rect 10446 35422 10498 35474
rect 10498 35422 10500 35474
rect 10444 35420 10500 35422
rect 10332 33516 10388 33572
rect 10444 34860 10500 34916
rect 9996 33458 10052 33460
rect 9996 33406 9998 33458
rect 9998 33406 10050 33458
rect 10050 33406 10052 33458
rect 9996 33404 10052 33406
rect 9436 31948 9492 32004
rect 9436 31666 9492 31668
rect 9436 31614 9438 31666
rect 9438 31614 9490 31666
rect 9490 31614 9492 31666
rect 9436 31612 9492 31614
rect 9548 30716 9604 30772
rect 9772 32396 9828 32452
rect 9884 32060 9940 32116
rect 9884 31836 9940 31892
rect 9436 30156 9492 30212
rect 9996 29932 10052 29988
rect 9660 29538 9716 29540
rect 9660 29486 9662 29538
rect 9662 29486 9714 29538
rect 9714 29486 9716 29538
rect 9660 29484 9716 29486
rect 9548 28866 9604 28868
rect 9548 28814 9550 28866
rect 9550 28814 9602 28866
rect 9602 28814 9604 28866
rect 9548 28812 9604 28814
rect 7084 26796 7140 26852
rect 9772 28642 9828 28644
rect 9772 28590 9774 28642
rect 9774 28590 9826 28642
rect 9826 28590 9828 28642
rect 9772 28588 9828 28590
rect 9660 28364 9716 28420
rect 9436 27916 9492 27972
rect 8652 27186 8708 27188
rect 8652 27134 8654 27186
rect 8654 27134 8706 27186
rect 8706 27134 8708 27186
rect 8652 27132 8708 27134
rect 7196 26572 7252 26628
rect 8652 26572 8708 26628
rect 6748 20972 6804 21028
rect 6860 24220 6916 24276
rect 6860 22204 6916 22260
rect 7196 24220 7252 24276
rect 7420 26124 7476 26180
rect 8092 25452 8148 25508
rect 7532 22988 7588 23044
rect 6300 19964 6356 20020
rect 6748 20748 6804 20804
rect 8428 25564 8484 25620
rect 8764 26290 8820 26292
rect 8764 26238 8766 26290
rect 8766 26238 8818 26290
rect 8818 26238 8820 26290
rect 8764 26236 8820 26238
rect 8428 23884 8484 23940
rect 8652 23938 8708 23940
rect 8652 23886 8654 23938
rect 8654 23886 8706 23938
rect 8706 23886 8708 23938
rect 8652 23884 8708 23886
rect 9436 26908 9492 26964
rect 9772 27858 9828 27860
rect 9772 27806 9774 27858
rect 9774 27806 9826 27858
rect 9826 27806 9828 27858
rect 9772 27804 9828 27806
rect 9884 27692 9940 27748
rect 10108 30044 10164 30100
rect 10556 34412 10612 34468
rect 10780 36428 10836 36484
rect 11228 38162 11284 38164
rect 11228 38110 11230 38162
rect 11230 38110 11282 38162
rect 11282 38110 11284 38162
rect 11228 38108 11284 38110
rect 11004 37884 11060 37940
rect 11004 36876 11060 36932
rect 10780 35308 10836 35364
rect 10556 33628 10612 33684
rect 10780 33346 10836 33348
rect 10780 33294 10782 33346
rect 10782 33294 10834 33346
rect 10834 33294 10836 33346
rect 10780 33292 10836 33294
rect 10780 33068 10836 33124
rect 11004 35138 11060 35140
rect 11004 35086 11006 35138
rect 11006 35086 11058 35138
rect 11058 35086 11060 35138
rect 11004 35084 11060 35086
rect 11788 40460 11844 40516
rect 11788 39564 11844 39620
rect 11788 39058 11844 39060
rect 11788 39006 11790 39058
rect 11790 39006 11842 39058
rect 11842 39006 11844 39058
rect 11788 39004 11844 39006
rect 11788 38834 11844 38836
rect 11788 38782 11790 38834
rect 11790 38782 11842 38834
rect 11842 38782 11844 38834
rect 11788 38780 11844 38782
rect 11452 35196 11508 35252
rect 11788 38220 11844 38276
rect 11676 36370 11732 36372
rect 11676 36318 11678 36370
rect 11678 36318 11730 36370
rect 11730 36318 11732 36370
rect 11676 36316 11732 36318
rect 11676 36092 11732 36148
rect 11340 34748 11396 34804
rect 11116 34636 11172 34692
rect 11676 34748 11732 34804
rect 12572 41970 12628 41972
rect 12572 41918 12574 41970
rect 12574 41918 12626 41970
rect 12626 41918 12628 41970
rect 12572 41916 12628 41918
rect 13132 43314 13188 43316
rect 13132 43262 13134 43314
rect 13134 43262 13186 43314
rect 13186 43262 13188 43314
rect 13132 43260 13188 43262
rect 12572 40012 12628 40068
rect 13020 39788 13076 39844
rect 13132 40796 13188 40852
rect 12908 39730 12964 39732
rect 12908 39678 12910 39730
rect 12910 39678 12962 39730
rect 12962 39678 12964 39730
rect 12908 39676 12964 39678
rect 12236 39618 12292 39620
rect 12236 39566 12238 39618
rect 12238 39566 12290 39618
rect 12290 39566 12292 39618
rect 12236 39564 12292 39566
rect 12572 39564 12628 39620
rect 12124 38780 12180 38836
rect 11900 37996 11956 38052
rect 12012 36988 12068 37044
rect 12796 39452 12852 39508
rect 12684 38892 12740 38948
rect 12348 37884 12404 37940
rect 12460 38780 12516 38836
rect 12348 37324 12404 37380
rect 12012 36764 12068 36820
rect 12012 36540 12068 36596
rect 11900 36428 11956 36484
rect 13132 39340 13188 39396
rect 12684 38050 12740 38052
rect 12684 37998 12686 38050
rect 12686 37998 12738 38050
rect 12738 37998 12740 38050
rect 12684 37996 12740 37998
rect 13132 37772 13188 37828
rect 12572 36540 12628 36596
rect 12684 37324 12740 37380
rect 11900 35644 11956 35700
rect 11452 33852 11508 33908
rect 10892 32674 10948 32676
rect 10892 32622 10894 32674
rect 10894 32622 10946 32674
rect 10946 32622 10948 32674
rect 10892 32620 10948 32622
rect 11004 32396 11060 32452
rect 10668 31388 10724 31444
rect 10556 30940 10612 30996
rect 10780 30380 10836 30436
rect 11116 31724 11172 31780
rect 11116 31164 11172 31220
rect 11228 31500 11284 31556
rect 11116 30322 11172 30324
rect 11116 30270 11118 30322
rect 11118 30270 11170 30322
rect 11170 30270 11172 30322
rect 11116 30268 11172 30270
rect 10332 29202 10388 29204
rect 10332 29150 10334 29202
rect 10334 29150 10386 29202
rect 10386 29150 10388 29202
rect 10332 29148 10388 29150
rect 10108 28924 10164 28980
rect 9996 26908 10052 26964
rect 10108 28700 10164 28756
rect 10556 28588 10612 28644
rect 10444 28418 10500 28420
rect 10444 28366 10446 28418
rect 10446 28366 10498 28418
rect 10498 28366 10500 28418
rect 10444 28364 10500 28366
rect 10108 26514 10164 26516
rect 10108 26462 10110 26514
rect 10110 26462 10162 26514
rect 10162 26462 10164 26514
rect 10108 26460 10164 26462
rect 9324 23660 9380 23716
rect 8316 23324 8372 23380
rect 8988 23548 9044 23604
rect 8316 22988 8372 23044
rect 8876 22876 8932 22932
rect 9436 22146 9492 22148
rect 9436 22094 9438 22146
rect 9438 22094 9490 22146
rect 9490 22094 9492 22146
rect 9436 22092 9492 22094
rect 8204 21644 8260 21700
rect 9100 21308 9156 21364
rect 7980 20748 8036 20804
rect 8764 20802 8820 20804
rect 8764 20750 8766 20802
rect 8766 20750 8818 20802
rect 8818 20750 8820 20802
rect 8764 20748 8820 20750
rect 9772 25228 9828 25284
rect 11452 30210 11508 30212
rect 11452 30158 11454 30210
rect 11454 30158 11506 30210
rect 11506 30158 11508 30210
rect 11452 30156 11508 30158
rect 10892 29484 10948 29540
rect 11676 33068 11732 33124
rect 11676 32450 11732 32452
rect 11676 32398 11678 32450
rect 11678 32398 11730 32450
rect 11730 32398 11732 32450
rect 11676 32396 11732 32398
rect 12796 36316 12852 36372
rect 12236 35196 12292 35252
rect 12124 34076 12180 34132
rect 12012 33516 12068 33572
rect 12236 34860 12292 34916
rect 12460 34412 12516 34468
rect 12124 33404 12180 33460
rect 12460 33404 12516 33460
rect 12012 32508 12068 32564
rect 12348 31836 12404 31892
rect 11900 31500 11956 31556
rect 11788 31164 11844 31220
rect 12348 30828 12404 30884
rect 12012 30380 12068 30436
rect 12348 30156 12404 30212
rect 12908 33234 12964 33236
rect 12908 33182 12910 33234
rect 12910 33182 12962 33234
rect 12962 33182 12964 33234
rect 12908 33180 12964 33182
rect 13132 33964 13188 34020
rect 13132 32674 13188 32676
rect 13132 32622 13134 32674
rect 13134 32622 13186 32674
rect 13186 32622 13188 32674
rect 13132 32620 13188 32622
rect 13020 32396 13076 32452
rect 12796 30994 12852 30996
rect 12796 30942 12798 30994
rect 12798 30942 12850 30994
rect 12850 30942 12852 30994
rect 12796 30940 12852 30942
rect 13020 31724 13076 31780
rect 12684 30322 12740 30324
rect 12684 30270 12686 30322
rect 12686 30270 12738 30322
rect 12738 30270 12740 30322
rect 12684 30268 12740 30270
rect 12460 30044 12516 30100
rect 11116 29260 11172 29316
rect 11228 29148 11284 29204
rect 10892 28812 10948 28868
rect 11004 29036 11060 29092
rect 10892 27580 10948 27636
rect 10220 23884 10276 23940
rect 9996 22988 10052 23044
rect 9884 21420 9940 21476
rect 10444 25228 10500 25284
rect 11340 28530 11396 28532
rect 11340 28478 11342 28530
rect 11342 28478 11394 28530
rect 11394 28478 11396 28530
rect 11340 28476 11396 28478
rect 12012 28476 12068 28532
rect 11452 28418 11508 28420
rect 11452 28366 11454 28418
rect 11454 28366 11506 28418
rect 11506 28366 11508 28418
rect 11452 28364 11508 28366
rect 11788 27692 11844 27748
rect 12236 28924 12292 28980
rect 12572 29596 12628 29652
rect 12572 28700 12628 28756
rect 12908 28700 12964 28756
rect 12796 28476 12852 28532
rect 12236 28364 12292 28420
rect 14364 50540 14420 50596
rect 13804 50092 13860 50148
rect 13916 50034 13972 50036
rect 13916 49982 13918 50034
rect 13918 49982 13970 50034
rect 13970 49982 13972 50034
rect 13916 49980 13972 49982
rect 14252 49532 14308 49588
rect 15148 51884 15204 51940
rect 14924 50706 14980 50708
rect 14924 50654 14926 50706
rect 14926 50654 14978 50706
rect 14978 50654 14980 50706
rect 14924 50652 14980 50654
rect 15372 51772 15428 51828
rect 16492 52946 16548 52948
rect 16492 52894 16494 52946
rect 16494 52894 16546 52946
rect 16546 52894 16548 52946
rect 16492 52892 16548 52894
rect 16828 52556 16884 52612
rect 17500 52556 17556 52612
rect 16156 51772 16212 51828
rect 16604 52108 16660 52164
rect 16044 50706 16100 50708
rect 16044 50654 16046 50706
rect 16046 50654 16098 50706
rect 16098 50654 16100 50706
rect 16044 50652 16100 50654
rect 17612 52162 17668 52164
rect 17612 52110 17614 52162
rect 17614 52110 17666 52162
rect 17666 52110 17668 52162
rect 17612 52108 17668 52110
rect 18508 55916 18564 55972
rect 18284 54402 18340 54404
rect 18284 54350 18286 54402
rect 18286 54350 18338 54402
rect 18338 54350 18340 54402
rect 18284 54348 18340 54350
rect 18284 53676 18340 53732
rect 19068 54514 19124 54516
rect 19068 54462 19070 54514
rect 19070 54462 19122 54514
rect 19122 54462 19124 54514
rect 19068 54460 19124 54462
rect 18732 54402 18788 54404
rect 18732 54350 18734 54402
rect 18734 54350 18786 54402
rect 18786 54350 18788 54402
rect 18732 54348 18788 54350
rect 18956 53676 19012 53732
rect 19836 56474 19892 56476
rect 19836 56422 19838 56474
rect 19838 56422 19890 56474
rect 19890 56422 19892 56474
rect 19836 56420 19892 56422
rect 19940 56474 19996 56476
rect 19940 56422 19942 56474
rect 19942 56422 19994 56474
rect 19994 56422 19996 56474
rect 19940 56420 19996 56422
rect 20044 56474 20100 56476
rect 20044 56422 20046 56474
rect 20046 56422 20098 56474
rect 20098 56422 20100 56474
rect 20044 56420 20100 56422
rect 20860 56252 20916 56308
rect 22092 56306 22148 56308
rect 22092 56254 22094 56306
rect 22094 56254 22146 56306
rect 22146 56254 22148 56306
rect 22092 56252 22148 56254
rect 22428 56140 22484 56196
rect 25564 56252 25620 56308
rect 27468 56306 27524 56308
rect 27468 56254 27470 56306
rect 27470 56254 27522 56306
rect 27522 56254 27524 56306
rect 27468 56252 27524 56254
rect 25340 56194 25396 56196
rect 25340 56142 25342 56194
rect 25342 56142 25394 56194
rect 25394 56142 25396 56194
rect 25340 56140 25396 56142
rect 21868 55186 21924 55188
rect 21868 55134 21870 55186
rect 21870 55134 21922 55186
rect 21922 55134 21924 55186
rect 21868 55132 21924 55134
rect 15372 50594 15428 50596
rect 15372 50542 15374 50594
rect 15374 50542 15426 50594
rect 15426 50542 15428 50594
rect 15372 50540 15428 50542
rect 15036 50034 15092 50036
rect 15036 49982 15038 50034
rect 15038 49982 15090 50034
rect 15090 49982 15092 50034
rect 15036 49980 15092 49982
rect 15708 48748 15764 48804
rect 15708 48412 15764 48468
rect 16380 48412 16436 48468
rect 16716 48860 16772 48916
rect 16828 48466 16884 48468
rect 16828 48414 16830 48466
rect 16830 48414 16882 48466
rect 16882 48414 16884 48466
rect 16828 48412 16884 48414
rect 13692 47068 13748 47124
rect 13580 45890 13636 45892
rect 13580 45838 13582 45890
rect 13582 45838 13634 45890
rect 13634 45838 13636 45890
rect 13580 45836 13636 45838
rect 16044 47516 16100 47572
rect 14364 46844 14420 46900
rect 13916 45724 13972 45780
rect 15932 46898 15988 46900
rect 15932 46846 15934 46898
rect 15934 46846 15986 46898
rect 15986 46846 15988 46898
rect 15932 46844 15988 46846
rect 13580 45052 13636 45108
rect 14476 45052 14532 45108
rect 13356 41858 13412 41860
rect 13356 41806 13358 41858
rect 13358 41806 13410 41858
rect 13410 41806 13412 41858
rect 13356 41804 13412 41806
rect 13580 40572 13636 40628
rect 13468 40460 13524 40516
rect 13356 39452 13412 39508
rect 13356 39004 13412 39060
rect 15148 46674 15204 46676
rect 15148 46622 15150 46674
rect 15150 46622 15202 46674
rect 15202 46622 15204 46674
rect 15148 46620 15204 46622
rect 15036 46002 15092 46004
rect 15036 45950 15038 46002
rect 15038 45950 15090 46002
rect 15090 45950 15092 46002
rect 15036 45948 15092 45950
rect 15148 45276 15204 45332
rect 15596 46620 15652 46676
rect 15820 46620 15876 46676
rect 15596 45890 15652 45892
rect 15596 45838 15598 45890
rect 15598 45838 15650 45890
rect 15650 45838 15652 45890
rect 15596 45836 15652 45838
rect 15372 45052 15428 45108
rect 15932 45052 15988 45108
rect 14700 43372 14756 43428
rect 16268 45276 16324 45332
rect 16492 45836 16548 45892
rect 15372 43650 15428 43652
rect 15372 43598 15374 43650
rect 15374 43598 15426 43650
rect 15426 43598 15428 43650
rect 15372 43596 15428 43598
rect 14924 43148 14980 43204
rect 15036 43484 15092 43540
rect 14700 42754 14756 42756
rect 14700 42702 14702 42754
rect 14702 42702 14754 42754
rect 14754 42702 14756 42754
rect 14700 42700 14756 42702
rect 15708 43538 15764 43540
rect 15708 43486 15710 43538
rect 15710 43486 15762 43538
rect 15762 43486 15764 43538
rect 15708 43484 15764 43486
rect 14812 42530 14868 42532
rect 14812 42478 14814 42530
rect 14814 42478 14866 42530
rect 14866 42478 14868 42530
rect 14812 42476 14868 42478
rect 16940 46620 16996 46676
rect 16716 45276 16772 45332
rect 16828 45106 16884 45108
rect 16828 45054 16830 45106
rect 16830 45054 16882 45106
rect 16882 45054 16884 45106
rect 16828 45052 16884 45054
rect 16268 43538 16324 43540
rect 16268 43486 16270 43538
rect 16270 43486 16322 43538
rect 16322 43486 16324 43538
rect 16268 43484 16324 43486
rect 16268 42476 16324 42532
rect 15148 41804 15204 41860
rect 14476 41356 14532 41412
rect 13804 41186 13860 41188
rect 13804 41134 13806 41186
rect 13806 41134 13858 41186
rect 13858 41134 13860 41186
rect 13804 41132 13860 41134
rect 15036 41244 15092 41300
rect 15260 41580 15316 41636
rect 15260 41244 15316 41300
rect 15260 40908 15316 40964
rect 16492 42754 16548 42756
rect 16492 42702 16494 42754
rect 16494 42702 16546 42754
rect 16546 42702 16548 42754
rect 16492 42700 16548 42702
rect 15820 41580 15876 41636
rect 14140 40796 14196 40852
rect 14028 40684 14084 40740
rect 15932 40962 15988 40964
rect 15932 40910 15934 40962
rect 15934 40910 15986 40962
rect 15986 40910 15988 40962
rect 15932 40908 15988 40910
rect 15372 40460 15428 40516
rect 16156 40460 16212 40516
rect 16716 43596 16772 43652
rect 16828 43148 16884 43204
rect 16716 41858 16772 41860
rect 16716 41806 16718 41858
rect 16718 41806 16770 41858
rect 16770 41806 16772 41858
rect 16716 41804 16772 41806
rect 16492 41468 16548 41524
rect 14028 39788 14084 39844
rect 13692 39340 13748 39396
rect 13692 38834 13748 38836
rect 13692 38782 13694 38834
rect 13694 38782 13746 38834
rect 13746 38782 13748 38834
rect 13692 38780 13748 38782
rect 14028 39618 14084 39620
rect 14028 39566 14030 39618
rect 14030 39566 14082 39618
rect 14082 39566 14084 39618
rect 14028 39564 14084 39566
rect 14028 39058 14084 39060
rect 14028 39006 14030 39058
rect 14030 39006 14082 39058
rect 14082 39006 14084 39058
rect 14028 39004 14084 39006
rect 13804 38556 13860 38612
rect 13692 38108 13748 38164
rect 13580 37996 13636 38052
rect 14252 38050 14308 38052
rect 14252 37998 14254 38050
rect 14254 37998 14306 38050
rect 14306 37998 14308 38050
rect 14252 37996 14308 37998
rect 13692 37938 13748 37940
rect 13692 37886 13694 37938
rect 13694 37886 13746 37938
rect 13746 37886 13748 37938
rect 13692 37884 13748 37886
rect 13580 36482 13636 36484
rect 13580 36430 13582 36482
rect 13582 36430 13634 36482
rect 13634 36430 13636 36482
rect 13580 36428 13636 36430
rect 15596 40348 15652 40404
rect 14812 38556 14868 38612
rect 15148 38556 15204 38612
rect 15372 39618 15428 39620
rect 15372 39566 15374 39618
rect 15374 39566 15426 39618
rect 15426 39566 15428 39618
rect 15372 39564 15428 39566
rect 15484 39506 15540 39508
rect 15484 39454 15486 39506
rect 15486 39454 15538 39506
rect 15538 39454 15540 39506
rect 15484 39452 15540 39454
rect 15372 39340 15428 39396
rect 15372 38892 15428 38948
rect 15820 39564 15876 39620
rect 16044 39340 16100 39396
rect 15820 39116 15876 39172
rect 13580 34860 13636 34916
rect 13804 35532 13860 35588
rect 13468 34412 13524 34468
rect 13804 34914 13860 34916
rect 13804 34862 13806 34914
rect 13806 34862 13858 34914
rect 13858 34862 13860 34914
rect 13804 34860 13860 34862
rect 13916 34748 13972 34804
rect 13468 34018 13524 34020
rect 13468 33966 13470 34018
rect 13470 33966 13522 34018
rect 13522 33966 13524 34018
rect 13468 33964 13524 33966
rect 14252 35698 14308 35700
rect 14252 35646 14254 35698
rect 14254 35646 14306 35698
rect 14306 35646 14308 35698
rect 14252 35644 14308 35646
rect 15148 37378 15204 37380
rect 15148 37326 15150 37378
rect 15150 37326 15202 37378
rect 15202 37326 15204 37378
rect 15148 37324 15204 37326
rect 14700 37266 14756 37268
rect 14700 37214 14702 37266
rect 14702 37214 14754 37266
rect 14754 37214 14756 37266
rect 14700 37212 14756 37214
rect 15372 37266 15428 37268
rect 15372 37214 15374 37266
rect 15374 37214 15426 37266
rect 15426 37214 15428 37266
rect 15372 37212 15428 37214
rect 16380 38668 16436 38724
rect 16604 39900 16660 39956
rect 16156 38050 16212 38052
rect 16156 37998 16158 38050
rect 16158 37998 16210 38050
rect 16210 37998 16212 38050
rect 16156 37996 16212 37998
rect 16604 37996 16660 38052
rect 16044 36988 16100 37044
rect 15708 35868 15764 35924
rect 15372 35420 15428 35476
rect 15260 35308 15316 35364
rect 15260 34972 15316 35028
rect 14140 34188 14196 34244
rect 14028 34076 14084 34132
rect 14140 33964 14196 34020
rect 14028 33740 14084 33796
rect 13804 33292 13860 33348
rect 13916 33516 13972 33572
rect 14028 33122 14084 33124
rect 14028 33070 14030 33122
rect 14030 33070 14082 33122
rect 14082 33070 14084 33122
rect 14028 33068 14084 33070
rect 13692 32284 13748 32340
rect 13356 31724 13412 31780
rect 13580 31836 13636 31892
rect 13468 31388 13524 31444
rect 13692 30940 13748 30996
rect 13916 32396 13972 32452
rect 13580 30380 13636 30436
rect 13804 30268 13860 30324
rect 13692 30210 13748 30212
rect 13692 30158 13694 30210
rect 13694 30158 13746 30210
rect 13746 30158 13748 30210
rect 13692 30156 13748 30158
rect 14364 33180 14420 33236
rect 14476 33852 14532 33908
rect 14364 31890 14420 31892
rect 14364 31838 14366 31890
rect 14366 31838 14418 31890
rect 14418 31838 14420 31890
rect 14364 31836 14420 31838
rect 14252 31612 14308 31668
rect 13916 29260 13972 29316
rect 12124 27244 12180 27300
rect 13804 27298 13860 27300
rect 13804 27246 13806 27298
rect 13806 27246 13858 27298
rect 13858 27246 13860 27298
rect 13804 27244 13860 27246
rect 14140 29372 14196 29428
rect 14140 28754 14196 28756
rect 14140 28702 14142 28754
rect 14142 28702 14194 28754
rect 14194 28702 14196 28754
rect 14140 28700 14196 28702
rect 11004 23996 11060 24052
rect 11340 23996 11396 24052
rect 11228 23100 11284 23156
rect 10332 22258 10388 22260
rect 10332 22206 10334 22258
rect 10334 22206 10386 22258
rect 10386 22206 10388 22258
rect 10332 22204 10388 22206
rect 10332 21980 10388 22036
rect 11116 22540 11172 22596
rect 11004 22092 11060 22148
rect 11228 22204 11284 22260
rect 11116 21980 11172 22036
rect 10444 21644 10500 21700
rect 9996 20860 10052 20916
rect 9548 20636 9604 20692
rect 9772 20188 9828 20244
rect 8652 20018 8708 20020
rect 8652 19966 8654 20018
rect 8654 19966 8706 20018
rect 8706 19966 8708 20018
rect 8652 19964 8708 19966
rect 6748 19740 6804 19796
rect 7868 19292 7924 19348
rect 7308 19234 7364 19236
rect 7308 19182 7310 19234
rect 7310 19182 7362 19234
rect 7362 19182 7364 19234
rect 7308 19180 7364 19182
rect 8316 19180 8372 19236
rect 9772 19794 9828 19796
rect 9772 19742 9774 19794
rect 9774 19742 9826 19794
rect 9826 19742 9828 19794
rect 9772 19740 9828 19742
rect 9548 19068 9604 19124
rect 8876 18674 8932 18676
rect 8876 18622 8878 18674
rect 8878 18622 8930 18674
rect 8930 18622 8932 18674
rect 8876 18620 8932 18622
rect 10668 21084 10724 21140
rect 10780 20972 10836 21028
rect 10668 20748 10724 20804
rect 10668 20018 10724 20020
rect 10668 19966 10670 20018
rect 10670 19966 10722 20018
rect 10722 19966 10724 20018
rect 10668 19964 10724 19966
rect 11116 21586 11172 21588
rect 11116 21534 11118 21586
rect 11118 21534 11170 21586
rect 11170 21534 11172 21586
rect 11116 21532 11172 21534
rect 11116 21196 11172 21252
rect 11004 20188 11060 20244
rect 11676 26460 11732 26516
rect 11788 25506 11844 25508
rect 11788 25454 11790 25506
rect 11790 25454 11842 25506
rect 11842 25454 11844 25506
rect 11788 25452 11844 25454
rect 11452 23548 11508 23604
rect 11452 21586 11508 21588
rect 11452 21534 11454 21586
rect 11454 21534 11506 21586
rect 11506 21534 11508 21586
rect 11452 21532 11508 21534
rect 12124 23884 12180 23940
rect 12348 23938 12404 23940
rect 12348 23886 12350 23938
rect 12350 23886 12402 23938
rect 12402 23886 12404 23938
rect 12348 23884 12404 23886
rect 11676 22876 11732 22932
rect 11788 23436 11844 23492
rect 11676 21698 11732 21700
rect 11676 21646 11678 21698
rect 11678 21646 11730 21698
rect 11730 21646 11732 21698
rect 11676 21644 11732 21646
rect 11452 21084 11508 21140
rect 11564 20690 11620 20692
rect 11564 20638 11566 20690
rect 11566 20638 11618 20690
rect 11618 20638 11620 20690
rect 11564 20636 11620 20638
rect 12124 23324 12180 23380
rect 12236 23212 12292 23268
rect 12908 26348 12964 26404
rect 12796 24162 12852 24164
rect 12796 24110 12798 24162
rect 12798 24110 12850 24162
rect 12850 24110 12852 24162
rect 12796 24108 12852 24110
rect 13132 26236 13188 26292
rect 12684 23548 12740 23604
rect 12572 23154 12628 23156
rect 12572 23102 12574 23154
rect 12574 23102 12626 23154
rect 12626 23102 12628 23154
rect 12572 23100 12628 23102
rect 12684 22988 12740 23044
rect 12796 23324 12852 23380
rect 12348 22258 12404 22260
rect 12348 22206 12350 22258
rect 12350 22206 12402 22258
rect 12402 22206 12404 22258
rect 12348 22204 12404 22206
rect 12572 21532 12628 21588
rect 11676 20300 11732 20356
rect 10892 19628 10948 19684
rect 10220 19180 10276 19236
rect 11452 19628 11508 19684
rect 11116 18956 11172 19012
rect 10892 17666 10948 17668
rect 10892 17614 10894 17666
rect 10894 17614 10946 17666
rect 10946 17614 10948 17666
rect 10892 17612 10948 17614
rect 11452 18620 11508 18676
rect 12012 20130 12068 20132
rect 12012 20078 12014 20130
rect 12014 20078 12066 20130
rect 12066 20078 12068 20130
rect 12012 20076 12068 20078
rect 12908 22428 12964 22484
rect 13132 22316 13188 22372
rect 13916 26908 13972 26964
rect 13692 25506 13748 25508
rect 13692 25454 13694 25506
rect 13694 25454 13746 25506
rect 13746 25454 13748 25506
rect 13692 25452 13748 25454
rect 13804 25228 13860 25284
rect 13804 24610 13860 24612
rect 13804 24558 13806 24610
rect 13806 24558 13858 24610
rect 13858 24558 13860 24610
rect 13804 24556 13860 24558
rect 13692 24220 13748 24276
rect 15036 33740 15092 33796
rect 15372 34802 15428 34804
rect 15372 34750 15374 34802
rect 15374 34750 15426 34802
rect 15426 34750 15428 34802
rect 15372 34748 15428 34750
rect 15260 34130 15316 34132
rect 15260 34078 15262 34130
rect 15262 34078 15314 34130
rect 15314 34078 15316 34130
rect 15260 34076 15316 34078
rect 15148 33628 15204 33684
rect 15260 33346 15316 33348
rect 15260 33294 15262 33346
rect 15262 33294 15314 33346
rect 15314 33294 15316 33346
rect 15260 33292 15316 33294
rect 14700 32620 14756 32676
rect 14588 31724 14644 31780
rect 15148 32508 15204 32564
rect 14924 31388 14980 31444
rect 15036 31276 15092 31332
rect 14588 29932 14644 29988
rect 14700 30268 14756 30324
rect 14924 30098 14980 30100
rect 14924 30046 14926 30098
rect 14926 30046 14978 30098
rect 14978 30046 14980 30098
rect 14924 30044 14980 30046
rect 14700 29596 14756 29652
rect 14476 29036 14532 29092
rect 14700 28364 14756 28420
rect 14252 26348 14308 26404
rect 14700 26290 14756 26292
rect 14700 26238 14702 26290
rect 14702 26238 14754 26290
rect 14754 26238 14756 26290
rect 14700 26236 14756 26238
rect 14364 26124 14420 26180
rect 14924 29314 14980 29316
rect 14924 29262 14926 29314
rect 14926 29262 14978 29314
rect 14978 29262 14980 29314
rect 14924 29260 14980 29262
rect 15148 30828 15204 30884
rect 15820 35532 15876 35588
rect 16156 35196 16212 35252
rect 15596 34636 15652 34692
rect 15708 34300 15764 34356
rect 16156 34300 16212 34356
rect 16716 37324 16772 37380
rect 16828 36988 16884 37044
rect 16604 36876 16660 36932
rect 17500 48972 17556 49028
rect 18060 48914 18116 48916
rect 18060 48862 18062 48914
rect 18062 48862 18114 48914
rect 18114 48862 18116 48914
rect 18060 48860 18116 48862
rect 18284 48748 18340 48804
rect 17612 47964 17668 48020
rect 17388 47516 17444 47572
rect 19292 53116 19348 53172
rect 19836 54906 19892 54908
rect 19836 54854 19838 54906
rect 19838 54854 19890 54906
rect 19890 54854 19892 54906
rect 19836 54852 19892 54854
rect 19940 54906 19996 54908
rect 19940 54854 19942 54906
rect 19942 54854 19994 54906
rect 19994 54854 19996 54906
rect 19940 54852 19996 54854
rect 20044 54906 20100 54908
rect 20044 54854 20046 54906
rect 20046 54854 20098 54906
rect 20098 54854 20100 54906
rect 20044 54852 20100 54854
rect 22540 55074 22596 55076
rect 22540 55022 22542 55074
rect 22542 55022 22594 55074
rect 22594 55022 22596 55074
rect 22540 55020 22596 55022
rect 25788 55356 25844 55412
rect 19852 53900 19908 53956
rect 21868 54348 21924 54404
rect 22204 54012 22260 54068
rect 21644 53564 21700 53620
rect 20972 53452 21028 53508
rect 19836 53338 19892 53340
rect 19836 53286 19838 53338
rect 19838 53286 19890 53338
rect 19890 53286 19892 53338
rect 19836 53284 19892 53286
rect 19940 53338 19996 53340
rect 19940 53286 19942 53338
rect 19942 53286 19994 53338
rect 19994 53286 19996 53338
rect 19940 53284 19996 53286
rect 20044 53338 20100 53340
rect 20044 53286 20046 53338
rect 20046 53286 20098 53338
rect 20098 53286 20100 53338
rect 20044 53284 20100 53286
rect 20524 53170 20580 53172
rect 20524 53118 20526 53170
rect 20526 53118 20578 53170
rect 20578 53118 20580 53170
rect 20524 53116 20580 53118
rect 18732 51212 18788 51268
rect 19180 50988 19236 51044
rect 19740 51884 19796 51940
rect 19836 51770 19892 51772
rect 19836 51718 19838 51770
rect 19838 51718 19890 51770
rect 19890 51718 19892 51770
rect 19836 51716 19892 51718
rect 19940 51770 19996 51772
rect 19940 51718 19942 51770
rect 19942 51718 19994 51770
rect 19994 51718 19996 51770
rect 19940 51716 19996 51718
rect 20044 51770 20100 51772
rect 20044 51718 20046 51770
rect 20046 51718 20098 51770
rect 20098 51718 20100 51770
rect 20044 51716 20100 51718
rect 20076 51436 20132 51492
rect 20412 51884 20468 51940
rect 20300 50988 20356 51044
rect 20860 51490 20916 51492
rect 20860 51438 20862 51490
rect 20862 51438 20914 51490
rect 20914 51438 20916 51490
rect 20860 51436 20916 51438
rect 20636 51266 20692 51268
rect 20636 51214 20638 51266
rect 20638 51214 20690 51266
rect 20690 51214 20692 51266
rect 20636 51212 20692 51214
rect 18732 50316 18788 50372
rect 18732 49026 18788 49028
rect 18732 48974 18734 49026
rect 18734 48974 18786 49026
rect 18786 48974 18788 49026
rect 18732 48972 18788 48974
rect 18620 48076 18676 48132
rect 17388 47068 17444 47124
rect 20524 50370 20580 50372
rect 20524 50318 20526 50370
rect 20526 50318 20578 50370
rect 20578 50318 20580 50370
rect 20524 50316 20580 50318
rect 19836 50202 19892 50204
rect 19836 50150 19838 50202
rect 19838 50150 19890 50202
rect 19890 50150 19892 50202
rect 19836 50148 19892 50150
rect 19940 50202 19996 50204
rect 19940 50150 19942 50202
rect 19942 50150 19994 50202
rect 19994 50150 19996 50202
rect 19940 50148 19996 50150
rect 20044 50202 20100 50204
rect 20044 50150 20046 50202
rect 20046 50150 20098 50202
rect 20098 50150 20100 50202
rect 20044 50148 20100 50150
rect 20300 48914 20356 48916
rect 20300 48862 20302 48914
rect 20302 48862 20354 48914
rect 20354 48862 20356 48914
rect 20300 48860 20356 48862
rect 19740 48802 19796 48804
rect 19740 48750 19742 48802
rect 19742 48750 19794 48802
rect 19794 48750 19796 48802
rect 19740 48748 19796 48750
rect 20412 48802 20468 48804
rect 20412 48750 20414 48802
rect 20414 48750 20466 48802
rect 20466 48750 20468 48802
rect 20412 48748 20468 48750
rect 19836 48634 19892 48636
rect 19836 48582 19838 48634
rect 19838 48582 19890 48634
rect 19890 48582 19892 48634
rect 19836 48580 19892 48582
rect 19940 48634 19996 48636
rect 19940 48582 19942 48634
rect 19942 48582 19994 48634
rect 19994 48582 19996 48634
rect 19940 48580 19996 48582
rect 20044 48634 20100 48636
rect 20044 48582 20046 48634
rect 20046 48582 20098 48634
rect 20098 48582 20100 48634
rect 20044 48580 20100 48582
rect 20300 48300 20356 48356
rect 20076 47458 20132 47460
rect 20076 47406 20078 47458
rect 20078 47406 20130 47458
rect 20130 47406 20132 47458
rect 20076 47404 20132 47406
rect 19836 47066 19892 47068
rect 19836 47014 19838 47066
rect 19838 47014 19890 47066
rect 19890 47014 19892 47066
rect 19836 47012 19892 47014
rect 19940 47066 19996 47068
rect 19940 47014 19942 47066
rect 19942 47014 19994 47066
rect 19994 47014 19996 47066
rect 19940 47012 19996 47014
rect 20044 47066 20100 47068
rect 20044 47014 20046 47066
rect 20046 47014 20098 47066
rect 20098 47014 20100 47066
rect 20044 47012 20100 47014
rect 20636 48130 20692 48132
rect 20636 48078 20638 48130
rect 20638 48078 20690 48130
rect 20690 48078 20692 48130
rect 20636 48076 20692 48078
rect 20860 47404 20916 47460
rect 22092 53618 22148 53620
rect 22092 53566 22094 53618
rect 22094 53566 22146 53618
rect 22146 53566 22148 53618
rect 22092 53564 22148 53566
rect 22988 53954 23044 53956
rect 22988 53902 22990 53954
rect 22990 53902 23042 53954
rect 23042 53902 23044 53954
rect 22988 53900 23044 53902
rect 23100 53788 23156 53844
rect 21644 52556 21700 52612
rect 21756 52892 21812 52948
rect 21308 51938 21364 51940
rect 21308 51886 21310 51938
rect 21310 51886 21362 51938
rect 21362 51886 21364 51938
rect 21308 51884 21364 51886
rect 21644 51938 21700 51940
rect 21644 51886 21646 51938
rect 21646 51886 21698 51938
rect 21698 51886 21700 51938
rect 21644 51884 21700 51886
rect 21308 51548 21364 51604
rect 21196 50764 21252 50820
rect 20972 46844 21028 46900
rect 17500 44044 17556 44100
rect 17948 44380 18004 44436
rect 17836 42082 17892 42084
rect 17836 42030 17838 42082
rect 17838 42030 17890 42082
rect 17890 42030 17892 42082
rect 17836 42028 17892 42030
rect 18620 46450 18676 46452
rect 18620 46398 18622 46450
rect 18622 46398 18674 46450
rect 18674 46398 18676 46450
rect 18620 46396 18676 46398
rect 18396 45724 18452 45780
rect 19292 45890 19348 45892
rect 19292 45838 19294 45890
rect 19294 45838 19346 45890
rect 19346 45838 19348 45890
rect 19292 45836 19348 45838
rect 21084 47964 21140 48020
rect 20188 46396 20244 46452
rect 20412 45836 20468 45892
rect 20188 45612 20244 45668
rect 20300 45778 20356 45780
rect 20300 45726 20302 45778
rect 20302 45726 20354 45778
rect 20354 45726 20356 45778
rect 20300 45724 20356 45726
rect 19836 45498 19892 45500
rect 19836 45446 19838 45498
rect 19838 45446 19890 45498
rect 19890 45446 19892 45498
rect 19836 45444 19892 45446
rect 19940 45498 19996 45500
rect 19940 45446 19942 45498
rect 19942 45446 19994 45498
rect 19994 45446 19996 45498
rect 19940 45444 19996 45446
rect 20044 45498 20100 45500
rect 20044 45446 20046 45498
rect 20046 45446 20098 45498
rect 20098 45446 20100 45498
rect 20044 45444 20100 45446
rect 19180 45052 19236 45108
rect 18620 44380 18676 44436
rect 20412 45388 20468 45444
rect 21420 51100 21476 51156
rect 22428 52946 22484 52948
rect 22428 52894 22430 52946
rect 22430 52894 22482 52946
rect 22482 52894 22484 52946
rect 22428 52892 22484 52894
rect 23100 53506 23156 53508
rect 23100 53454 23102 53506
rect 23102 53454 23154 53506
rect 23154 53454 23156 53506
rect 23100 53452 23156 53454
rect 23772 55186 23828 55188
rect 23772 55134 23774 55186
rect 23774 55134 23826 55186
rect 23826 55134 23828 55186
rect 23772 55132 23828 55134
rect 23660 55074 23716 55076
rect 23660 55022 23662 55074
rect 23662 55022 23714 55074
rect 23714 55022 23716 55074
rect 23660 55020 23716 55022
rect 23436 54460 23492 54516
rect 23324 54236 23380 54292
rect 23884 54514 23940 54516
rect 23884 54462 23886 54514
rect 23886 54462 23938 54514
rect 23938 54462 23940 54514
rect 23884 54460 23940 54462
rect 22092 51884 22148 51940
rect 21980 51548 22036 51604
rect 21868 51100 21924 51156
rect 21980 50876 22036 50932
rect 21644 47458 21700 47460
rect 21644 47406 21646 47458
rect 21646 47406 21698 47458
rect 21698 47406 21700 47458
rect 21644 47404 21700 47406
rect 21420 46620 21476 46676
rect 21308 46508 21364 46564
rect 21308 45948 21364 46004
rect 21868 45724 21924 45780
rect 21084 45052 21140 45108
rect 21196 45388 21252 45444
rect 19852 44434 19908 44436
rect 19852 44382 19854 44434
rect 19854 44382 19906 44434
rect 19906 44382 19908 44434
rect 19852 44380 19908 44382
rect 19292 44156 19348 44212
rect 18284 43708 18340 43764
rect 19404 44098 19460 44100
rect 19404 44046 19406 44098
rect 19406 44046 19458 44098
rect 19458 44046 19460 44098
rect 19404 44044 19460 44046
rect 19836 43930 19892 43932
rect 19836 43878 19838 43930
rect 19838 43878 19890 43930
rect 19890 43878 19892 43930
rect 19836 43876 19892 43878
rect 19940 43930 19996 43932
rect 19940 43878 19942 43930
rect 19942 43878 19994 43930
rect 19994 43878 19996 43930
rect 19940 43876 19996 43878
rect 20044 43930 20100 43932
rect 20044 43878 20046 43930
rect 20046 43878 20098 43930
rect 20098 43878 20100 43930
rect 20044 43876 20100 43878
rect 20300 44098 20356 44100
rect 20300 44046 20302 44098
rect 20302 44046 20354 44098
rect 20354 44046 20356 44098
rect 20300 44044 20356 44046
rect 20748 44156 20804 44212
rect 20188 43596 20244 43652
rect 20300 43708 20356 43764
rect 18508 42588 18564 42644
rect 19292 42642 19348 42644
rect 19292 42590 19294 42642
rect 19294 42590 19346 42642
rect 19346 42590 19348 42642
rect 19292 42588 19348 42590
rect 19068 42082 19124 42084
rect 19068 42030 19070 42082
rect 19070 42030 19122 42082
rect 19122 42030 19124 42082
rect 19068 42028 19124 42030
rect 17612 41746 17668 41748
rect 17612 41694 17614 41746
rect 17614 41694 17666 41746
rect 17666 41694 17668 41746
rect 17612 41692 17668 41694
rect 17164 39004 17220 39060
rect 17612 40514 17668 40516
rect 17612 40462 17614 40514
rect 17614 40462 17666 40514
rect 17666 40462 17668 40514
rect 17612 40460 17668 40462
rect 17948 41020 18004 41076
rect 17612 39394 17668 39396
rect 17612 39342 17614 39394
rect 17614 39342 17666 39394
rect 17666 39342 17668 39394
rect 17612 39340 17668 39342
rect 17388 38892 17444 38948
rect 17948 40012 18004 40068
rect 17948 39228 18004 39284
rect 17948 39058 18004 39060
rect 17948 39006 17950 39058
rect 17950 39006 18002 39058
rect 18002 39006 18004 39058
rect 17948 39004 18004 39006
rect 20860 42754 20916 42756
rect 20860 42702 20862 42754
rect 20862 42702 20914 42754
rect 20914 42702 20916 42754
rect 20860 42700 20916 42702
rect 20524 42642 20580 42644
rect 20524 42590 20526 42642
rect 20526 42590 20578 42642
rect 20578 42590 20580 42642
rect 20524 42588 20580 42590
rect 20748 42588 20804 42644
rect 19836 42362 19892 42364
rect 19836 42310 19838 42362
rect 19838 42310 19890 42362
rect 19890 42310 19892 42362
rect 19836 42308 19892 42310
rect 19940 42362 19996 42364
rect 19940 42310 19942 42362
rect 19942 42310 19994 42362
rect 19994 42310 19996 42362
rect 19940 42308 19996 42310
rect 20044 42362 20100 42364
rect 20044 42310 20046 42362
rect 20046 42310 20098 42362
rect 20098 42310 20100 42362
rect 20044 42308 20100 42310
rect 20524 42028 20580 42084
rect 18396 41020 18452 41076
rect 19180 41692 19236 41748
rect 19180 40908 19236 40964
rect 20636 41916 20692 41972
rect 19628 40962 19684 40964
rect 19628 40910 19630 40962
rect 19630 40910 19682 40962
rect 19682 40910 19684 40962
rect 19628 40908 19684 40910
rect 20524 40908 20580 40964
rect 19836 40794 19892 40796
rect 19836 40742 19838 40794
rect 19838 40742 19890 40794
rect 19890 40742 19892 40794
rect 19836 40740 19892 40742
rect 19940 40794 19996 40796
rect 19940 40742 19942 40794
rect 19942 40742 19994 40794
rect 19994 40742 19996 40794
rect 19940 40740 19996 40742
rect 20044 40794 20100 40796
rect 20044 40742 20046 40794
rect 20046 40742 20098 40794
rect 20098 40742 20100 40794
rect 20044 40740 20100 40742
rect 19404 40348 19460 40404
rect 19516 40012 19572 40068
rect 21756 45106 21812 45108
rect 21756 45054 21758 45106
rect 21758 45054 21810 45106
rect 21810 45054 21812 45106
rect 21756 45052 21812 45054
rect 22204 50988 22260 51044
rect 22092 50818 22148 50820
rect 22092 50766 22094 50818
rect 22094 50766 22146 50818
rect 22146 50766 22148 50818
rect 22092 50764 22148 50766
rect 22652 52162 22708 52164
rect 22652 52110 22654 52162
rect 22654 52110 22706 52162
rect 22706 52110 22708 52162
rect 22652 52108 22708 52110
rect 22540 51212 22596 51268
rect 22764 51212 22820 51268
rect 22876 51938 22932 51940
rect 22876 51886 22878 51938
rect 22878 51886 22930 51938
rect 22930 51886 22932 51938
rect 22876 51884 22932 51886
rect 23548 52162 23604 52164
rect 23548 52110 23550 52162
rect 23550 52110 23602 52162
rect 23602 52110 23604 52162
rect 23548 52108 23604 52110
rect 23324 51884 23380 51940
rect 24332 55020 24388 55076
rect 24108 54290 24164 54292
rect 24108 54238 24110 54290
rect 24110 54238 24162 54290
rect 24162 54238 24164 54290
rect 24108 54236 24164 54238
rect 24220 53842 24276 53844
rect 24220 53790 24222 53842
rect 24222 53790 24274 53842
rect 24274 53790 24276 53842
rect 24220 53788 24276 53790
rect 25452 55132 25508 55188
rect 27020 55410 27076 55412
rect 27020 55358 27022 55410
rect 27022 55358 27074 55410
rect 27074 55358 27076 55410
rect 27020 55356 27076 55358
rect 27132 55244 27188 55300
rect 25788 55020 25844 55076
rect 27132 54514 27188 54516
rect 27132 54462 27134 54514
rect 27134 54462 27186 54514
rect 27186 54462 27188 54514
rect 27132 54460 27188 54462
rect 24780 53730 24836 53732
rect 24780 53678 24782 53730
rect 24782 53678 24834 53730
rect 24834 53678 24836 53730
rect 24780 53676 24836 53678
rect 25340 53730 25396 53732
rect 25340 53678 25342 53730
rect 25342 53678 25394 53730
rect 25394 53678 25396 53730
rect 25340 53676 25396 53678
rect 24220 53452 24276 53508
rect 25004 53452 25060 53508
rect 24220 53170 24276 53172
rect 24220 53118 24222 53170
rect 24222 53118 24274 53170
rect 24274 53118 24276 53170
rect 24220 53116 24276 53118
rect 25228 53116 25284 53172
rect 24108 52892 24164 52948
rect 26124 53730 26180 53732
rect 26124 53678 26126 53730
rect 26126 53678 26178 53730
rect 26178 53678 26180 53730
rect 26124 53676 26180 53678
rect 25900 53506 25956 53508
rect 25900 53454 25902 53506
rect 25902 53454 25954 53506
rect 25954 53454 25956 53506
rect 25900 53452 25956 53454
rect 27244 54012 27300 54068
rect 27132 53564 27188 53620
rect 25788 53170 25844 53172
rect 25788 53118 25790 53170
rect 25790 53118 25842 53170
rect 25842 53118 25844 53170
rect 25788 53116 25844 53118
rect 25340 52946 25396 52948
rect 25340 52894 25342 52946
rect 25342 52894 25394 52946
rect 25394 52894 25396 52946
rect 25340 52892 25396 52894
rect 23660 51154 23716 51156
rect 23660 51102 23662 51154
rect 23662 51102 23714 51154
rect 23714 51102 23716 51154
rect 23660 51100 23716 51102
rect 23324 50876 23380 50932
rect 23100 50594 23156 50596
rect 23100 50542 23102 50594
rect 23102 50542 23154 50594
rect 23154 50542 23156 50594
rect 23100 50540 23156 50542
rect 23772 50594 23828 50596
rect 23772 50542 23774 50594
rect 23774 50542 23826 50594
rect 23826 50542 23828 50594
rect 23772 50540 23828 50542
rect 24220 52162 24276 52164
rect 24220 52110 24222 52162
rect 24222 52110 24274 52162
rect 24274 52110 24276 52162
rect 24220 52108 24276 52110
rect 23884 50428 23940 50484
rect 23772 49868 23828 49924
rect 23996 49922 24052 49924
rect 23996 49870 23998 49922
rect 23998 49870 24050 49922
rect 24050 49870 24052 49922
rect 23996 49868 24052 49870
rect 23436 49644 23492 49700
rect 24220 49868 24276 49924
rect 22092 48412 22148 48468
rect 22764 48748 22820 48804
rect 22204 48354 22260 48356
rect 22204 48302 22206 48354
rect 22206 48302 22258 48354
rect 22258 48302 22260 48354
rect 22204 48300 22260 48302
rect 22428 48076 22484 48132
rect 23324 48130 23380 48132
rect 23324 48078 23326 48130
rect 23326 48078 23378 48130
rect 23378 48078 23380 48130
rect 23324 48076 23380 48078
rect 23996 47964 24052 48020
rect 24332 48802 24388 48804
rect 24332 48750 24334 48802
rect 24334 48750 24386 48802
rect 24386 48750 24388 48802
rect 24332 48748 24388 48750
rect 24444 48188 24500 48244
rect 23548 47458 23604 47460
rect 23548 47406 23550 47458
rect 23550 47406 23602 47458
rect 23602 47406 23604 47458
rect 23548 47404 23604 47406
rect 21980 45500 22036 45556
rect 22092 45836 22148 45892
rect 21980 44044 22036 44100
rect 21868 43650 21924 43652
rect 21868 43598 21870 43650
rect 21870 43598 21922 43650
rect 21922 43598 21924 43650
rect 21868 43596 21924 43598
rect 21756 42866 21812 42868
rect 21756 42814 21758 42866
rect 21758 42814 21810 42866
rect 21810 42814 21812 42866
rect 21756 42812 21812 42814
rect 21980 42754 22036 42756
rect 21980 42702 21982 42754
rect 21982 42702 22034 42754
rect 22034 42702 22036 42754
rect 21980 42700 22036 42702
rect 21420 42642 21476 42644
rect 21420 42590 21422 42642
rect 21422 42590 21474 42642
rect 21474 42590 21476 42642
rect 21420 42588 21476 42590
rect 21644 41916 21700 41972
rect 18396 38892 18452 38948
rect 18508 39340 18564 39396
rect 16940 36876 16996 36932
rect 16492 36652 16548 36708
rect 16380 35980 16436 36036
rect 16492 35756 16548 35812
rect 16268 34636 16324 34692
rect 15932 34076 15988 34132
rect 15484 32172 15540 32228
rect 15708 32172 15764 32228
rect 15372 31948 15428 32004
rect 16044 33234 16100 33236
rect 16044 33182 16046 33234
rect 16046 33182 16098 33234
rect 16098 33182 16100 33234
rect 16044 33180 16100 33182
rect 16044 32172 16100 32228
rect 15932 31724 15988 31780
rect 16044 31948 16100 32004
rect 17612 37884 17668 37940
rect 17388 36540 17444 36596
rect 17276 36092 17332 36148
rect 18844 37826 18900 37828
rect 18844 37774 18846 37826
rect 18846 37774 18898 37826
rect 18898 37774 18900 37826
rect 18844 37772 18900 37774
rect 19180 38834 19236 38836
rect 19180 38782 19182 38834
rect 19182 38782 19234 38834
rect 19234 38782 19236 38834
rect 19180 38780 19236 38782
rect 20748 40124 20804 40180
rect 20076 39788 20132 39844
rect 19516 39116 19572 39172
rect 19836 39226 19892 39228
rect 19836 39174 19838 39226
rect 19838 39174 19890 39226
rect 19890 39174 19892 39226
rect 19836 39172 19892 39174
rect 19940 39226 19996 39228
rect 19940 39174 19942 39226
rect 19942 39174 19994 39226
rect 19994 39174 19996 39226
rect 19940 39172 19996 39174
rect 20044 39226 20100 39228
rect 20044 39174 20046 39226
rect 20046 39174 20098 39226
rect 20098 39174 20100 39226
rect 20044 39172 20100 39174
rect 19628 38892 19684 38948
rect 21196 40290 21252 40292
rect 21196 40238 21198 40290
rect 21198 40238 21250 40290
rect 21250 40238 21252 40290
rect 21196 40236 21252 40238
rect 21980 40124 22036 40180
rect 21084 38892 21140 38948
rect 20076 38444 20132 38500
rect 19180 38108 19236 38164
rect 19292 38220 19348 38276
rect 19180 37938 19236 37940
rect 19180 37886 19182 37938
rect 19182 37886 19234 37938
rect 19234 37886 19236 37938
rect 19180 37884 19236 37886
rect 18172 37436 18228 37492
rect 18284 37266 18340 37268
rect 18284 37214 18286 37266
rect 18286 37214 18338 37266
rect 18338 37214 18340 37266
rect 18284 37212 18340 37214
rect 18172 37100 18228 37156
rect 17500 35810 17556 35812
rect 17500 35758 17502 35810
rect 17502 35758 17554 35810
rect 17554 35758 17556 35810
rect 17500 35756 17556 35758
rect 18060 36988 18116 37044
rect 18060 36540 18116 36596
rect 18396 36988 18452 37044
rect 18284 36764 18340 36820
rect 19628 38108 19684 38164
rect 18844 37100 18900 37156
rect 18844 36876 18900 36932
rect 17276 34860 17332 34916
rect 16604 33852 16660 33908
rect 16716 34242 16772 34244
rect 16716 34190 16718 34242
rect 16718 34190 16770 34242
rect 16770 34190 16772 34242
rect 16716 34188 16772 34190
rect 16492 32450 16548 32452
rect 16492 32398 16494 32450
rect 16494 32398 16546 32450
rect 16546 32398 16548 32450
rect 16492 32396 16548 32398
rect 17052 33346 17108 33348
rect 17052 33294 17054 33346
rect 17054 33294 17106 33346
rect 17106 33294 17108 33346
rect 17052 33292 17108 33294
rect 17388 32620 17444 32676
rect 17164 32396 17220 32452
rect 16604 31724 16660 31780
rect 15484 30210 15540 30212
rect 15484 30158 15486 30210
rect 15486 30158 15538 30210
rect 15538 30158 15540 30210
rect 15484 30156 15540 30158
rect 16044 30210 16100 30212
rect 16044 30158 16046 30210
rect 16046 30158 16098 30210
rect 16098 30158 16100 30210
rect 16044 30156 16100 30158
rect 15596 29708 15652 29764
rect 14924 26460 14980 26516
rect 14812 26012 14868 26068
rect 15148 25788 15204 25844
rect 14364 25228 14420 25284
rect 14700 24556 14756 24612
rect 14924 24108 14980 24164
rect 14028 23884 14084 23940
rect 14140 23772 14196 23828
rect 13580 23660 13636 23716
rect 13468 23154 13524 23156
rect 13468 23102 13470 23154
rect 13470 23102 13522 23154
rect 13522 23102 13524 23154
rect 13468 23100 13524 23102
rect 13916 22540 13972 22596
rect 14028 22316 14084 22372
rect 13580 22204 13636 22260
rect 12908 21420 12964 21476
rect 14252 21980 14308 22036
rect 13916 21644 13972 21700
rect 14140 21698 14196 21700
rect 14140 21646 14142 21698
rect 14142 21646 14194 21698
rect 14194 21646 14196 21698
rect 14140 21644 14196 21646
rect 15372 26236 15428 26292
rect 15148 25228 15204 25284
rect 15148 24108 15204 24164
rect 16044 29426 16100 29428
rect 16044 29374 16046 29426
rect 16046 29374 16098 29426
rect 16098 29374 16100 29426
rect 16044 29372 16100 29374
rect 16044 27692 16100 27748
rect 15708 27132 15764 27188
rect 15596 26684 15652 26740
rect 16604 31388 16660 31444
rect 16268 29596 16324 29652
rect 16492 30828 16548 30884
rect 16380 28754 16436 28756
rect 16380 28702 16382 28754
rect 16382 28702 16434 28754
rect 16434 28702 16436 28754
rect 16380 28700 16436 28702
rect 16156 27244 16212 27300
rect 16268 28588 16324 28644
rect 16044 27020 16100 27076
rect 15820 26962 15876 26964
rect 15820 26910 15822 26962
rect 15822 26910 15874 26962
rect 15874 26910 15876 26962
rect 15820 26908 15876 26910
rect 15932 26460 15988 26516
rect 16268 26236 16324 26292
rect 16156 26178 16212 26180
rect 16156 26126 16158 26178
rect 16158 26126 16210 26178
rect 16210 26126 16212 26178
rect 16156 26124 16212 26126
rect 15820 26012 15876 26068
rect 15484 23884 15540 23940
rect 15036 23324 15092 23380
rect 15708 25228 15764 25284
rect 14812 22316 14868 22372
rect 14588 22204 14644 22260
rect 14476 21644 14532 21700
rect 13244 21308 13300 21364
rect 12460 20690 12516 20692
rect 12460 20638 12462 20690
rect 12462 20638 12514 20690
rect 12514 20638 12516 20690
rect 12460 20636 12516 20638
rect 12012 19740 12068 19796
rect 12124 19346 12180 19348
rect 12124 19294 12126 19346
rect 12126 19294 12178 19346
rect 12178 19294 12180 19346
rect 12124 19292 12180 19294
rect 12572 20076 12628 20132
rect 12684 20188 12740 20244
rect 12348 19964 12404 20020
rect 11788 19068 11844 19124
rect 12908 20578 12964 20580
rect 12908 20526 12910 20578
rect 12910 20526 12962 20578
rect 12962 20526 12964 20578
rect 12908 20524 12964 20526
rect 13692 21586 13748 21588
rect 13692 21534 13694 21586
rect 13694 21534 13746 21586
rect 13746 21534 13748 21586
rect 13692 21532 13748 21534
rect 14028 21308 14084 21364
rect 14364 21308 14420 21364
rect 13468 21084 13524 21140
rect 14252 20972 14308 21028
rect 14140 20914 14196 20916
rect 14140 20862 14142 20914
rect 14142 20862 14194 20914
rect 14194 20862 14196 20914
rect 14140 20860 14196 20862
rect 13020 19852 13076 19908
rect 12908 19628 12964 19684
rect 11788 18508 11844 18564
rect 10556 17052 10612 17108
rect 12460 18508 12516 18564
rect 12796 17724 12852 17780
rect 12012 17106 12068 17108
rect 12012 17054 12014 17106
rect 12014 17054 12066 17106
rect 12066 17054 12068 17106
rect 12012 17052 12068 17054
rect 13020 17612 13076 17668
rect 13244 20636 13300 20692
rect 13468 20690 13524 20692
rect 13468 20638 13470 20690
rect 13470 20638 13522 20690
rect 13522 20638 13524 20690
rect 13468 20636 13524 20638
rect 13244 20130 13300 20132
rect 13244 20078 13246 20130
rect 13246 20078 13298 20130
rect 13298 20078 13300 20130
rect 13244 20076 13300 20078
rect 13804 20076 13860 20132
rect 13580 19180 13636 19236
rect 14028 19906 14084 19908
rect 14028 19854 14030 19906
rect 14030 19854 14082 19906
rect 14082 19854 14084 19906
rect 14028 19852 14084 19854
rect 14140 19234 14196 19236
rect 14140 19182 14142 19234
rect 14142 19182 14194 19234
rect 14194 19182 14196 19234
rect 14140 19180 14196 19182
rect 13132 18396 13188 18452
rect 13580 19010 13636 19012
rect 13580 18958 13582 19010
rect 13582 18958 13634 19010
rect 13634 18958 13636 19010
rect 13580 18956 13636 18958
rect 13692 17948 13748 18004
rect 13580 17778 13636 17780
rect 13580 17726 13582 17778
rect 13582 17726 13634 17778
rect 13634 17726 13636 17778
rect 13580 17724 13636 17726
rect 13580 17106 13636 17108
rect 13580 17054 13582 17106
rect 13582 17054 13634 17106
rect 13634 17054 13636 17106
rect 13580 17052 13636 17054
rect 11564 16882 11620 16884
rect 11564 16830 11566 16882
rect 11566 16830 11618 16882
rect 11618 16830 11620 16882
rect 11564 16828 11620 16830
rect 14028 16882 14084 16884
rect 14028 16830 14030 16882
rect 14030 16830 14082 16882
rect 14082 16830 14084 16882
rect 14028 16828 14084 16830
rect 14028 16268 14084 16324
rect 15148 21868 15204 21924
rect 15596 21810 15652 21812
rect 15596 21758 15598 21810
rect 15598 21758 15650 21810
rect 15650 21758 15652 21810
rect 15596 21756 15652 21758
rect 14588 21420 14644 21476
rect 14700 21308 14756 21364
rect 14700 20636 14756 20692
rect 14476 20524 14532 20580
rect 14588 20412 14644 20468
rect 15484 21532 15540 21588
rect 15036 20412 15092 20468
rect 15372 21308 15428 21364
rect 14924 20300 14980 20356
rect 14700 20076 14756 20132
rect 15148 20076 15204 20132
rect 14700 19740 14756 19796
rect 14924 19852 14980 19908
rect 16268 26012 16324 26068
rect 16156 25116 16212 25172
rect 15932 24780 15988 24836
rect 16492 27468 16548 27524
rect 16492 27244 16548 27300
rect 17052 31724 17108 31780
rect 17052 31276 17108 31332
rect 16828 30268 16884 30324
rect 16828 29932 16884 29988
rect 17052 30156 17108 30212
rect 17052 28642 17108 28644
rect 17052 28590 17054 28642
rect 17054 28590 17106 28642
rect 17106 28590 17108 28642
rect 17052 28588 17108 28590
rect 17724 33628 17780 33684
rect 17836 33404 17892 33460
rect 18172 35586 18228 35588
rect 18172 35534 18174 35586
rect 18174 35534 18226 35586
rect 18226 35534 18228 35586
rect 18172 35532 18228 35534
rect 18172 33292 18228 33348
rect 17500 31724 17556 31780
rect 17500 31388 17556 31444
rect 17388 30994 17444 30996
rect 17388 30942 17390 30994
rect 17390 30942 17442 30994
rect 17442 30942 17444 30994
rect 17388 30940 17444 30942
rect 18956 35980 19012 36036
rect 18620 35196 18676 35252
rect 19292 36988 19348 37044
rect 19180 36876 19236 36932
rect 19404 36764 19460 36820
rect 19404 35922 19460 35924
rect 19404 35870 19406 35922
rect 19406 35870 19458 35922
rect 19458 35870 19460 35922
rect 19404 35868 19460 35870
rect 20188 38108 20244 38164
rect 19836 37658 19892 37660
rect 19836 37606 19838 37658
rect 19838 37606 19890 37658
rect 19890 37606 19892 37658
rect 19836 37604 19892 37606
rect 19940 37658 19996 37660
rect 19940 37606 19942 37658
rect 19942 37606 19994 37658
rect 19994 37606 19996 37658
rect 19940 37604 19996 37606
rect 20044 37658 20100 37660
rect 20044 37606 20046 37658
rect 20046 37606 20098 37658
rect 20098 37606 20100 37658
rect 20044 37604 20100 37606
rect 19852 37490 19908 37492
rect 19852 37438 19854 37490
rect 19854 37438 19906 37490
rect 19906 37438 19908 37490
rect 19852 37436 19908 37438
rect 19740 37266 19796 37268
rect 19740 37214 19742 37266
rect 19742 37214 19794 37266
rect 19794 37214 19796 37266
rect 19740 37212 19796 37214
rect 19964 37100 20020 37156
rect 20076 36876 20132 36932
rect 20748 37938 20804 37940
rect 20748 37886 20750 37938
rect 20750 37886 20802 37938
rect 20802 37886 20804 37938
rect 20748 37884 20804 37886
rect 22204 45500 22260 45556
rect 22540 46620 22596 46676
rect 22876 47234 22932 47236
rect 22876 47182 22878 47234
rect 22878 47182 22930 47234
rect 22930 47182 22932 47234
rect 22876 47180 22932 47182
rect 23100 46674 23156 46676
rect 23100 46622 23102 46674
rect 23102 46622 23154 46674
rect 23154 46622 23156 46674
rect 23100 46620 23156 46622
rect 23212 46562 23268 46564
rect 23212 46510 23214 46562
rect 23214 46510 23266 46562
rect 23266 46510 23268 46562
rect 23212 46508 23268 46510
rect 22988 45836 23044 45892
rect 22876 45666 22932 45668
rect 22876 45614 22878 45666
rect 22878 45614 22930 45666
rect 22930 45614 22932 45666
rect 22876 45612 22932 45614
rect 23436 45164 23492 45220
rect 22540 44994 22596 44996
rect 22540 44942 22542 44994
rect 22542 44942 22594 44994
rect 22594 44942 22596 44994
rect 22540 44940 22596 44942
rect 22428 40124 22484 40180
rect 22204 39730 22260 39732
rect 22204 39678 22206 39730
rect 22206 39678 22258 39730
rect 22258 39678 22260 39730
rect 22204 39676 22260 39678
rect 21308 38722 21364 38724
rect 21308 38670 21310 38722
rect 21310 38670 21362 38722
rect 21362 38670 21364 38722
rect 21308 38668 21364 38670
rect 20860 37378 20916 37380
rect 20860 37326 20862 37378
rect 20862 37326 20914 37378
rect 20914 37326 20916 37378
rect 20860 37324 20916 37326
rect 19836 36090 19892 36092
rect 19836 36038 19838 36090
rect 19838 36038 19890 36090
rect 19890 36038 19892 36090
rect 19836 36036 19892 36038
rect 19940 36090 19996 36092
rect 19940 36038 19942 36090
rect 19942 36038 19994 36090
rect 19994 36038 19996 36090
rect 19940 36036 19996 36038
rect 20044 36090 20100 36092
rect 20044 36038 20046 36090
rect 20046 36038 20098 36090
rect 20098 36038 20100 36090
rect 20044 36036 20100 36038
rect 19516 35756 19572 35812
rect 19964 35868 20020 35924
rect 19404 34972 19460 35028
rect 19628 34914 19684 34916
rect 19628 34862 19630 34914
rect 19630 34862 19682 34914
rect 19682 34862 19684 34914
rect 19628 34860 19684 34862
rect 20076 35196 20132 35252
rect 20412 36428 20468 36484
rect 20636 36092 20692 36148
rect 20636 35308 20692 35364
rect 20860 36988 20916 37044
rect 20972 37212 21028 37268
rect 20524 35196 20580 35252
rect 19292 34802 19348 34804
rect 19292 34750 19294 34802
rect 19294 34750 19346 34802
rect 19346 34750 19348 34802
rect 19292 34748 19348 34750
rect 20300 34860 20356 34916
rect 18508 34188 18564 34244
rect 18508 33516 18564 33572
rect 18060 32338 18116 32340
rect 18060 32286 18062 32338
rect 18062 32286 18114 32338
rect 18114 32286 18116 32338
rect 18060 32284 18116 32286
rect 18284 31948 18340 32004
rect 18284 31778 18340 31780
rect 18284 31726 18286 31778
rect 18286 31726 18338 31778
rect 18338 31726 18340 31778
rect 18284 31724 18340 31726
rect 19068 33852 19124 33908
rect 19180 33740 19236 33796
rect 18620 32284 18676 32340
rect 18060 30940 18116 30996
rect 17388 29426 17444 29428
rect 17388 29374 17390 29426
rect 17390 29374 17442 29426
rect 17442 29374 17444 29426
rect 17388 29372 17444 29374
rect 17388 28476 17444 28532
rect 16828 27244 16884 27300
rect 16604 26012 16660 26068
rect 16716 24780 16772 24836
rect 16716 23548 16772 23604
rect 16156 23100 16212 23156
rect 15820 22204 15876 22260
rect 15932 22652 15988 22708
rect 15484 20188 15540 20244
rect 15260 19964 15316 20020
rect 15148 19122 15204 19124
rect 15148 19070 15150 19122
rect 15150 19070 15202 19122
rect 15202 19070 15204 19122
rect 15148 19068 15204 19070
rect 14812 18956 14868 19012
rect 14700 18284 14756 18340
rect 15820 20636 15876 20692
rect 15708 19906 15764 19908
rect 15708 19854 15710 19906
rect 15710 19854 15762 19906
rect 15762 19854 15764 19906
rect 15708 19852 15764 19854
rect 15596 19180 15652 19236
rect 15596 18450 15652 18452
rect 15596 18398 15598 18450
rect 15598 18398 15650 18450
rect 15650 18398 15652 18450
rect 15596 18396 15652 18398
rect 15148 17724 15204 17780
rect 14924 16268 14980 16324
rect 16828 22764 16884 22820
rect 17836 28700 17892 28756
rect 17724 27692 17780 27748
rect 17388 26460 17444 26516
rect 17948 26514 18004 26516
rect 17948 26462 17950 26514
rect 17950 26462 18002 26514
rect 18002 26462 18004 26514
rect 17948 26460 18004 26462
rect 19836 34522 19892 34524
rect 19836 34470 19838 34522
rect 19838 34470 19890 34522
rect 19890 34470 19892 34522
rect 19836 34468 19892 34470
rect 19940 34522 19996 34524
rect 19940 34470 19942 34522
rect 19942 34470 19994 34522
rect 19994 34470 19996 34522
rect 19940 34468 19996 34470
rect 20044 34522 20100 34524
rect 20044 34470 20046 34522
rect 20046 34470 20098 34522
rect 20098 34470 20100 34522
rect 20044 34468 20100 34470
rect 19628 33628 19684 33684
rect 20524 33740 20580 33796
rect 20972 36316 21028 36372
rect 21980 38444 22036 38500
rect 21756 37884 21812 37940
rect 21868 38220 21924 38276
rect 21644 37772 21700 37828
rect 21868 37660 21924 37716
rect 21868 37266 21924 37268
rect 21868 37214 21870 37266
rect 21870 37214 21922 37266
rect 21922 37214 21924 37266
rect 21868 37212 21924 37214
rect 21532 36876 21588 36932
rect 21420 36764 21476 36820
rect 21644 36764 21700 36820
rect 21308 36204 21364 36260
rect 21084 35698 21140 35700
rect 21084 35646 21086 35698
rect 21086 35646 21138 35698
rect 21138 35646 21140 35698
rect 21084 35644 21140 35646
rect 21532 36428 21588 36484
rect 21532 35810 21588 35812
rect 21532 35758 21534 35810
rect 21534 35758 21586 35810
rect 21586 35758 21588 35810
rect 21532 35756 21588 35758
rect 21420 35308 21476 35364
rect 21420 35026 21476 35028
rect 21420 34974 21422 35026
rect 21422 34974 21474 35026
rect 21474 34974 21476 35026
rect 21420 34972 21476 34974
rect 21308 34802 21364 34804
rect 21308 34750 21310 34802
rect 21310 34750 21362 34802
rect 21362 34750 21364 34802
rect 21308 34748 21364 34750
rect 22316 39452 22372 39508
rect 22428 39116 22484 39172
rect 23548 44940 23604 44996
rect 23660 44322 23716 44324
rect 23660 44270 23662 44322
rect 23662 44270 23714 44322
rect 23714 44270 23716 44322
rect 23660 44268 23716 44270
rect 22764 44098 22820 44100
rect 22764 44046 22766 44098
rect 22766 44046 22818 44098
rect 22818 44046 22820 44098
rect 22764 44044 22820 44046
rect 22652 42866 22708 42868
rect 22652 42814 22654 42866
rect 22654 42814 22706 42866
rect 22706 42814 22708 42866
rect 22652 42812 22708 42814
rect 22652 41916 22708 41972
rect 22652 37772 22708 37828
rect 22316 37660 22372 37716
rect 22316 37266 22372 37268
rect 22316 37214 22318 37266
rect 22318 37214 22370 37266
rect 22370 37214 22372 37266
rect 22316 37212 22372 37214
rect 22204 37100 22260 37156
rect 21868 36092 21924 36148
rect 22316 36092 22372 36148
rect 22764 37436 22820 37492
rect 22540 36988 22596 37044
rect 19628 33180 19684 33236
rect 19068 31724 19124 31780
rect 18620 30882 18676 30884
rect 18620 30830 18622 30882
rect 18622 30830 18674 30882
rect 18674 30830 18676 30882
rect 18620 30828 18676 30830
rect 18732 31500 18788 31556
rect 18396 29596 18452 29652
rect 18172 28812 18228 28868
rect 18396 28588 18452 28644
rect 18620 28028 18676 28084
rect 19180 30044 19236 30100
rect 18956 28364 19012 28420
rect 18732 27580 18788 27636
rect 18620 27244 18676 27300
rect 18172 27132 18228 27188
rect 18396 26852 18452 26908
rect 17388 26012 17444 26068
rect 17724 25004 17780 25060
rect 18172 25228 18228 25284
rect 18620 26402 18676 26404
rect 18620 26350 18622 26402
rect 18622 26350 18674 26402
rect 18674 26350 18676 26402
rect 18620 26348 18676 26350
rect 18620 25452 18676 25508
rect 18732 25394 18788 25396
rect 18732 25342 18734 25394
rect 18734 25342 18786 25394
rect 18786 25342 18788 25394
rect 18732 25340 18788 25342
rect 18284 24220 18340 24276
rect 17612 23660 17668 23716
rect 17948 23884 18004 23940
rect 17612 23212 17668 23268
rect 17836 23548 17892 23604
rect 17724 22764 17780 22820
rect 17612 22540 17668 22596
rect 17612 22370 17668 22372
rect 17612 22318 17614 22370
rect 17614 22318 17666 22370
rect 17666 22318 17668 22370
rect 17612 22316 17668 22318
rect 16716 21868 16772 21924
rect 16156 21532 16212 21588
rect 16268 20690 16324 20692
rect 16268 20638 16270 20690
rect 16270 20638 16322 20690
rect 16322 20638 16324 20690
rect 16268 20636 16324 20638
rect 16268 19964 16324 20020
rect 16492 20130 16548 20132
rect 16492 20078 16494 20130
rect 16494 20078 16546 20130
rect 16546 20078 16548 20130
rect 16492 20076 16548 20078
rect 16044 19346 16100 19348
rect 16044 19294 16046 19346
rect 16046 19294 16098 19346
rect 16098 19294 16100 19346
rect 16044 19292 16100 19294
rect 16492 19010 16548 19012
rect 16492 18958 16494 19010
rect 16494 18958 16546 19010
rect 16546 18958 16548 19010
rect 16492 18956 16548 18958
rect 16940 21532 16996 21588
rect 17724 21308 17780 21364
rect 16940 19964 16996 20020
rect 16716 19404 16772 19460
rect 16380 18338 16436 18340
rect 16380 18286 16382 18338
rect 16382 18286 16434 18338
rect 16434 18286 16436 18338
rect 16380 18284 16436 18286
rect 16604 16156 16660 16212
rect 16044 15820 16100 15876
rect 14700 15148 14756 15204
rect 4476 14922 4532 14924
rect 4476 14870 4478 14922
rect 4478 14870 4530 14922
rect 4530 14870 4532 14922
rect 4476 14868 4532 14870
rect 4580 14922 4636 14924
rect 4580 14870 4582 14922
rect 4582 14870 4634 14922
rect 4634 14870 4636 14922
rect 4580 14868 4636 14870
rect 4684 14922 4740 14924
rect 4684 14870 4686 14922
rect 4686 14870 4738 14922
rect 4738 14870 4740 14922
rect 4684 14868 4740 14870
rect 4476 13354 4532 13356
rect 4476 13302 4478 13354
rect 4478 13302 4530 13354
rect 4530 13302 4532 13354
rect 4476 13300 4532 13302
rect 4580 13354 4636 13356
rect 4580 13302 4582 13354
rect 4582 13302 4634 13354
rect 4634 13302 4636 13354
rect 4580 13300 4636 13302
rect 4684 13354 4740 13356
rect 4684 13302 4686 13354
rect 4686 13302 4738 13354
rect 4738 13302 4740 13354
rect 4684 13300 4740 13302
rect 4476 11786 4532 11788
rect 4476 11734 4478 11786
rect 4478 11734 4530 11786
rect 4530 11734 4532 11786
rect 4476 11732 4532 11734
rect 4580 11786 4636 11788
rect 4580 11734 4582 11786
rect 4582 11734 4634 11786
rect 4634 11734 4636 11786
rect 4580 11732 4636 11734
rect 4684 11786 4740 11788
rect 4684 11734 4686 11786
rect 4686 11734 4738 11786
rect 4738 11734 4740 11786
rect 4684 11732 4740 11734
rect 4476 10218 4532 10220
rect 4476 10166 4478 10218
rect 4478 10166 4530 10218
rect 4530 10166 4532 10218
rect 4476 10164 4532 10166
rect 4580 10218 4636 10220
rect 4580 10166 4582 10218
rect 4582 10166 4634 10218
rect 4634 10166 4636 10218
rect 4580 10164 4636 10166
rect 4684 10218 4740 10220
rect 4684 10166 4686 10218
rect 4686 10166 4738 10218
rect 4738 10166 4740 10218
rect 4684 10164 4740 10166
rect 16268 15314 16324 15316
rect 16268 15262 16270 15314
rect 16270 15262 16322 15314
rect 16322 15262 16324 15314
rect 16268 15260 16324 15262
rect 16380 15202 16436 15204
rect 16380 15150 16382 15202
rect 16382 15150 16434 15202
rect 16434 15150 16436 15202
rect 16380 15148 16436 15150
rect 16940 18956 16996 19012
rect 16940 18396 16996 18452
rect 16940 17612 16996 17668
rect 18284 23772 18340 23828
rect 18620 24668 18676 24724
rect 18396 23378 18452 23380
rect 18396 23326 18398 23378
rect 18398 23326 18450 23378
rect 18450 23326 18452 23378
rect 18396 23324 18452 23326
rect 18060 22988 18116 23044
rect 18060 21868 18116 21924
rect 18172 22876 18228 22932
rect 18508 22764 18564 22820
rect 17948 21756 18004 21812
rect 17948 20914 18004 20916
rect 17948 20862 17950 20914
rect 17950 20862 18002 20914
rect 18002 20862 18004 20914
rect 17948 20860 18004 20862
rect 17724 20802 17780 20804
rect 17724 20750 17726 20802
rect 17726 20750 17778 20802
rect 17778 20750 17780 20802
rect 17724 20748 17780 20750
rect 17388 20130 17444 20132
rect 17388 20078 17390 20130
rect 17390 20078 17442 20130
rect 17442 20078 17444 20130
rect 17388 20076 17444 20078
rect 17164 19292 17220 19348
rect 17836 20076 17892 20132
rect 17612 19964 17668 20020
rect 17500 19906 17556 19908
rect 17500 19854 17502 19906
rect 17502 19854 17554 19906
rect 17554 19854 17556 19906
rect 17500 19852 17556 19854
rect 17388 19010 17444 19012
rect 17388 18958 17390 19010
rect 17390 18958 17442 19010
rect 17442 18958 17444 19010
rect 17388 18956 17444 18958
rect 17500 18508 17556 18564
rect 17724 18450 17780 18452
rect 17724 18398 17726 18450
rect 17726 18398 17778 18450
rect 17778 18398 17780 18450
rect 17724 18396 17780 18398
rect 17052 17052 17108 17108
rect 16828 16940 16884 16996
rect 17500 18284 17556 18340
rect 17164 16268 17220 16324
rect 17836 17500 17892 17556
rect 16716 15148 16772 15204
rect 17276 15874 17332 15876
rect 17276 15822 17278 15874
rect 17278 15822 17330 15874
rect 17330 15822 17332 15874
rect 17276 15820 17332 15822
rect 17164 15260 17220 15316
rect 14028 13580 14084 13636
rect 15260 13580 15316 13636
rect 18060 20018 18116 20020
rect 18060 19966 18062 20018
rect 18062 19966 18114 20018
rect 18114 19966 18116 20018
rect 18060 19964 18116 19966
rect 18284 21532 18340 21588
rect 18956 27020 19012 27076
rect 20524 33122 20580 33124
rect 20524 33070 20526 33122
rect 20526 33070 20578 33122
rect 20578 33070 20580 33122
rect 20524 33068 20580 33070
rect 19836 32954 19892 32956
rect 19836 32902 19838 32954
rect 19838 32902 19890 32954
rect 19890 32902 19892 32954
rect 19836 32900 19892 32902
rect 19940 32954 19996 32956
rect 19940 32902 19942 32954
rect 19942 32902 19994 32954
rect 19994 32902 19996 32954
rect 19940 32900 19996 32902
rect 20044 32954 20100 32956
rect 20044 32902 20046 32954
rect 20046 32902 20098 32954
rect 20098 32902 20100 32954
rect 20044 32900 20100 32902
rect 20188 32396 20244 32452
rect 19836 31386 19892 31388
rect 19836 31334 19838 31386
rect 19838 31334 19890 31386
rect 19890 31334 19892 31386
rect 19836 31332 19892 31334
rect 19940 31386 19996 31388
rect 19940 31334 19942 31386
rect 19942 31334 19994 31386
rect 19994 31334 19996 31386
rect 19940 31332 19996 31334
rect 20044 31386 20100 31388
rect 20044 31334 20046 31386
rect 20046 31334 20098 31386
rect 20098 31334 20100 31386
rect 20044 31332 20100 31334
rect 19628 30882 19684 30884
rect 19628 30830 19630 30882
rect 19630 30830 19682 30882
rect 19682 30830 19684 30882
rect 19628 30828 19684 30830
rect 20076 30492 20132 30548
rect 19404 29596 19460 29652
rect 19628 30210 19684 30212
rect 19628 30158 19630 30210
rect 19630 30158 19682 30210
rect 19682 30158 19684 30210
rect 19628 30156 19684 30158
rect 19180 28028 19236 28084
rect 19180 27356 19236 27412
rect 19836 29818 19892 29820
rect 19836 29766 19838 29818
rect 19838 29766 19890 29818
rect 19890 29766 19892 29818
rect 19836 29764 19892 29766
rect 19940 29818 19996 29820
rect 19940 29766 19942 29818
rect 19942 29766 19994 29818
rect 19994 29766 19996 29818
rect 19940 29764 19996 29766
rect 20044 29818 20100 29820
rect 20044 29766 20046 29818
rect 20046 29766 20098 29818
rect 20098 29766 20100 29818
rect 20044 29764 20100 29766
rect 19740 29596 19796 29652
rect 20412 31890 20468 31892
rect 20412 31838 20414 31890
rect 20414 31838 20466 31890
rect 20466 31838 20468 31890
rect 20412 31836 20468 31838
rect 21308 33628 21364 33684
rect 20972 33516 21028 33572
rect 20748 32060 20804 32116
rect 21308 33068 21364 33124
rect 21196 31948 21252 32004
rect 20636 31778 20692 31780
rect 20636 31726 20638 31778
rect 20638 31726 20690 31778
rect 20690 31726 20692 31778
rect 20636 31724 20692 31726
rect 20748 31612 20804 31668
rect 20636 31164 20692 31220
rect 20524 30994 20580 30996
rect 20524 30942 20526 30994
rect 20526 30942 20578 30994
rect 20578 30942 20580 30994
rect 20524 30940 20580 30942
rect 20972 31612 21028 31668
rect 20412 30210 20468 30212
rect 20412 30158 20414 30210
rect 20414 30158 20466 30210
rect 20466 30158 20468 30210
rect 20412 30156 20468 30158
rect 20300 29036 20356 29092
rect 19852 28754 19908 28756
rect 19852 28702 19854 28754
rect 19854 28702 19906 28754
rect 19906 28702 19908 28754
rect 19852 28700 19908 28702
rect 19836 28250 19892 28252
rect 19836 28198 19838 28250
rect 19838 28198 19890 28250
rect 19890 28198 19892 28250
rect 19836 28196 19892 28198
rect 19940 28250 19996 28252
rect 19940 28198 19942 28250
rect 19942 28198 19994 28250
rect 19994 28198 19996 28250
rect 19940 28196 19996 28198
rect 20044 28250 20100 28252
rect 20044 28198 20046 28250
rect 20046 28198 20098 28250
rect 20098 28198 20100 28250
rect 20044 28196 20100 28198
rect 19068 26908 19124 26964
rect 19068 26684 19124 26740
rect 18956 26402 19012 26404
rect 18956 26350 18958 26402
rect 18958 26350 19010 26402
rect 19010 26350 19012 26402
rect 18956 26348 19012 26350
rect 19516 27356 19572 27412
rect 20188 27074 20244 27076
rect 20188 27022 20190 27074
rect 20190 27022 20242 27074
rect 20242 27022 20244 27074
rect 20188 27020 20244 27022
rect 19516 26796 19572 26852
rect 20300 26796 20356 26852
rect 19836 26682 19892 26684
rect 19836 26630 19838 26682
rect 19838 26630 19890 26682
rect 19890 26630 19892 26682
rect 19836 26628 19892 26630
rect 19940 26682 19996 26684
rect 19940 26630 19942 26682
rect 19942 26630 19994 26682
rect 19994 26630 19996 26682
rect 19940 26628 19996 26630
rect 20044 26682 20100 26684
rect 20044 26630 20046 26682
rect 20046 26630 20098 26682
rect 20098 26630 20100 26682
rect 20044 26628 20100 26630
rect 20188 26684 20244 26740
rect 20300 26514 20356 26516
rect 20300 26462 20302 26514
rect 20302 26462 20354 26514
rect 20354 26462 20356 26514
rect 20300 26460 20356 26462
rect 19068 25452 19124 25508
rect 19292 25394 19348 25396
rect 19292 25342 19294 25394
rect 19294 25342 19346 25394
rect 19346 25342 19348 25394
rect 19292 25340 19348 25342
rect 19740 26012 19796 26068
rect 18844 24892 18900 24948
rect 18956 24722 19012 24724
rect 18956 24670 18958 24722
rect 18958 24670 19010 24722
rect 19010 24670 19012 24722
rect 18956 24668 19012 24670
rect 19404 25116 19460 25172
rect 19516 25004 19572 25060
rect 18956 23996 19012 24052
rect 18508 21308 18564 21364
rect 18844 22540 18900 22596
rect 18732 21810 18788 21812
rect 18732 21758 18734 21810
rect 18734 21758 18786 21810
rect 18786 21758 18788 21810
rect 18732 21756 18788 21758
rect 18284 20412 18340 20468
rect 18396 19964 18452 20020
rect 18396 19516 18452 19572
rect 18060 18284 18116 18340
rect 17948 17388 18004 17444
rect 18284 17836 18340 17892
rect 17500 17106 17556 17108
rect 17500 17054 17502 17106
rect 17502 17054 17554 17106
rect 17554 17054 17556 17106
rect 17500 17052 17556 17054
rect 18172 16940 18228 16996
rect 17612 16268 17668 16324
rect 17500 16156 17556 16212
rect 20300 26124 20356 26180
rect 20860 30604 20916 30660
rect 20748 30210 20804 30212
rect 20748 30158 20750 30210
rect 20750 30158 20802 30210
rect 20802 30158 20804 30210
rect 20748 30156 20804 30158
rect 20748 29650 20804 29652
rect 20748 29598 20750 29650
rect 20750 29598 20802 29650
rect 20802 29598 20804 29650
rect 20748 29596 20804 29598
rect 21532 33906 21588 33908
rect 21532 33854 21534 33906
rect 21534 33854 21586 33906
rect 21586 33854 21588 33906
rect 21532 33852 21588 33854
rect 22204 35308 22260 35364
rect 21644 33292 21700 33348
rect 22092 33740 22148 33796
rect 22092 33346 22148 33348
rect 22092 33294 22094 33346
rect 22094 33294 22146 33346
rect 22146 33294 22148 33346
rect 22092 33292 22148 33294
rect 21420 31500 21476 31556
rect 21532 31724 21588 31780
rect 21420 30044 21476 30100
rect 20636 29148 20692 29204
rect 21420 29148 21476 29204
rect 22092 32562 22148 32564
rect 22092 32510 22094 32562
rect 22094 32510 22146 32562
rect 22146 32510 22148 32562
rect 22092 32508 22148 32510
rect 21644 29036 21700 29092
rect 21756 32060 21812 32116
rect 21868 31836 21924 31892
rect 21980 31778 22036 31780
rect 21980 31726 21982 31778
rect 21982 31726 22034 31778
rect 22034 31726 22036 31778
rect 21980 31724 22036 31726
rect 21980 31164 22036 31220
rect 21868 30210 21924 30212
rect 21868 30158 21870 30210
rect 21870 30158 21922 30210
rect 21922 30158 21924 30210
rect 21868 30156 21924 30158
rect 21756 30044 21812 30100
rect 23996 47570 24052 47572
rect 23996 47518 23998 47570
rect 23998 47518 24050 47570
rect 24050 47518 24052 47570
rect 23996 47516 24052 47518
rect 24108 47404 24164 47460
rect 24668 48130 24724 48132
rect 24668 48078 24670 48130
rect 24670 48078 24722 48130
rect 24722 48078 24724 48130
rect 24668 48076 24724 48078
rect 24556 47964 24612 48020
rect 24668 47404 24724 47460
rect 24444 47068 24500 47124
rect 24668 47180 24724 47236
rect 23884 46562 23940 46564
rect 23884 46510 23886 46562
rect 23886 46510 23938 46562
rect 23938 46510 23940 46562
rect 23884 46508 23940 46510
rect 25788 52332 25844 52388
rect 26348 52332 26404 52388
rect 27020 53506 27076 53508
rect 27020 53454 27022 53506
rect 27022 53454 27074 53506
rect 27074 53454 27076 53506
rect 27020 53452 27076 53454
rect 26908 52332 26964 52388
rect 25340 49138 25396 49140
rect 25340 49086 25342 49138
rect 25342 49086 25394 49138
rect 25394 49086 25396 49138
rect 25340 49084 25396 49086
rect 25676 51100 25732 51156
rect 26236 50428 26292 50484
rect 25676 49644 25732 49700
rect 25564 48972 25620 49028
rect 25900 49586 25956 49588
rect 25900 49534 25902 49586
rect 25902 49534 25954 49586
rect 25954 49534 25956 49586
rect 25900 49532 25956 49534
rect 27468 54684 27524 54740
rect 27468 54460 27524 54516
rect 28252 55074 28308 55076
rect 28252 55022 28254 55074
rect 28254 55022 28306 55074
rect 28306 55022 28308 55074
rect 28252 55020 28308 55022
rect 27356 53228 27412 53284
rect 27804 53676 27860 53732
rect 27916 54684 27972 54740
rect 28028 54460 28084 54516
rect 27692 53564 27748 53620
rect 30716 55186 30772 55188
rect 30716 55134 30718 55186
rect 30718 55134 30770 55186
rect 30770 55134 30772 55186
rect 30716 55132 30772 55134
rect 30156 55020 30212 55076
rect 30044 54348 30100 54404
rect 30940 54348 30996 54404
rect 31388 54402 31444 54404
rect 31388 54350 31390 54402
rect 31390 54350 31442 54402
rect 31442 54350 31444 54402
rect 31388 54348 31444 54350
rect 32172 55468 32228 55524
rect 31836 55356 31892 55412
rect 32508 55132 32564 55188
rect 31836 53900 31892 53956
rect 32508 53788 32564 53844
rect 29148 53730 29204 53732
rect 29148 53678 29150 53730
rect 29150 53678 29202 53730
rect 29202 53678 29204 53730
rect 29148 53676 29204 53678
rect 32956 53730 33012 53732
rect 32956 53678 32958 53730
rect 32958 53678 33010 53730
rect 33010 53678 33012 53730
rect 32956 53676 33012 53678
rect 28476 53228 28532 53284
rect 28588 53564 28644 53620
rect 26796 51548 26852 51604
rect 27020 51490 27076 51492
rect 27020 51438 27022 51490
rect 27022 51438 27074 51490
rect 27074 51438 27076 51490
rect 27020 51436 27076 51438
rect 28028 51602 28084 51604
rect 28028 51550 28030 51602
rect 28030 51550 28082 51602
rect 28082 51550 28084 51602
rect 28028 51548 28084 51550
rect 28140 51490 28196 51492
rect 28140 51438 28142 51490
rect 28142 51438 28194 51490
rect 28194 51438 28196 51490
rect 28140 51436 28196 51438
rect 26796 50428 26852 50484
rect 28028 51212 28084 51268
rect 30828 53618 30884 53620
rect 30828 53566 30830 53618
rect 30830 53566 30882 53618
rect 30882 53566 30884 53618
rect 30828 53564 30884 53566
rect 29596 53506 29652 53508
rect 29596 53454 29598 53506
rect 29598 53454 29650 53506
rect 29650 53454 29652 53506
rect 29596 53452 29652 53454
rect 30268 53506 30324 53508
rect 30268 53454 30270 53506
rect 30270 53454 30322 53506
rect 30322 53454 30324 53506
rect 30268 53452 30324 53454
rect 29260 53228 29316 53284
rect 29260 52162 29316 52164
rect 29260 52110 29262 52162
rect 29262 52110 29314 52162
rect 29314 52110 29316 52162
rect 29260 52108 29316 52110
rect 28028 50706 28084 50708
rect 28028 50654 28030 50706
rect 28030 50654 28082 50706
rect 28082 50654 28084 50706
rect 28028 50652 28084 50654
rect 28700 50652 28756 50708
rect 26460 49756 26516 49812
rect 26460 48972 26516 49028
rect 26460 48802 26516 48804
rect 26460 48750 26462 48802
rect 26462 48750 26514 48802
rect 26514 48750 26516 48802
rect 26460 48748 26516 48750
rect 25564 48242 25620 48244
rect 25564 48190 25566 48242
rect 25566 48190 25618 48242
rect 25618 48190 25620 48242
rect 25564 48188 25620 48190
rect 25340 48130 25396 48132
rect 25340 48078 25342 48130
rect 25342 48078 25394 48130
rect 25394 48078 25396 48130
rect 25340 48076 25396 48078
rect 23996 45778 24052 45780
rect 23996 45726 23998 45778
rect 23998 45726 24050 45778
rect 24050 45726 24052 45778
rect 23996 45724 24052 45726
rect 25004 47404 25060 47460
rect 24332 45164 24388 45220
rect 24556 45666 24612 45668
rect 24556 45614 24558 45666
rect 24558 45614 24610 45666
rect 24610 45614 24612 45666
rect 24556 45612 24612 45614
rect 24668 44994 24724 44996
rect 24668 44942 24670 44994
rect 24670 44942 24722 44994
rect 24722 44942 24724 44994
rect 24668 44940 24724 44942
rect 24556 44268 24612 44324
rect 24668 44492 24724 44548
rect 23996 43596 24052 43652
rect 23996 42812 24052 42868
rect 23884 42028 23940 42084
rect 24556 42866 24612 42868
rect 24556 42814 24558 42866
rect 24558 42814 24610 42866
rect 24610 42814 24612 42866
rect 24556 42812 24612 42814
rect 25340 47346 25396 47348
rect 25340 47294 25342 47346
rect 25342 47294 25394 47346
rect 25394 47294 25396 47346
rect 25340 47292 25396 47294
rect 25004 46844 25060 46900
rect 25340 46898 25396 46900
rect 25340 46846 25342 46898
rect 25342 46846 25394 46898
rect 25394 46846 25396 46898
rect 25340 46844 25396 46846
rect 27356 49084 27412 49140
rect 26796 47964 26852 48020
rect 27020 48130 27076 48132
rect 27020 48078 27022 48130
rect 27022 48078 27074 48130
rect 27074 48078 27076 48130
rect 27020 48076 27076 48078
rect 26908 47404 26964 47460
rect 27580 49810 27636 49812
rect 27580 49758 27582 49810
rect 27582 49758 27634 49810
rect 27634 49758 27636 49810
rect 27580 49756 27636 49758
rect 27132 47740 27188 47796
rect 27132 47180 27188 47236
rect 25004 45500 25060 45556
rect 25340 45666 25396 45668
rect 25340 45614 25342 45666
rect 25342 45614 25394 45666
rect 25394 45614 25396 45666
rect 25340 45612 25396 45614
rect 25452 45500 25508 45556
rect 25004 45164 25060 45220
rect 25004 44940 25060 44996
rect 24892 44322 24948 44324
rect 24892 44270 24894 44322
rect 24894 44270 24946 44322
rect 24946 44270 24948 44322
rect 24892 44268 24948 44270
rect 25452 45106 25508 45108
rect 25452 45054 25454 45106
rect 25454 45054 25506 45106
rect 25506 45054 25508 45106
rect 25452 45052 25508 45054
rect 25452 44492 25508 44548
rect 25452 44268 25508 44324
rect 24892 43596 24948 43652
rect 24668 41970 24724 41972
rect 24668 41918 24670 41970
rect 24670 41918 24722 41970
rect 24722 41918 24724 41970
rect 24668 41916 24724 41918
rect 23884 40514 23940 40516
rect 23884 40462 23886 40514
rect 23886 40462 23938 40514
rect 23938 40462 23940 40514
rect 23884 40460 23940 40462
rect 24444 40402 24500 40404
rect 24444 40350 24446 40402
rect 24446 40350 24498 40402
rect 24498 40350 24500 40402
rect 24444 40348 24500 40350
rect 23548 39506 23604 39508
rect 23548 39454 23550 39506
rect 23550 39454 23602 39506
rect 23602 39454 23604 39506
rect 23548 39452 23604 39454
rect 23324 39340 23380 39396
rect 22988 38834 23044 38836
rect 22988 38782 22990 38834
rect 22990 38782 23042 38834
rect 23042 38782 23044 38834
rect 22988 38780 23044 38782
rect 23212 38834 23268 38836
rect 23212 38782 23214 38834
rect 23214 38782 23266 38834
rect 23266 38782 23268 38834
rect 23212 38780 23268 38782
rect 23100 37884 23156 37940
rect 23772 38780 23828 38836
rect 22988 37042 23044 37044
rect 22988 36990 22990 37042
rect 22990 36990 23042 37042
rect 23042 36990 23044 37042
rect 22988 36988 23044 36990
rect 22652 35308 22708 35364
rect 22876 35644 22932 35700
rect 22764 35196 22820 35252
rect 23772 37436 23828 37492
rect 23436 37100 23492 37156
rect 23212 34748 23268 34804
rect 23212 34188 23268 34244
rect 22540 34018 22596 34020
rect 22540 33966 22542 34018
rect 22542 33966 22594 34018
rect 22594 33966 22596 34018
rect 22540 33964 22596 33966
rect 23212 33740 23268 33796
rect 22316 33516 22372 33572
rect 22652 33516 22708 33572
rect 22316 32732 22372 32788
rect 22876 33234 22932 33236
rect 22876 33182 22878 33234
rect 22878 33182 22930 33234
rect 22930 33182 22932 33234
rect 22876 33180 22932 33182
rect 22988 32396 23044 32452
rect 23548 35196 23604 35252
rect 23436 35084 23492 35140
rect 23772 35196 23828 35252
rect 23548 33628 23604 33684
rect 23436 33180 23492 33236
rect 23772 33122 23828 33124
rect 23772 33070 23774 33122
rect 23774 33070 23826 33122
rect 23826 33070 23828 33122
rect 23772 33068 23828 33070
rect 22316 30044 22372 30100
rect 22092 29596 22148 29652
rect 22764 31164 22820 31220
rect 22988 30380 23044 30436
rect 25788 45388 25844 45444
rect 25340 41970 25396 41972
rect 25340 41918 25342 41970
rect 25342 41918 25394 41970
rect 25394 41918 25396 41970
rect 25340 41916 25396 41918
rect 25228 41804 25284 41860
rect 25116 41244 25172 41300
rect 24668 40460 24724 40516
rect 24108 39564 24164 39620
rect 23996 39452 24052 39508
rect 24332 38668 24388 38724
rect 23996 37996 24052 38052
rect 24220 37996 24276 38052
rect 24108 37436 24164 37492
rect 24556 39394 24612 39396
rect 24556 39342 24558 39394
rect 24558 39342 24610 39394
rect 24610 39342 24612 39394
rect 24556 39340 24612 39342
rect 24668 38946 24724 38948
rect 24668 38894 24670 38946
rect 24670 38894 24722 38946
rect 24722 38894 24724 38946
rect 24668 38892 24724 38894
rect 24556 38834 24612 38836
rect 24556 38782 24558 38834
rect 24558 38782 24610 38834
rect 24610 38782 24612 38834
rect 24556 38780 24612 38782
rect 25004 39618 25060 39620
rect 25004 39566 25006 39618
rect 25006 39566 25058 39618
rect 25058 39566 25060 39618
rect 25004 39564 25060 39566
rect 24780 38332 24836 38388
rect 24556 37212 24612 37268
rect 24780 37212 24836 37268
rect 25564 41804 25620 41860
rect 25228 40348 25284 40404
rect 25228 38722 25284 38724
rect 25228 38670 25230 38722
rect 25230 38670 25282 38722
rect 25282 38670 25284 38722
rect 25228 38668 25284 38670
rect 25676 41410 25732 41412
rect 25676 41358 25678 41410
rect 25678 41358 25730 41410
rect 25730 41358 25732 41410
rect 25676 41356 25732 41358
rect 25452 41298 25508 41300
rect 25452 41246 25454 41298
rect 25454 41246 25506 41298
rect 25506 41246 25508 41298
rect 25452 41244 25508 41246
rect 26012 45052 26068 45108
rect 26124 45276 26180 45332
rect 26236 44546 26292 44548
rect 26236 44494 26238 44546
rect 26238 44494 26290 44546
rect 26290 44494 26292 44546
rect 26236 44492 26292 44494
rect 25900 44268 25956 44324
rect 28252 50594 28308 50596
rect 28252 50542 28254 50594
rect 28254 50542 28306 50594
rect 28306 50542 28308 50594
rect 28252 50540 28308 50542
rect 28924 50540 28980 50596
rect 28476 50428 28532 50484
rect 31276 53506 31332 53508
rect 31276 53454 31278 53506
rect 31278 53454 31330 53506
rect 31330 53454 31332 53506
rect 31276 53452 31332 53454
rect 29596 51996 29652 52052
rect 29708 52780 29764 52836
rect 30828 52834 30884 52836
rect 30828 52782 30830 52834
rect 30830 52782 30882 52834
rect 30882 52782 30884 52834
rect 30828 52780 30884 52782
rect 30156 52162 30212 52164
rect 30156 52110 30158 52162
rect 30158 52110 30210 52162
rect 30210 52110 30212 52162
rect 30156 52108 30212 52110
rect 30604 51996 30660 52052
rect 30268 51324 30324 51380
rect 29596 50818 29652 50820
rect 29596 50766 29598 50818
rect 29598 50766 29650 50818
rect 29650 50766 29652 50818
rect 29596 50764 29652 50766
rect 30156 50706 30212 50708
rect 30156 50654 30158 50706
rect 30158 50654 30210 50706
rect 30210 50654 30212 50706
rect 30156 50652 30212 50654
rect 29484 50482 29540 50484
rect 29484 50430 29486 50482
rect 29486 50430 29538 50482
rect 29538 50430 29540 50482
rect 29484 50428 29540 50430
rect 29596 50540 29652 50596
rect 28700 49810 28756 49812
rect 28700 49758 28702 49810
rect 28702 49758 28754 49810
rect 28754 49758 28756 49810
rect 28700 49756 28756 49758
rect 29372 49756 29428 49812
rect 27916 49532 27972 49588
rect 30828 51996 30884 52052
rect 32060 53452 32116 53508
rect 31724 53228 31780 53284
rect 31388 52780 31444 52836
rect 30828 50876 30884 50932
rect 31612 51996 31668 52052
rect 31276 50988 31332 51044
rect 31388 51100 31444 51156
rect 31164 50764 31220 50820
rect 30268 50594 30324 50596
rect 30268 50542 30270 50594
rect 30270 50542 30322 50594
rect 30322 50542 30324 50594
rect 30268 50540 30324 50542
rect 29932 50482 29988 50484
rect 29932 50430 29934 50482
rect 29934 50430 29986 50482
rect 29986 50430 29988 50482
rect 29932 50428 29988 50430
rect 30380 50428 30436 50484
rect 29708 49084 29764 49140
rect 28028 48972 28084 49028
rect 27804 47740 27860 47796
rect 27916 48354 27972 48356
rect 27916 48302 27918 48354
rect 27918 48302 27970 48354
rect 27970 48302 27972 48354
rect 27916 48300 27972 48302
rect 28588 48972 28644 49028
rect 29260 49026 29316 49028
rect 29260 48974 29262 49026
rect 29262 48974 29314 49026
rect 29314 48974 29316 49026
rect 29260 48972 29316 48974
rect 29484 48300 29540 48356
rect 27916 47516 27972 47572
rect 28364 48076 28420 48132
rect 28028 47458 28084 47460
rect 28028 47406 28030 47458
rect 28030 47406 28082 47458
rect 28082 47406 28084 47458
rect 28028 47404 28084 47406
rect 28700 47964 28756 48020
rect 27916 47346 27972 47348
rect 27916 47294 27918 47346
rect 27918 47294 27970 47346
rect 27970 47294 27972 47346
rect 27916 47292 27972 47294
rect 29484 47628 29540 47684
rect 29372 47404 29428 47460
rect 29260 46732 29316 46788
rect 29820 47068 29876 47124
rect 31052 50482 31108 50484
rect 31052 50430 31054 50482
rect 31054 50430 31106 50482
rect 31106 50430 31108 50482
rect 31052 50428 31108 50430
rect 30268 47628 30324 47684
rect 30716 47404 30772 47460
rect 29932 46786 29988 46788
rect 29932 46734 29934 46786
rect 29934 46734 29986 46786
rect 29986 46734 29988 46786
rect 29932 46732 29988 46734
rect 30380 46956 30436 47012
rect 29596 46508 29652 46564
rect 29708 46674 29764 46676
rect 29708 46622 29710 46674
rect 29710 46622 29762 46674
rect 29762 46622 29764 46674
rect 29708 46620 29764 46622
rect 28140 45500 28196 45556
rect 30940 46844 30996 46900
rect 31276 46620 31332 46676
rect 26908 43820 26964 43876
rect 26572 43484 26628 43540
rect 26236 42754 26292 42756
rect 26236 42702 26238 42754
rect 26238 42702 26290 42754
rect 26290 42702 26292 42754
rect 26236 42700 26292 42702
rect 25900 41356 25956 41412
rect 26684 43596 26740 43652
rect 27580 44492 27636 44548
rect 27356 43596 27412 43652
rect 26460 43148 26516 43204
rect 25788 41244 25844 41300
rect 26348 39394 26404 39396
rect 26348 39342 26350 39394
rect 26350 39342 26402 39394
rect 26402 39342 26404 39394
rect 26348 39340 26404 39342
rect 26124 38892 26180 38948
rect 26572 37996 26628 38052
rect 25452 37490 25508 37492
rect 25452 37438 25454 37490
rect 25454 37438 25506 37490
rect 25506 37438 25508 37490
rect 25452 37436 25508 37438
rect 25340 37378 25396 37380
rect 25340 37326 25342 37378
rect 25342 37326 25394 37378
rect 25394 37326 25396 37378
rect 25340 37324 25396 37326
rect 25228 37266 25284 37268
rect 25228 37214 25230 37266
rect 25230 37214 25282 37266
rect 25282 37214 25284 37266
rect 25228 37212 25284 37214
rect 25564 37212 25620 37268
rect 24108 35474 24164 35476
rect 24108 35422 24110 35474
rect 24110 35422 24162 35474
rect 24162 35422 24164 35474
rect 24108 35420 24164 35422
rect 23996 34972 24052 35028
rect 24668 36370 24724 36372
rect 24668 36318 24670 36370
rect 24670 36318 24722 36370
rect 24722 36318 24724 36370
rect 24668 36316 24724 36318
rect 24780 34748 24836 34804
rect 23996 33852 24052 33908
rect 24332 34130 24388 34132
rect 24332 34078 24334 34130
rect 24334 34078 24386 34130
rect 24386 34078 24388 34130
rect 24332 34076 24388 34078
rect 24668 34130 24724 34132
rect 24668 34078 24670 34130
rect 24670 34078 24722 34130
rect 24722 34078 24724 34130
rect 24668 34076 24724 34078
rect 23996 32396 24052 32452
rect 24220 32338 24276 32340
rect 24220 32286 24222 32338
rect 24222 32286 24274 32338
rect 24274 32286 24276 32338
rect 24220 32284 24276 32286
rect 23548 31836 23604 31892
rect 23660 30940 23716 30996
rect 21756 28700 21812 28756
rect 21196 26460 21252 26516
rect 20524 26348 20580 26404
rect 20860 26402 20916 26404
rect 20860 26350 20862 26402
rect 20862 26350 20914 26402
rect 20914 26350 20916 26402
rect 20860 26348 20916 26350
rect 20860 26066 20916 26068
rect 20860 26014 20862 26066
rect 20862 26014 20914 26066
rect 20914 26014 20916 26066
rect 20860 26012 20916 26014
rect 20188 25452 20244 25508
rect 19964 25340 20020 25396
rect 20076 25282 20132 25284
rect 20076 25230 20078 25282
rect 20078 25230 20130 25282
rect 20130 25230 20132 25282
rect 20076 25228 20132 25230
rect 20412 25394 20468 25396
rect 20412 25342 20414 25394
rect 20414 25342 20466 25394
rect 20466 25342 20468 25394
rect 20412 25340 20468 25342
rect 21868 26796 21924 26852
rect 22988 28754 23044 28756
rect 22988 28702 22990 28754
rect 22990 28702 23042 28754
rect 23042 28702 23044 28754
rect 22988 28700 23044 28702
rect 22316 28364 22372 28420
rect 21980 26460 22036 26516
rect 21420 26124 21476 26180
rect 21196 25452 21252 25508
rect 19836 25114 19892 25116
rect 19836 25062 19838 25114
rect 19838 25062 19890 25114
rect 19890 25062 19892 25114
rect 19836 25060 19892 25062
rect 19940 25114 19996 25116
rect 19940 25062 19942 25114
rect 19942 25062 19994 25114
rect 19994 25062 19996 25114
rect 19940 25060 19996 25062
rect 20044 25114 20100 25116
rect 20044 25062 20046 25114
rect 20046 25062 20098 25114
rect 20098 25062 20100 25114
rect 20044 25060 20100 25062
rect 20076 24722 20132 24724
rect 20076 24670 20078 24722
rect 20078 24670 20130 24722
rect 20130 24670 20132 24722
rect 20076 24668 20132 24670
rect 19516 24332 19572 24388
rect 19516 23996 19572 24052
rect 20188 23996 20244 24052
rect 20300 23884 20356 23940
rect 19516 23826 19572 23828
rect 19516 23774 19518 23826
rect 19518 23774 19570 23826
rect 19570 23774 19572 23826
rect 19516 23772 19572 23774
rect 19964 23714 20020 23716
rect 19964 23662 19966 23714
rect 19966 23662 20018 23714
rect 20018 23662 20020 23714
rect 19964 23660 20020 23662
rect 19068 23378 19124 23380
rect 19068 23326 19070 23378
rect 19070 23326 19122 23378
rect 19122 23326 19124 23378
rect 19068 23324 19124 23326
rect 18956 21644 19012 21700
rect 19068 23100 19124 23156
rect 19836 23546 19892 23548
rect 19836 23494 19838 23546
rect 19838 23494 19890 23546
rect 19890 23494 19892 23546
rect 19836 23492 19892 23494
rect 19940 23546 19996 23548
rect 19940 23494 19942 23546
rect 19942 23494 19994 23546
rect 19994 23494 19996 23546
rect 19940 23492 19996 23494
rect 20044 23546 20100 23548
rect 20044 23494 20046 23546
rect 20046 23494 20098 23546
rect 20098 23494 20100 23546
rect 20044 23492 20100 23494
rect 19740 23154 19796 23156
rect 19740 23102 19742 23154
rect 19742 23102 19794 23154
rect 19794 23102 19796 23154
rect 19740 23100 19796 23102
rect 19180 21644 19236 21700
rect 20188 22370 20244 22372
rect 20188 22318 20190 22370
rect 20190 22318 20242 22370
rect 20242 22318 20244 22370
rect 20188 22316 20244 22318
rect 19852 22146 19908 22148
rect 19852 22094 19854 22146
rect 19854 22094 19906 22146
rect 19906 22094 19908 22146
rect 19852 22092 19908 22094
rect 19180 21084 19236 21140
rect 19068 20578 19124 20580
rect 19068 20526 19070 20578
rect 19070 20526 19122 20578
rect 19122 20526 19124 20578
rect 19068 20524 19124 20526
rect 19180 20412 19236 20468
rect 18956 19964 19012 20020
rect 18844 19852 18900 19908
rect 18732 19234 18788 19236
rect 18732 19182 18734 19234
rect 18734 19182 18786 19234
rect 18786 19182 18788 19234
rect 18732 19180 18788 19182
rect 18844 19068 18900 19124
rect 18620 18508 18676 18564
rect 18844 17836 18900 17892
rect 18732 17554 18788 17556
rect 18732 17502 18734 17554
rect 18734 17502 18786 17554
rect 18786 17502 18788 17554
rect 18732 17500 18788 17502
rect 18620 16994 18676 16996
rect 18620 16942 18622 16994
rect 18622 16942 18674 16994
rect 18674 16942 18676 16994
rect 18620 16940 18676 16942
rect 18732 16882 18788 16884
rect 18732 16830 18734 16882
rect 18734 16830 18786 16882
rect 18786 16830 18788 16882
rect 18732 16828 18788 16830
rect 18508 15986 18564 15988
rect 18508 15934 18510 15986
rect 18510 15934 18562 15986
rect 18562 15934 18564 15986
rect 18508 15932 18564 15934
rect 18396 15820 18452 15876
rect 16940 13804 16996 13860
rect 16828 13692 16884 13748
rect 16716 13580 16772 13636
rect 16604 12348 16660 12404
rect 16940 12124 16996 12180
rect 16492 11116 16548 11172
rect 16044 10892 16100 10948
rect 15036 10780 15092 10836
rect 5964 9884 6020 9940
rect 4476 8650 4532 8652
rect 4476 8598 4478 8650
rect 4478 8598 4530 8650
rect 4530 8598 4532 8650
rect 4476 8596 4532 8598
rect 4580 8650 4636 8652
rect 4580 8598 4582 8650
rect 4582 8598 4634 8650
rect 4634 8598 4636 8650
rect 4580 8596 4636 8598
rect 4684 8650 4740 8652
rect 4684 8598 4686 8650
rect 4686 8598 4738 8650
rect 4738 8598 4740 8650
rect 4684 8596 4740 8598
rect 16604 10892 16660 10948
rect 18060 14476 18116 14532
rect 17836 13858 17892 13860
rect 17836 13806 17838 13858
rect 17838 13806 17890 13858
rect 17890 13806 17892 13858
rect 17836 13804 17892 13806
rect 18172 13916 18228 13972
rect 17948 13746 18004 13748
rect 17948 13694 17950 13746
rect 17950 13694 18002 13746
rect 18002 13694 18004 13746
rect 17948 13692 18004 13694
rect 18844 15874 18900 15876
rect 18844 15822 18846 15874
rect 18846 15822 18898 15874
rect 18898 15822 18900 15874
rect 18844 15820 18900 15822
rect 18844 15596 18900 15652
rect 19180 19628 19236 19684
rect 19404 20972 19460 21028
rect 19836 21978 19892 21980
rect 19836 21926 19838 21978
rect 19838 21926 19890 21978
rect 19890 21926 19892 21978
rect 19836 21924 19892 21926
rect 19940 21978 19996 21980
rect 19940 21926 19942 21978
rect 19942 21926 19994 21978
rect 19994 21926 19996 21978
rect 19940 21924 19996 21926
rect 20044 21978 20100 21980
rect 20044 21926 20046 21978
rect 20046 21926 20098 21978
rect 20098 21926 20100 21978
rect 20044 21924 20100 21926
rect 20076 21810 20132 21812
rect 20076 21758 20078 21810
rect 20078 21758 20130 21810
rect 20130 21758 20132 21810
rect 20076 21756 20132 21758
rect 19740 21644 19796 21700
rect 19516 20748 19572 20804
rect 19404 20636 19460 20692
rect 19404 17724 19460 17780
rect 19180 17442 19236 17444
rect 19180 17390 19182 17442
rect 19182 17390 19234 17442
rect 19234 17390 19236 17442
rect 19180 17388 19236 17390
rect 19180 15874 19236 15876
rect 19180 15822 19182 15874
rect 19182 15822 19234 15874
rect 19234 15822 19236 15874
rect 19180 15820 19236 15822
rect 19404 17500 19460 17556
rect 19740 20636 19796 20692
rect 20188 21084 20244 21140
rect 20188 20802 20244 20804
rect 20188 20750 20190 20802
rect 20190 20750 20242 20802
rect 20242 20750 20244 20802
rect 20188 20748 20244 20750
rect 19836 20410 19892 20412
rect 19836 20358 19838 20410
rect 19838 20358 19890 20410
rect 19890 20358 19892 20410
rect 19836 20356 19892 20358
rect 19940 20410 19996 20412
rect 19940 20358 19942 20410
rect 19942 20358 19994 20410
rect 19994 20358 19996 20410
rect 19940 20356 19996 20358
rect 20044 20410 20100 20412
rect 20044 20358 20046 20410
rect 20046 20358 20098 20410
rect 20098 20358 20100 20410
rect 20044 20356 20100 20358
rect 19628 20188 19684 20244
rect 19628 19906 19684 19908
rect 19628 19854 19630 19906
rect 19630 19854 19682 19906
rect 19682 19854 19684 19906
rect 19628 19852 19684 19854
rect 20188 20018 20244 20020
rect 20188 19966 20190 20018
rect 20190 19966 20242 20018
rect 20242 19966 20244 20018
rect 20188 19964 20244 19966
rect 20188 19516 20244 19572
rect 19836 18842 19892 18844
rect 19836 18790 19838 18842
rect 19838 18790 19890 18842
rect 19890 18790 19892 18842
rect 19836 18788 19892 18790
rect 19940 18842 19996 18844
rect 19940 18790 19942 18842
rect 19942 18790 19994 18842
rect 19994 18790 19996 18842
rect 19940 18788 19996 18790
rect 20044 18842 20100 18844
rect 20044 18790 20046 18842
rect 20046 18790 20098 18842
rect 20098 18790 20100 18842
rect 20044 18788 20100 18790
rect 19740 17778 19796 17780
rect 19740 17726 19742 17778
rect 19742 17726 19794 17778
rect 19794 17726 19796 17778
rect 19740 17724 19796 17726
rect 20524 24834 20580 24836
rect 20524 24782 20526 24834
rect 20526 24782 20578 24834
rect 20578 24782 20580 24834
rect 20524 24780 20580 24782
rect 20972 24556 21028 24612
rect 20636 23772 20692 23828
rect 20860 24220 20916 24276
rect 20524 22876 20580 22932
rect 20860 22428 20916 22484
rect 20412 22146 20468 22148
rect 20412 22094 20414 22146
rect 20414 22094 20466 22146
rect 20466 22094 20468 22146
rect 20412 22092 20468 22094
rect 23436 28866 23492 28868
rect 23436 28814 23438 28866
rect 23438 28814 23490 28866
rect 23490 28814 23492 28866
rect 23436 28812 23492 28814
rect 24556 32562 24612 32564
rect 24556 32510 24558 32562
rect 24558 32510 24610 32562
rect 24610 32510 24612 32562
rect 24556 32508 24612 32510
rect 25900 37826 25956 37828
rect 25900 37774 25902 37826
rect 25902 37774 25954 37826
rect 25954 37774 25956 37826
rect 25900 37772 25956 37774
rect 26012 37490 26068 37492
rect 26012 37438 26014 37490
rect 26014 37438 26066 37490
rect 26066 37438 26068 37490
rect 26012 37436 26068 37438
rect 26460 37266 26516 37268
rect 26460 37214 26462 37266
rect 26462 37214 26514 37266
rect 26514 37214 26516 37266
rect 26460 37212 26516 37214
rect 25340 35420 25396 35476
rect 25340 35084 25396 35140
rect 25116 35026 25172 35028
rect 25116 34974 25118 35026
rect 25118 34974 25170 35026
rect 25170 34974 25172 35026
rect 25116 34972 25172 34974
rect 25564 34972 25620 35028
rect 26012 34242 26068 34244
rect 26012 34190 26014 34242
rect 26014 34190 26066 34242
rect 26066 34190 26068 34242
rect 26012 34188 26068 34190
rect 25900 34076 25956 34132
rect 25788 33404 25844 33460
rect 25340 32396 25396 32452
rect 25116 32284 25172 32340
rect 24444 31612 24500 31668
rect 24668 31164 24724 31220
rect 24444 31052 24500 31108
rect 23884 30044 23940 30100
rect 23548 28700 23604 28756
rect 23996 29484 24052 29540
rect 24220 30492 24276 30548
rect 25228 31052 25284 31108
rect 25116 30828 25172 30884
rect 24220 30044 24276 30100
rect 24556 30156 24612 30212
rect 24108 28700 24164 28756
rect 23772 28642 23828 28644
rect 23772 28590 23774 28642
rect 23774 28590 23826 28642
rect 23826 28590 23828 28642
rect 23772 28588 23828 28590
rect 24780 29484 24836 29540
rect 24556 29260 24612 29316
rect 23660 28364 23716 28420
rect 24668 28364 24724 28420
rect 23324 28140 23380 28196
rect 24332 28140 24388 28196
rect 22764 28082 22820 28084
rect 22764 28030 22766 28082
rect 22766 28030 22818 28082
rect 22818 28030 22820 28082
rect 22764 28028 22820 28030
rect 23324 27970 23380 27972
rect 23324 27918 23326 27970
rect 23326 27918 23378 27970
rect 23378 27918 23380 27970
rect 23324 27916 23380 27918
rect 22204 26236 22260 26292
rect 21644 25116 21700 25172
rect 21308 24668 21364 24724
rect 21420 24892 21476 24948
rect 21308 23154 21364 23156
rect 21308 23102 21310 23154
rect 21310 23102 21362 23154
rect 21362 23102 21364 23154
rect 21308 23100 21364 23102
rect 20972 21868 21028 21924
rect 21084 22092 21140 22148
rect 20524 21756 20580 21812
rect 21980 25564 22036 25620
rect 21868 25394 21924 25396
rect 21868 25342 21870 25394
rect 21870 25342 21922 25394
rect 21922 25342 21924 25394
rect 21868 25340 21924 25342
rect 21756 24892 21812 24948
rect 21644 23996 21700 24052
rect 21532 23660 21588 23716
rect 21868 23154 21924 23156
rect 21868 23102 21870 23154
rect 21870 23102 21922 23154
rect 21922 23102 21924 23154
rect 21868 23100 21924 23102
rect 22652 25564 22708 25620
rect 23212 25900 23268 25956
rect 22652 25116 22708 25172
rect 22316 24220 22372 24276
rect 22764 24780 22820 24836
rect 22204 23660 22260 23716
rect 22316 23548 22372 23604
rect 22988 25116 23044 25172
rect 23100 25228 23156 25284
rect 22764 23548 22820 23604
rect 22876 23772 22932 23828
rect 24332 27186 24388 27188
rect 24332 27134 24334 27186
rect 24334 27134 24386 27186
rect 24386 27134 24388 27186
rect 24332 27132 24388 27134
rect 23884 26908 23940 26964
rect 23548 26514 23604 26516
rect 23548 26462 23550 26514
rect 23550 26462 23602 26514
rect 23602 26462 23604 26514
rect 23548 26460 23604 26462
rect 23548 25394 23604 25396
rect 23548 25342 23550 25394
rect 23550 25342 23602 25394
rect 23602 25342 23604 25394
rect 23548 25340 23604 25342
rect 24668 26178 24724 26180
rect 24668 26126 24670 26178
rect 24670 26126 24722 26178
rect 24722 26126 24724 26178
rect 24668 26124 24724 26126
rect 23436 25116 23492 25172
rect 24556 25394 24612 25396
rect 24556 25342 24558 25394
rect 24558 25342 24610 25394
rect 24610 25342 24612 25394
rect 24556 25340 24612 25342
rect 25452 32002 25508 32004
rect 25452 31950 25454 32002
rect 25454 31950 25506 32002
rect 25506 31950 25508 32002
rect 25452 31948 25508 31950
rect 25228 26684 25284 26740
rect 25340 27132 25396 27188
rect 24892 26124 24948 26180
rect 24892 25452 24948 25508
rect 24780 25282 24836 25284
rect 24780 25230 24782 25282
rect 24782 25230 24834 25282
rect 24834 25230 24836 25282
rect 24780 25228 24836 25230
rect 26572 34188 26628 34244
rect 27916 44322 27972 44324
rect 27916 44270 27918 44322
rect 27918 44270 27970 44322
rect 27970 44270 27972 44322
rect 27916 44268 27972 44270
rect 28028 43538 28084 43540
rect 28028 43486 28030 43538
rect 28030 43486 28082 43538
rect 28082 43486 28084 43538
rect 28028 43484 28084 43486
rect 29596 45106 29652 45108
rect 29596 45054 29598 45106
rect 29598 45054 29650 45106
rect 29650 45054 29652 45106
rect 29596 45052 29652 45054
rect 29372 44268 29428 44324
rect 27692 43260 27748 43316
rect 29484 43708 29540 43764
rect 29148 43148 29204 43204
rect 27356 42754 27412 42756
rect 27356 42702 27358 42754
rect 27358 42702 27410 42754
rect 27410 42702 27412 42754
rect 27356 42700 27412 42702
rect 27692 41916 27748 41972
rect 28364 42476 28420 42532
rect 27356 40236 27412 40292
rect 27804 41132 27860 41188
rect 27916 40460 27972 40516
rect 28028 40348 28084 40404
rect 27468 39788 27524 39844
rect 27132 39676 27188 39732
rect 30380 45500 30436 45556
rect 30604 43820 30660 43876
rect 29596 43148 29652 43204
rect 30492 43260 30548 43316
rect 29260 41970 29316 41972
rect 29260 41918 29262 41970
rect 29262 41918 29314 41970
rect 29314 41918 29316 41970
rect 29260 41916 29316 41918
rect 28588 41858 28644 41860
rect 28588 41806 28590 41858
rect 28590 41806 28642 41858
rect 28642 41806 28644 41858
rect 28588 41804 28644 41806
rect 29820 41804 29876 41860
rect 28700 41244 28756 41300
rect 28364 40012 28420 40068
rect 28476 40572 28532 40628
rect 27916 39506 27972 39508
rect 27916 39454 27918 39506
rect 27918 39454 27970 39506
rect 27970 39454 27972 39506
rect 27916 39452 27972 39454
rect 27356 39340 27412 39396
rect 28588 39618 28644 39620
rect 28588 39566 28590 39618
rect 28590 39566 28642 39618
rect 28642 39566 28644 39618
rect 28588 39564 28644 39566
rect 28028 39116 28084 39172
rect 26908 37884 26964 37940
rect 26796 37212 26852 37268
rect 27020 36092 27076 36148
rect 27132 34972 27188 35028
rect 26908 33628 26964 33684
rect 26684 33404 26740 33460
rect 26572 33292 26628 33348
rect 26796 32620 26852 32676
rect 26572 32396 26628 32452
rect 26348 31948 26404 32004
rect 26796 31778 26852 31780
rect 26796 31726 26798 31778
rect 26798 31726 26850 31778
rect 26850 31726 26852 31778
rect 26796 31724 26852 31726
rect 25564 30044 25620 30100
rect 27244 30044 27300 30100
rect 25564 28588 25620 28644
rect 26796 29426 26852 29428
rect 26796 29374 26798 29426
rect 26798 29374 26850 29426
rect 26850 29374 26852 29426
rect 26796 29372 26852 29374
rect 26012 29260 26068 29316
rect 28364 38556 28420 38612
rect 28252 38108 28308 38164
rect 28028 37996 28084 38052
rect 27804 37378 27860 37380
rect 27804 37326 27806 37378
rect 27806 37326 27858 37378
rect 27858 37326 27860 37378
rect 27804 37324 27860 37326
rect 27468 37154 27524 37156
rect 27468 37102 27470 37154
rect 27470 37102 27522 37154
rect 27522 37102 27524 37154
rect 27468 37100 27524 37102
rect 27580 34914 27636 34916
rect 27580 34862 27582 34914
rect 27582 34862 27634 34914
rect 27634 34862 27636 34914
rect 27580 34860 27636 34862
rect 28364 36988 28420 37044
rect 28364 36092 28420 36148
rect 28588 35698 28644 35700
rect 28588 35646 28590 35698
rect 28590 35646 28642 35698
rect 28642 35646 28644 35698
rect 28588 35644 28644 35646
rect 29036 41186 29092 41188
rect 29036 41134 29038 41186
rect 29038 41134 29090 41186
rect 29090 41134 29092 41186
rect 29036 41132 29092 41134
rect 28924 40572 28980 40628
rect 29036 40460 29092 40516
rect 29820 40572 29876 40628
rect 29932 41020 29988 41076
rect 29708 40460 29764 40516
rect 30044 40402 30100 40404
rect 30044 40350 30046 40402
rect 30046 40350 30098 40402
rect 30098 40350 30100 40402
rect 30044 40348 30100 40350
rect 28812 39900 28868 39956
rect 29260 39900 29316 39956
rect 30380 39900 30436 39956
rect 28924 39564 28980 39620
rect 29036 39452 29092 39508
rect 30380 39058 30436 39060
rect 30380 39006 30382 39058
rect 30382 39006 30434 39058
rect 30434 39006 30436 39058
rect 30380 39004 30436 39006
rect 29148 38050 29204 38052
rect 29148 37998 29150 38050
rect 29150 37998 29202 38050
rect 29202 37998 29204 38050
rect 29148 37996 29204 37998
rect 29260 36092 29316 36148
rect 29484 37100 29540 37156
rect 29484 36204 29540 36260
rect 28812 35756 28868 35812
rect 28252 33852 28308 33908
rect 27916 33628 27972 33684
rect 27804 33516 27860 33572
rect 27468 31836 27524 31892
rect 27692 32508 27748 32564
rect 27580 29372 27636 29428
rect 27132 28700 27188 28756
rect 25900 28028 25956 28084
rect 25788 26908 25844 26964
rect 25564 26402 25620 26404
rect 25564 26350 25566 26402
rect 25566 26350 25618 26402
rect 25618 26350 25620 26402
rect 25564 26348 25620 26350
rect 25676 25564 25732 25620
rect 23884 24780 23940 24836
rect 24444 24834 24500 24836
rect 24444 24782 24446 24834
rect 24446 24782 24498 24834
rect 24498 24782 24500 24834
rect 24444 24780 24500 24782
rect 24556 24668 24612 24724
rect 23212 24220 23268 24276
rect 23324 23884 23380 23940
rect 23996 24332 24052 24388
rect 23100 23548 23156 23604
rect 23212 23436 23268 23492
rect 23436 23714 23492 23716
rect 23436 23662 23438 23714
rect 23438 23662 23490 23714
rect 23490 23662 23492 23714
rect 23436 23660 23492 23662
rect 21980 22988 22036 23044
rect 21980 21980 22036 22036
rect 25788 25116 25844 25172
rect 26124 27858 26180 27860
rect 26124 27806 26126 27858
rect 26126 27806 26178 27858
rect 26178 27806 26180 27858
rect 26124 27804 26180 27806
rect 26236 27746 26292 27748
rect 26236 27694 26238 27746
rect 26238 27694 26290 27746
rect 26290 27694 26292 27746
rect 26236 27692 26292 27694
rect 26124 27020 26180 27076
rect 26012 26514 26068 26516
rect 26012 26462 26014 26514
rect 26014 26462 26066 26514
rect 26066 26462 26068 26514
rect 26012 26460 26068 26462
rect 26012 25788 26068 25844
rect 26796 26908 26852 26964
rect 26684 26796 26740 26852
rect 27356 28252 27412 28308
rect 27468 28028 27524 28084
rect 26572 26572 26628 26628
rect 27132 26572 27188 26628
rect 26796 25788 26852 25844
rect 24556 23772 24612 23828
rect 24220 23548 24276 23604
rect 22988 22092 23044 22148
rect 22876 21980 22932 22036
rect 23436 21980 23492 22036
rect 21084 21698 21140 21700
rect 21084 21646 21086 21698
rect 21086 21646 21138 21698
rect 21138 21646 21140 21698
rect 21084 21644 21140 21646
rect 20412 20972 20468 21028
rect 20636 21362 20692 21364
rect 20636 21310 20638 21362
rect 20638 21310 20690 21362
rect 20690 21310 20692 21362
rect 20636 21308 20692 21310
rect 21308 21308 21364 21364
rect 20636 21084 20692 21140
rect 20412 20802 20468 20804
rect 20412 20750 20414 20802
rect 20414 20750 20466 20802
rect 20466 20750 20468 20802
rect 20412 20748 20468 20750
rect 21420 21026 21476 21028
rect 21420 20974 21422 21026
rect 21422 20974 21474 21026
rect 21474 20974 21476 21026
rect 21420 20972 21476 20974
rect 21308 20748 21364 20804
rect 21644 21084 21700 21140
rect 21532 20860 21588 20916
rect 20748 20636 20804 20692
rect 21420 20690 21476 20692
rect 21420 20638 21422 20690
rect 21422 20638 21474 20690
rect 21474 20638 21476 20690
rect 21420 20636 21476 20638
rect 23100 21698 23156 21700
rect 23100 21646 23102 21698
rect 23102 21646 23154 21698
rect 23154 21646 23156 21698
rect 23100 21644 23156 21646
rect 22764 21586 22820 21588
rect 22764 21534 22766 21586
rect 22766 21534 22818 21586
rect 22818 21534 22820 21586
rect 22764 21532 22820 21534
rect 22092 20690 22148 20692
rect 22092 20638 22094 20690
rect 22094 20638 22146 20690
rect 22146 20638 22148 20690
rect 22092 20636 22148 20638
rect 21868 20300 21924 20356
rect 20972 20188 21028 20244
rect 20300 19346 20356 19348
rect 20300 19294 20302 19346
rect 20302 19294 20354 19346
rect 20354 19294 20356 19346
rect 20300 19292 20356 19294
rect 20524 17778 20580 17780
rect 20524 17726 20526 17778
rect 20526 17726 20578 17778
rect 20578 17726 20580 17778
rect 20524 17724 20580 17726
rect 19836 17274 19892 17276
rect 19836 17222 19838 17274
rect 19838 17222 19890 17274
rect 19890 17222 19892 17274
rect 19836 17220 19892 17222
rect 19940 17274 19996 17276
rect 19940 17222 19942 17274
rect 19942 17222 19994 17274
rect 19994 17222 19996 17274
rect 19940 17220 19996 17222
rect 20044 17274 20100 17276
rect 20044 17222 20046 17274
rect 20046 17222 20098 17274
rect 20098 17222 20100 17274
rect 20044 17220 20100 17222
rect 20076 17052 20132 17108
rect 20412 16044 20468 16100
rect 21420 19180 21476 19236
rect 22764 20412 22820 20468
rect 21868 20076 21924 20132
rect 21980 19628 22036 19684
rect 22652 20130 22708 20132
rect 22652 20078 22654 20130
rect 22654 20078 22706 20130
rect 22706 20078 22708 20130
rect 22652 20076 22708 20078
rect 22204 19964 22260 20020
rect 22652 19794 22708 19796
rect 22652 19742 22654 19794
rect 22654 19742 22706 19794
rect 22706 19742 22708 19794
rect 22652 19740 22708 19742
rect 21756 19292 21812 19348
rect 22092 19234 22148 19236
rect 22092 19182 22094 19234
rect 22094 19182 22146 19234
rect 22146 19182 22148 19234
rect 22092 19180 22148 19182
rect 21532 18284 21588 18340
rect 21644 17500 21700 17556
rect 21756 17836 21812 17892
rect 21196 16044 21252 16100
rect 21644 16716 21700 16772
rect 21644 16156 21700 16212
rect 20748 15986 20804 15988
rect 20748 15934 20750 15986
rect 20750 15934 20802 15986
rect 20802 15934 20804 15986
rect 20748 15932 20804 15934
rect 19628 15708 19684 15764
rect 19836 15706 19892 15708
rect 19836 15654 19838 15706
rect 19838 15654 19890 15706
rect 19890 15654 19892 15706
rect 19836 15652 19892 15654
rect 19940 15706 19996 15708
rect 19940 15654 19942 15706
rect 19942 15654 19994 15706
rect 19994 15654 19996 15706
rect 19940 15652 19996 15654
rect 20044 15706 20100 15708
rect 20044 15654 20046 15706
rect 20046 15654 20098 15706
rect 20098 15654 20100 15706
rect 20044 15652 20100 15654
rect 20412 15820 20468 15876
rect 19740 15260 19796 15316
rect 19292 15148 19348 15204
rect 17500 12402 17556 12404
rect 17500 12350 17502 12402
rect 17502 12350 17554 12402
rect 17554 12350 17556 12402
rect 17500 12348 17556 12350
rect 18172 12850 18228 12852
rect 18172 12798 18174 12850
rect 18174 12798 18226 12850
rect 18226 12798 18228 12850
rect 18172 12796 18228 12798
rect 17948 12348 18004 12404
rect 17724 11506 17780 11508
rect 17724 11454 17726 11506
rect 17726 11454 17778 11506
rect 17778 11454 17780 11506
rect 17724 11452 17780 11454
rect 17164 10892 17220 10948
rect 17052 10780 17108 10836
rect 17612 10834 17668 10836
rect 17612 10782 17614 10834
rect 17614 10782 17666 10834
rect 17666 10782 17668 10834
rect 17612 10780 17668 10782
rect 16940 10556 16996 10612
rect 16492 9100 16548 9156
rect 4476 7082 4532 7084
rect 4476 7030 4478 7082
rect 4478 7030 4530 7082
rect 4530 7030 4532 7082
rect 4476 7028 4532 7030
rect 4580 7082 4636 7084
rect 4580 7030 4582 7082
rect 4582 7030 4634 7082
rect 4634 7030 4636 7082
rect 4580 7028 4636 7030
rect 4684 7082 4740 7084
rect 4684 7030 4686 7082
rect 4686 7030 4738 7082
rect 4738 7030 4740 7082
rect 4684 7028 4740 7030
rect 17948 12178 18004 12180
rect 17948 12126 17950 12178
rect 17950 12126 18002 12178
rect 18002 12126 18004 12178
rect 17948 12124 18004 12126
rect 18060 11452 18116 11508
rect 18732 13634 18788 13636
rect 18732 13582 18734 13634
rect 18734 13582 18786 13634
rect 18786 13582 18788 13634
rect 18732 13580 18788 13582
rect 18956 13580 19012 13636
rect 20748 15484 20804 15540
rect 21308 15260 21364 15316
rect 22204 18450 22260 18452
rect 22204 18398 22206 18450
rect 22206 18398 22258 18450
rect 22258 18398 22260 18450
rect 22204 18396 22260 18398
rect 22204 17612 22260 17668
rect 21868 17052 21924 17108
rect 22652 19292 22708 19348
rect 23548 21868 23604 21924
rect 25676 23826 25732 23828
rect 25676 23774 25678 23826
rect 25678 23774 25730 23826
rect 25730 23774 25732 23826
rect 25676 23772 25732 23774
rect 25452 23660 25508 23716
rect 25340 23548 25396 23604
rect 25340 23042 25396 23044
rect 25340 22990 25342 23042
rect 25342 22990 25394 23042
rect 25394 22990 25396 23042
rect 25340 22988 25396 22990
rect 25228 22876 25284 22932
rect 23884 22092 23940 22148
rect 24444 22204 24500 22260
rect 23660 21308 23716 21364
rect 23884 21084 23940 21140
rect 23996 21420 24052 21476
rect 23436 20690 23492 20692
rect 23436 20638 23438 20690
rect 23438 20638 23490 20690
rect 23490 20638 23492 20690
rect 23436 20636 23492 20638
rect 23660 20188 23716 20244
rect 22764 17612 22820 17668
rect 22316 16828 22372 16884
rect 21980 16604 22036 16660
rect 21868 15484 21924 15540
rect 19836 14138 19892 14140
rect 19836 14086 19838 14138
rect 19838 14086 19890 14138
rect 19890 14086 19892 14138
rect 19836 14084 19892 14086
rect 19940 14138 19996 14140
rect 19940 14086 19942 14138
rect 19942 14086 19994 14138
rect 19994 14086 19996 14138
rect 19940 14084 19996 14086
rect 20044 14138 20100 14140
rect 20044 14086 20046 14138
rect 20046 14086 20098 14138
rect 20098 14086 20100 14138
rect 20044 14084 20100 14086
rect 19628 13746 19684 13748
rect 19628 13694 19630 13746
rect 19630 13694 19682 13746
rect 19682 13694 19684 13746
rect 19628 13692 19684 13694
rect 19404 13468 19460 13524
rect 19068 12796 19124 12852
rect 18732 12402 18788 12404
rect 18732 12350 18734 12402
rect 18734 12350 18786 12402
rect 18786 12350 18788 12402
rect 18732 12348 18788 12350
rect 20188 13580 20244 13636
rect 19740 12796 19796 12852
rect 20188 13356 20244 13412
rect 19836 12570 19892 12572
rect 19836 12518 19838 12570
rect 19838 12518 19890 12570
rect 19890 12518 19892 12570
rect 19836 12516 19892 12518
rect 19940 12570 19996 12572
rect 19940 12518 19942 12570
rect 19942 12518 19994 12570
rect 19994 12518 19996 12570
rect 19940 12516 19996 12518
rect 20044 12570 20100 12572
rect 20044 12518 20046 12570
rect 20046 12518 20098 12570
rect 20098 12518 20100 12570
rect 20044 12516 20100 12518
rect 19740 12290 19796 12292
rect 19740 12238 19742 12290
rect 19742 12238 19794 12290
rect 19794 12238 19796 12290
rect 19740 12236 19796 12238
rect 18060 11170 18116 11172
rect 18060 11118 18062 11170
rect 18062 11118 18114 11170
rect 18114 11118 18116 11170
rect 18060 11116 18116 11118
rect 18284 10780 18340 10836
rect 18060 10610 18116 10612
rect 18060 10558 18062 10610
rect 18062 10558 18114 10610
rect 18114 10558 18116 10610
rect 18060 10556 18116 10558
rect 18732 11340 18788 11396
rect 17836 8988 17892 9044
rect 17948 9100 18004 9156
rect 17948 8204 18004 8260
rect 17052 7644 17108 7700
rect 18060 7698 18116 7700
rect 18060 7646 18062 7698
rect 18062 7646 18114 7698
rect 18114 7646 18116 7698
rect 18060 7644 18116 7646
rect 18172 7474 18228 7476
rect 18172 7422 18174 7474
rect 18174 7422 18226 7474
rect 18226 7422 18228 7474
rect 18172 7420 18228 7422
rect 16604 7308 16660 7364
rect 17500 7362 17556 7364
rect 17500 7310 17502 7362
rect 17502 7310 17554 7362
rect 17554 7310 17556 7362
rect 17500 7308 17556 7310
rect 18396 9154 18452 9156
rect 18396 9102 18398 9154
rect 18398 9102 18450 9154
rect 18450 9102 18452 9154
rect 18396 9100 18452 9102
rect 18620 10892 18676 10948
rect 18844 12124 18900 12180
rect 19740 11900 19796 11956
rect 20524 14418 20580 14420
rect 20524 14366 20526 14418
rect 20526 14366 20578 14418
rect 20578 14366 20580 14418
rect 20524 14364 20580 14366
rect 20636 13692 20692 13748
rect 21308 13020 21364 13076
rect 20524 12402 20580 12404
rect 20524 12350 20526 12402
rect 20526 12350 20578 12402
rect 20578 12350 20580 12402
rect 20524 12348 20580 12350
rect 20300 12178 20356 12180
rect 20300 12126 20302 12178
rect 20302 12126 20354 12178
rect 20354 12126 20356 12178
rect 20300 12124 20356 12126
rect 20300 11900 20356 11956
rect 18844 11116 18900 11172
rect 19404 11170 19460 11172
rect 19404 11118 19406 11170
rect 19406 11118 19458 11170
rect 19458 11118 19460 11170
rect 19404 11116 19460 11118
rect 19180 10780 19236 10836
rect 19836 11002 19892 11004
rect 19836 10950 19838 11002
rect 19838 10950 19890 11002
rect 19890 10950 19892 11002
rect 19836 10948 19892 10950
rect 19940 11002 19996 11004
rect 19940 10950 19942 11002
rect 19942 10950 19994 11002
rect 19994 10950 19996 11002
rect 19940 10948 19996 10950
rect 20044 11002 20100 11004
rect 20044 10950 20046 11002
rect 20046 10950 20098 11002
rect 20098 10950 20100 11002
rect 20044 10948 20100 10950
rect 18620 9212 18676 9268
rect 19068 9548 19124 9604
rect 19068 9100 19124 9156
rect 19068 8540 19124 8596
rect 18732 8258 18788 8260
rect 18732 8206 18734 8258
rect 18734 8206 18786 8258
rect 18786 8206 18788 8258
rect 18732 8204 18788 8206
rect 18956 8258 19012 8260
rect 18956 8206 18958 8258
rect 18958 8206 19010 8258
rect 19010 8206 19012 8258
rect 18956 8204 19012 8206
rect 18396 7308 18452 7364
rect 15372 6636 15428 6692
rect 16492 6690 16548 6692
rect 16492 6638 16494 6690
rect 16494 6638 16546 6690
rect 16546 6638 16548 6690
rect 16492 6636 16548 6638
rect 4476 5514 4532 5516
rect 4476 5462 4478 5514
rect 4478 5462 4530 5514
rect 4530 5462 4532 5514
rect 4476 5460 4532 5462
rect 4580 5514 4636 5516
rect 4580 5462 4582 5514
rect 4582 5462 4634 5514
rect 4634 5462 4636 5514
rect 4580 5460 4636 5462
rect 4684 5514 4740 5516
rect 4684 5462 4686 5514
rect 4686 5462 4738 5514
rect 4738 5462 4740 5514
rect 4684 5460 4740 5462
rect 19628 10108 19684 10164
rect 19836 9434 19892 9436
rect 19836 9382 19838 9434
rect 19838 9382 19890 9434
rect 19890 9382 19892 9434
rect 19836 9380 19892 9382
rect 19940 9434 19996 9436
rect 19940 9382 19942 9434
rect 19942 9382 19994 9434
rect 19994 9382 19996 9434
rect 19940 9380 19996 9382
rect 20044 9434 20100 9436
rect 20044 9382 20046 9434
rect 20046 9382 20098 9434
rect 20098 9382 20100 9434
rect 20044 9380 20100 9382
rect 19852 9266 19908 9268
rect 19852 9214 19854 9266
rect 19854 9214 19906 9266
rect 19906 9214 19908 9266
rect 19852 9212 19908 9214
rect 19404 6636 19460 6692
rect 19836 7866 19892 7868
rect 19836 7814 19838 7866
rect 19838 7814 19890 7866
rect 19890 7814 19892 7866
rect 19836 7812 19892 7814
rect 19940 7866 19996 7868
rect 19940 7814 19942 7866
rect 19942 7814 19994 7866
rect 19994 7814 19996 7866
rect 19940 7812 19996 7814
rect 20044 7866 20100 7868
rect 20044 7814 20046 7866
rect 20046 7814 20098 7866
rect 20098 7814 20100 7866
rect 20044 7812 20100 7814
rect 20636 11282 20692 11284
rect 20636 11230 20638 11282
rect 20638 11230 20690 11282
rect 20690 11230 20692 11282
rect 20636 11228 20692 11230
rect 21308 12348 21364 12404
rect 21420 11282 21476 11284
rect 21420 11230 21422 11282
rect 21422 11230 21474 11282
rect 21474 11230 21476 11282
rect 21420 11228 21476 11230
rect 20972 10108 21028 10164
rect 20412 9212 20468 9268
rect 21308 9154 21364 9156
rect 21308 9102 21310 9154
rect 21310 9102 21362 9154
rect 21362 9102 21364 9154
rect 21308 9100 21364 9102
rect 20300 8540 20356 8596
rect 19740 6690 19796 6692
rect 19740 6638 19742 6690
rect 19742 6638 19794 6690
rect 19794 6638 19796 6690
rect 19740 6636 19796 6638
rect 19836 6298 19892 6300
rect 19836 6246 19838 6298
rect 19838 6246 19890 6298
rect 19890 6246 19892 6298
rect 19836 6244 19892 6246
rect 19940 6298 19996 6300
rect 19940 6246 19942 6298
rect 19942 6246 19994 6298
rect 19994 6246 19996 6298
rect 19940 6244 19996 6246
rect 20044 6298 20100 6300
rect 20044 6246 20046 6298
rect 20046 6246 20098 6298
rect 20098 6246 20100 6298
rect 20044 6244 20100 6246
rect 18396 5852 18452 5908
rect 18844 5906 18900 5908
rect 18844 5854 18846 5906
rect 18846 5854 18898 5906
rect 18898 5854 18900 5906
rect 18844 5852 18900 5854
rect 18620 5404 18676 5460
rect 16492 5068 16548 5124
rect 17948 5122 18004 5124
rect 17948 5070 17950 5122
rect 17950 5070 18002 5122
rect 18002 5070 18004 5122
rect 17948 5068 18004 5070
rect 19964 5906 20020 5908
rect 19964 5854 19966 5906
rect 19966 5854 20018 5906
rect 20018 5854 20020 5906
rect 19964 5852 20020 5854
rect 21532 10220 21588 10276
rect 21756 11788 21812 11844
rect 21868 11394 21924 11396
rect 21868 11342 21870 11394
rect 21870 11342 21922 11394
rect 21922 11342 21924 11394
rect 21868 11340 21924 11342
rect 22204 16098 22260 16100
rect 22204 16046 22206 16098
rect 22206 16046 22258 16098
rect 22258 16046 22260 16098
rect 22204 16044 22260 16046
rect 22540 17388 22596 17444
rect 23212 18450 23268 18452
rect 23212 18398 23214 18450
rect 23214 18398 23266 18450
rect 23266 18398 23268 18450
rect 23212 18396 23268 18398
rect 23548 18284 23604 18340
rect 23660 18620 23716 18676
rect 23548 17836 23604 17892
rect 22988 16716 23044 16772
rect 23100 17052 23156 17108
rect 23660 17052 23716 17108
rect 24668 21586 24724 21588
rect 24668 21534 24670 21586
rect 24670 21534 24722 21586
rect 24722 21534 24724 21586
rect 24668 21532 24724 21534
rect 24892 20860 24948 20916
rect 23884 20690 23940 20692
rect 23884 20638 23886 20690
rect 23886 20638 23938 20690
rect 23938 20638 23940 20690
rect 23884 20636 23940 20638
rect 24332 20690 24388 20692
rect 24332 20638 24334 20690
rect 24334 20638 24386 20690
rect 24386 20638 24388 20690
rect 24332 20636 24388 20638
rect 25452 22652 25508 22708
rect 26124 24722 26180 24724
rect 26124 24670 26126 24722
rect 26126 24670 26178 24722
rect 26178 24670 26180 24722
rect 26124 24668 26180 24670
rect 28364 33180 28420 33236
rect 28476 33292 28532 33348
rect 28364 32562 28420 32564
rect 28364 32510 28366 32562
rect 28366 32510 28418 32562
rect 28418 32510 28420 32562
rect 28364 32508 28420 32510
rect 27916 31724 27972 31780
rect 28028 31666 28084 31668
rect 28028 31614 28030 31666
rect 28030 31614 28082 31666
rect 28082 31614 28084 31666
rect 28028 31612 28084 31614
rect 28028 30716 28084 30772
rect 27916 30604 27972 30660
rect 28364 31612 28420 31668
rect 28700 34690 28756 34692
rect 28700 34638 28702 34690
rect 28702 34638 28754 34690
rect 28754 34638 28756 34690
rect 28700 34636 28756 34638
rect 29372 35644 29428 35700
rect 29596 35810 29652 35812
rect 29596 35758 29598 35810
rect 29598 35758 29650 35810
rect 29650 35758 29652 35810
rect 29596 35756 29652 35758
rect 29148 35026 29204 35028
rect 29148 34974 29150 35026
rect 29150 34974 29202 35026
rect 29202 34974 29204 35026
rect 29148 34972 29204 34974
rect 30828 43708 30884 43764
rect 31052 44044 31108 44100
rect 32956 53452 33012 53508
rect 33068 53004 33124 53060
rect 33292 54348 33348 54404
rect 32508 51378 32564 51380
rect 32508 51326 32510 51378
rect 32510 51326 32562 51378
rect 32562 51326 32564 51378
rect 32508 51324 32564 51326
rect 32732 50988 32788 51044
rect 32620 50876 32676 50932
rect 32508 50540 32564 50596
rect 33180 50876 33236 50932
rect 33628 55468 33684 55524
rect 33404 53452 33460 53508
rect 33516 53788 33572 53844
rect 34188 55410 34244 55412
rect 34188 55358 34190 55410
rect 34190 55358 34242 55410
rect 34242 55358 34244 55410
rect 34188 55356 34244 55358
rect 33740 53900 33796 53956
rect 32844 49138 32900 49140
rect 32844 49086 32846 49138
rect 32846 49086 32898 49138
rect 32898 49086 32900 49138
rect 32844 49084 32900 49086
rect 31500 49026 31556 49028
rect 31500 48974 31502 49026
rect 31502 48974 31554 49026
rect 31554 48974 31556 49026
rect 31500 48972 31556 48974
rect 31500 47458 31556 47460
rect 31500 47406 31502 47458
rect 31502 47406 31554 47458
rect 31554 47406 31556 47458
rect 31500 47404 31556 47406
rect 32172 47458 32228 47460
rect 32172 47406 32174 47458
rect 32174 47406 32226 47458
rect 32226 47406 32228 47458
rect 32172 47404 32228 47406
rect 33628 52050 33684 52052
rect 33628 51998 33630 52050
rect 33630 51998 33682 52050
rect 33682 51998 33684 52050
rect 33628 51996 33684 51998
rect 33516 50594 33572 50596
rect 33516 50542 33518 50594
rect 33518 50542 33570 50594
rect 33570 50542 33572 50594
rect 33516 50540 33572 50542
rect 34636 53506 34692 53508
rect 34636 53454 34638 53506
rect 34638 53454 34690 53506
rect 34690 53454 34692 53506
rect 34636 53452 34692 53454
rect 34300 53058 34356 53060
rect 34300 53006 34302 53058
rect 34302 53006 34354 53058
rect 34354 53006 34356 53058
rect 34300 53004 34356 53006
rect 34300 52668 34356 52724
rect 38108 57036 38164 57092
rect 36540 56252 36596 56308
rect 35084 56082 35140 56084
rect 35084 56030 35086 56082
rect 35086 56030 35138 56082
rect 35138 56030 35140 56082
rect 35084 56028 35140 56030
rect 35868 56028 35924 56084
rect 35196 55690 35252 55692
rect 35196 55638 35198 55690
rect 35198 55638 35250 55690
rect 35250 55638 35252 55690
rect 35196 55636 35252 55638
rect 35300 55690 35356 55692
rect 35300 55638 35302 55690
rect 35302 55638 35354 55690
rect 35354 55638 35356 55690
rect 35300 55636 35356 55638
rect 35404 55690 35460 55692
rect 35404 55638 35406 55690
rect 35406 55638 35458 55690
rect 35458 55638 35460 55690
rect 35404 55636 35460 55638
rect 34972 54572 35028 54628
rect 38780 56082 38836 56084
rect 38780 56030 38782 56082
rect 38782 56030 38834 56082
rect 38834 56030 38836 56082
rect 38780 56028 38836 56030
rect 38108 55970 38164 55972
rect 38108 55918 38110 55970
rect 38110 55918 38162 55970
rect 38162 55918 38164 55970
rect 38108 55916 38164 55918
rect 35980 55468 36036 55524
rect 37548 55468 37604 55524
rect 35868 54514 35924 54516
rect 35868 54462 35870 54514
rect 35870 54462 35922 54514
rect 35922 54462 35924 54514
rect 35868 54460 35924 54462
rect 35196 54122 35252 54124
rect 35196 54070 35198 54122
rect 35198 54070 35250 54122
rect 35250 54070 35252 54122
rect 35196 54068 35252 54070
rect 35300 54122 35356 54124
rect 35300 54070 35302 54122
rect 35302 54070 35354 54122
rect 35354 54070 35356 54122
rect 35300 54068 35356 54070
rect 35404 54122 35460 54124
rect 35404 54070 35406 54122
rect 35406 54070 35458 54122
rect 35458 54070 35460 54122
rect 35404 54068 35460 54070
rect 35084 53116 35140 53172
rect 34748 52274 34804 52276
rect 34748 52222 34750 52274
rect 34750 52222 34802 52274
rect 34802 52222 34804 52274
rect 34748 52220 34804 52222
rect 34972 52892 35028 52948
rect 34300 52108 34356 52164
rect 35084 52780 35140 52836
rect 35868 52834 35924 52836
rect 35868 52782 35870 52834
rect 35870 52782 35922 52834
rect 35922 52782 35924 52834
rect 35868 52780 35924 52782
rect 35196 52668 35252 52724
rect 35196 52554 35252 52556
rect 35196 52502 35198 52554
rect 35198 52502 35250 52554
rect 35250 52502 35252 52554
rect 35196 52500 35252 52502
rect 35300 52554 35356 52556
rect 35300 52502 35302 52554
rect 35302 52502 35354 52554
rect 35354 52502 35356 52554
rect 35300 52500 35356 52502
rect 35404 52554 35460 52556
rect 35404 52502 35406 52554
rect 35406 52502 35458 52554
rect 35458 52502 35460 52554
rect 35404 52500 35460 52502
rect 35532 52274 35588 52276
rect 35532 52222 35534 52274
rect 35534 52222 35586 52274
rect 35586 52222 35588 52274
rect 35532 52220 35588 52222
rect 36540 54348 36596 54404
rect 37100 54626 37156 54628
rect 37100 54574 37102 54626
rect 37102 54574 37154 54626
rect 37154 54574 37156 54626
rect 37100 54572 37156 54574
rect 37996 55468 38052 55524
rect 38556 55468 38612 55524
rect 37100 53506 37156 53508
rect 37100 53454 37102 53506
rect 37102 53454 37154 53506
rect 37154 53454 37156 53506
rect 37100 53452 37156 53454
rect 36204 52946 36260 52948
rect 36204 52894 36206 52946
rect 36206 52894 36258 52946
rect 36258 52894 36260 52946
rect 36204 52892 36260 52894
rect 37436 53788 37492 53844
rect 38444 54684 38500 54740
rect 37772 54572 37828 54628
rect 37324 53228 37380 53284
rect 37884 54460 37940 54516
rect 38332 54348 38388 54404
rect 37212 53004 37268 53060
rect 37996 53788 38052 53844
rect 37324 52892 37380 52948
rect 36204 52220 36260 52276
rect 35420 51938 35476 51940
rect 35420 51886 35422 51938
rect 35422 51886 35474 51938
rect 35474 51886 35476 51938
rect 35420 51884 35476 51886
rect 35532 51602 35588 51604
rect 35532 51550 35534 51602
rect 35534 51550 35586 51602
rect 35586 51550 35588 51602
rect 35532 51548 35588 51550
rect 35980 52108 36036 52164
rect 36092 51884 36148 51940
rect 35196 50986 35252 50988
rect 35196 50934 35198 50986
rect 35198 50934 35250 50986
rect 35250 50934 35252 50986
rect 35196 50932 35252 50934
rect 35300 50986 35356 50988
rect 35300 50934 35302 50986
rect 35302 50934 35354 50986
rect 35354 50934 35356 50986
rect 35300 50932 35356 50934
rect 35404 50986 35460 50988
rect 35404 50934 35406 50986
rect 35406 50934 35458 50986
rect 35458 50934 35460 50986
rect 35404 50932 35460 50934
rect 33964 50652 34020 50708
rect 35756 50652 35812 50708
rect 33852 50540 33908 50596
rect 33516 49868 33572 49924
rect 34412 50482 34468 50484
rect 34412 50430 34414 50482
rect 34414 50430 34466 50482
rect 34466 50430 34468 50482
rect 34412 50428 34468 50430
rect 34300 50204 34356 50260
rect 34636 50204 34692 50260
rect 33740 49138 33796 49140
rect 33740 49086 33742 49138
rect 33742 49086 33794 49138
rect 33794 49086 33796 49138
rect 33740 49084 33796 49086
rect 34972 50204 35028 50260
rect 35084 50316 35140 50372
rect 34188 49026 34244 49028
rect 34188 48974 34190 49026
rect 34190 48974 34242 49026
rect 34242 48974 34244 49026
rect 34188 48972 34244 48974
rect 35532 49756 35588 49812
rect 35196 49418 35252 49420
rect 35196 49366 35198 49418
rect 35198 49366 35250 49418
rect 35250 49366 35252 49418
rect 35196 49364 35252 49366
rect 35300 49418 35356 49420
rect 35300 49366 35302 49418
rect 35302 49366 35354 49418
rect 35354 49366 35356 49418
rect 35300 49364 35356 49366
rect 35404 49418 35460 49420
rect 35404 49366 35406 49418
rect 35406 49366 35458 49418
rect 35458 49366 35460 49418
rect 35404 49364 35460 49366
rect 35420 49196 35476 49252
rect 33404 48748 33460 48804
rect 35196 47850 35252 47852
rect 35196 47798 35198 47850
rect 35198 47798 35250 47850
rect 35250 47798 35252 47850
rect 35196 47796 35252 47798
rect 35300 47850 35356 47852
rect 35300 47798 35302 47850
rect 35302 47798 35354 47850
rect 35354 47798 35356 47850
rect 35300 47796 35356 47798
rect 35404 47850 35460 47852
rect 35404 47798 35406 47850
rect 35406 47798 35458 47850
rect 35458 47798 35460 47850
rect 35404 47796 35460 47798
rect 34972 47458 35028 47460
rect 34972 47406 34974 47458
rect 34974 47406 35026 47458
rect 35026 47406 35028 47458
rect 34972 47404 35028 47406
rect 33740 47292 33796 47348
rect 33292 46844 33348 46900
rect 32396 45164 32452 45220
rect 31948 45106 32004 45108
rect 31948 45054 31950 45106
rect 31950 45054 32002 45106
rect 32002 45054 32004 45106
rect 31948 45052 32004 45054
rect 31500 44434 31556 44436
rect 31500 44382 31502 44434
rect 31502 44382 31554 44434
rect 31554 44382 31556 44434
rect 31500 44380 31556 44382
rect 33404 45218 33460 45220
rect 33404 45166 33406 45218
rect 33406 45166 33458 45218
rect 33458 45166 33460 45218
rect 33404 45164 33460 45166
rect 32956 44268 33012 44324
rect 31836 44098 31892 44100
rect 31836 44046 31838 44098
rect 31838 44046 31890 44098
rect 31890 44046 31892 44098
rect 31836 44044 31892 44046
rect 34412 46620 34468 46676
rect 34524 46956 34580 47012
rect 33740 45330 33796 45332
rect 33740 45278 33742 45330
rect 33742 45278 33794 45330
rect 33794 45278 33796 45330
rect 33740 45276 33796 45278
rect 33964 45276 34020 45332
rect 33068 43260 33124 43316
rect 30716 41804 30772 41860
rect 32060 42754 32116 42756
rect 32060 42702 32062 42754
rect 32062 42702 32114 42754
rect 32114 42702 32116 42754
rect 32060 42700 32116 42702
rect 33068 42754 33124 42756
rect 33068 42702 33070 42754
rect 33070 42702 33122 42754
rect 33122 42702 33124 42754
rect 33068 42700 33124 42702
rect 33292 42754 33348 42756
rect 33292 42702 33294 42754
rect 33294 42702 33346 42754
rect 33346 42702 33348 42754
rect 33292 42700 33348 42702
rect 32956 42476 33012 42532
rect 31500 41356 31556 41412
rect 31836 42140 31892 42196
rect 31724 40684 31780 40740
rect 30940 40012 30996 40068
rect 30716 39452 30772 39508
rect 33068 41746 33124 41748
rect 33068 41694 33070 41746
rect 33070 41694 33122 41746
rect 33122 41694 33124 41746
rect 33068 41692 33124 41694
rect 32508 41298 32564 41300
rect 32508 41246 32510 41298
rect 32510 41246 32562 41298
rect 32562 41246 32564 41298
rect 32508 41244 32564 41246
rect 32844 41186 32900 41188
rect 32844 41134 32846 41186
rect 32846 41134 32898 41186
rect 32898 41134 32900 41186
rect 32844 41132 32900 41134
rect 33628 42588 33684 42644
rect 33404 41916 33460 41972
rect 33404 41132 33460 41188
rect 33068 41074 33124 41076
rect 33068 41022 33070 41074
rect 33070 41022 33122 41074
rect 33122 41022 33124 41074
rect 33068 41020 33124 41022
rect 33180 40684 33236 40740
rect 30044 37266 30100 37268
rect 30044 37214 30046 37266
rect 30046 37214 30098 37266
rect 30098 37214 30100 37266
rect 30044 37212 30100 37214
rect 31276 39452 31332 39508
rect 31276 39004 31332 39060
rect 30380 36428 30436 36484
rect 29708 34914 29764 34916
rect 29708 34862 29710 34914
rect 29710 34862 29762 34914
rect 29762 34862 29764 34914
rect 29708 34860 29764 34862
rect 29484 34748 29540 34804
rect 29484 33516 29540 33572
rect 29148 33234 29204 33236
rect 29148 33182 29150 33234
rect 29150 33182 29202 33234
rect 29202 33182 29204 33234
rect 29148 33180 29204 33182
rect 29820 33516 29876 33572
rect 29036 32562 29092 32564
rect 29036 32510 29038 32562
rect 29038 32510 29090 32562
rect 29090 32510 29092 32562
rect 29036 32508 29092 32510
rect 29372 32396 29428 32452
rect 30156 33516 30212 33572
rect 29148 31890 29204 31892
rect 29148 31838 29150 31890
rect 29150 31838 29202 31890
rect 29202 31838 29204 31890
rect 29148 31836 29204 31838
rect 29484 31500 29540 31556
rect 28252 30268 28308 30324
rect 28588 30210 28644 30212
rect 28588 30158 28590 30210
rect 28590 30158 28642 30210
rect 28642 30158 28644 30210
rect 28588 30156 28644 30158
rect 28476 30098 28532 30100
rect 28476 30046 28478 30098
rect 28478 30046 28530 30098
rect 28530 30046 28532 30098
rect 28476 30044 28532 30046
rect 27916 29148 27972 29204
rect 28588 29596 28644 29652
rect 27804 28642 27860 28644
rect 27804 28590 27806 28642
rect 27806 28590 27858 28642
rect 27858 28590 27860 28642
rect 27804 28588 27860 28590
rect 27692 28028 27748 28084
rect 27916 28476 27972 28532
rect 27804 27916 27860 27972
rect 27916 27804 27972 27860
rect 28364 27804 28420 27860
rect 28476 27692 28532 27748
rect 28476 27020 28532 27076
rect 28812 28252 28868 28308
rect 28588 26684 28644 26740
rect 27468 25618 27524 25620
rect 27468 25566 27470 25618
rect 27470 25566 27522 25618
rect 27522 25566 27524 25618
rect 27468 25564 27524 25566
rect 27916 26178 27972 26180
rect 27916 26126 27918 26178
rect 27918 26126 27970 26178
rect 27970 26126 27972 26178
rect 27916 26124 27972 26126
rect 28700 26348 28756 26404
rect 27020 25340 27076 25396
rect 26796 25116 26852 25172
rect 27692 24892 27748 24948
rect 26236 23324 26292 23380
rect 25900 22428 25956 22484
rect 25340 21586 25396 21588
rect 25340 21534 25342 21586
rect 25342 21534 25394 21586
rect 25394 21534 25396 21586
rect 25340 21532 25396 21534
rect 25340 20972 25396 21028
rect 25676 21084 25732 21140
rect 24220 19516 24276 19572
rect 25564 19404 25620 19460
rect 25116 19292 25172 19348
rect 23996 18450 24052 18452
rect 23996 18398 23998 18450
rect 23998 18398 24050 18450
rect 24050 18398 24052 18450
rect 23996 18396 24052 18398
rect 23884 18284 23940 18340
rect 24108 17612 24164 17668
rect 24220 19180 24276 19236
rect 23548 15484 23604 15540
rect 22988 15372 23044 15428
rect 22876 14364 22932 14420
rect 24108 15314 24164 15316
rect 24108 15262 24110 15314
rect 24110 15262 24162 15314
rect 24162 15262 24164 15314
rect 24108 15260 24164 15262
rect 23884 15202 23940 15204
rect 23884 15150 23886 15202
rect 23886 15150 23938 15202
rect 23938 15150 23940 15202
rect 23884 15148 23940 15150
rect 25340 19068 25396 19124
rect 24668 18674 24724 18676
rect 24668 18622 24670 18674
rect 24670 18622 24722 18674
rect 24722 18622 24724 18674
rect 24668 18620 24724 18622
rect 25228 18620 25284 18676
rect 24668 18396 24724 18452
rect 25004 18172 25060 18228
rect 25452 18508 25508 18564
rect 28588 24946 28644 24948
rect 28588 24894 28590 24946
rect 28590 24894 28642 24946
rect 28642 24894 28644 24946
rect 28588 24892 28644 24894
rect 28140 23996 28196 24052
rect 28476 24108 28532 24164
rect 28140 23714 28196 23716
rect 28140 23662 28142 23714
rect 28142 23662 28194 23714
rect 28194 23662 28196 23714
rect 28140 23660 28196 23662
rect 27916 23378 27972 23380
rect 27916 23326 27918 23378
rect 27918 23326 27970 23378
rect 27970 23326 27972 23378
rect 27916 23324 27972 23326
rect 27804 22988 27860 23044
rect 28140 22988 28196 23044
rect 28028 22540 28084 22596
rect 26236 22146 26292 22148
rect 26236 22094 26238 22146
rect 26238 22094 26290 22146
rect 26290 22094 26292 22146
rect 26236 22092 26292 22094
rect 26124 21868 26180 21924
rect 27020 21868 27076 21924
rect 26684 21586 26740 21588
rect 26684 21534 26686 21586
rect 26686 21534 26738 21586
rect 26738 21534 26740 21586
rect 26684 21532 26740 21534
rect 26348 21420 26404 21476
rect 26460 21026 26516 21028
rect 26460 20974 26462 21026
rect 26462 20974 26514 21026
rect 26514 20974 26516 21026
rect 26460 20972 26516 20974
rect 27692 21532 27748 21588
rect 28028 21756 28084 21812
rect 28140 21362 28196 21364
rect 28140 21310 28142 21362
rect 28142 21310 28194 21362
rect 28194 21310 28196 21362
rect 28140 21308 28196 21310
rect 27356 20914 27412 20916
rect 27356 20862 27358 20914
rect 27358 20862 27410 20914
rect 27410 20862 27412 20914
rect 27356 20860 27412 20862
rect 26572 20690 26628 20692
rect 26572 20638 26574 20690
rect 26574 20638 26626 20690
rect 26626 20638 26628 20690
rect 26572 20636 26628 20638
rect 26908 20300 26964 20356
rect 25900 19628 25956 19684
rect 26236 19852 26292 19908
rect 25788 19404 25844 19460
rect 26236 19234 26292 19236
rect 26236 19182 26238 19234
rect 26238 19182 26290 19234
rect 26290 19182 26292 19234
rect 26236 19180 26292 19182
rect 25900 18508 25956 18564
rect 26572 18620 26628 18676
rect 26796 19628 26852 19684
rect 26796 18620 26852 18676
rect 28588 22540 28644 22596
rect 28476 21868 28532 21924
rect 28364 20578 28420 20580
rect 28364 20526 28366 20578
rect 28366 20526 28418 20578
rect 28418 20526 28420 20578
rect 28364 20524 28420 20526
rect 27916 19628 27972 19684
rect 27916 19068 27972 19124
rect 26012 17666 26068 17668
rect 26012 17614 26014 17666
rect 26014 17614 26066 17666
rect 26066 17614 26068 17666
rect 26012 17612 26068 17614
rect 26236 17666 26292 17668
rect 26236 17614 26238 17666
rect 26238 17614 26290 17666
rect 26290 17614 26292 17666
rect 26236 17612 26292 17614
rect 26460 17442 26516 17444
rect 26460 17390 26462 17442
rect 26462 17390 26514 17442
rect 26514 17390 26516 17442
rect 26460 17388 26516 17390
rect 26908 17164 26964 17220
rect 25676 16604 25732 16660
rect 23996 13916 24052 13972
rect 23884 13858 23940 13860
rect 23884 13806 23886 13858
rect 23886 13806 23938 13858
rect 23938 13806 23940 13858
rect 23884 13804 23940 13806
rect 22092 13020 22148 13076
rect 22876 13244 22932 13300
rect 22092 12850 22148 12852
rect 22092 12798 22094 12850
rect 22094 12798 22146 12850
rect 22146 12798 22148 12850
rect 22092 12796 22148 12798
rect 22092 10220 22148 10276
rect 22652 9884 22708 9940
rect 21980 9548 22036 9604
rect 21308 6636 21364 6692
rect 20636 6188 20692 6244
rect 20524 5906 20580 5908
rect 20524 5854 20526 5906
rect 20526 5854 20578 5906
rect 20578 5854 20580 5906
rect 20524 5852 20580 5854
rect 20972 6076 21028 6132
rect 21532 6188 21588 6244
rect 22092 9100 22148 9156
rect 22092 7756 22148 7812
rect 22764 7980 22820 8036
rect 22204 7196 22260 7252
rect 21980 6748 22036 6804
rect 21644 6076 21700 6132
rect 21420 5404 21476 5460
rect 21532 5010 21588 5012
rect 21532 4958 21534 5010
rect 21534 4958 21586 5010
rect 21586 4958 21588 5010
rect 21532 4956 21588 4958
rect 19836 4730 19892 4732
rect 19836 4678 19838 4730
rect 19838 4678 19890 4730
rect 19890 4678 19892 4730
rect 19836 4676 19892 4678
rect 19940 4730 19996 4732
rect 19940 4678 19942 4730
rect 19942 4678 19994 4730
rect 19994 4678 19996 4730
rect 19940 4676 19996 4678
rect 20044 4730 20100 4732
rect 20044 4678 20046 4730
rect 20046 4678 20098 4730
rect 20098 4678 20100 4730
rect 20044 4676 20100 4678
rect 24332 13746 24388 13748
rect 24332 13694 24334 13746
rect 24334 13694 24386 13746
rect 24386 13694 24388 13746
rect 24332 13692 24388 13694
rect 24220 13468 24276 13524
rect 25788 15932 25844 15988
rect 25228 15538 25284 15540
rect 25228 15486 25230 15538
rect 25230 15486 25282 15538
rect 25282 15486 25284 15538
rect 25228 15484 25284 15486
rect 24780 15148 24836 15204
rect 25564 15202 25620 15204
rect 25564 15150 25566 15202
rect 25566 15150 25618 15202
rect 25618 15150 25620 15202
rect 25564 15148 25620 15150
rect 24556 13132 24612 13188
rect 24108 12236 24164 12292
rect 23772 12012 23828 12068
rect 23660 11564 23716 11620
rect 23212 11506 23268 11508
rect 23212 11454 23214 11506
rect 23214 11454 23266 11506
rect 23266 11454 23268 11506
rect 23212 11452 23268 11454
rect 22988 11394 23044 11396
rect 22988 11342 22990 11394
rect 22990 11342 23042 11394
rect 23042 11342 23044 11394
rect 22988 11340 23044 11342
rect 23100 10108 23156 10164
rect 24556 12236 24612 12292
rect 24220 11452 24276 11508
rect 25004 14530 25060 14532
rect 25004 14478 25006 14530
rect 25006 14478 25058 14530
rect 25058 14478 25060 14530
rect 25004 14476 25060 14478
rect 25004 14306 25060 14308
rect 25004 14254 25006 14306
rect 25006 14254 25058 14306
rect 25058 14254 25060 14306
rect 25004 14252 25060 14254
rect 25564 13916 25620 13972
rect 25116 13132 25172 13188
rect 25452 13580 25508 13636
rect 26236 15260 26292 15316
rect 26236 15036 26292 15092
rect 26012 14252 26068 14308
rect 25676 13468 25732 13524
rect 25116 12012 25172 12068
rect 25788 13356 25844 13412
rect 24892 11564 24948 11620
rect 25116 11788 25172 11844
rect 23884 11116 23940 11172
rect 23884 10610 23940 10612
rect 23884 10558 23886 10610
rect 23886 10558 23938 10610
rect 23938 10558 23940 10610
rect 23884 10556 23940 10558
rect 23772 9042 23828 9044
rect 23772 8990 23774 9042
rect 23774 8990 23826 9042
rect 23826 8990 23828 9042
rect 23772 8988 23828 8990
rect 24444 9996 24500 10052
rect 24556 10108 24612 10164
rect 24668 9938 24724 9940
rect 24668 9886 24670 9938
rect 24670 9886 24722 9938
rect 24722 9886 24724 9938
rect 24668 9884 24724 9886
rect 24892 8876 24948 8932
rect 22988 8316 23044 8372
rect 23772 8316 23828 8372
rect 23996 8258 24052 8260
rect 23996 8206 23998 8258
rect 23998 8206 24050 8258
rect 24050 8206 24052 8258
rect 23996 8204 24052 8206
rect 23884 8034 23940 8036
rect 23884 7982 23886 8034
rect 23886 7982 23938 8034
rect 23938 7982 23940 8034
rect 23884 7980 23940 7982
rect 23884 7474 23940 7476
rect 23884 7422 23886 7474
rect 23886 7422 23938 7474
rect 23938 7422 23940 7474
rect 23884 7420 23940 7422
rect 22876 7308 22932 7364
rect 24332 8258 24388 8260
rect 24332 8206 24334 8258
rect 24334 8206 24386 8258
rect 24386 8206 24388 8258
rect 24332 8204 24388 8206
rect 25340 12066 25396 12068
rect 25340 12014 25342 12066
rect 25342 12014 25394 12066
rect 25394 12014 25396 12066
rect 25340 12012 25396 12014
rect 25676 13074 25732 13076
rect 25676 13022 25678 13074
rect 25678 13022 25730 13074
rect 25730 13022 25732 13074
rect 25676 13020 25732 13022
rect 25676 12236 25732 12292
rect 26012 13580 26068 13636
rect 26124 13356 26180 13412
rect 25676 11900 25732 11956
rect 25788 11788 25844 11844
rect 25900 12236 25956 12292
rect 25788 11394 25844 11396
rect 25788 11342 25790 11394
rect 25790 11342 25842 11394
rect 25842 11342 25844 11394
rect 25788 11340 25844 11342
rect 25676 11170 25732 11172
rect 25676 11118 25678 11170
rect 25678 11118 25730 11170
rect 25730 11118 25732 11170
rect 25676 11116 25732 11118
rect 25452 10610 25508 10612
rect 25452 10558 25454 10610
rect 25454 10558 25506 10610
rect 25506 10558 25508 10610
rect 25452 10556 25508 10558
rect 26012 11394 26068 11396
rect 26012 11342 26014 11394
rect 26014 11342 26066 11394
rect 26066 11342 26068 11394
rect 26012 11340 26068 11342
rect 26572 15932 26628 15988
rect 26908 16604 26964 16660
rect 27244 16940 27300 16996
rect 27132 16044 27188 16100
rect 26572 15148 26628 15204
rect 26572 13916 26628 13972
rect 27468 15148 27524 15204
rect 27132 15036 27188 15092
rect 26908 14924 26964 14980
rect 26460 13692 26516 13748
rect 26572 13356 26628 13412
rect 26796 12348 26852 12404
rect 26796 11954 26852 11956
rect 26796 11902 26798 11954
rect 26798 11902 26850 11954
rect 26850 11902 26852 11954
rect 26796 11900 26852 11902
rect 26684 11394 26740 11396
rect 26684 11342 26686 11394
rect 26686 11342 26738 11394
rect 26738 11342 26740 11394
rect 26684 11340 26740 11342
rect 26684 11004 26740 11060
rect 26012 10780 26068 10836
rect 26684 10722 26740 10724
rect 26684 10670 26686 10722
rect 26686 10670 26738 10722
rect 26738 10670 26740 10722
rect 26684 10668 26740 10670
rect 25452 10050 25508 10052
rect 25452 9998 25454 10050
rect 25454 9998 25506 10050
rect 25506 9998 25508 10050
rect 25452 9996 25508 9998
rect 25452 9660 25508 9716
rect 26012 9660 26068 9716
rect 25788 8930 25844 8932
rect 25788 8878 25790 8930
rect 25790 8878 25842 8930
rect 25842 8878 25844 8930
rect 25788 8876 25844 8878
rect 25004 7980 25060 8036
rect 24220 7474 24276 7476
rect 24220 7422 24222 7474
rect 24222 7422 24274 7474
rect 24274 7422 24276 7474
rect 24220 7420 24276 7422
rect 22540 6636 22596 6692
rect 22428 6300 22484 6356
rect 22988 6690 23044 6692
rect 22988 6638 22990 6690
rect 22990 6638 23042 6690
rect 23042 6638 23044 6690
rect 22988 6636 23044 6638
rect 22540 6076 22596 6132
rect 22876 5180 22932 5236
rect 22204 4956 22260 5012
rect 4476 3946 4532 3948
rect 4476 3894 4478 3946
rect 4478 3894 4530 3946
rect 4530 3894 4532 3946
rect 4476 3892 4532 3894
rect 4580 3946 4636 3948
rect 4580 3894 4582 3946
rect 4582 3894 4634 3946
rect 4634 3894 4636 3946
rect 4580 3892 4636 3894
rect 4684 3946 4740 3948
rect 4684 3894 4686 3946
rect 4686 3894 4738 3946
rect 4738 3894 4740 3946
rect 4684 3892 4740 3894
rect 23772 6860 23828 6916
rect 23324 6636 23380 6692
rect 23436 6466 23492 6468
rect 23436 6414 23438 6466
rect 23438 6414 23490 6466
rect 23490 6414 23492 6466
rect 23436 6412 23492 6414
rect 24332 6636 24388 6692
rect 24892 7308 24948 7364
rect 24668 6578 24724 6580
rect 24668 6526 24670 6578
rect 24670 6526 24722 6578
rect 24722 6526 24724 6578
rect 24668 6524 24724 6526
rect 23660 6300 23716 6356
rect 23324 5740 23380 5796
rect 23324 5122 23380 5124
rect 23324 5070 23326 5122
rect 23326 5070 23378 5122
rect 23378 5070 23380 5122
rect 23324 5068 23380 5070
rect 24108 5122 24164 5124
rect 24108 5070 24110 5122
rect 24110 5070 24162 5122
rect 24162 5070 24164 5122
rect 24108 5068 24164 5070
rect 25452 8258 25508 8260
rect 25452 8206 25454 8258
rect 25454 8206 25506 8258
rect 25506 8206 25508 8258
rect 25452 8204 25508 8206
rect 25228 7420 25284 7476
rect 25116 6802 25172 6804
rect 25116 6750 25118 6802
rect 25118 6750 25170 6802
rect 25170 6750 25172 6802
rect 25116 6748 25172 6750
rect 25900 7532 25956 7588
rect 25340 7308 25396 7364
rect 25788 6914 25844 6916
rect 25788 6862 25790 6914
rect 25790 6862 25842 6914
rect 25842 6862 25844 6914
rect 25788 6860 25844 6862
rect 27916 15202 27972 15204
rect 27916 15150 27918 15202
rect 27918 15150 27970 15202
rect 27970 15150 27972 15202
rect 27916 15148 27972 15150
rect 28140 17612 28196 17668
rect 28140 17442 28196 17444
rect 28140 17390 28142 17442
rect 28142 17390 28194 17442
rect 28194 17390 28196 17442
rect 28140 17388 28196 17390
rect 28364 18284 28420 18340
rect 28700 21474 28756 21476
rect 28700 21422 28702 21474
rect 28702 21422 28754 21474
rect 28754 21422 28756 21474
rect 28700 21420 28756 21422
rect 29036 30322 29092 30324
rect 29036 30270 29038 30322
rect 29038 30270 29090 30322
rect 29090 30270 29092 30322
rect 29036 30268 29092 30270
rect 29596 31164 29652 31220
rect 30380 31276 30436 31332
rect 29820 30156 29876 30212
rect 29148 29708 29204 29764
rect 29708 29932 29764 29988
rect 29372 29372 29428 29428
rect 29148 29148 29204 29204
rect 29372 28588 29428 28644
rect 29036 27692 29092 27748
rect 29372 27244 29428 27300
rect 29708 29538 29764 29540
rect 29708 29486 29710 29538
rect 29710 29486 29762 29538
rect 29762 29486 29764 29538
rect 29708 29484 29764 29486
rect 29932 29932 29988 29988
rect 29932 29708 29988 29764
rect 30044 29484 30100 29540
rect 30716 37154 30772 37156
rect 30716 37102 30718 37154
rect 30718 37102 30770 37154
rect 30770 37102 30772 37154
rect 30716 37100 30772 37102
rect 30716 36258 30772 36260
rect 30716 36206 30718 36258
rect 30718 36206 30770 36258
rect 30770 36206 30772 36258
rect 30716 36204 30772 36206
rect 31164 38556 31220 38612
rect 30940 37996 30996 38052
rect 30940 36540 30996 36596
rect 30604 33516 30660 33572
rect 30492 30210 30548 30212
rect 30492 30158 30494 30210
rect 30494 30158 30546 30210
rect 30546 30158 30548 30210
rect 30492 30156 30548 30158
rect 30604 31052 30660 31108
rect 31724 39228 31780 39284
rect 31836 39004 31892 39060
rect 32060 40460 32116 40516
rect 32172 40124 32228 40180
rect 31948 38780 32004 38836
rect 32060 39340 32116 39396
rect 31836 38556 31892 38612
rect 32396 40236 32452 40292
rect 33852 44322 33908 44324
rect 33852 44270 33854 44322
rect 33854 44270 33906 44322
rect 33906 44270 33908 44322
rect 33852 44268 33908 44270
rect 34748 46898 34804 46900
rect 34748 46846 34750 46898
rect 34750 46846 34802 46898
rect 34802 46846 34804 46898
rect 34748 46844 34804 46846
rect 34636 46732 34692 46788
rect 34300 45388 34356 45444
rect 34412 45330 34468 45332
rect 34412 45278 34414 45330
rect 34414 45278 34466 45330
rect 34466 45278 34468 45330
rect 34412 45276 34468 45278
rect 35196 47068 35252 47124
rect 35308 46786 35364 46788
rect 35308 46734 35310 46786
rect 35310 46734 35362 46786
rect 35362 46734 35364 46786
rect 35308 46732 35364 46734
rect 34748 45948 34804 46004
rect 34860 46060 34916 46116
rect 35532 47404 35588 47460
rect 35420 46450 35476 46452
rect 35420 46398 35422 46450
rect 35422 46398 35474 46450
rect 35474 46398 35476 46450
rect 35420 46396 35476 46398
rect 37100 52780 37156 52836
rect 36988 51490 37044 51492
rect 36988 51438 36990 51490
rect 36990 51438 37042 51490
rect 37042 51438 37044 51490
rect 36988 51436 37044 51438
rect 37660 52946 37716 52948
rect 37660 52894 37662 52946
rect 37662 52894 37714 52946
rect 37714 52894 37716 52946
rect 37660 52892 37716 52894
rect 37436 52162 37492 52164
rect 37436 52110 37438 52162
rect 37438 52110 37490 52162
rect 37490 52110 37492 52162
rect 37436 52108 37492 52110
rect 38444 53730 38500 53732
rect 38444 53678 38446 53730
rect 38446 53678 38498 53730
rect 38498 53678 38500 53730
rect 38444 53676 38500 53678
rect 38892 54684 38948 54740
rect 38668 53788 38724 53844
rect 38332 52892 38388 52948
rect 38220 52220 38276 52276
rect 38108 52108 38164 52164
rect 39340 55692 39396 55748
rect 40796 56306 40852 56308
rect 40796 56254 40798 56306
rect 40798 56254 40850 56306
rect 40850 56254 40852 56306
rect 40796 56252 40852 56254
rect 41132 56028 41188 56084
rect 39452 54572 39508 54628
rect 39676 54514 39732 54516
rect 39676 54462 39678 54514
rect 39678 54462 39730 54514
rect 39730 54462 39732 54514
rect 39676 54460 39732 54462
rect 39228 54348 39284 54404
rect 39116 53676 39172 53732
rect 39004 52556 39060 52612
rect 39116 52162 39172 52164
rect 39116 52110 39118 52162
rect 39118 52110 39170 52162
rect 39170 52110 39172 52162
rect 39116 52108 39172 52110
rect 38556 51996 38612 52052
rect 37660 51602 37716 51604
rect 37660 51550 37662 51602
rect 37662 51550 37714 51602
rect 37714 51550 37716 51602
rect 37660 51548 37716 51550
rect 37100 50818 37156 50820
rect 37100 50766 37102 50818
rect 37102 50766 37154 50818
rect 37154 50766 37156 50818
rect 37100 50764 37156 50766
rect 36876 50652 36932 50708
rect 37548 50706 37604 50708
rect 37548 50654 37550 50706
rect 37550 50654 37602 50706
rect 37602 50654 37604 50706
rect 37548 50652 37604 50654
rect 36316 50482 36372 50484
rect 36316 50430 36318 50482
rect 36318 50430 36370 50482
rect 36370 50430 36372 50482
rect 36316 50428 36372 50430
rect 38108 51490 38164 51492
rect 38108 51438 38110 51490
rect 38110 51438 38162 51490
rect 38162 51438 38164 51490
rect 38108 51436 38164 51438
rect 36988 50482 37044 50484
rect 36988 50430 36990 50482
rect 36990 50430 37042 50482
rect 37042 50430 37044 50482
rect 36988 50428 37044 50430
rect 35980 50204 36036 50260
rect 36764 50204 36820 50260
rect 35868 49980 35924 50036
rect 36652 50034 36708 50036
rect 36652 49982 36654 50034
rect 36654 49982 36706 50034
rect 36706 49982 36708 50034
rect 36652 49980 36708 49982
rect 36316 49810 36372 49812
rect 36316 49758 36318 49810
rect 36318 49758 36370 49810
rect 36370 49758 36372 49810
rect 36316 49756 36372 49758
rect 35980 49698 36036 49700
rect 35980 49646 35982 49698
rect 35982 49646 36034 49698
rect 36034 49646 36036 49698
rect 35980 49644 36036 49646
rect 35980 49250 36036 49252
rect 35980 49198 35982 49250
rect 35982 49198 36034 49250
rect 36034 49198 36036 49250
rect 35980 49196 36036 49198
rect 36988 49084 37044 49140
rect 37100 49532 37156 49588
rect 37436 49420 37492 49476
rect 35756 47292 35812 47348
rect 36764 48972 36820 49028
rect 36092 48914 36148 48916
rect 36092 48862 36094 48914
rect 36094 48862 36146 48914
rect 36146 48862 36148 48914
rect 36092 48860 36148 48862
rect 37100 48860 37156 48916
rect 38108 50204 38164 50260
rect 38220 49698 38276 49700
rect 38220 49646 38222 49698
rect 38222 49646 38274 49698
rect 38274 49646 38276 49698
rect 38220 49644 38276 49646
rect 37772 49084 37828 49140
rect 35196 46282 35252 46284
rect 35196 46230 35198 46282
rect 35198 46230 35250 46282
rect 35250 46230 35252 46282
rect 35196 46228 35252 46230
rect 35300 46282 35356 46284
rect 35300 46230 35302 46282
rect 35302 46230 35354 46282
rect 35354 46230 35356 46282
rect 35300 46228 35356 46230
rect 35404 46282 35460 46284
rect 35404 46230 35406 46282
rect 35406 46230 35458 46282
rect 35458 46230 35460 46282
rect 35404 46228 35460 46230
rect 35196 45948 35252 46004
rect 37212 48748 37268 48804
rect 36316 47068 36372 47124
rect 36428 47292 36484 47348
rect 35868 46060 35924 46116
rect 36092 46396 36148 46452
rect 35756 45276 35812 45332
rect 35196 44714 35252 44716
rect 35196 44662 35198 44714
rect 35198 44662 35250 44714
rect 35250 44662 35252 44714
rect 35196 44660 35252 44662
rect 35300 44714 35356 44716
rect 35300 44662 35302 44714
rect 35302 44662 35354 44714
rect 35354 44662 35356 44714
rect 35300 44660 35356 44662
rect 35404 44714 35460 44716
rect 35404 44662 35406 44714
rect 35406 44662 35458 44714
rect 35458 44662 35460 44714
rect 35404 44660 35460 44662
rect 34748 44380 34804 44436
rect 37212 47346 37268 47348
rect 37212 47294 37214 47346
rect 37214 47294 37266 47346
rect 37266 47294 37268 47346
rect 37212 47292 37268 47294
rect 37100 46956 37156 47012
rect 36988 46562 37044 46564
rect 36988 46510 36990 46562
rect 36990 46510 37042 46562
rect 37042 46510 37044 46562
rect 36988 46508 37044 46510
rect 36876 45948 36932 46004
rect 36316 45836 36372 45892
rect 36764 45836 36820 45892
rect 36316 43650 36372 43652
rect 36316 43598 36318 43650
rect 36318 43598 36370 43650
rect 36370 43598 36372 43650
rect 36316 43596 36372 43598
rect 34076 42754 34132 42756
rect 34076 42702 34078 42754
rect 34078 42702 34130 42754
rect 34130 42702 34132 42754
rect 34076 42700 34132 42702
rect 34300 42530 34356 42532
rect 34300 42478 34302 42530
rect 34302 42478 34354 42530
rect 34354 42478 34356 42530
rect 34300 42476 34356 42478
rect 34524 42252 34580 42308
rect 33852 41804 33908 41860
rect 33852 41244 33908 41300
rect 33852 40908 33908 40964
rect 33516 40572 33572 40628
rect 33628 40460 33684 40516
rect 33292 39676 33348 39732
rect 32396 39340 32452 39396
rect 33292 39228 33348 39284
rect 33516 39228 33572 39284
rect 33180 39058 33236 39060
rect 33180 39006 33182 39058
rect 33182 39006 33234 39058
rect 33234 39006 33236 39058
rect 33180 39004 33236 39006
rect 33964 40460 34020 40516
rect 33740 39340 33796 39396
rect 33068 38780 33124 38836
rect 31164 36428 31220 36484
rect 34412 40572 34468 40628
rect 34524 41692 34580 41748
rect 34748 42028 34804 42084
rect 35196 43146 35252 43148
rect 35196 43094 35198 43146
rect 35198 43094 35250 43146
rect 35250 43094 35252 43146
rect 35196 43092 35252 43094
rect 35300 43146 35356 43148
rect 35300 43094 35302 43146
rect 35302 43094 35354 43146
rect 35354 43094 35356 43146
rect 35300 43092 35356 43094
rect 35404 43146 35460 43148
rect 35404 43094 35406 43146
rect 35406 43094 35458 43146
rect 35458 43094 35460 43146
rect 35404 43092 35460 43094
rect 36316 42476 36372 42532
rect 35196 41970 35252 41972
rect 35196 41918 35198 41970
rect 35198 41918 35250 41970
rect 35250 41918 35252 41970
rect 35196 41916 35252 41918
rect 35196 41578 35252 41580
rect 35196 41526 35198 41578
rect 35198 41526 35250 41578
rect 35250 41526 35252 41578
rect 35196 41524 35252 41526
rect 35300 41578 35356 41580
rect 35300 41526 35302 41578
rect 35302 41526 35354 41578
rect 35354 41526 35356 41578
rect 35300 41524 35356 41526
rect 35404 41578 35460 41580
rect 35404 41526 35406 41578
rect 35406 41526 35458 41578
rect 35458 41526 35460 41578
rect 35404 41524 35460 41526
rect 37212 46060 37268 46116
rect 36988 43596 37044 43652
rect 36876 43538 36932 43540
rect 36876 43486 36878 43538
rect 36878 43486 36930 43538
rect 36930 43486 36932 43538
rect 36876 43484 36932 43486
rect 37548 47682 37604 47684
rect 37548 47630 37550 47682
rect 37550 47630 37602 47682
rect 37602 47630 37604 47682
rect 37548 47628 37604 47630
rect 38332 48972 38388 49028
rect 38444 47628 38500 47684
rect 38220 46956 38276 47012
rect 39452 53228 39508 53284
rect 40460 55020 40516 55076
rect 39788 53116 39844 53172
rect 40012 54460 40068 54516
rect 40124 53676 40180 53732
rect 38780 51266 38836 51268
rect 38780 51214 38782 51266
rect 38782 51214 38834 51266
rect 38834 51214 38836 51266
rect 38780 51212 38836 51214
rect 38668 49532 38724 49588
rect 39340 51660 39396 51716
rect 39228 51602 39284 51604
rect 39228 51550 39230 51602
rect 39230 51550 39282 51602
rect 39282 51550 39284 51602
rect 39228 51548 39284 51550
rect 39228 50764 39284 50820
rect 40236 53564 40292 53620
rect 41020 54626 41076 54628
rect 41020 54574 41022 54626
rect 41022 54574 41074 54626
rect 41074 54574 41076 54626
rect 41020 54572 41076 54574
rect 41468 55356 41524 55412
rect 42364 55132 42420 55188
rect 41468 54402 41524 54404
rect 41468 54350 41470 54402
rect 41470 54350 41522 54402
rect 41522 54350 41524 54402
rect 41468 54348 41524 54350
rect 42364 54796 42420 54852
rect 40908 53340 40964 53396
rect 41692 53564 41748 53620
rect 41468 53452 41524 53508
rect 41916 53170 41972 53172
rect 41916 53118 41918 53170
rect 41918 53118 41970 53170
rect 41970 53118 41972 53170
rect 41916 53116 41972 53118
rect 39004 49756 39060 49812
rect 39788 51378 39844 51380
rect 39788 51326 39790 51378
rect 39790 51326 39842 51378
rect 39842 51326 39844 51378
rect 39788 51324 39844 51326
rect 39676 51212 39732 51268
rect 40124 50316 40180 50372
rect 39116 49532 39172 49588
rect 39452 49420 39508 49476
rect 39004 49138 39060 49140
rect 39004 49086 39006 49138
rect 39006 49086 39058 49138
rect 39058 49086 39060 49138
rect 39004 49084 39060 49086
rect 38892 47964 38948 48020
rect 38780 46956 38836 47012
rect 38332 45164 38388 45220
rect 38556 46508 38612 46564
rect 38108 45052 38164 45108
rect 38220 44940 38276 44996
rect 39564 48018 39620 48020
rect 39564 47966 39566 48018
rect 39566 47966 39618 48018
rect 39618 47966 39620 48018
rect 39564 47964 39620 47966
rect 39564 47404 39620 47460
rect 39116 46508 39172 46564
rect 39228 46284 39284 46340
rect 40460 51660 40516 51716
rect 41692 52220 41748 52276
rect 42588 55074 42644 55076
rect 42588 55022 42590 55074
rect 42590 55022 42642 55074
rect 42642 55022 42644 55074
rect 42588 55020 42644 55022
rect 42476 54460 42532 54516
rect 41468 51660 41524 51716
rect 41356 51548 41412 51604
rect 41244 51490 41300 51492
rect 41244 51438 41246 51490
rect 41246 51438 41298 51490
rect 41298 51438 41300 51490
rect 41244 51436 41300 51438
rect 40796 51324 40852 51380
rect 40460 50428 40516 50484
rect 40236 49084 40292 49140
rect 40012 48354 40068 48356
rect 40012 48302 40014 48354
rect 40014 48302 40066 48354
rect 40066 48302 40068 48354
rect 40012 48300 40068 48302
rect 39788 47516 39844 47572
rect 39564 46284 39620 46340
rect 38668 45330 38724 45332
rect 38668 45278 38670 45330
rect 38670 45278 38722 45330
rect 38722 45278 38724 45330
rect 38668 45276 38724 45278
rect 38556 45218 38612 45220
rect 38556 45166 38558 45218
rect 38558 45166 38610 45218
rect 38610 45166 38612 45218
rect 38556 45164 38612 45166
rect 38780 45164 38836 45220
rect 39116 45106 39172 45108
rect 39116 45054 39118 45106
rect 39118 45054 39170 45106
rect 39170 45054 39172 45106
rect 39116 45052 39172 45054
rect 37324 43650 37380 43652
rect 37324 43598 37326 43650
rect 37326 43598 37378 43650
rect 37378 43598 37380 43650
rect 37324 43596 37380 43598
rect 37548 43708 37604 43764
rect 37100 42530 37156 42532
rect 37100 42478 37102 42530
rect 37102 42478 37154 42530
rect 37154 42478 37156 42530
rect 37100 42476 37156 42478
rect 37212 42140 37268 42196
rect 36764 41804 36820 41860
rect 36540 41692 36596 41748
rect 37212 41356 37268 41412
rect 34636 40684 34692 40740
rect 34972 40908 35028 40964
rect 34748 40460 34804 40516
rect 34188 39788 34244 39844
rect 34076 39676 34132 39732
rect 33964 38946 34020 38948
rect 33964 38894 33966 38946
rect 33966 38894 34018 38946
rect 34018 38894 34020 38946
rect 33964 38892 34020 38894
rect 32396 38050 32452 38052
rect 32396 37998 32398 38050
rect 32398 37998 32450 38050
rect 32450 37998 32452 38050
rect 32396 37996 32452 37998
rect 33628 38050 33684 38052
rect 33628 37998 33630 38050
rect 33630 37998 33682 38050
rect 33682 37998 33684 38050
rect 33628 37996 33684 37998
rect 33068 37772 33124 37828
rect 32172 37212 32228 37268
rect 32508 37266 32564 37268
rect 32508 37214 32510 37266
rect 32510 37214 32562 37266
rect 32562 37214 32564 37266
rect 32508 37212 32564 37214
rect 32956 36988 33012 37044
rect 32172 36540 32228 36596
rect 31164 35698 31220 35700
rect 31164 35646 31166 35698
rect 31166 35646 31218 35698
rect 31218 35646 31220 35698
rect 31164 35644 31220 35646
rect 30828 34860 30884 34916
rect 31276 34300 31332 34356
rect 30828 34188 30884 34244
rect 31948 34354 32004 34356
rect 31948 34302 31950 34354
rect 31950 34302 32002 34354
rect 32002 34302 32004 34354
rect 31948 34300 32004 34302
rect 31836 34242 31892 34244
rect 31836 34190 31838 34242
rect 31838 34190 31890 34242
rect 31890 34190 31892 34242
rect 31836 34188 31892 34190
rect 30828 33852 30884 33908
rect 31052 33852 31108 33908
rect 31948 33906 32004 33908
rect 31948 33854 31950 33906
rect 31950 33854 32002 33906
rect 32002 33854 32004 33906
rect 31948 33852 32004 33854
rect 31164 33404 31220 33460
rect 30940 31724 30996 31780
rect 31836 32620 31892 32676
rect 33404 37826 33460 37828
rect 33404 37774 33406 37826
rect 33406 37774 33458 37826
rect 33458 37774 33460 37826
rect 33404 37772 33460 37774
rect 33404 36988 33460 37044
rect 33964 37772 34020 37828
rect 34076 37996 34132 38052
rect 33852 37212 33908 37268
rect 33180 36540 33236 36596
rect 33628 36428 33684 36484
rect 33628 35532 33684 35588
rect 33180 34300 33236 34356
rect 33292 34076 33348 34132
rect 32508 33628 32564 33684
rect 32284 33346 32340 33348
rect 32284 33294 32286 33346
rect 32286 33294 32338 33346
rect 32338 33294 32340 33346
rect 32284 33292 32340 33294
rect 32396 32562 32452 32564
rect 32396 32510 32398 32562
rect 32398 32510 32450 32562
rect 32450 32510 32452 32562
rect 32396 32508 32452 32510
rect 31164 31388 31220 31444
rect 30380 29596 30436 29652
rect 30156 28924 30212 28980
rect 30380 29260 30436 29316
rect 30380 28700 30436 28756
rect 30156 28530 30212 28532
rect 30156 28478 30158 28530
rect 30158 28478 30210 28530
rect 30210 28478 30212 28530
rect 30156 28476 30212 28478
rect 30156 28028 30212 28084
rect 29708 27858 29764 27860
rect 29708 27806 29710 27858
rect 29710 27806 29762 27858
rect 29762 27806 29764 27858
rect 29708 27804 29764 27806
rect 29148 27074 29204 27076
rect 29148 27022 29150 27074
rect 29150 27022 29202 27074
rect 29202 27022 29204 27074
rect 29148 27020 29204 27022
rect 29260 26290 29316 26292
rect 29260 26238 29262 26290
rect 29262 26238 29314 26290
rect 29314 26238 29316 26290
rect 29260 26236 29316 26238
rect 30044 26012 30100 26068
rect 29036 24668 29092 24724
rect 29596 24722 29652 24724
rect 29596 24670 29598 24722
rect 29598 24670 29650 24722
rect 29650 24670 29652 24722
rect 29596 24668 29652 24670
rect 29260 24556 29316 24612
rect 29036 23042 29092 23044
rect 29036 22990 29038 23042
rect 29038 22990 29090 23042
rect 29090 22990 29092 23042
rect 29036 22988 29092 22990
rect 29708 24556 29764 24612
rect 29708 24108 29764 24164
rect 29484 22988 29540 23044
rect 29148 22428 29204 22484
rect 29372 22540 29428 22596
rect 30604 28642 30660 28644
rect 30604 28590 30606 28642
rect 30606 28590 30658 28642
rect 30658 28590 30660 28642
rect 30604 28588 30660 28590
rect 30716 27804 30772 27860
rect 31388 31276 31444 31332
rect 31164 30268 31220 30324
rect 31276 30044 31332 30100
rect 31052 29986 31108 29988
rect 31052 29934 31054 29986
rect 31054 29934 31106 29986
rect 31106 29934 31108 29986
rect 31052 29932 31108 29934
rect 30940 29372 30996 29428
rect 31052 29596 31108 29652
rect 30940 29148 30996 29204
rect 31164 29484 31220 29540
rect 31500 30268 31556 30324
rect 31836 29596 31892 29652
rect 31948 30210 32004 30212
rect 31948 30158 31950 30210
rect 31950 30158 32002 30210
rect 32002 30158 32004 30210
rect 31948 30156 32004 30158
rect 31500 29314 31556 29316
rect 31500 29262 31502 29314
rect 31502 29262 31554 29314
rect 31554 29262 31556 29314
rect 31500 29260 31556 29262
rect 31948 29148 32004 29204
rect 32060 29036 32116 29092
rect 32172 31948 32228 32004
rect 33180 33458 33236 33460
rect 33180 33406 33182 33458
rect 33182 33406 33234 33458
rect 33234 33406 33236 33458
rect 33180 33404 33236 33406
rect 32732 33346 32788 33348
rect 32732 33294 32734 33346
rect 32734 33294 32786 33346
rect 32786 33294 32788 33346
rect 32732 33292 32788 33294
rect 33404 33516 33460 33572
rect 34524 37100 34580 37156
rect 34748 36370 34804 36372
rect 34748 36318 34750 36370
rect 34750 36318 34802 36370
rect 34802 36318 34804 36370
rect 34748 36316 34804 36318
rect 34412 35586 34468 35588
rect 34412 35534 34414 35586
rect 34414 35534 34466 35586
rect 34466 35534 34468 35586
rect 34412 35532 34468 35534
rect 33852 34188 33908 34244
rect 33404 32338 33460 32340
rect 33404 32286 33406 32338
rect 33406 32286 33458 32338
rect 33458 32286 33460 32338
rect 33404 32284 33460 32286
rect 33180 31948 33236 32004
rect 34524 34130 34580 34132
rect 34524 34078 34526 34130
rect 34526 34078 34578 34130
rect 34578 34078 34580 34130
rect 34524 34076 34580 34078
rect 33740 33292 33796 33348
rect 33740 32732 33796 32788
rect 33852 33404 33908 33460
rect 34748 33404 34804 33460
rect 33964 33292 34020 33348
rect 33516 31948 33572 32004
rect 33628 32396 33684 32452
rect 34076 32396 34132 32452
rect 34860 32396 34916 32452
rect 34524 32338 34580 32340
rect 34524 32286 34526 32338
rect 34526 32286 34578 32338
rect 34578 32286 34580 32338
rect 34524 32284 34580 32286
rect 32508 31164 32564 31220
rect 32396 31106 32452 31108
rect 32396 31054 32398 31106
rect 32398 31054 32450 31106
rect 32450 31054 32452 31106
rect 32396 31052 32452 31054
rect 33404 30828 33460 30884
rect 32396 30770 32452 30772
rect 32396 30718 32398 30770
rect 32398 30718 32450 30770
rect 32450 30718 32452 30770
rect 32396 30716 32452 30718
rect 32396 30044 32452 30100
rect 32284 29708 32340 29764
rect 32508 29426 32564 29428
rect 32508 29374 32510 29426
rect 32510 29374 32562 29426
rect 32562 29374 32564 29426
rect 32508 29372 32564 29374
rect 33516 30380 33572 30436
rect 33964 31554 34020 31556
rect 33964 31502 33966 31554
rect 33966 31502 34018 31554
rect 34018 31502 34020 31554
rect 33964 31500 34020 31502
rect 34188 31276 34244 31332
rect 33964 31052 34020 31108
rect 32844 30210 32900 30212
rect 32844 30158 32846 30210
rect 32846 30158 32898 30210
rect 32898 30158 32900 30210
rect 32844 30156 32900 30158
rect 33964 30156 34020 30212
rect 33180 29820 33236 29876
rect 33516 29708 33572 29764
rect 32956 29484 33012 29540
rect 31276 28140 31332 28196
rect 31836 27970 31892 27972
rect 31836 27918 31838 27970
rect 31838 27918 31890 27970
rect 31890 27918 31892 27970
rect 31836 27916 31892 27918
rect 31164 27692 31220 27748
rect 31276 27186 31332 27188
rect 31276 27134 31278 27186
rect 31278 27134 31330 27186
rect 31330 27134 31332 27186
rect 31276 27132 31332 27134
rect 32508 27858 32564 27860
rect 32508 27806 32510 27858
rect 32510 27806 32562 27858
rect 32562 27806 32564 27858
rect 32508 27804 32564 27806
rect 32508 27580 32564 27636
rect 32172 27356 32228 27412
rect 30492 26572 30548 26628
rect 30492 24722 30548 24724
rect 30492 24670 30494 24722
rect 30494 24670 30546 24722
rect 30546 24670 30548 24722
rect 30492 24668 30548 24670
rect 32172 26572 32228 26628
rect 32508 26402 32564 26404
rect 32508 26350 32510 26402
rect 32510 26350 32562 26402
rect 32562 26350 32564 26402
rect 32508 26348 32564 26350
rect 30716 26236 30772 26292
rect 32620 26236 32676 26292
rect 32396 26066 32452 26068
rect 32396 26014 32398 26066
rect 32398 26014 32450 26066
rect 32450 26014 32452 26066
rect 32396 26012 32452 26014
rect 31612 25676 31668 25732
rect 30156 22988 30212 23044
rect 30940 24220 30996 24276
rect 29932 22092 29988 22148
rect 30940 23772 30996 23828
rect 30828 23714 30884 23716
rect 30828 23662 30830 23714
rect 30830 23662 30882 23714
rect 30882 23662 30884 23714
rect 30828 23660 30884 23662
rect 30604 22988 30660 23044
rect 30492 22146 30548 22148
rect 30492 22094 30494 22146
rect 30494 22094 30546 22146
rect 30546 22094 30548 22146
rect 30492 22092 30548 22094
rect 30828 21868 30884 21924
rect 30268 21644 30324 21700
rect 29596 21084 29652 21140
rect 29260 20636 29316 20692
rect 28924 19852 28980 19908
rect 29036 20524 29092 20580
rect 29036 18732 29092 18788
rect 29148 18620 29204 18676
rect 28476 17836 28532 17892
rect 28588 17724 28644 17780
rect 28924 17724 28980 17780
rect 28476 17554 28532 17556
rect 28476 17502 28478 17554
rect 28478 17502 28530 17554
rect 28530 17502 28532 17554
rect 28476 17500 28532 17502
rect 28364 16940 28420 16996
rect 29148 17554 29204 17556
rect 29148 17502 29150 17554
rect 29150 17502 29202 17554
rect 29202 17502 29204 17554
rect 29148 17500 29204 17502
rect 29260 17388 29316 17444
rect 29708 19740 29764 19796
rect 31276 23996 31332 24052
rect 32396 24610 32452 24612
rect 32396 24558 32398 24610
rect 32398 24558 32450 24610
rect 32450 24558 32452 24610
rect 32396 24556 32452 24558
rect 31836 23996 31892 24052
rect 31612 23938 31668 23940
rect 31612 23886 31614 23938
rect 31614 23886 31666 23938
rect 31666 23886 31668 23938
rect 31612 23884 31668 23886
rect 32060 23826 32116 23828
rect 32060 23774 32062 23826
rect 32062 23774 32114 23826
rect 32114 23774 32116 23826
rect 32060 23772 32116 23774
rect 31164 23042 31220 23044
rect 31164 22990 31166 23042
rect 31166 22990 31218 23042
rect 31218 22990 31220 23042
rect 31164 22988 31220 22990
rect 31052 21698 31108 21700
rect 31052 21646 31054 21698
rect 31054 21646 31106 21698
rect 31106 21646 31108 21698
rect 31052 21644 31108 21646
rect 32284 23884 32340 23940
rect 31388 21868 31444 21924
rect 31612 21756 31668 21812
rect 31388 21532 31444 21588
rect 31500 20636 31556 20692
rect 30156 19740 30212 19796
rect 30380 19404 30436 19460
rect 30268 18732 30324 18788
rect 29820 17724 29876 17780
rect 30044 18284 30100 18340
rect 29372 17276 29428 17332
rect 29708 17276 29764 17332
rect 27692 13634 27748 13636
rect 27692 13582 27694 13634
rect 27694 13582 27746 13634
rect 27746 13582 27748 13634
rect 27692 13580 27748 13582
rect 27020 13468 27076 13524
rect 27580 13468 27636 13524
rect 27132 13356 27188 13412
rect 27132 11228 27188 11284
rect 27132 10108 27188 10164
rect 27468 10444 27524 10500
rect 26572 9714 26628 9716
rect 26572 9662 26574 9714
rect 26574 9662 26626 9714
rect 26626 9662 26628 9714
rect 26572 9660 26628 9662
rect 26124 6690 26180 6692
rect 26124 6638 26126 6690
rect 26126 6638 26178 6690
rect 26178 6638 26180 6690
rect 26124 6636 26180 6638
rect 26012 6524 26068 6580
rect 24668 6130 24724 6132
rect 24668 6078 24670 6130
rect 24670 6078 24722 6130
rect 24722 6078 24724 6130
rect 24668 6076 24724 6078
rect 24780 5628 24836 5684
rect 25004 5234 25060 5236
rect 25004 5182 25006 5234
rect 25006 5182 25058 5234
rect 25058 5182 25060 5234
rect 25004 5180 25060 5182
rect 25564 6300 25620 6356
rect 25340 6076 25396 6132
rect 26012 5906 26068 5908
rect 26012 5854 26014 5906
rect 26014 5854 26066 5906
rect 26066 5854 26068 5906
rect 26012 5852 26068 5854
rect 26236 5852 26292 5908
rect 25452 5794 25508 5796
rect 25452 5742 25454 5794
rect 25454 5742 25506 5794
rect 25506 5742 25508 5794
rect 25452 5740 25508 5742
rect 26348 5794 26404 5796
rect 26348 5742 26350 5794
rect 26350 5742 26402 5794
rect 26402 5742 26404 5794
rect 26348 5740 26404 5742
rect 25452 5516 25508 5572
rect 26460 5516 26516 5572
rect 25564 4956 25620 5012
rect 26684 8316 26740 8372
rect 27020 7698 27076 7700
rect 27020 7646 27022 7698
rect 27022 7646 27074 7698
rect 27074 7646 27076 7698
rect 27020 7644 27076 7646
rect 27804 13356 27860 13412
rect 27692 13132 27748 13188
rect 28252 13468 28308 13524
rect 27916 12236 27972 12292
rect 27804 11394 27860 11396
rect 27804 11342 27806 11394
rect 27806 11342 27858 11394
rect 27858 11342 27860 11394
rect 27804 11340 27860 11342
rect 27804 10108 27860 10164
rect 29596 14642 29652 14644
rect 29596 14590 29598 14642
rect 29598 14590 29650 14642
rect 29650 14590 29652 14642
rect 29596 14588 29652 14590
rect 29372 12796 29428 12852
rect 29596 12572 29652 12628
rect 28476 12290 28532 12292
rect 28476 12238 28478 12290
rect 28478 12238 28530 12290
rect 28530 12238 28532 12290
rect 28476 12236 28532 12238
rect 28364 11394 28420 11396
rect 28364 11342 28366 11394
rect 28366 11342 28418 11394
rect 28418 11342 28420 11394
rect 28364 11340 28420 11342
rect 29148 11788 29204 11844
rect 30156 16882 30212 16884
rect 30156 16830 30158 16882
rect 30158 16830 30210 16882
rect 30210 16830 30212 16882
rect 30156 16828 30212 16830
rect 30492 19292 30548 19348
rect 31052 19292 31108 19348
rect 31276 19292 31332 19348
rect 31388 17554 31444 17556
rect 31388 17502 31390 17554
rect 31390 17502 31442 17554
rect 31442 17502 31444 17554
rect 31388 17500 31444 17502
rect 31164 17442 31220 17444
rect 31164 17390 31166 17442
rect 31166 17390 31218 17442
rect 31218 17390 31220 17442
rect 31164 17388 31220 17390
rect 30492 16716 30548 16772
rect 31724 20018 31780 20020
rect 31724 19966 31726 20018
rect 31726 19966 31778 20018
rect 31778 19966 31780 20018
rect 31724 19964 31780 19966
rect 32172 22204 32228 22260
rect 32060 21644 32116 21700
rect 32172 19964 32228 20020
rect 32060 19346 32116 19348
rect 32060 19294 32062 19346
rect 32062 19294 32114 19346
rect 32114 19294 32116 19346
rect 32060 19292 32116 19294
rect 32508 20636 32564 20692
rect 32060 18732 32116 18788
rect 33292 29426 33348 29428
rect 33292 29374 33294 29426
rect 33294 29374 33346 29426
rect 33346 29374 33348 29426
rect 33292 29372 33348 29374
rect 33404 29036 33460 29092
rect 32956 28924 33012 28980
rect 33068 28252 33124 28308
rect 33180 27692 33236 27748
rect 33292 27580 33348 27636
rect 32956 27356 33012 27412
rect 33628 29932 33684 29988
rect 33740 29372 33796 29428
rect 33964 29986 34020 29988
rect 33964 29934 33966 29986
rect 33966 29934 34018 29986
rect 34018 29934 34020 29986
rect 33964 29932 34020 29934
rect 34076 29426 34132 29428
rect 34076 29374 34078 29426
rect 34078 29374 34130 29426
rect 34130 29374 34132 29426
rect 34076 29372 34132 29374
rect 33516 28812 33572 28868
rect 34188 28754 34244 28756
rect 34188 28702 34190 28754
rect 34190 28702 34242 28754
rect 34242 28702 34244 28754
rect 34188 28700 34244 28702
rect 34076 28140 34132 28196
rect 33628 27916 33684 27972
rect 36988 41186 37044 41188
rect 36988 41134 36990 41186
rect 36990 41134 37042 41186
rect 37042 41134 37044 41186
rect 36988 41132 37044 41134
rect 35756 41020 35812 41076
rect 37100 41074 37156 41076
rect 37100 41022 37102 41074
rect 37102 41022 37154 41074
rect 37154 41022 37156 41074
rect 37100 41020 37156 41022
rect 39228 44828 39284 44884
rect 37772 43650 37828 43652
rect 37772 43598 37774 43650
rect 37774 43598 37826 43650
rect 37826 43598 37828 43650
rect 37772 43596 37828 43598
rect 40012 45164 40068 45220
rect 39564 44994 39620 44996
rect 39564 44942 39566 44994
rect 39566 44942 39618 44994
rect 39618 44942 39620 44994
rect 39564 44940 39620 44942
rect 39676 44380 39732 44436
rect 38444 43372 38500 43428
rect 38220 42754 38276 42756
rect 38220 42702 38222 42754
rect 38222 42702 38274 42754
rect 38274 42702 38276 42754
rect 38220 42700 38276 42702
rect 38108 42530 38164 42532
rect 38108 42478 38110 42530
rect 38110 42478 38162 42530
rect 38162 42478 38164 42530
rect 38108 42476 38164 42478
rect 38780 43484 38836 43540
rect 39004 43538 39060 43540
rect 39004 43486 39006 43538
rect 39006 43486 39058 43538
rect 39058 43486 39060 43538
rect 39004 43484 39060 43486
rect 38556 43260 38612 43316
rect 38780 42924 38836 42980
rect 38556 42476 38612 42532
rect 37660 41074 37716 41076
rect 37660 41022 37662 41074
rect 37662 41022 37714 41074
rect 37714 41022 37716 41074
rect 37660 41020 37716 41022
rect 35756 40514 35812 40516
rect 35756 40462 35758 40514
rect 35758 40462 35810 40514
rect 35810 40462 35812 40514
rect 35756 40460 35812 40462
rect 36428 40572 36484 40628
rect 35308 40348 35364 40404
rect 35756 40236 35812 40292
rect 35196 40010 35252 40012
rect 35196 39958 35198 40010
rect 35198 39958 35250 40010
rect 35250 39958 35252 40010
rect 35196 39956 35252 39958
rect 35300 40010 35356 40012
rect 35300 39958 35302 40010
rect 35302 39958 35354 40010
rect 35354 39958 35356 40010
rect 35300 39956 35356 39958
rect 35404 40010 35460 40012
rect 35404 39958 35406 40010
rect 35406 39958 35458 40010
rect 35458 39958 35460 40010
rect 35404 39956 35460 39958
rect 35644 39842 35700 39844
rect 35644 39790 35646 39842
rect 35646 39790 35698 39842
rect 35698 39790 35700 39842
rect 35644 39788 35700 39790
rect 35308 39730 35364 39732
rect 35308 39678 35310 39730
rect 35310 39678 35362 39730
rect 35362 39678 35364 39730
rect 35308 39676 35364 39678
rect 36540 40402 36596 40404
rect 36540 40350 36542 40402
rect 36542 40350 36594 40402
rect 36594 40350 36596 40402
rect 36540 40348 36596 40350
rect 35196 38442 35252 38444
rect 35196 38390 35198 38442
rect 35198 38390 35250 38442
rect 35250 38390 35252 38442
rect 35196 38388 35252 38390
rect 35300 38442 35356 38444
rect 35300 38390 35302 38442
rect 35302 38390 35354 38442
rect 35354 38390 35356 38442
rect 35300 38388 35356 38390
rect 35404 38442 35460 38444
rect 35404 38390 35406 38442
rect 35406 38390 35458 38442
rect 35458 38390 35460 38442
rect 35404 38388 35460 38390
rect 35084 37100 35140 37156
rect 35196 36874 35252 36876
rect 35196 36822 35198 36874
rect 35198 36822 35250 36874
rect 35250 36822 35252 36874
rect 35196 36820 35252 36822
rect 35300 36874 35356 36876
rect 35300 36822 35302 36874
rect 35302 36822 35354 36874
rect 35354 36822 35356 36874
rect 35300 36820 35356 36822
rect 35404 36874 35460 36876
rect 35404 36822 35406 36874
rect 35406 36822 35458 36874
rect 35458 36822 35460 36874
rect 35404 36820 35460 36822
rect 35644 37100 35700 37156
rect 35980 39228 36036 39284
rect 36428 39394 36484 39396
rect 36428 39342 36430 39394
rect 36430 39342 36482 39394
rect 36482 39342 36484 39394
rect 36428 39340 36484 39342
rect 37100 40290 37156 40292
rect 37100 40238 37102 40290
rect 37102 40238 37154 40290
rect 37154 40238 37156 40290
rect 37100 40236 37156 40238
rect 36988 37548 37044 37604
rect 35308 36370 35364 36372
rect 35308 36318 35310 36370
rect 35310 36318 35362 36370
rect 35362 36318 35364 36370
rect 35308 36316 35364 36318
rect 35868 36316 35924 36372
rect 36316 36370 36372 36372
rect 36316 36318 36318 36370
rect 36318 36318 36370 36370
rect 36370 36318 36372 36370
rect 36316 36316 36372 36318
rect 36204 36258 36260 36260
rect 36204 36206 36206 36258
rect 36206 36206 36258 36258
rect 36258 36206 36260 36258
rect 36204 36204 36260 36206
rect 36540 35644 36596 35700
rect 35196 35306 35252 35308
rect 35196 35254 35198 35306
rect 35198 35254 35250 35306
rect 35250 35254 35252 35306
rect 35196 35252 35252 35254
rect 35300 35306 35356 35308
rect 35300 35254 35302 35306
rect 35302 35254 35354 35306
rect 35354 35254 35356 35306
rect 35300 35252 35356 35254
rect 35404 35306 35460 35308
rect 35404 35254 35406 35306
rect 35406 35254 35458 35306
rect 35458 35254 35460 35306
rect 35404 35252 35460 35254
rect 36092 34636 36148 34692
rect 35084 34130 35140 34132
rect 35084 34078 35086 34130
rect 35086 34078 35138 34130
rect 35138 34078 35140 34130
rect 35084 34076 35140 34078
rect 35196 33738 35252 33740
rect 35196 33686 35198 33738
rect 35198 33686 35250 33738
rect 35250 33686 35252 33738
rect 35196 33684 35252 33686
rect 35300 33738 35356 33740
rect 35300 33686 35302 33738
rect 35302 33686 35354 33738
rect 35354 33686 35356 33738
rect 35300 33684 35356 33686
rect 35404 33738 35460 33740
rect 35404 33686 35406 33738
rect 35406 33686 35458 33738
rect 35458 33686 35460 33738
rect 35404 33684 35460 33686
rect 35756 32786 35812 32788
rect 35756 32734 35758 32786
rect 35758 32734 35810 32786
rect 35810 32734 35812 32786
rect 35756 32732 35812 32734
rect 35532 32508 35588 32564
rect 35196 32170 35252 32172
rect 35196 32118 35198 32170
rect 35198 32118 35250 32170
rect 35250 32118 35252 32170
rect 35196 32116 35252 32118
rect 35300 32170 35356 32172
rect 35300 32118 35302 32170
rect 35302 32118 35354 32170
rect 35354 32118 35356 32170
rect 35300 32116 35356 32118
rect 35404 32170 35460 32172
rect 35404 32118 35406 32170
rect 35406 32118 35458 32170
rect 35458 32118 35460 32170
rect 35404 32116 35460 32118
rect 36540 32172 36596 32228
rect 35756 31948 35812 32004
rect 34636 31052 34692 31108
rect 35308 31724 35364 31780
rect 34524 30098 34580 30100
rect 34524 30046 34526 30098
rect 34526 30046 34578 30098
rect 34578 30046 34580 30098
rect 34524 30044 34580 30046
rect 34972 31554 35028 31556
rect 34972 31502 34974 31554
rect 34974 31502 35026 31554
rect 35026 31502 35028 31554
rect 34972 31500 35028 31502
rect 36652 31948 36708 32004
rect 36988 36316 37044 36372
rect 38444 41074 38500 41076
rect 38444 41022 38446 41074
rect 38446 41022 38498 41074
rect 38498 41022 38500 41074
rect 38444 41020 38500 41022
rect 38332 40962 38388 40964
rect 38332 40910 38334 40962
rect 38334 40910 38386 40962
rect 38386 40910 38388 40962
rect 38332 40908 38388 40910
rect 37436 40402 37492 40404
rect 37436 40350 37438 40402
rect 37438 40350 37490 40402
rect 37490 40350 37492 40402
rect 37436 40348 37492 40350
rect 37548 39506 37604 39508
rect 37548 39454 37550 39506
rect 37550 39454 37602 39506
rect 37602 39454 37604 39506
rect 37548 39452 37604 39454
rect 37996 39506 38052 39508
rect 37996 39454 37998 39506
rect 37998 39454 38050 39506
rect 38050 39454 38052 39506
rect 37996 39452 38052 39454
rect 39004 42754 39060 42756
rect 39004 42702 39006 42754
rect 39006 42702 39058 42754
rect 39058 42702 39060 42754
rect 39004 42700 39060 42702
rect 39228 42924 39284 42980
rect 39340 42140 39396 42196
rect 38780 41468 38836 41524
rect 39116 41804 39172 41860
rect 38780 41186 38836 41188
rect 38780 41134 38782 41186
rect 38782 41134 38834 41186
rect 38834 41134 38836 41186
rect 38780 41132 38836 41134
rect 38668 40908 38724 40964
rect 39340 41468 39396 41524
rect 38892 40348 38948 40404
rect 38556 38892 38612 38948
rect 39004 39900 39060 39956
rect 40348 48242 40404 48244
rect 40348 48190 40350 48242
rect 40350 48190 40402 48242
rect 40402 48190 40404 48242
rect 40348 48188 40404 48190
rect 42028 51436 42084 51492
rect 42028 50706 42084 50708
rect 42028 50654 42030 50706
rect 42030 50654 42082 50706
rect 42082 50654 42084 50706
rect 42028 50652 42084 50654
rect 42252 54348 42308 54404
rect 42924 55970 42980 55972
rect 42924 55918 42926 55970
rect 42926 55918 42978 55970
rect 42978 55918 42980 55970
rect 42924 55916 42980 55918
rect 43260 55468 43316 55524
rect 44604 57036 44660 57092
rect 42812 54572 42868 54628
rect 42812 53788 42868 53844
rect 43036 55186 43092 55188
rect 43036 55134 43038 55186
rect 43038 55134 43090 55186
rect 43090 55134 43092 55186
rect 43036 55132 43092 55134
rect 42700 53506 42756 53508
rect 42700 53454 42702 53506
rect 42702 53454 42754 53506
rect 42754 53454 42756 53506
rect 42700 53452 42756 53454
rect 42364 52220 42420 52276
rect 43260 55356 43316 55412
rect 43372 54796 43428 54852
rect 43596 55468 43652 55524
rect 43708 55132 43764 55188
rect 43484 54684 43540 54740
rect 43596 55020 43652 55076
rect 43148 53228 43204 53284
rect 44044 55916 44100 55972
rect 44940 55186 44996 55188
rect 44940 55134 44942 55186
rect 44942 55134 44994 55186
rect 44994 55134 44996 55186
rect 44940 55132 44996 55134
rect 44828 55074 44884 55076
rect 44828 55022 44830 55074
rect 44830 55022 44882 55074
rect 44882 55022 44884 55074
rect 44828 55020 44884 55022
rect 44268 54796 44324 54852
rect 44716 54514 44772 54516
rect 44716 54462 44718 54514
rect 44718 54462 44770 54514
rect 44770 54462 44772 54514
rect 44716 54460 44772 54462
rect 44268 53676 44324 53732
rect 44828 54012 44884 54068
rect 44044 53452 44100 53508
rect 43820 53004 43876 53060
rect 44156 53340 44212 53396
rect 43596 52780 43652 52836
rect 43484 52050 43540 52052
rect 43484 51998 43486 52050
rect 43486 51998 43538 52050
rect 43538 51998 43540 52050
rect 43484 51996 43540 51998
rect 42924 51938 42980 51940
rect 42924 51886 42926 51938
rect 42926 51886 42978 51938
rect 42978 51886 42980 51938
rect 42924 51884 42980 51886
rect 42364 51212 42420 51268
rect 41580 50316 41636 50372
rect 41468 50204 41524 50260
rect 42140 49922 42196 49924
rect 42140 49870 42142 49922
rect 42142 49870 42194 49922
rect 42194 49870 42196 49922
rect 42140 49868 42196 49870
rect 40572 48802 40628 48804
rect 40572 48750 40574 48802
rect 40574 48750 40626 48802
rect 40626 48750 40628 48802
rect 40572 48748 40628 48750
rect 40460 48076 40516 48132
rect 41244 49532 41300 49588
rect 41356 49084 41412 49140
rect 43036 50428 43092 50484
rect 42924 49868 42980 49924
rect 41916 48748 41972 48804
rect 42028 49084 42084 49140
rect 41468 48242 41524 48244
rect 41468 48190 41470 48242
rect 41470 48190 41522 48242
rect 41522 48190 41524 48242
rect 41468 48188 41524 48190
rect 41244 48076 41300 48132
rect 41020 47570 41076 47572
rect 41020 47518 41022 47570
rect 41022 47518 41074 47570
rect 41074 47518 41076 47570
rect 41020 47516 41076 47518
rect 41020 46956 41076 47012
rect 40348 45890 40404 45892
rect 40348 45838 40350 45890
rect 40350 45838 40402 45890
rect 40402 45838 40404 45890
rect 40348 45836 40404 45838
rect 40236 45276 40292 45332
rect 40908 45330 40964 45332
rect 40908 45278 40910 45330
rect 40910 45278 40962 45330
rect 40962 45278 40964 45330
rect 40908 45276 40964 45278
rect 40348 45106 40404 45108
rect 40348 45054 40350 45106
rect 40350 45054 40402 45106
rect 40402 45054 40404 45106
rect 40348 45052 40404 45054
rect 41692 48354 41748 48356
rect 41692 48302 41694 48354
rect 41694 48302 41746 48354
rect 41746 48302 41748 48354
rect 41692 48300 41748 48302
rect 41468 47292 41524 47348
rect 41356 47234 41412 47236
rect 41356 47182 41358 47234
rect 41358 47182 41410 47234
rect 41410 47182 41412 47234
rect 41356 47180 41412 47182
rect 41244 47068 41300 47124
rect 41692 47404 41748 47460
rect 42476 48636 42532 48692
rect 45052 53788 45108 53844
rect 44940 53730 44996 53732
rect 44940 53678 44942 53730
rect 44942 53678 44994 53730
rect 44994 53678 44996 53730
rect 44940 53676 44996 53678
rect 44156 52220 44212 52276
rect 44380 53004 44436 53060
rect 44044 51436 44100 51492
rect 44268 51884 44324 51940
rect 43932 51266 43988 51268
rect 43932 51214 43934 51266
rect 43934 51214 43986 51266
rect 43986 51214 43988 51266
rect 43932 51212 43988 51214
rect 43708 50204 43764 50260
rect 42364 48354 42420 48356
rect 42364 48302 42366 48354
rect 42366 48302 42418 48354
rect 42418 48302 42420 48354
rect 42364 48300 42420 48302
rect 44604 51996 44660 52052
rect 44604 50428 44660 50484
rect 44828 53228 44884 53284
rect 44828 52108 44884 52164
rect 45276 55410 45332 55412
rect 45276 55358 45278 55410
rect 45278 55358 45330 55410
rect 45330 55358 45332 55410
rect 45276 55356 45332 55358
rect 45500 54796 45556 54852
rect 45276 53842 45332 53844
rect 45276 53790 45278 53842
rect 45278 53790 45330 53842
rect 45330 53790 45332 53842
rect 45276 53788 45332 53790
rect 45724 54738 45780 54740
rect 45724 54686 45726 54738
rect 45726 54686 45778 54738
rect 45778 54686 45780 54738
rect 45724 54684 45780 54686
rect 45164 52220 45220 52276
rect 45612 52162 45668 52164
rect 45612 52110 45614 52162
rect 45614 52110 45666 52162
rect 45666 52110 45668 52162
rect 45612 52108 45668 52110
rect 45052 50428 45108 50484
rect 45276 51266 45332 51268
rect 45276 51214 45278 51266
rect 45278 51214 45330 51266
rect 45330 51214 45332 51266
rect 45276 51212 45332 51214
rect 44716 50092 44772 50148
rect 44492 49756 44548 49812
rect 45052 49698 45108 49700
rect 45052 49646 45054 49698
rect 45054 49646 45106 49698
rect 45106 49646 45108 49698
rect 45052 49644 45108 49646
rect 44380 49532 44436 49588
rect 45388 49250 45444 49252
rect 45388 49198 45390 49250
rect 45390 49198 45442 49250
rect 45442 49198 45444 49250
rect 45388 49196 45444 49198
rect 44268 48636 44324 48692
rect 44940 48636 44996 48692
rect 43372 48466 43428 48468
rect 43372 48414 43374 48466
rect 43374 48414 43426 48466
rect 43426 48414 43428 48466
rect 43372 48412 43428 48414
rect 44044 48466 44100 48468
rect 44044 48414 44046 48466
rect 44046 48414 44098 48466
rect 44098 48414 44100 48466
rect 44044 48412 44100 48414
rect 42028 46956 42084 47012
rect 41580 45106 41636 45108
rect 41580 45054 41582 45106
rect 41582 45054 41634 45106
rect 41634 45054 41636 45106
rect 41580 45052 41636 45054
rect 42364 47180 42420 47236
rect 42476 47068 42532 47124
rect 42028 44828 42084 44884
rect 40236 44380 40292 44436
rect 41916 44380 41972 44436
rect 40236 43820 40292 43876
rect 41132 44322 41188 44324
rect 41132 44270 41134 44322
rect 41134 44270 41186 44322
rect 41186 44270 41188 44322
rect 41132 44268 41188 44270
rect 41580 44322 41636 44324
rect 41580 44270 41582 44322
rect 41582 44270 41634 44322
rect 41634 44270 41636 44322
rect 41580 44268 41636 44270
rect 41020 43708 41076 43764
rect 40124 43260 40180 43316
rect 40236 42924 40292 42980
rect 40124 41746 40180 41748
rect 40124 41694 40126 41746
rect 40126 41694 40178 41746
rect 40178 41694 40180 41746
rect 40124 41692 40180 41694
rect 39564 41132 39620 41188
rect 40348 40908 40404 40964
rect 38892 38668 38948 38724
rect 37548 37548 37604 37604
rect 37436 37436 37492 37492
rect 38220 37826 38276 37828
rect 38220 37774 38222 37826
rect 38222 37774 38274 37826
rect 38274 37774 38276 37826
rect 38220 37772 38276 37774
rect 38220 37490 38276 37492
rect 38220 37438 38222 37490
rect 38222 37438 38274 37490
rect 38274 37438 38276 37490
rect 38220 37436 38276 37438
rect 38556 37490 38612 37492
rect 38556 37438 38558 37490
rect 38558 37438 38610 37490
rect 38610 37438 38612 37490
rect 38556 37436 38612 37438
rect 38780 38108 38836 38164
rect 39228 37490 39284 37492
rect 39228 37438 39230 37490
rect 39230 37438 39282 37490
rect 39282 37438 39284 37490
rect 39228 37436 39284 37438
rect 37772 36204 37828 36260
rect 38556 35196 38612 35252
rect 38556 34860 38612 34916
rect 37436 34636 37492 34692
rect 37884 34690 37940 34692
rect 37884 34638 37886 34690
rect 37886 34638 37938 34690
rect 37938 34638 37940 34690
rect 37884 34636 37940 34638
rect 37324 34242 37380 34244
rect 37324 34190 37326 34242
rect 37326 34190 37378 34242
rect 37378 34190 37380 34242
rect 37324 34188 37380 34190
rect 36988 33628 37044 33684
rect 36092 31778 36148 31780
rect 36092 31726 36094 31778
rect 36094 31726 36146 31778
rect 36146 31726 36148 31778
rect 36092 31724 36148 31726
rect 35420 30716 35476 30772
rect 35196 30602 35252 30604
rect 35196 30550 35198 30602
rect 35198 30550 35250 30602
rect 35250 30550 35252 30602
rect 35196 30548 35252 30550
rect 35300 30602 35356 30604
rect 35300 30550 35302 30602
rect 35302 30550 35354 30602
rect 35354 30550 35356 30602
rect 35300 30548 35356 30550
rect 35404 30602 35460 30604
rect 35404 30550 35406 30602
rect 35406 30550 35458 30602
rect 35458 30550 35460 30602
rect 35404 30548 35460 30550
rect 35084 30044 35140 30100
rect 34524 29484 34580 29540
rect 34748 29372 34804 29428
rect 36092 30716 36148 30772
rect 35980 30380 36036 30436
rect 35756 30322 35812 30324
rect 35756 30270 35758 30322
rect 35758 30270 35810 30322
rect 35810 30270 35812 30322
rect 35756 30268 35812 30270
rect 35532 30044 35588 30100
rect 34972 28252 35028 28308
rect 34412 27916 34468 27972
rect 35196 29034 35252 29036
rect 35196 28982 35198 29034
rect 35198 28982 35250 29034
rect 35250 28982 35252 29034
rect 35196 28980 35252 28982
rect 35300 29034 35356 29036
rect 35300 28982 35302 29034
rect 35302 28982 35354 29034
rect 35354 28982 35356 29034
rect 35300 28980 35356 28982
rect 35404 29034 35460 29036
rect 35404 28982 35406 29034
rect 35406 28982 35458 29034
rect 35458 28982 35460 29034
rect 35404 28980 35460 28982
rect 35420 28754 35476 28756
rect 35420 28702 35422 28754
rect 35422 28702 35474 28754
rect 35474 28702 35476 28754
rect 35420 28700 35476 28702
rect 35644 28866 35700 28868
rect 35644 28814 35646 28866
rect 35646 28814 35698 28866
rect 35698 28814 35700 28866
rect 35644 28812 35700 28814
rect 35532 28028 35588 28084
rect 35644 28140 35700 28196
rect 34412 27746 34468 27748
rect 34412 27694 34414 27746
rect 34414 27694 34466 27746
rect 34466 27694 34468 27746
rect 34412 27692 34468 27694
rect 34748 27634 34804 27636
rect 34748 27582 34750 27634
rect 34750 27582 34802 27634
rect 34802 27582 34804 27634
rect 34748 27580 34804 27582
rect 34636 27244 34692 27300
rect 33180 26236 33236 26292
rect 33180 25564 33236 25620
rect 35084 27634 35140 27636
rect 35084 27582 35086 27634
rect 35086 27582 35138 27634
rect 35138 27582 35140 27634
rect 35084 27580 35140 27582
rect 35868 27580 35924 27636
rect 35196 27466 35252 27468
rect 35196 27414 35198 27466
rect 35198 27414 35250 27466
rect 35250 27414 35252 27466
rect 35196 27412 35252 27414
rect 35300 27466 35356 27468
rect 35300 27414 35302 27466
rect 35302 27414 35354 27466
rect 35354 27414 35356 27466
rect 35300 27412 35356 27414
rect 35404 27466 35460 27468
rect 35404 27414 35406 27466
rect 35406 27414 35458 27466
rect 35458 27414 35460 27466
rect 35404 27412 35460 27414
rect 35196 27244 35252 27300
rect 35196 27020 35252 27076
rect 35532 26796 35588 26852
rect 33068 23884 33124 23940
rect 33628 25676 33684 25732
rect 34076 25618 34132 25620
rect 34076 25566 34078 25618
rect 34078 25566 34130 25618
rect 34130 25566 34132 25618
rect 34076 25564 34132 25566
rect 34524 25340 34580 25396
rect 33516 23660 33572 23716
rect 34188 22316 34244 22372
rect 33964 21532 34020 21588
rect 33852 20524 33908 20580
rect 33628 20300 33684 20356
rect 33292 19292 33348 19348
rect 33292 18450 33348 18452
rect 33292 18398 33294 18450
rect 33294 18398 33346 18450
rect 33346 18398 33348 18450
rect 33292 18396 33348 18398
rect 33740 20130 33796 20132
rect 33740 20078 33742 20130
rect 33742 20078 33794 20130
rect 33794 20078 33796 20130
rect 33740 20076 33796 20078
rect 34188 20300 34244 20356
rect 34748 26012 34804 26068
rect 34636 23938 34692 23940
rect 34636 23886 34638 23938
rect 34638 23886 34690 23938
rect 34690 23886 34692 23938
rect 34636 23884 34692 23886
rect 36092 26908 36148 26964
rect 36988 31612 37044 31668
rect 36540 30882 36596 30884
rect 36540 30830 36542 30882
rect 36542 30830 36594 30882
rect 36594 30830 36596 30882
rect 36540 30828 36596 30830
rect 36428 29986 36484 29988
rect 36428 29934 36430 29986
rect 36430 29934 36482 29986
rect 36482 29934 36484 29986
rect 36428 29932 36484 29934
rect 35756 26850 35812 26852
rect 35756 26798 35758 26850
rect 35758 26798 35810 26850
rect 35810 26798 35812 26850
rect 35756 26796 35812 26798
rect 35196 25898 35252 25900
rect 35196 25846 35198 25898
rect 35198 25846 35250 25898
rect 35250 25846 35252 25898
rect 35196 25844 35252 25846
rect 35300 25898 35356 25900
rect 35300 25846 35302 25898
rect 35302 25846 35354 25898
rect 35354 25846 35356 25898
rect 35300 25844 35356 25846
rect 35404 25898 35460 25900
rect 35404 25846 35406 25898
rect 35406 25846 35458 25898
rect 35458 25846 35460 25898
rect 35404 25844 35460 25846
rect 35532 25506 35588 25508
rect 35532 25454 35534 25506
rect 35534 25454 35586 25506
rect 35586 25454 35588 25506
rect 35532 25452 35588 25454
rect 35980 25564 36036 25620
rect 34860 25004 34916 25060
rect 35868 25116 35924 25172
rect 35196 24330 35252 24332
rect 35196 24278 35198 24330
rect 35198 24278 35250 24330
rect 35250 24278 35252 24330
rect 35196 24276 35252 24278
rect 35300 24330 35356 24332
rect 35300 24278 35302 24330
rect 35302 24278 35354 24330
rect 35354 24278 35356 24330
rect 35300 24276 35356 24278
rect 35404 24330 35460 24332
rect 35404 24278 35406 24330
rect 35406 24278 35458 24330
rect 35458 24278 35460 24330
rect 35404 24276 35460 24278
rect 36428 25394 36484 25396
rect 36428 25342 36430 25394
rect 36430 25342 36482 25394
rect 36482 25342 36484 25394
rect 36428 25340 36484 25342
rect 36316 24610 36372 24612
rect 36316 24558 36318 24610
rect 36318 24558 36370 24610
rect 36370 24558 36372 24610
rect 36316 24556 36372 24558
rect 34972 23548 35028 23604
rect 35196 23772 35252 23828
rect 34860 22652 34916 22708
rect 35532 23548 35588 23604
rect 35196 22762 35252 22764
rect 35196 22710 35198 22762
rect 35198 22710 35250 22762
rect 35250 22710 35252 22762
rect 35196 22708 35252 22710
rect 35300 22762 35356 22764
rect 35300 22710 35302 22762
rect 35302 22710 35354 22762
rect 35354 22710 35356 22762
rect 35300 22708 35356 22710
rect 35404 22762 35460 22764
rect 35404 22710 35406 22762
rect 35406 22710 35458 22762
rect 35458 22710 35460 22762
rect 35404 22708 35460 22710
rect 34748 22204 34804 22260
rect 34636 21756 34692 21812
rect 35084 22370 35140 22372
rect 35084 22318 35086 22370
rect 35086 22318 35138 22370
rect 35138 22318 35140 22370
rect 35084 22316 35140 22318
rect 36092 23938 36148 23940
rect 36092 23886 36094 23938
rect 36094 23886 36146 23938
rect 36146 23886 36148 23938
rect 36092 23884 36148 23886
rect 35868 22652 35924 22708
rect 36316 23436 36372 23492
rect 35756 22316 35812 22372
rect 34860 21532 34916 21588
rect 35196 21194 35252 21196
rect 35196 21142 35198 21194
rect 35198 21142 35250 21194
rect 35250 21142 35252 21194
rect 35196 21140 35252 21142
rect 35300 21194 35356 21196
rect 35300 21142 35302 21194
rect 35302 21142 35354 21194
rect 35354 21142 35356 21194
rect 35300 21140 35356 21142
rect 35404 21194 35460 21196
rect 35404 21142 35406 21194
rect 35406 21142 35458 21194
rect 35458 21142 35460 21194
rect 35404 21140 35460 21142
rect 36428 22428 36484 22484
rect 36316 22316 36372 22372
rect 35868 22146 35924 22148
rect 35868 22094 35870 22146
rect 35870 22094 35922 22146
rect 35922 22094 35924 22146
rect 35868 22092 35924 22094
rect 35756 21026 35812 21028
rect 35756 20974 35758 21026
rect 35758 20974 35810 21026
rect 35810 20974 35812 21026
rect 35756 20972 35812 20974
rect 34860 20690 34916 20692
rect 34860 20638 34862 20690
rect 34862 20638 34914 20690
rect 34914 20638 34916 20690
rect 34860 20636 34916 20638
rect 34972 20188 35028 20244
rect 31724 17948 31780 18004
rect 30940 15372 30996 15428
rect 30044 14028 30100 14084
rect 30492 14642 30548 14644
rect 30492 14590 30494 14642
rect 30494 14590 30546 14642
rect 30546 14590 30548 14642
rect 30492 14588 30548 14590
rect 30268 13244 30324 13300
rect 29820 12572 29876 12628
rect 29932 12796 29988 12852
rect 28140 10668 28196 10724
rect 28028 10556 28084 10612
rect 29596 11170 29652 11172
rect 29596 11118 29598 11170
rect 29598 11118 29650 11170
rect 29650 11118 29652 11170
rect 29596 11116 29652 11118
rect 29148 10610 29204 10612
rect 29148 10558 29150 10610
rect 29150 10558 29202 10610
rect 29202 10558 29204 10610
rect 29148 10556 29204 10558
rect 29260 10498 29316 10500
rect 29260 10446 29262 10498
rect 29262 10446 29314 10498
rect 29314 10446 29316 10498
rect 29260 10444 29316 10446
rect 29820 10780 29876 10836
rect 28588 10108 28644 10164
rect 30156 12572 30212 12628
rect 30044 12460 30100 12516
rect 31388 16882 31444 16884
rect 31388 16830 31390 16882
rect 31390 16830 31442 16882
rect 31442 16830 31444 16882
rect 31388 16828 31444 16830
rect 31164 16716 31220 16772
rect 30828 14364 30884 14420
rect 30828 14028 30884 14084
rect 30380 12290 30436 12292
rect 30380 12238 30382 12290
rect 30382 12238 30434 12290
rect 30434 12238 30436 12290
rect 30380 12236 30436 12238
rect 30604 12124 30660 12180
rect 30044 11788 30100 11844
rect 30156 10834 30212 10836
rect 30156 10782 30158 10834
rect 30158 10782 30210 10834
rect 30210 10782 30212 10834
rect 30156 10780 30212 10782
rect 30268 9714 30324 9716
rect 30268 9662 30270 9714
rect 30270 9662 30322 9714
rect 30322 9662 30324 9714
rect 30268 9660 30324 9662
rect 29036 7644 29092 7700
rect 28924 7586 28980 7588
rect 28924 7534 28926 7586
rect 28926 7534 28978 7586
rect 28978 7534 28980 7586
rect 28924 7532 28980 7534
rect 27356 6748 27412 6804
rect 26684 6524 26740 6580
rect 27020 6188 27076 6244
rect 27692 6748 27748 6804
rect 28476 6748 28532 6804
rect 28364 6690 28420 6692
rect 28364 6638 28366 6690
rect 28366 6638 28418 6690
rect 28418 6638 28420 6690
rect 28364 6636 28420 6638
rect 27020 5628 27076 5684
rect 27916 6130 27972 6132
rect 27916 6078 27918 6130
rect 27918 6078 27970 6130
rect 27970 6078 27972 6130
rect 27916 6076 27972 6078
rect 28364 6412 28420 6468
rect 27356 5852 27412 5908
rect 27692 5906 27748 5908
rect 27692 5854 27694 5906
rect 27694 5854 27746 5906
rect 27746 5854 27748 5906
rect 27692 5852 27748 5854
rect 27804 5794 27860 5796
rect 27804 5742 27806 5794
rect 27806 5742 27858 5794
rect 27858 5742 27860 5794
rect 27804 5740 27860 5742
rect 29260 6690 29316 6692
rect 29260 6638 29262 6690
rect 29262 6638 29314 6690
rect 29314 6638 29316 6690
rect 29260 6636 29316 6638
rect 30716 11170 30772 11172
rect 30716 11118 30718 11170
rect 30718 11118 30770 11170
rect 30770 11118 30772 11170
rect 30716 11116 30772 11118
rect 30716 10668 30772 10724
rect 30940 11900 30996 11956
rect 32284 17836 32340 17892
rect 31948 16268 32004 16324
rect 32284 17388 32340 17444
rect 32284 16716 32340 16772
rect 33516 18284 33572 18340
rect 33404 18172 33460 18228
rect 33180 17890 33236 17892
rect 33180 17838 33182 17890
rect 33182 17838 33234 17890
rect 33234 17838 33236 17890
rect 33180 17836 33236 17838
rect 32956 17778 33012 17780
rect 32956 17726 32958 17778
rect 32958 17726 33010 17778
rect 33010 17726 33012 17778
rect 32956 17724 33012 17726
rect 33516 17164 33572 17220
rect 32508 16604 32564 16660
rect 32172 15932 32228 15988
rect 32396 15484 32452 15540
rect 31164 12124 31220 12180
rect 31052 11676 31108 11732
rect 31948 14588 32004 14644
rect 31948 14364 32004 14420
rect 31836 13916 31892 13972
rect 31724 12460 31780 12516
rect 31612 12290 31668 12292
rect 31612 12238 31614 12290
rect 31614 12238 31666 12290
rect 31666 12238 31668 12290
rect 31612 12236 31668 12238
rect 32172 12460 32228 12516
rect 32172 12290 32228 12292
rect 32172 12238 32174 12290
rect 32174 12238 32226 12290
rect 32226 12238 32228 12290
rect 32172 12236 32228 12238
rect 31164 11788 31220 11844
rect 30828 10610 30884 10612
rect 30828 10558 30830 10610
rect 30830 10558 30882 10610
rect 30882 10558 30884 10610
rect 30828 10556 30884 10558
rect 31276 10610 31332 10612
rect 31276 10558 31278 10610
rect 31278 10558 31330 10610
rect 31330 10558 31332 10610
rect 31276 10556 31332 10558
rect 31164 9996 31220 10052
rect 31052 9660 31108 9716
rect 31500 9100 31556 9156
rect 31948 11676 32004 11732
rect 32732 14588 32788 14644
rect 32396 11452 32452 11508
rect 31948 10610 32004 10612
rect 31948 10558 31950 10610
rect 31950 10558 32002 10610
rect 32002 10558 32004 10610
rect 31948 10556 32004 10558
rect 32508 10220 32564 10276
rect 31612 8316 31668 8372
rect 31948 9996 32004 10052
rect 30268 7644 30324 7700
rect 30044 7474 30100 7476
rect 30044 7422 30046 7474
rect 30046 7422 30098 7474
rect 30098 7422 30100 7474
rect 30044 7420 30100 7422
rect 30380 6748 30436 6804
rect 30044 6690 30100 6692
rect 30044 6638 30046 6690
rect 30046 6638 30098 6690
rect 30098 6638 30100 6690
rect 30044 6636 30100 6638
rect 28588 6524 28644 6580
rect 29260 6188 29316 6244
rect 29596 6018 29652 6020
rect 29596 5966 29598 6018
rect 29598 5966 29650 6018
rect 29650 5966 29652 6018
rect 29596 5964 29652 5966
rect 29036 5906 29092 5908
rect 29036 5854 29038 5906
rect 29038 5854 29090 5906
rect 29090 5854 29092 5906
rect 29036 5852 29092 5854
rect 30268 6578 30324 6580
rect 30268 6526 30270 6578
rect 30270 6526 30322 6578
rect 30322 6526 30324 6578
rect 30268 6524 30324 6526
rect 29708 5852 29764 5908
rect 29820 6076 29876 6132
rect 30492 6466 30548 6468
rect 30492 6414 30494 6466
rect 30494 6414 30546 6466
rect 30546 6414 30548 6466
rect 30492 6412 30548 6414
rect 30268 5852 30324 5908
rect 30828 7250 30884 7252
rect 30828 7198 30830 7250
rect 30830 7198 30882 7250
rect 30882 7198 30884 7250
rect 30828 7196 30884 7198
rect 31612 7644 31668 7700
rect 31500 7474 31556 7476
rect 31500 7422 31502 7474
rect 31502 7422 31554 7474
rect 31554 7422 31556 7474
rect 31500 7420 31556 7422
rect 32396 9996 32452 10052
rect 33628 16604 33684 16660
rect 33740 19628 33796 19684
rect 33292 15932 33348 15988
rect 33516 16098 33572 16100
rect 33516 16046 33518 16098
rect 33518 16046 33570 16098
rect 33570 16046 33572 16098
rect 33516 16044 33572 16046
rect 33292 15538 33348 15540
rect 33292 15486 33294 15538
rect 33294 15486 33346 15538
rect 33346 15486 33348 15538
rect 33292 15484 33348 15486
rect 34412 19906 34468 19908
rect 34412 19854 34414 19906
rect 34414 19854 34466 19906
rect 34466 19854 34468 19906
rect 34412 19852 34468 19854
rect 35084 20130 35140 20132
rect 35084 20078 35086 20130
rect 35086 20078 35138 20130
rect 35138 20078 35140 20130
rect 35084 20076 35140 20078
rect 36204 20690 36260 20692
rect 36204 20638 36206 20690
rect 36206 20638 36258 20690
rect 36258 20638 36260 20690
rect 36204 20636 36260 20638
rect 35980 20524 36036 20580
rect 35532 20300 35588 20356
rect 35868 20300 35924 20356
rect 35756 20188 35812 20244
rect 35644 20130 35700 20132
rect 35644 20078 35646 20130
rect 35646 20078 35698 20130
rect 35698 20078 35700 20130
rect 35644 20076 35700 20078
rect 34748 19628 34804 19684
rect 35196 19626 35252 19628
rect 35196 19574 35198 19626
rect 35198 19574 35250 19626
rect 35250 19574 35252 19626
rect 35196 19572 35252 19574
rect 35300 19626 35356 19628
rect 35300 19574 35302 19626
rect 35302 19574 35354 19626
rect 35354 19574 35356 19626
rect 35300 19572 35356 19574
rect 35404 19626 35460 19628
rect 35404 19574 35406 19626
rect 35406 19574 35458 19626
rect 35458 19574 35460 19626
rect 35404 19572 35460 19574
rect 34524 19346 34580 19348
rect 34524 19294 34526 19346
rect 34526 19294 34578 19346
rect 34578 19294 34580 19346
rect 34524 19292 34580 19294
rect 34412 18844 34468 18900
rect 34636 19068 34692 19124
rect 34636 18338 34692 18340
rect 34636 18286 34638 18338
rect 34638 18286 34690 18338
rect 34690 18286 34692 18338
rect 34636 18284 34692 18286
rect 34300 18172 34356 18228
rect 35084 19068 35140 19124
rect 35420 19122 35476 19124
rect 35420 19070 35422 19122
rect 35422 19070 35474 19122
rect 35474 19070 35476 19122
rect 35420 19068 35476 19070
rect 35196 18844 35252 18900
rect 35196 18620 35252 18676
rect 35084 18450 35140 18452
rect 35084 18398 35086 18450
rect 35086 18398 35138 18450
rect 35138 18398 35140 18450
rect 35084 18396 35140 18398
rect 35308 18396 35364 18452
rect 35532 18450 35588 18452
rect 35532 18398 35534 18450
rect 35534 18398 35586 18450
rect 35586 18398 35588 18450
rect 35532 18396 35588 18398
rect 33964 17836 34020 17892
rect 34188 17724 34244 17780
rect 34300 17554 34356 17556
rect 34300 17502 34302 17554
rect 34302 17502 34354 17554
rect 34354 17502 34356 17554
rect 34300 17500 34356 17502
rect 35196 18058 35252 18060
rect 35196 18006 35198 18058
rect 35198 18006 35250 18058
rect 35250 18006 35252 18058
rect 35196 18004 35252 18006
rect 35300 18058 35356 18060
rect 35300 18006 35302 18058
rect 35302 18006 35354 18058
rect 35354 18006 35356 18058
rect 35300 18004 35356 18006
rect 35404 18058 35460 18060
rect 35404 18006 35406 18058
rect 35406 18006 35458 18058
rect 35458 18006 35460 18058
rect 35404 18004 35460 18006
rect 35756 19852 35812 19908
rect 35980 19852 36036 19908
rect 35868 18674 35924 18676
rect 35868 18622 35870 18674
rect 35870 18622 35922 18674
rect 35922 18622 35924 18674
rect 35868 18620 35924 18622
rect 35868 18396 35924 18452
rect 36092 20076 36148 20132
rect 36092 19404 36148 19460
rect 36316 20076 36372 20132
rect 36316 19740 36372 19796
rect 36092 18620 36148 18676
rect 36204 18844 36260 18900
rect 34636 17724 34692 17780
rect 34972 17724 35028 17780
rect 34860 17666 34916 17668
rect 34860 17614 34862 17666
rect 34862 17614 34914 17666
rect 34914 17614 34916 17666
rect 34860 17612 34916 17614
rect 34524 17554 34580 17556
rect 34524 17502 34526 17554
rect 34526 17502 34578 17554
rect 34578 17502 34580 17554
rect 34524 17500 34580 17502
rect 34188 17164 34244 17220
rect 34412 17106 34468 17108
rect 34412 17054 34414 17106
rect 34414 17054 34466 17106
rect 34466 17054 34468 17106
rect 34412 17052 34468 17054
rect 34300 15986 34356 15988
rect 34300 15934 34302 15986
rect 34302 15934 34354 15986
rect 34354 15934 34356 15986
rect 34300 15932 34356 15934
rect 33964 15820 34020 15876
rect 33852 15538 33908 15540
rect 33852 15486 33854 15538
rect 33854 15486 33906 15538
rect 33906 15486 33908 15538
rect 33852 15484 33908 15486
rect 33964 15260 34020 15316
rect 34188 15260 34244 15316
rect 33404 14588 33460 14644
rect 33740 13858 33796 13860
rect 33740 13806 33742 13858
rect 33742 13806 33794 13858
rect 33794 13806 33796 13858
rect 33740 13804 33796 13806
rect 33628 13692 33684 13748
rect 33740 13580 33796 13636
rect 33628 12124 33684 12180
rect 33068 11394 33124 11396
rect 33068 11342 33070 11394
rect 33070 11342 33122 11394
rect 33122 11342 33124 11394
rect 33068 11340 33124 11342
rect 34188 14924 34244 14980
rect 34076 14700 34132 14756
rect 34076 13580 34132 13636
rect 34188 13468 34244 13524
rect 34636 16044 34692 16100
rect 34860 16828 34916 16884
rect 36316 17948 36372 18004
rect 36092 17666 36148 17668
rect 36092 17614 36094 17666
rect 36094 17614 36146 17666
rect 36146 17614 36148 17666
rect 36092 17612 36148 17614
rect 36428 17836 36484 17892
rect 35420 17106 35476 17108
rect 35420 17054 35422 17106
rect 35422 17054 35474 17106
rect 35474 17054 35476 17106
rect 35420 17052 35476 17054
rect 35196 16490 35252 16492
rect 35196 16438 35198 16490
rect 35198 16438 35250 16490
rect 35250 16438 35252 16490
rect 35196 16436 35252 16438
rect 35300 16490 35356 16492
rect 35300 16438 35302 16490
rect 35302 16438 35354 16490
rect 35354 16438 35356 16490
rect 35300 16436 35356 16438
rect 35404 16490 35460 16492
rect 35404 16438 35406 16490
rect 35406 16438 35458 16490
rect 35458 16438 35460 16490
rect 35404 16436 35460 16438
rect 35420 16156 35476 16212
rect 36316 17106 36372 17108
rect 36316 17054 36318 17106
rect 36318 17054 36370 17106
rect 36370 17054 36372 17106
rect 36316 17052 36372 17054
rect 35980 16828 36036 16884
rect 35868 16268 35924 16324
rect 36428 16994 36484 16996
rect 36428 16942 36430 16994
rect 36430 16942 36482 16994
rect 36482 16942 36484 16994
rect 36428 16940 36484 16942
rect 36428 16604 36484 16660
rect 37436 33516 37492 33572
rect 37548 33180 37604 33236
rect 37548 31612 37604 31668
rect 37436 31388 37492 31444
rect 37212 31218 37268 31220
rect 37212 31166 37214 31218
rect 37214 31166 37266 31218
rect 37266 31166 37268 31218
rect 37212 31164 37268 31166
rect 37100 30268 37156 30324
rect 37548 30380 37604 30436
rect 38108 31218 38164 31220
rect 38108 31166 38110 31218
rect 38110 31166 38162 31218
rect 38162 31166 38164 31218
rect 38108 31164 38164 31166
rect 38332 31052 38388 31108
rect 38220 30994 38276 30996
rect 38220 30942 38222 30994
rect 38222 30942 38274 30994
rect 38274 30942 38276 30994
rect 38220 30940 38276 30942
rect 38108 30380 38164 30436
rect 37996 27692 38052 27748
rect 36988 27074 37044 27076
rect 36988 27022 36990 27074
rect 36990 27022 37042 27074
rect 37042 27022 37044 27074
rect 36988 27020 37044 27022
rect 36876 26908 36932 26964
rect 37996 26908 38052 26964
rect 36988 26796 37044 26852
rect 36764 25676 36820 25732
rect 37212 26850 37268 26852
rect 37212 26798 37214 26850
rect 37214 26798 37266 26850
rect 37266 26798 37268 26850
rect 37212 26796 37268 26798
rect 36988 25506 37044 25508
rect 36988 25454 36990 25506
rect 36990 25454 37042 25506
rect 37042 25454 37044 25506
rect 36988 25452 37044 25454
rect 37436 26460 37492 26516
rect 38220 26572 38276 26628
rect 37996 26514 38052 26516
rect 37996 26462 37998 26514
rect 37998 26462 38050 26514
rect 38050 26462 38052 26514
rect 37996 26460 38052 26462
rect 37212 25228 37268 25284
rect 38780 34802 38836 34804
rect 38780 34750 38782 34802
rect 38782 34750 38834 34802
rect 38834 34750 38836 34802
rect 38780 34748 38836 34750
rect 39116 33516 39172 33572
rect 39116 33234 39172 33236
rect 39116 33182 39118 33234
rect 39118 33182 39170 33234
rect 39170 33182 39172 33234
rect 39116 33180 39172 33182
rect 39900 38220 39956 38276
rect 41468 43762 41524 43764
rect 41468 43710 41470 43762
rect 41470 43710 41522 43762
rect 41522 43710 41524 43762
rect 41468 43708 41524 43710
rect 42588 47292 42644 47348
rect 42476 45836 42532 45892
rect 42364 44940 42420 44996
rect 42364 44380 42420 44436
rect 42028 43484 42084 43540
rect 40684 43260 40740 43316
rect 40908 40402 40964 40404
rect 40908 40350 40910 40402
rect 40910 40350 40962 40402
rect 40962 40350 40964 40402
rect 40908 40348 40964 40350
rect 41132 40348 41188 40404
rect 41356 42028 41412 42084
rect 41468 41692 41524 41748
rect 41916 40514 41972 40516
rect 41916 40462 41918 40514
rect 41918 40462 41970 40514
rect 41970 40462 41972 40514
rect 41916 40460 41972 40462
rect 40460 38668 40516 38724
rect 40124 38108 40180 38164
rect 39676 37772 39732 37828
rect 40236 37772 40292 37828
rect 39788 37324 39844 37380
rect 42252 40348 42308 40404
rect 42700 47180 42756 47236
rect 43484 47068 43540 47124
rect 43596 47180 43652 47236
rect 44828 47292 44884 47348
rect 43708 46620 43764 46676
rect 42812 45948 42868 46004
rect 43260 45890 43316 45892
rect 43260 45838 43262 45890
rect 43262 45838 43314 45890
rect 43314 45838 43316 45890
rect 43260 45836 43316 45838
rect 43596 45890 43652 45892
rect 43596 45838 43598 45890
rect 43598 45838 43650 45890
rect 43650 45838 43652 45890
rect 43596 45836 43652 45838
rect 43372 45164 43428 45220
rect 42812 45106 42868 45108
rect 42812 45054 42814 45106
rect 42814 45054 42866 45106
rect 42866 45054 42868 45106
rect 42812 45052 42868 45054
rect 42700 44882 42756 44884
rect 42700 44830 42702 44882
rect 42702 44830 42754 44882
rect 42754 44830 42756 44882
rect 42700 44828 42756 44830
rect 42924 44546 42980 44548
rect 42924 44494 42926 44546
rect 42926 44494 42978 44546
rect 42978 44494 42980 44546
rect 42924 44492 42980 44494
rect 43596 44994 43652 44996
rect 43596 44942 43598 44994
rect 43598 44942 43650 44994
rect 43650 44942 43652 44994
rect 43596 44940 43652 44942
rect 44268 46674 44324 46676
rect 44268 46622 44270 46674
rect 44270 46622 44322 46674
rect 44322 46622 44324 46674
rect 44268 46620 44324 46622
rect 43932 44492 43988 44548
rect 44044 45948 44100 46004
rect 43372 43820 43428 43876
rect 44828 46002 44884 46004
rect 44828 45950 44830 46002
rect 44830 45950 44882 46002
rect 44882 45950 44884 46002
rect 44828 45948 44884 45950
rect 45052 47458 45108 47460
rect 45052 47406 45054 47458
rect 45054 47406 45106 47458
rect 45106 47406 45108 47458
rect 45052 47404 45108 47406
rect 45388 47234 45444 47236
rect 45388 47182 45390 47234
rect 45390 47182 45442 47234
rect 45442 47182 45444 47234
rect 45388 47180 45444 47182
rect 44156 45666 44212 45668
rect 44156 45614 44158 45666
rect 44158 45614 44210 45666
rect 44210 45614 44212 45666
rect 44156 45612 44212 45614
rect 45052 45500 45108 45556
rect 44044 44268 44100 44324
rect 43596 43538 43652 43540
rect 43596 43486 43598 43538
rect 43598 43486 43650 43538
rect 43650 43486 43652 43538
rect 43596 43484 43652 43486
rect 43820 44210 43876 44212
rect 43820 44158 43822 44210
rect 43822 44158 43874 44210
rect 43874 44158 43876 44210
rect 43820 44156 43876 44158
rect 43484 41692 43540 41748
rect 42812 41356 42868 41412
rect 44268 44322 44324 44324
rect 44268 44270 44270 44322
rect 44270 44270 44322 44322
rect 44322 44270 44324 44322
rect 44268 44268 44324 44270
rect 44044 44098 44100 44100
rect 44044 44046 44046 44098
rect 44046 44046 44098 44098
rect 44098 44046 44100 44098
rect 44044 44044 44100 44046
rect 44044 43820 44100 43876
rect 44940 45276 44996 45332
rect 44940 44210 44996 44212
rect 44940 44158 44942 44210
rect 44942 44158 44994 44210
rect 44994 44158 44996 44210
rect 44940 44156 44996 44158
rect 45388 45330 45444 45332
rect 45388 45278 45390 45330
rect 45390 45278 45442 45330
rect 45442 45278 45444 45330
rect 45388 45276 45444 45278
rect 45612 45164 45668 45220
rect 45164 45106 45220 45108
rect 45164 45054 45166 45106
rect 45166 45054 45218 45106
rect 45218 45054 45220 45106
rect 45164 45052 45220 45054
rect 45276 44434 45332 44436
rect 45276 44382 45278 44434
rect 45278 44382 45330 44434
rect 45330 44382 45332 44434
rect 45276 44380 45332 44382
rect 45164 44268 45220 44324
rect 45052 43484 45108 43540
rect 43820 40460 43876 40516
rect 42700 40402 42756 40404
rect 42700 40350 42702 40402
rect 42702 40350 42754 40402
rect 42754 40350 42756 40402
rect 42700 40348 42756 40350
rect 42476 39900 42532 39956
rect 41580 37996 41636 38052
rect 40348 37324 40404 37380
rect 40460 36988 40516 37044
rect 40124 36316 40180 36372
rect 38668 30994 38724 30996
rect 38668 30942 38670 30994
rect 38670 30942 38722 30994
rect 38722 30942 38724 30994
rect 38668 30940 38724 30942
rect 38780 30380 38836 30436
rect 39900 33346 39956 33348
rect 39900 33294 39902 33346
rect 39902 33294 39954 33346
rect 39954 33294 39956 33346
rect 39900 33292 39956 33294
rect 40012 33180 40068 33236
rect 40348 33346 40404 33348
rect 40348 33294 40350 33346
rect 40350 33294 40402 33346
rect 40402 33294 40404 33346
rect 40348 33292 40404 33294
rect 39564 31724 39620 31780
rect 39900 31836 39956 31892
rect 39004 31164 39060 31220
rect 40012 32284 40068 32340
rect 39228 31106 39284 31108
rect 39228 31054 39230 31106
rect 39230 31054 39282 31106
rect 39282 31054 39284 31106
rect 39228 31052 39284 31054
rect 39564 30882 39620 30884
rect 39564 30830 39566 30882
rect 39566 30830 39618 30882
rect 39618 30830 39620 30882
rect 39564 30828 39620 30830
rect 39228 29372 39284 29428
rect 39900 28530 39956 28532
rect 39900 28478 39902 28530
rect 39902 28478 39954 28530
rect 39954 28478 39956 28530
rect 39900 28476 39956 28478
rect 39564 27746 39620 27748
rect 39564 27694 39566 27746
rect 39566 27694 39618 27746
rect 39618 27694 39620 27746
rect 39564 27692 39620 27694
rect 38892 26460 38948 26516
rect 39340 26402 39396 26404
rect 39340 26350 39342 26402
rect 39342 26350 39394 26402
rect 39394 26350 39396 26402
rect 39340 26348 39396 26350
rect 39452 25452 39508 25508
rect 39228 24556 39284 24612
rect 39676 24610 39732 24612
rect 39676 24558 39678 24610
rect 39678 24558 39730 24610
rect 39730 24558 39732 24610
rect 39676 24556 39732 24558
rect 37436 23436 37492 23492
rect 37100 22146 37156 22148
rect 37100 22094 37102 22146
rect 37102 22094 37154 22146
rect 37154 22094 37156 22146
rect 37100 22092 37156 22094
rect 37548 21756 37604 21812
rect 36988 20690 37044 20692
rect 36988 20638 36990 20690
rect 36990 20638 37042 20690
rect 37042 20638 37044 20690
rect 36988 20636 37044 20638
rect 36652 20524 36708 20580
rect 36988 20412 37044 20468
rect 37100 20076 37156 20132
rect 37660 20972 37716 21028
rect 37884 21756 37940 21812
rect 37100 19906 37156 19908
rect 37100 19854 37102 19906
rect 37102 19854 37154 19906
rect 37154 19854 37156 19906
rect 37100 19852 37156 19854
rect 37212 19234 37268 19236
rect 37212 19182 37214 19234
rect 37214 19182 37266 19234
rect 37266 19182 37268 19234
rect 37212 19180 37268 19182
rect 36876 18844 36932 18900
rect 37212 18396 37268 18452
rect 36876 17948 36932 18004
rect 36652 17164 36708 17220
rect 36652 16882 36708 16884
rect 36652 16830 36654 16882
rect 36654 16830 36706 16882
rect 36706 16830 36708 16882
rect 36652 16828 36708 16830
rect 36316 16156 36372 16212
rect 35084 15314 35140 15316
rect 35084 15262 35086 15314
rect 35086 15262 35138 15314
rect 35138 15262 35140 15314
rect 35084 15260 35140 15262
rect 34188 13074 34244 13076
rect 34188 13022 34190 13074
rect 34190 13022 34242 13074
rect 34242 13022 34244 13074
rect 34188 13020 34244 13022
rect 33964 12908 34020 12964
rect 33852 12348 33908 12404
rect 34076 12850 34132 12852
rect 34076 12798 34078 12850
rect 34078 12798 34130 12850
rect 34130 12798 34132 12850
rect 34076 12796 34132 12798
rect 35644 15708 35700 15764
rect 35980 15708 36036 15764
rect 35868 15596 35924 15652
rect 35420 15036 35476 15092
rect 35868 15202 35924 15204
rect 35868 15150 35870 15202
rect 35870 15150 35922 15202
rect 35922 15150 35924 15202
rect 35868 15148 35924 15150
rect 35196 14922 35252 14924
rect 35196 14870 35198 14922
rect 35198 14870 35250 14922
rect 35250 14870 35252 14922
rect 35196 14868 35252 14870
rect 35300 14922 35356 14924
rect 35300 14870 35302 14922
rect 35302 14870 35354 14922
rect 35354 14870 35356 14922
rect 35300 14868 35356 14870
rect 35404 14922 35460 14924
rect 35404 14870 35406 14922
rect 35406 14870 35458 14922
rect 35458 14870 35460 14922
rect 35404 14868 35460 14870
rect 34748 14140 34804 14196
rect 35196 13916 35252 13972
rect 34412 13746 34468 13748
rect 34412 13694 34414 13746
rect 34414 13694 34466 13746
rect 34466 13694 34468 13746
rect 34412 13692 34468 13694
rect 34748 13522 34804 13524
rect 34748 13470 34750 13522
rect 34750 13470 34802 13522
rect 34802 13470 34804 13522
rect 34748 13468 34804 13470
rect 34412 12962 34468 12964
rect 34412 12910 34414 12962
rect 34414 12910 34466 12962
rect 34466 12910 34468 12962
rect 34412 12908 34468 12910
rect 34300 12684 34356 12740
rect 35532 13916 35588 13972
rect 35196 13354 35252 13356
rect 35196 13302 35198 13354
rect 35198 13302 35250 13354
rect 35250 13302 35252 13354
rect 35196 13300 35252 13302
rect 35300 13354 35356 13356
rect 35300 13302 35302 13354
rect 35302 13302 35354 13354
rect 35354 13302 35356 13354
rect 35300 13300 35356 13302
rect 35404 13354 35460 13356
rect 35404 13302 35406 13354
rect 35406 13302 35458 13354
rect 35458 13302 35460 13354
rect 35404 13300 35460 13302
rect 35084 13020 35140 13076
rect 35084 12850 35140 12852
rect 35084 12798 35086 12850
rect 35086 12798 35138 12850
rect 35138 12798 35140 12850
rect 35084 12796 35140 12798
rect 35756 13858 35812 13860
rect 35756 13806 35758 13858
rect 35758 13806 35810 13858
rect 35810 13806 35812 13858
rect 35756 13804 35812 13806
rect 35644 12796 35700 12852
rect 34636 12684 34692 12740
rect 33180 9996 33236 10052
rect 32732 8204 32788 8260
rect 33180 7586 33236 7588
rect 33180 7534 33182 7586
rect 33182 7534 33234 7586
rect 33234 7534 33236 7586
rect 33180 7532 33236 7534
rect 32172 7196 32228 7252
rect 31276 6748 31332 6804
rect 32172 6748 32228 6804
rect 33068 6748 33124 6804
rect 33852 9996 33908 10052
rect 34076 12066 34132 12068
rect 34076 12014 34078 12066
rect 34078 12014 34130 12066
rect 34130 12014 34132 12066
rect 34076 12012 34132 12014
rect 34300 11340 34356 11396
rect 34636 12012 34692 12068
rect 34636 11004 34692 11060
rect 34748 11228 34804 11284
rect 33516 9324 33572 9380
rect 33404 9042 33460 9044
rect 33404 8990 33406 9042
rect 33406 8990 33458 9042
rect 33458 8990 33460 9042
rect 33404 8988 33460 8990
rect 33852 9042 33908 9044
rect 33852 8990 33854 9042
rect 33854 8990 33906 9042
rect 33906 8990 33908 9042
rect 33852 8988 33908 8990
rect 33740 7586 33796 7588
rect 33740 7534 33742 7586
rect 33742 7534 33794 7586
rect 33794 7534 33796 7586
rect 33740 7532 33796 7534
rect 34188 9212 34244 9268
rect 34076 9154 34132 9156
rect 34076 9102 34078 9154
rect 34078 9102 34130 9154
rect 34130 9102 34132 9154
rect 34076 9100 34132 9102
rect 34636 10332 34692 10388
rect 34524 9996 34580 10052
rect 35196 11786 35252 11788
rect 35196 11734 35198 11786
rect 35198 11734 35250 11786
rect 35250 11734 35252 11786
rect 35196 11732 35252 11734
rect 35300 11786 35356 11788
rect 35300 11734 35302 11786
rect 35302 11734 35354 11786
rect 35354 11734 35356 11786
rect 35300 11732 35356 11734
rect 35404 11786 35460 11788
rect 35404 11734 35406 11786
rect 35406 11734 35458 11786
rect 35458 11734 35460 11786
rect 35404 11732 35460 11734
rect 35644 11394 35700 11396
rect 35644 11342 35646 11394
rect 35646 11342 35698 11394
rect 35698 11342 35700 11394
rect 35644 11340 35700 11342
rect 34972 11228 35028 11284
rect 35532 11116 35588 11172
rect 35196 10218 35252 10220
rect 35196 10166 35198 10218
rect 35198 10166 35250 10218
rect 35250 10166 35252 10218
rect 35196 10164 35252 10166
rect 35300 10218 35356 10220
rect 35300 10166 35302 10218
rect 35302 10166 35354 10218
rect 35354 10166 35356 10218
rect 35300 10164 35356 10166
rect 35404 10218 35460 10220
rect 35404 10166 35406 10218
rect 35406 10166 35458 10218
rect 35458 10166 35460 10218
rect 35404 10164 35460 10166
rect 35420 9996 35476 10052
rect 35084 9826 35140 9828
rect 35084 9774 35086 9826
rect 35086 9774 35138 9826
rect 35138 9774 35140 9826
rect 35084 9772 35140 9774
rect 35868 11004 35924 11060
rect 35868 10444 35924 10500
rect 35756 10332 35812 10388
rect 36540 16044 36596 16100
rect 36204 15036 36260 15092
rect 36204 14700 36260 14756
rect 36204 13804 36260 13860
rect 36092 11282 36148 11284
rect 36092 11230 36094 11282
rect 36094 11230 36146 11282
rect 36146 11230 36148 11282
rect 36092 11228 36148 11230
rect 36092 10892 36148 10948
rect 36092 10108 36148 10164
rect 36316 10332 36372 10388
rect 34636 8258 34692 8260
rect 34636 8206 34638 8258
rect 34638 8206 34690 8258
rect 34690 8206 34692 8258
rect 34636 8204 34692 8206
rect 34412 7980 34468 8036
rect 34412 7474 34468 7476
rect 34412 7422 34414 7474
rect 34414 7422 34466 7474
rect 34466 7422 34468 7474
rect 34412 7420 34468 7422
rect 34412 6802 34468 6804
rect 34412 6750 34414 6802
rect 34414 6750 34466 6802
rect 34466 6750 34468 6802
rect 34412 6748 34468 6750
rect 34300 6636 34356 6692
rect 31052 6578 31108 6580
rect 31052 6526 31054 6578
rect 31054 6526 31106 6578
rect 31106 6526 31108 6578
rect 31052 6524 31108 6526
rect 31724 6524 31780 6580
rect 31276 6076 31332 6132
rect 31500 6018 31556 6020
rect 31500 5966 31502 6018
rect 31502 5966 31554 6018
rect 31554 5966 31556 6018
rect 31500 5964 31556 5966
rect 26572 4956 26628 5012
rect 28140 5068 28196 5124
rect 27356 4956 27412 5012
rect 29036 5068 29092 5124
rect 29932 5122 29988 5124
rect 29932 5070 29934 5122
rect 29934 5070 29986 5122
rect 29986 5070 29988 5122
rect 29932 5068 29988 5070
rect 31052 5180 31108 5236
rect 32844 6466 32900 6468
rect 32844 6414 32846 6466
rect 32846 6414 32898 6466
rect 32898 6414 32900 6466
rect 32844 6412 32900 6414
rect 32620 6188 32676 6244
rect 33068 6130 33124 6132
rect 33068 6078 33070 6130
rect 33070 6078 33122 6130
rect 33122 6078 33124 6130
rect 33068 6076 33124 6078
rect 32396 5292 32452 5348
rect 34076 6188 34132 6244
rect 33740 6018 33796 6020
rect 33740 5966 33742 6018
rect 33742 5966 33794 6018
rect 33794 5966 33796 6018
rect 33740 5964 33796 5966
rect 32732 5234 32788 5236
rect 32732 5182 32734 5234
rect 32734 5182 32786 5234
rect 32786 5182 32788 5234
rect 32732 5180 32788 5182
rect 33180 5122 33236 5124
rect 33180 5070 33182 5122
rect 33182 5070 33234 5122
rect 33234 5070 33236 5122
rect 33180 5068 33236 5070
rect 33516 5852 33572 5908
rect 34748 7586 34804 7588
rect 34748 7534 34750 7586
rect 34750 7534 34802 7586
rect 34802 7534 34804 7586
rect 34748 7532 34804 7534
rect 35084 9266 35140 9268
rect 35084 9214 35086 9266
rect 35086 9214 35138 9266
rect 35138 9214 35140 9266
rect 35084 9212 35140 9214
rect 35196 8650 35252 8652
rect 35196 8598 35198 8650
rect 35198 8598 35250 8650
rect 35250 8598 35252 8650
rect 35196 8596 35252 8598
rect 35300 8650 35356 8652
rect 35300 8598 35302 8650
rect 35302 8598 35354 8650
rect 35354 8598 35356 8650
rect 35300 8596 35356 8598
rect 35404 8650 35460 8652
rect 35404 8598 35406 8650
rect 35406 8598 35458 8650
rect 35458 8598 35460 8650
rect 35404 8596 35460 8598
rect 35644 8204 35700 8260
rect 35084 7756 35140 7812
rect 35308 7756 35364 7812
rect 35420 7586 35476 7588
rect 35420 7534 35422 7586
rect 35422 7534 35474 7586
rect 35474 7534 35476 7586
rect 35420 7532 35476 7534
rect 34860 7420 34916 7476
rect 35196 7082 35252 7084
rect 35196 7030 35198 7082
rect 35198 7030 35250 7082
rect 35250 7030 35252 7082
rect 35196 7028 35252 7030
rect 35300 7082 35356 7084
rect 35300 7030 35302 7082
rect 35302 7030 35354 7082
rect 35354 7030 35356 7082
rect 35300 7028 35356 7030
rect 35404 7082 35460 7084
rect 35404 7030 35406 7082
rect 35406 7030 35458 7082
rect 35458 7030 35460 7082
rect 35404 7028 35460 7030
rect 34748 6748 34804 6804
rect 34860 6636 34916 6692
rect 35308 6690 35364 6692
rect 35308 6638 35310 6690
rect 35310 6638 35362 6690
rect 35362 6638 35364 6690
rect 35308 6636 35364 6638
rect 34972 6018 35028 6020
rect 34972 5966 34974 6018
rect 34974 5966 35026 6018
rect 35026 5966 35028 6018
rect 34972 5964 35028 5966
rect 35420 5906 35476 5908
rect 35420 5854 35422 5906
rect 35422 5854 35474 5906
rect 35474 5854 35476 5906
rect 35420 5852 35476 5854
rect 35308 5740 35364 5796
rect 35532 5628 35588 5684
rect 35868 9324 35924 9380
rect 35756 7644 35812 7700
rect 36092 7532 36148 7588
rect 36204 7980 36260 8036
rect 35756 7474 35812 7476
rect 35756 7422 35758 7474
rect 35758 7422 35810 7474
rect 35810 7422 35812 7474
rect 35756 7420 35812 7422
rect 35196 5514 35252 5516
rect 35196 5462 35198 5514
rect 35198 5462 35250 5514
rect 35250 5462 35252 5514
rect 35196 5460 35252 5462
rect 35300 5514 35356 5516
rect 35300 5462 35302 5514
rect 35302 5462 35354 5514
rect 35354 5462 35356 5514
rect 35300 5460 35356 5462
rect 35404 5514 35460 5516
rect 35404 5462 35406 5514
rect 35406 5462 35458 5514
rect 35458 5462 35460 5514
rect 35404 5460 35460 5462
rect 35980 6636 36036 6692
rect 35868 6076 35924 6132
rect 36092 6524 36148 6580
rect 35308 5292 35364 5348
rect 33516 4956 33572 5012
rect 36092 5628 36148 5684
rect 35868 5180 35924 5236
rect 37100 17052 37156 17108
rect 37100 16658 37156 16660
rect 37100 16606 37102 16658
rect 37102 16606 37154 16658
rect 37154 16606 37156 16658
rect 37100 16604 37156 16606
rect 36988 16268 37044 16324
rect 37212 16156 37268 16212
rect 36876 15596 36932 15652
rect 37548 19516 37604 19572
rect 37548 18956 37604 19012
rect 37660 17724 37716 17780
rect 37772 20076 37828 20132
rect 37772 19068 37828 19124
rect 38556 23826 38612 23828
rect 38556 23774 38558 23826
rect 38558 23774 38610 23826
rect 38610 23774 38612 23826
rect 38556 23772 38612 23774
rect 39564 23378 39620 23380
rect 39564 23326 39566 23378
rect 39566 23326 39618 23378
rect 39618 23326 39620 23378
rect 39564 23324 39620 23326
rect 38556 23212 38612 23268
rect 38332 21532 38388 21588
rect 40012 22876 40068 22932
rect 40124 32172 40180 32228
rect 38220 21308 38276 21364
rect 38556 21308 38612 21364
rect 38668 21532 38724 21588
rect 38668 21196 38724 21252
rect 40012 21644 40068 21700
rect 39228 21532 39284 21588
rect 38556 20690 38612 20692
rect 38556 20638 38558 20690
rect 38558 20638 38610 20690
rect 38610 20638 38612 20690
rect 38556 20636 38612 20638
rect 39228 21196 39284 21252
rect 39788 21586 39844 21588
rect 39788 21534 39790 21586
rect 39790 21534 39842 21586
rect 39842 21534 39844 21586
rect 39788 21532 39844 21534
rect 41580 37266 41636 37268
rect 41580 37214 41582 37266
rect 41582 37214 41634 37266
rect 41634 37214 41636 37266
rect 41580 37212 41636 37214
rect 42028 38274 42084 38276
rect 42028 38222 42030 38274
rect 42030 38222 42082 38274
rect 42082 38222 42084 38274
rect 42028 38220 42084 38222
rect 42364 38220 42420 38276
rect 41916 37490 41972 37492
rect 41916 37438 41918 37490
rect 41918 37438 41970 37490
rect 41970 37438 41972 37490
rect 41916 37436 41972 37438
rect 44156 40124 44212 40180
rect 43372 39730 43428 39732
rect 43372 39678 43374 39730
rect 43374 39678 43426 39730
rect 43426 39678 43428 39730
rect 43372 39676 43428 39678
rect 43260 39564 43316 39620
rect 42476 37996 42532 38052
rect 42140 37100 42196 37156
rect 42252 37212 42308 37268
rect 41356 35196 41412 35252
rect 41804 36594 41860 36596
rect 41804 36542 41806 36594
rect 41806 36542 41858 36594
rect 41858 36542 41860 36594
rect 41804 36540 41860 36542
rect 42924 38668 42980 38724
rect 42812 38050 42868 38052
rect 42812 37998 42814 38050
rect 42814 37998 42866 38050
rect 42866 37998 42868 38050
rect 42812 37996 42868 37998
rect 42700 37436 42756 37492
rect 42924 37154 42980 37156
rect 42924 37102 42926 37154
rect 42926 37102 42978 37154
rect 42978 37102 42980 37154
rect 42924 37100 42980 37102
rect 42140 36370 42196 36372
rect 42140 36318 42142 36370
rect 42142 36318 42194 36370
rect 42194 36318 42196 36370
rect 42140 36316 42196 36318
rect 42812 36540 42868 36596
rect 43932 38722 43988 38724
rect 43932 38670 43934 38722
rect 43934 38670 43986 38722
rect 43986 38670 43988 38722
rect 43932 38668 43988 38670
rect 43820 38274 43876 38276
rect 43820 38222 43822 38274
rect 43822 38222 43874 38274
rect 43874 38222 43876 38274
rect 43820 38220 43876 38222
rect 44156 39676 44212 39732
rect 46508 54012 46564 54068
rect 47852 56082 47908 56084
rect 47852 56030 47854 56082
rect 47854 56030 47906 56082
rect 47906 56030 47908 56082
rect 47852 56028 47908 56030
rect 47628 55858 47684 55860
rect 47628 55806 47630 55858
rect 47630 55806 47682 55858
rect 47682 55806 47684 55858
rect 47628 55804 47684 55806
rect 47516 52834 47572 52836
rect 47516 52782 47518 52834
rect 47518 52782 47570 52834
rect 47570 52782 47572 52834
rect 47516 52780 47572 52782
rect 47740 52556 47796 52612
rect 47404 51490 47460 51492
rect 47404 51438 47406 51490
rect 47406 51438 47458 51490
rect 47458 51438 47460 51490
rect 47404 51436 47460 51438
rect 46844 50482 46900 50484
rect 46844 50430 46846 50482
rect 46846 50430 46898 50482
rect 46898 50430 46900 50482
rect 46844 50428 46900 50430
rect 46396 49922 46452 49924
rect 46396 49870 46398 49922
rect 46398 49870 46450 49922
rect 46450 49870 46452 49922
rect 46396 49868 46452 49870
rect 46732 49810 46788 49812
rect 46732 49758 46734 49810
rect 46734 49758 46786 49810
rect 46786 49758 46788 49810
rect 46732 49756 46788 49758
rect 48076 53452 48132 53508
rect 47964 52556 48020 52612
rect 47852 50428 47908 50484
rect 46284 49698 46340 49700
rect 46284 49646 46286 49698
rect 46286 49646 46338 49698
rect 46338 49646 46340 49698
rect 46284 49644 46340 49646
rect 47404 49196 47460 49252
rect 45836 48802 45892 48804
rect 45836 48750 45838 48802
rect 45838 48750 45890 48802
rect 45890 48750 45892 48802
rect 45836 48748 45892 48750
rect 46396 48972 46452 49028
rect 45948 48524 46004 48580
rect 46060 47180 46116 47236
rect 45836 45890 45892 45892
rect 45836 45838 45838 45890
rect 45838 45838 45890 45890
rect 45890 45838 45892 45890
rect 45836 45836 45892 45838
rect 46172 45276 46228 45332
rect 46284 45164 46340 45220
rect 46172 44044 46228 44100
rect 47628 49026 47684 49028
rect 47628 48974 47630 49026
rect 47630 48974 47682 49026
rect 47682 48974 47684 49026
rect 47628 48972 47684 48974
rect 48300 50204 48356 50260
rect 46620 48300 46676 48356
rect 47404 48802 47460 48804
rect 47404 48750 47406 48802
rect 47406 48750 47458 48802
rect 47458 48750 47460 48802
rect 47404 48748 47460 48750
rect 48188 48802 48244 48804
rect 48188 48750 48190 48802
rect 48190 48750 48242 48802
rect 48242 48750 48244 48802
rect 48188 48748 48244 48750
rect 48076 48636 48132 48692
rect 47404 48354 47460 48356
rect 47404 48302 47406 48354
rect 47406 48302 47458 48354
rect 47458 48302 47460 48354
rect 47404 48300 47460 48302
rect 46844 47570 46900 47572
rect 46844 47518 46846 47570
rect 46846 47518 46898 47570
rect 46898 47518 46900 47570
rect 46844 47516 46900 47518
rect 47964 47516 48020 47572
rect 47404 47458 47460 47460
rect 47404 47406 47406 47458
rect 47406 47406 47458 47458
rect 47458 47406 47460 47458
rect 47404 47404 47460 47406
rect 46620 47292 46676 47348
rect 47628 47346 47684 47348
rect 47628 47294 47630 47346
rect 47630 47294 47682 47346
rect 47682 47294 47684 47346
rect 47628 47292 47684 47294
rect 46508 45106 46564 45108
rect 46508 45054 46510 45106
rect 46510 45054 46562 45106
rect 46562 45054 46564 45106
rect 46508 45052 46564 45054
rect 45724 41916 45780 41972
rect 46060 42028 46116 42084
rect 45724 41746 45780 41748
rect 45724 41694 45726 41746
rect 45726 41694 45778 41746
rect 45778 41694 45780 41746
rect 45724 41692 45780 41694
rect 45388 40348 45444 40404
rect 45612 40460 45668 40516
rect 45500 40290 45556 40292
rect 45500 40238 45502 40290
rect 45502 40238 45554 40290
rect 45554 40238 45556 40290
rect 45500 40236 45556 40238
rect 45836 40178 45892 40180
rect 45836 40126 45838 40178
rect 45838 40126 45890 40178
rect 45890 40126 45892 40178
rect 45836 40124 45892 40126
rect 46172 40460 46228 40516
rect 47628 45500 47684 45556
rect 46732 44940 46788 44996
rect 47516 44994 47572 44996
rect 47516 44942 47518 44994
rect 47518 44942 47570 44994
rect 47570 44942 47572 44994
rect 47516 44940 47572 44942
rect 46620 44380 46676 44436
rect 47180 44828 47236 44884
rect 47292 44380 47348 44436
rect 47180 44044 47236 44100
rect 47740 44882 47796 44884
rect 47740 44830 47742 44882
rect 47742 44830 47794 44882
rect 47794 44830 47796 44882
rect 47740 44828 47796 44830
rect 48188 44380 48244 44436
rect 47180 42530 47236 42532
rect 47180 42478 47182 42530
rect 47182 42478 47234 42530
rect 47234 42478 47236 42530
rect 47180 42476 47236 42478
rect 47068 42082 47124 42084
rect 47068 42030 47070 42082
rect 47070 42030 47122 42082
rect 47122 42030 47124 42082
rect 47068 42028 47124 42030
rect 46396 40236 46452 40292
rect 48076 41970 48132 41972
rect 48076 41918 48078 41970
rect 48078 41918 48130 41970
rect 48130 41918 48132 41970
rect 48076 41916 48132 41918
rect 46956 40124 47012 40180
rect 47068 40012 47124 40068
rect 45500 39452 45556 39508
rect 43372 37324 43428 37380
rect 43596 37378 43652 37380
rect 43596 37326 43598 37378
rect 43598 37326 43650 37378
rect 43650 37326 43652 37378
rect 43596 37324 43652 37326
rect 42700 35308 42756 35364
rect 41468 34188 41524 34244
rect 40796 33516 40852 33572
rect 40236 27186 40292 27188
rect 40236 27134 40238 27186
rect 40238 27134 40290 27186
rect 40290 27134 40292 27186
rect 40236 27132 40292 27134
rect 41244 33404 41300 33460
rect 41020 33234 41076 33236
rect 41020 33182 41022 33234
rect 41022 33182 41074 33234
rect 41074 33182 41076 33234
rect 41020 33180 41076 33182
rect 41692 34018 41748 34020
rect 41692 33966 41694 34018
rect 41694 33966 41746 34018
rect 41746 33966 41748 34018
rect 41692 33964 41748 33966
rect 41356 33292 41412 33348
rect 41692 33404 41748 33460
rect 41468 31836 41524 31892
rect 41580 31724 41636 31780
rect 42028 31666 42084 31668
rect 42028 31614 42030 31666
rect 42030 31614 42082 31666
rect 42082 31614 42084 31666
rect 42028 31612 42084 31614
rect 41804 31164 41860 31220
rect 42476 31218 42532 31220
rect 42476 31166 42478 31218
rect 42478 31166 42530 31218
rect 42530 31166 42532 31218
rect 42476 31164 42532 31166
rect 41356 29986 41412 29988
rect 41356 29934 41358 29986
rect 41358 29934 41410 29986
rect 41410 29934 41412 29986
rect 41356 29932 41412 29934
rect 40348 26908 40404 26964
rect 40348 25900 40404 25956
rect 40908 28476 40964 28532
rect 41020 27132 41076 27188
rect 41356 27692 41412 27748
rect 42812 31106 42868 31108
rect 42812 31054 42814 31106
rect 42814 31054 42866 31106
rect 42866 31054 42868 31106
rect 42812 31052 42868 31054
rect 42252 29932 42308 29988
rect 43260 35420 43316 35476
rect 43260 35084 43316 35140
rect 43820 35196 43876 35252
rect 43484 34690 43540 34692
rect 43484 34638 43486 34690
rect 43486 34638 43538 34690
rect 43538 34638 43540 34690
rect 43484 34636 43540 34638
rect 43260 34076 43316 34132
rect 43148 33458 43204 33460
rect 43148 33406 43150 33458
rect 43150 33406 43202 33458
rect 43202 33406 43204 33458
rect 43148 33404 43204 33406
rect 43260 33292 43316 33348
rect 44380 34636 44436 34692
rect 43820 34076 43876 34132
rect 43484 32674 43540 32676
rect 43484 32622 43486 32674
rect 43486 32622 43538 32674
rect 43538 32622 43540 32674
rect 43484 32620 43540 32622
rect 43596 32172 43652 32228
rect 43372 31724 43428 31780
rect 43260 31052 43316 31108
rect 44268 34018 44324 34020
rect 44268 33966 44270 34018
rect 44270 33966 44322 34018
rect 44322 33966 44324 34018
rect 44268 33964 44324 33966
rect 44716 33292 44772 33348
rect 44940 33234 44996 33236
rect 44940 33182 44942 33234
rect 44942 33182 44994 33234
rect 44994 33182 44996 33234
rect 44940 33180 44996 33182
rect 44604 33068 44660 33124
rect 44044 32674 44100 32676
rect 44044 32622 44046 32674
rect 44046 32622 44098 32674
rect 44098 32622 44100 32674
rect 44044 32620 44100 32622
rect 44604 32172 44660 32228
rect 44268 32060 44324 32116
rect 43596 31052 43652 31108
rect 43820 31612 43876 31668
rect 44940 32674 44996 32676
rect 44940 32622 44942 32674
rect 44942 32622 44994 32674
rect 44994 32622 44996 32674
rect 44940 32620 44996 32622
rect 44604 31164 44660 31220
rect 44828 31106 44884 31108
rect 44828 31054 44830 31106
rect 44830 31054 44882 31106
rect 44882 31054 44884 31106
rect 44828 31052 44884 31054
rect 43036 29708 43092 29764
rect 42364 29260 42420 29316
rect 42924 29314 42980 29316
rect 42924 29262 42926 29314
rect 42926 29262 42978 29314
rect 42978 29262 42980 29314
rect 42924 29260 42980 29262
rect 42588 28588 42644 28644
rect 42140 27970 42196 27972
rect 42140 27918 42142 27970
rect 42142 27918 42194 27970
rect 42194 27918 42196 27970
rect 42140 27916 42196 27918
rect 42476 27916 42532 27972
rect 41916 26796 41972 26852
rect 41132 26460 41188 26516
rect 41244 26684 41300 26740
rect 41132 25900 41188 25956
rect 41356 25452 41412 25508
rect 41916 25506 41972 25508
rect 41916 25454 41918 25506
rect 41918 25454 41970 25506
rect 41970 25454 41972 25506
rect 41916 25452 41972 25454
rect 41580 24556 41636 24612
rect 40908 22988 40964 23044
rect 40460 22652 40516 22708
rect 41580 22988 41636 23044
rect 39004 20748 39060 20804
rect 39564 20748 39620 20804
rect 39228 20578 39284 20580
rect 39228 20526 39230 20578
rect 39230 20526 39282 20578
rect 39282 20526 39284 20578
rect 39228 20524 39284 20526
rect 38892 20188 38948 20244
rect 38108 20076 38164 20132
rect 38892 19852 38948 19908
rect 37996 18956 38052 19012
rect 38220 18396 38276 18452
rect 38668 19010 38724 19012
rect 38668 18958 38670 19010
rect 38670 18958 38722 19010
rect 38722 18958 38724 19010
rect 38668 18956 38724 18958
rect 37884 17836 37940 17892
rect 37548 16098 37604 16100
rect 37548 16046 37550 16098
rect 37550 16046 37602 16098
rect 37602 16046 37604 16098
rect 37548 16044 37604 16046
rect 37660 15708 37716 15764
rect 38444 17164 38500 17220
rect 37884 16882 37940 16884
rect 37884 16830 37886 16882
rect 37886 16830 37938 16882
rect 37938 16830 37940 16882
rect 37884 16828 37940 16830
rect 37436 15484 37492 15540
rect 38556 16716 38612 16772
rect 38780 18396 38836 18452
rect 39228 19628 39284 19684
rect 39676 20076 39732 20132
rect 39116 19516 39172 19572
rect 41020 22204 41076 22260
rect 40348 21810 40404 21812
rect 40348 21758 40350 21810
rect 40350 21758 40402 21810
rect 40402 21758 40404 21810
rect 40348 21756 40404 21758
rect 40236 20524 40292 20580
rect 40796 21644 40852 21700
rect 41916 22204 41972 22260
rect 41580 22146 41636 22148
rect 41580 22094 41582 22146
rect 41582 22094 41634 22146
rect 41634 22094 41636 22146
rect 41580 22092 41636 22094
rect 41804 22146 41860 22148
rect 41804 22094 41806 22146
rect 41806 22094 41858 22146
rect 41858 22094 41860 22146
rect 41804 22092 41860 22094
rect 42364 26514 42420 26516
rect 42364 26462 42366 26514
rect 42366 26462 42418 26514
rect 42418 26462 42420 26514
rect 42364 26460 42420 26462
rect 42924 28476 42980 28532
rect 42812 27970 42868 27972
rect 42812 27918 42814 27970
rect 42814 27918 42866 27970
rect 42866 27918 42868 27970
rect 42812 27916 42868 27918
rect 43484 29708 43540 29764
rect 43484 28588 43540 28644
rect 44044 30044 44100 30100
rect 43596 28476 43652 28532
rect 42924 26460 42980 26516
rect 43596 27692 43652 27748
rect 43148 26796 43204 26852
rect 43036 25452 43092 25508
rect 43372 25506 43428 25508
rect 43372 25454 43374 25506
rect 43374 25454 43426 25506
rect 43426 25454 43428 25506
rect 43372 25452 43428 25454
rect 43708 25452 43764 25508
rect 43932 24892 43988 24948
rect 43708 23324 43764 23380
rect 43148 22988 43204 23044
rect 42140 21980 42196 22036
rect 40796 20636 40852 20692
rect 41244 20524 41300 20580
rect 40012 19906 40068 19908
rect 40012 19854 40014 19906
rect 40014 19854 40066 19906
rect 40066 19854 40068 19906
rect 40012 19852 40068 19854
rect 40236 19852 40292 19908
rect 41020 19906 41076 19908
rect 41020 19854 41022 19906
rect 41022 19854 41074 19906
rect 41074 19854 41076 19906
rect 41020 19852 41076 19854
rect 41132 19740 41188 19796
rect 40460 19516 40516 19572
rect 40012 18396 40068 18452
rect 38892 17554 38948 17556
rect 38892 17502 38894 17554
rect 38894 17502 38946 17554
rect 38946 17502 38948 17554
rect 38892 17500 38948 17502
rect 38780 16882 38836 16884
rect 38780 16830 38782 16882
rect 38782 16830 38834 16882
rect 38834 16830 38836 16882
rect 38780 16828 38836 16830
rect 38556 15708 38612 15764
rect 38108 15372 38164 15428
rect 36764 13468 36820 13524
rect 38332 15202 38388 15204
rect 38332 15150 38334 15202
rect 38334 15150 38386 15202
rect 38386 15150 38388 15202
rect 38332 15148 38388 15150
rect 38668 15372 38724 15428
rect 38556 15148 38612 15204
rect 37772 13020 37828 13076
rect 37436 12908 37492 12964
rect 39452 18060 39508 18116
rect 40348 18284 40404 18340
rect 39116 17666 39172 17668
rect 39116 17614 39118 17666
rect 39118 17614 39170 17666
rect 39170 17614 39172 17666
rect 39116 17612 39172 17614
rect 39788 16940 39844 16996
rect 39564 16882 39620 16884
rect 39564 16830 39566 16882
rect 39566 16830 39618 16882
rect 39618 16830 39620 16882
rect 39564 16828 39620 16830
rect 39116 16492 39172 16548
rect 39004 16044 39060 16100
rect 39564 16156 39620 16212
rect 39228 15484 39284 15540
rect 39452 15820 39508 15876
rect 38892 15426 38948 15428
rect 38892 15374 38894 15426
rect 38894 15374 38946 15426
rect 38946 15374 38948 15426
rect 38892 15372 38948 15374
rect 38780 13580 38836 13636
rect 38892 14924 38948 14980
rect 37772 12178 37828 12180
rect 37772 12126 37774 12178
rect 37774 12126 37826 12178
rect 37826 12126 37828 12178
rect 37772 12124 37828 12126
rect 38556 13468 38612 13524
rect 36988 11170 37044 11172
rect 36988 11118 36990 11170
rect 36990 11118 37042 11170
rect 37042 11118 37044 11170
rect 36988 11116 37044 11118
rect 36540 9772 36596 9828
rect 36428 8034 36484 8036
rect 36428 7982 36430 8034
rect 36430 7982 36482 8034
rect 36482 7982 36484 8034
rect 36428 7980 36484 7982
rect 36540 7756 36596 7812
rect 36876 6636 36932 6692
rect 36540 6524 36596 6580
rect 36540 6300 36596 6356
rect 36316 6018 36372 6020
rect 36316 5966 36318 6018
rect 36318 5966 36370 6018
rect 36370 5966 36372 6018
rect 36316 5964 36372 5966
rect 36652 5740 36708 5796
rect 37324 10332 37380 10388
rect 37212 10108 37268 10164
rect 37324 9324 37380 9380
rect 38108 11564 38164 11620
rect 37660 11452 37716 11508
rect 38780 11676 38836 11732
rect 38780 11452 38836 11508
rect 38556 11282 38612 11284
rect 38556 11230 38558 11282
rect 38558 11230 38610 11282
rect 38610 11230 38612 11282
rect 38556 11228 38612 11230
rect 37660 10722 37716 10724
rect 37660 10670 37662 10722
rect 37662 10670 37714 10722
rect 37714 10670 37716 10722
rect 37660 10668 37716 10670
rect 39900 16098 39956 16100
rect 39900 16046 39902 16098
rect 39902 16046 39954 16098
rect 39954 16046 39956 16098
rect 39900 16044 39956 16046
rect 39788 15596 39844 15652
rect 40236 15538 40292 15540
rect 40236 15486 40238 15538
rect 40238 15486 40290 15538
rect 40290 15486 40292 15538
rect 40236 15484 40292 15486
rect 39116 15148 39172 15204
rect 41356 20018 41412 20020
rect 41356 19966 41358 20018
rect 41358 19966 41410 20018
rect 41410 19966 41412 20018
rect 41356 19964 41412 19966
rect 42140 20076 42196 20132
rect 42476 22258 42532 22260
rect 42476 22206 42478 22258
rect 42478 22206 42530 22258
rect 42530 22206 42532 22258
rect 42476 22204 42532 22206
rect 42588 21980 42644 22036
rect 41916 20018 41972 20020
rect 41916 19966 41918 20018
rect 41918 19966 41970 20018
rect 41970 19966 41972 20018
rect 41916 19964 41972 19966
rect 41804 19628 41860 19684
rect 42252 19516 42308 19572
rect 42700 20690 42756 20692
rect 42700 20638 42702 20690
rect 42702 20638 42754 20690
rect 42754 20638 42756 20690
rect 42700 20636 42756 20638
rect 43148 20690 43204 20692
rect 43148 20638 43150 20690
rect 43150 20638 43202 20690
rect 43202 20638 43204 20690
rect 43148 20636 43204 20638
rect 43596 21420 43652 21476
rect 43708 22092 43764 22148
rect 43260 20130 43316 20132
rect 43260 20078 43262 20130
rect 43262 20078 43314 20130
rect 43314 20078 43316 20130
rect 43260 20076 43316 20078
rect 42812 19740 42868 19796
rect 42140 18956 42196 19012
rect 41804 18732 41860 18788
rect 40908 18450 40964 18452
rect 40908 18398 40910 18450
rect 40910 18398 40962 18450
rect 40962 18398 40964 18450
rect 40908 18396 40964 18398
rect 41020 17276 41076 17332
rect 41356 17164 41412 17220
rect 41132 16994 41188 16996
rect 41132 16942 41134 16994
rect 41134 16942 41186 16994
rect 41186 16942 41188 16994
rect 41132 16940 41188 16942
rect 40908 16882 40964 16884
rect 40908 16830 40910 16882
rect 40910 16830 40962 16882
rect 40962 16830 40964 16882
rect 40908 16828 40964 16830
rect 41020 15596 41076 15652
rect 41692 18396 41748 18452
rect 41468 16604 41524 16660
rect 41804 17554 41860 17556
rect 41804 17502 41806 17554
rect 41806 17502 41858 17554
rect 41858 17502 41860 17554
rect 41804 17500 41860 17502
rect 41580 16380 41636 16436
rect 41692 16492 41748 16548
rect 41580 15538 41636 15540
rect 41580 15486 41582 15538
rect 41582 15486 41634 15538
rect 41634 15486 41636 15538
rect 41580 15484 41636 15486
rect 41020 15148 41076 15204
rect 39340 14140 39396 14196
rect 39116 11564 39172 11620
rect 38892 11394 38948 11396
rect 38892 11342 38894 11394
rect 38894 11342 38946 11394
rect 38946 11342 38948 11394
rect 38892 11340 38948 11342
rect 40012 11394 40068 11396
rect 40012 11342 40014 11394
rect 40014 11342 40066 11394
rect 40066 11342 40068 11394
rect 40012 11340 40068 11342
rect 42700 18956 42756 19012
rect 42476 18562 42532 18564
rect 42476 18510 42478 18562
rect 42478 18510 42530 18562
rect 42530 18510 42532 18562
rect 42476 18508 42532 18510
rect 42252 17164 42308 17220
rect 42140 16044 42196 16100
rect 42252 16940 42308 16996
rect 41916 15372 41972 15428
rect 42028 15820 42084 15876
rect 42252 15314 42308 15316
rect 42252 15262 42254 15314
rect 42254 15262 42306 15314
rect 42306 15262 42308 15314
rect 42252 15260 42308 15262
rect 42364 15932 42420 15988
rect 41916 15148 41972 15204
rect 42588 18338 42644 18340
rect 42588 18286 42590 18338
rect 42590 18286 42642 18338
rect 42642 18286 42644 18338
rect 42588 18284 42644 18286
rect 42924 18450 42980 18452
rect 42924 18398 42926 18450
rect 42926 18398 42978 18450
rect 42978 18398 42980 18450
rect 42924 18396 42980 18398
rect 43932 20690 43988 20692
rect 43932 20638 43934 20690
rect 43934 20638 43986 20690
rect 43986 20638 43988 20690
rect 43932 20636 43988 20638
rect 44604 28476 44660 28532
rect 44268 27746 44324 27748
rect 44268 27694 44270 27746
rect 44270 27694 44322 27746
rect 44322 27694 44324 27746
rect 44268 27692 44324 27694
rect 44940 27020 44996 27076
rect 45276 38220 45332 38276
rect 46732 39676 46788 39732
rect 45948 38834 46004 38836
rect 45948 38782 45950 38834
rect 45950 38782 46002 38834
rect 46002 38782 46004 38834
rect 45948 38780 46004 38782
rect 46172 37996 46228 38052
rect 45388 37938 45444 37940
rect 45388 37886 45390 37938
rect 45390 37886 45442 37938
rect 45442 37886 45444 37938
rect 45388 37884 45444 37886
rect 45388 35196 45444 35252
rect 45388 33180 45444 33236
rect 45276 33068 45332 33124
rect 45276 32674 45332 32676
rect 45276 32622 45278 32674
rect 45278 32622 45330 32674
rect 45330 32622 45332 32674
rect 45276 32620 45332 32622
rect 45724 35420 45780 35476
rect 45612 33180 45668 33236
rect 45164 31164 45220 31220
rect 45388 30156 45444 30212
rect 45388 29932 45444 29988
rect 45612 29932 45668 29988
rect 45724 29708 45780 29764
rect 45276 27746 45332 27748
rect 45276 27694 45278 27746
rect 45278 27694 45330 27746
rect 45330 27694 45332 27746
rect 45276 27692 45332 27694
rect 45052 26124 45108 26180
rect 45052 25116 45108 25172
rect 44828 24946 44884 24948
rect 44828 24894 44830 24946
rect 44830 24894 44882 24946
rect 44882 24894 44884 24946
rect 44828 24892 44884 24894
rect 45164 24892 45220 24948
rect 45052 24834 45108 24836
rect 45052 24782 45054 24834
rect 45054 24782 45106 24834
rect 45106 24782 45108 24834
rect 45052 24780 45108 24782
rect 44604 24668 44660 24724
rect 45276 24668 45332 24724
rect 45388 25116 45444 25172
rect 45612 24834 45668 24836
rect 45612 24782 45614 24834
rect 45614 24782 45666 24834
rect 45666 24782 45668 24834
rect 45612 24780 45668 24782
rect 45724 24722 45780 24724
rect 45724 24670 45726 24722
rect 45726 24670 45778 24722
rect 45778 24670 45780 24722
rect 45724 24668 45780 24670
rect 45388 24556 45444 24612
rect 46284 37324 46340 37380
rect 46508 37212 46564 37268
rect 47180 39900 47236 39956
rect 47068 39676 47124 39732
rect 47516 40460 47572 40516
rect 47964 40460 48020 40516
rect 47404 40124 47460 40180
rect 46732 39506 46788 39508
rect 46732 39454 46734 39506
rect 46734 39454 46786 39506
rect 46786 39454 46788 39506
rect 46732 39452 46788 39454
rect 46732 38780 46788 38836
rect 47628 39618 47684 39620
rect 47628 39566 47630 39618
rect 47630 39566 47682 39618
rect 47682 39566 47684 39618
rect 47628 39564 47684 39566
rect 47404 38780 47460 38836
rect 46844 38050 46900 38052
rect 46844 37998 46846 38050
rect 46846 37998 46898 38050
rect 46898 37998 46900 38050
rect 46844 37996 46900 37998
rect 47292 37884 47348 37940
rect 47180 37378 47236 37380
rect 47180 37326 47182 37378
rect 47182 37326 47234 37378
rect 47234 37326 47236 37378
rect 47180 37324 47236 37326
rect 46844 36988 46900 37044
rect 47068 37266 47124 37268
rect 47068 37214 47070 37266
rect 47070 37214 47122 37266
rect 47122 37214 47124 37266
rect 47068 37212 47124 37214
rect 46956 36258 47012 36260
rect 46956 36206 46958 36258
rect 46958 36206 47010 36258
rect 47010 36206 47012 36258
rect 46956 36204 47012 36206
rect 45948 35474 46004 35476
rect 45948 35422 45950 35474
rect 45950 35422 46002 35474
rect 46002 35422 46004 35474
rect 45948 35420 46004 35422
rect 47180 37154 47236 37156
rect 47180 37102 47182 37154
rect 47182 37102 47234 37154
rect 47234 37102 47236 37154
rect 47180 37100 47236 37102
rect 48188 40514 48244 40516
rect 48188 40462 48190 40514
rect 48190 40462 48242 40514
rect 48242 40462 48244 40514
rect 48188 40460 48244 40462
rect 47964 40012 48020 40068
rect 48412 42476 48468 42532
rect 48076 38834 48132 38836
rect 48076 38782 48078 38834
rect 48078 38782 48130 38834
rect 48130 38782 48132 38834
rect 48076 38780 48132 38782
rect 47516 36204 47572 36260
rect 48188 38668 48244 38724
rect 47852 36988 47908 37044
rect 48188 36204 48244 36260
rect 46844 33964 46900 34020
rect 46284 33068 46340 33124
rect 48188 34018 48244 34020
rect 48188 33966 48190 34018
rect 48190 33966 48242 34018
rect 48242 33966 48244 34018
rect 48188 33964 48244 33966
rect 46396 32620 46452 32676
rect 46060 31666 46116 31668
rect 46060 31614 46062 31666
rect 46062 31614 46114 31666
rect 46114 31614 46116 31666
rect 46060 31612 46116 31614
rect 46060 30156 46116 30212
rect 47852 32844 47908 32900
rect 47628 32732 47684 32788
rect 48188 32732 48244 32788
rect 47404 32674 47460 32676
rect 47404 32622 47406 32674
rect 47406 32622 47458 32674
rect 47458 32622 47460 32674
rect 47404 32620 47460 32622
rect 46844 31612 46900 31668
rect 47180 31106 47236 31108
rect 47180 31054 47182 31106
rect 47182 31054 47234 31106
rect 47234 31054 47236 31106
rect 47180 31052 47236 31054
rect 47628 31052 47684 31108
rect 47068 30940 47124 30996
rect 46396 30828 46452 30884
rect 47740 30994 47796 30996
rect 47740 30942 47742 30994
rect 47742 30942 47794 30994
rect 47794 30942 47796 30994
rect 47740 30940 47796 30942
rect 47292 30828 47348 30884
rect 46396 28364 46452 28420
rect 47180 29986 47236 29988
rect 47180 29934 47182 29986
rect 47182 29934 47234 29986
rect 47234 29934 47236 29986
rect 47180 29932 47236 29934
rect 46508 27692 46564 27748
rect 46284 27074 46340 27076
rect 46284 27022 46286 27074
rect 46286 27022 46338 27074
rect 46338 27022 46340 27074
rect 46284 27020 46340 27022
rect 44940 23436 44996 23492
rect 45164 23324 45220 23380
rect 44716 23266 44772 23268
rect 44716 23214 44718 23266
rect 44718 23214 44770 23266
rect 44770 23214 44772 23266
rect 44716 23212 44772 23214
rect 44268 23042 44324 23044
rect 44268 22990 44270 23042
rect 44270 22990 44322 23042
rect 44322 22990 44324 23042
rect 44268 22988 44324 22990
rect 45948 26908 46004 26964
rect 45612 23772 45668 23828
rect 44940 22988 44996 23044
rect 44156 21980 44212 22036
rect 44716 21474 44772 21476
rect 44716 21422 44718 21474
rect 44718 21422 44770 21474
rect 44770 21422 44772 21474
rect 44716 21420 44772 21422
rect 44380 20860 44436 20916
rect 44268 20300 44324 20356
rect 44940 20914 44996 20916
rect 44940 20862 44942 20914
rect 44942 20862 44994 20914
rect 44994 20862 44996 20914
rect 44940 20860 44996 20862
rect 45276 21756 45332 21812
rect 45500 21308 45556 21364
rect 45388 20860 45444 20916
rect 44380 20076 44436 20132
rect 43708 20018 43764 20020
rect 43708 19966 43710 20018
rect 43710 19966 43762 20018
rect 43762 19966 43764 20018
rect 43708 19964 43764 19966
rect 43708 19404 43764 19460
rect 44268 19906 44324 19908
rect 44268 19854 44270 19906
rect 44270 19854 44322 19906
rect 44322 19854 44324 19906
rect 44268 19852 44324 19854
rect 43372 19122 43428 19124
rect 43372 19070 43374 19122
rect 43374 19070 43426 19122
rect 43426 19070 43428 19122
rect 43372 19068 43428 19070
rect 43372 18396 43428 18452
rect 42924 17276 42980 17332
rect 42700 17052 42756 17108
rect 43036 16940 43092 16996
rect 43596 18450 43652 18452
rect 43596 18398 43598 18450
rect 43598 18398 43650 18450
rect 43650 18398 43652 18450
rect 43596 18396 43652 18398
rect 44268 19180 44324 19236
rect 43596 17612 43652 17668
rect 43932 18338 43988 18340
rect 43932 18286 43934 18338
rect 43934 18286 43986 18338
rect 43986 18286 43988 18338
rect 43932 18284 43988 18286
rect 44828 19068 44884 19124
rect 45276 20300 45332 20356
rect 45052 20018 45108 20020
rect 45052 19966 45054 20018
rect 45054 19966 45106 20018
rect 45106 19966 45108 20018
rect 45052 19964 45108 19966
rect 44940 18620 44996 18676
rect 44380 18284 44436 18340
rect 44044 18226 44100 18228
rect 44044 18174 44046 18226
rect 44046 18174 44098 18226
rect 44098 18174 44100 18226
rect 44044 18172 44100 18174
rect 44828 18450 44884 18452
rect 44828 18398 44830 18450
rect 44830 18398 44882 18450
rect 44882 18398 44884 18450
rect 44828 18396 44884 18398
rect 45164 18508 45220 18564
rect 43708 17724 43764 17780
rect 45052 18172 45108 18228
rect 43484 17388 43540 17444
rect 43372 17052 43428 17108
rect 43596 17276 43652 17332
rect 43820 17106 43876 17108
rect 43820 17054 43822 17106
rect 43822 17054 43874 17106
rect 43874 17054 43876 17106
rect 43820 17052 43876 17054
rect 43260 16828 43316 16884
rect 43148 16716 43204 16772
rect 42924 16604 42980 16660
rect 43148 16492 43204 16548
rect 43036 15596 43092 15652
rect 42588 15484 42644 15540
rect 41132 13020 41188 13076
rect 41916 12572 41972 12628
rect 42028 12684 42084 12740
rect 40236 11676 40292 11732
rect 38892 10834 38948 10836
rect 38892 10782 38894 10834
rect 38894 10782 38946 10834
rect 38946 10782 38948 10834
rect 38892 10780 38948 10782
rect 39564 11004 39620 11060
rect 39676 11116 39732 11172
rect 37548 10108 37604 10164
rect 39564 10556 39620 10612
rect 38108 9324 38164 9380
rect 37772 8930 37828 8932
rect 37772 8878 37774 8930
rect 37774 8878 37826 8930
rect 37826 8878 37828 8930
rect 37772 8876 37828 8878
rect 37660 8316 37716 8372
rect 37100 7980 37156 8036
rect 37548 7980 37604 8036
rect 37548 6578 37604 6580
rect 37548 6526 37550 6578
rect 37550 6526 37602 6578
rect 37602 6526 37604 6578
rect 37548 6524 37604 6526
rect 37772 6578 37828 6580
rect 37772 6526 37774 6578
rect 37774 6526 37826 6578
rect 37826 6526 37828 6578
rect 37772 6524 37828 6526
rect 37996 7532 38052 7588
rect 40236 11004 40292 11060
rect 40572 10780 40628 10836
rect 42028 12236 42084 12292
rect 41132 11452 41188 11508
rect 41132 11228 41188 11284
rect 41468 11340 41524 11396
rect 40796 10668 40852 10724
rect 40012 10610 40068 10612
rect 40012 10558 40014 10610
rect 40014 10558 40066 10610
rect 40066 10558 40068 10610
rect 40012 10556 40068 10558
rect 40236 10610 40292 10612
rect 40236 10558 40238 10610
rect 40238 10558 40290 10610
rect 40290 10558 40292 10610
rect 40236 10556 40292 10558
rect 39788 9100 39844 9156
rect 39676 8258 39732 8260
rect 39676 8206 39678 8258
rect 39678 8206 39730 8258
rect 39730 8206 39732 8258
rect 39676 8204 39732 8206
rect 39004 7980 39060 8036
rect 38892 7698 38948 7700
rect 38892 7646 38894 7698
rect 38894 7646 38946 7698
rect 38946 7646 38948 7698
rect 38892 7644 38948 7646
rect 38668 7532 38724 7588
rect 39564 7532 39620 7588
rect 41132 10780 41188 10836
rect 41692 11282 41748 11284
rect 41692 11230 41694 11282
rect 41694 11230 41746 11282
rect 41746 11230 41748 11282
rect 41692 11228 41748 11230
rect 42028 10722 42084 10724
rect 42028 10670 42030 10722
rect 42030 10670 42082 10722
rect 42082 10670 42084 10722
rect 42028 10668 42084 10670
rect 41356 10610 41412 10612
rect 41356 10558 41358 10610
rect 41358 10558 41410 10610
rect 41410 10558 41412 10610
rect 41356 10556 41412 10558
rect 43036 15372 43092 15428
rect 42700 15314 42756 15316
rect 42700 15262 42702 15314
rect 42702 15262 42754 15314
rect 42754 15262 42756 15314
rect 42700 15260 42756 15262
rect 44044 17724 44100 17780
rect 44156 17666 44212 17668
rect 44156 17614 44158 17666
rect 44158 17614 44210 17666
rect 44210 17614 44212 17666
rect 44156 17612 44212 17614
rect 44380 17500 44436 17556
rect 43932 16492 43988 16548
rect 44156 16492 44212 16548
rect 44044 16156 44100 16212
rect 43372 16044 43428 16100
rect 43708 16098 43764 16100
rect 43708 16046 43710 16098
rect 43710 16046 43762 16098
rect 43762 16046 43764 16098
rect 43708 16044 43764 16046
rect 43372 15874 43428 15876
rect 43372 15822 43374 15874
rect 43374 15822 43426 15874
rect 43426 15822 43428 15874
rect 43372 15820 43428 15822
rect 43596 15596 43652 15652
rect 43708 15314 43764 15316
rect 43708 15262 43710 15314
rect 43710 15262 43762 15314
rect 43762 15262 43764 15314
rect 43708 15260 43764 15262
rect 44156 15148 44212 15204
rect 42924 14812 42980 14868
rect 42364 12738 42420 12740
rect 42364 12686 42366 12738
rect 42366 12686 42418 12738
rect 42418 12686 42420 12738
rect 42364 12684 42420 12686
rect 42700 12572 42756 12628
rect 42252 11452 42308 11508
rect 42476 11170 42532 11172
rect 42476 11118 42478 11170
rect 42478 11118 42530 11170
rect 42530 11118 42532 11170
rect 42476 11116 42532 11118
rect 43036 14364 43092 14420
rect 44940 17554 44996 17556
rect 44940 17502 44942 17554
rect 44942 17502 44994 17554
rect 44994 17502 44996 17554
rect 44940 17500 44996 17502
rect 44380 15820 44436 15876
rect 44716 17276 44772 17332
rect 45164 17276 45220 17332
rect 45052 17164 45108 17220
rect 44716 16770 44772 16772
rect 44716 16718 44718 16770
rect 44718 16718 44770 16770
rect 44770 16718 44772 16770
rect 44716 16716 44772 16718
rect 45164 16268 45220 16324
rect 45052 16098 45108 16100
rect 45052 16046 45054 16098
rect 45054 16046 45106 16098
rect 45106 16046 45108 16098
rect 45052 16044 45108 16046
rect 44940 15986 44996 15988
rect 44940 15934 44942 15986
rect 44942 15934 44994 15986
rect 44994 15934 44996 15986
rect 44940 15932 44996 15934
rect 44828 15708 44884 15764
rect 44604 15260 44660 15316
rect 44268 14364 44324 14420
rect 44940 15148 44996 15204
rect 45164 15372 45220 15428
rect 45500 20076 45556 20132
rect 47180 28364 47236 28420
rect 47740 27020 47796 27076
rect 47852 26962 47908 26964
rect 47852 26910 47854 26962
rect 47854 26910 47906 26962
rect 47906 26910 47908 26962
rect 47852 26908 47908 26910
rect 48300 26908 48356 26964
rect 46284 24892 46340 24948
rect 46172 24610 46228 24612
rect 46172 24558 46174 24610
rect 46174 24558 46226 24610
rect 46226 24558 46228 24610
rect 46172 24556 46228 24558
rect 46172 23266 46228 23268
rect 46172 23214 46174 23266
rect 46174 23214 46226 23266
rect 46226 23214 46228 23266
rect 46172 23212 46228 23214
rect 46732 24668 46788 24724
rect 47516 24722 47572 24724
rect 47516 24670 47518 24722
rect 47518 24670 47570 24722
rect 47570 24670 47572 24722
rect 47516 24668 47572 24670
rect 46620 23324 46676 23380
rect 46060 21644 46116 21700
rect 46620 21810 46676 21812
rect 46620 21758 46622 21810
rect 46622 21758 46674 21810
rect 46674 21758 46676 21810
rect 46620 21756 46676 21758
rect 48300 24556 48356 24612
rect 46956 23826 47012 23828
rect 46956 23774 46958 23826
rect 46958 23774 47010 23826
rect 47010 23774 47012 23826
rect 46956 23772 47012 23774
rect 46844 23100 46900 23156
rect 46732 21644 46788 21700
rect 47740 23436 47796 23492
rect 47404 23154 47460 23156
rect 47404 23102 47406 23154
rect 47406 23102 47458 23154
rect 47458 23102 47460 23154
rect 47404 23100 47460 23102
rect 48076 23324 48132 23380
rect 47180 21810 47236 21812
rect 47180 21758 47182 21810
rect 47182 21758 47234 21810
rect 47234 21758 47236 21810
rect 47180 21756 47236 21758
rect 47068 21698 47124 21700
rect 47068 21646 47070 21698
rect 47070 21646 47122 21698
rect 47122 21646 47124 21698
rect 47068 21644 47124 21646
rect 46284 21084 46340 21140
rect 46844 20860 46900 20916
rect 45724 20018 45780 20020
rect 45724 19966 45726 20018
rect 45726 19966 45778 20018
rect 45778 19966 45780 20018
rect 45724 19964 45780 19966
rect 46172 20018 46228 20020
rect 46172 19966 46174 20018
rect 46174 19966 46226 20018
rect 46226 19966 46228 20018
rect 46172 19964 46228 19966
rect 46620 19852 46676 19908
rect 45388 17388 45444 17444
rect 45612 17164 45668 17220
rect 45500 16828 45556 16884
rect 45388 16604 45444 16660
rect 45388 16380 45444 16436
rect 45724 16268 45780 16324
rect 46396 18620 46452 18676
rect 46060 17554 46116 17556
rect 46060 17502 46062 17554
rect 46062 17502 46114 17554
rect 46114 17502 46116 17554
rect 46060 17500 46116 17502
rect 46060 17164 46116 17220
rect 45948 16604 46004 16660
rect 46284 16882 46340 16884
rect 46284 16830 46286 16882
rect 46286 16830 46338 16882
rect 46338 16830 46340 16882
rect 46284 16828 46340 16830
rect 46508 16828 46564 16884
rect 46060 16492 46116 16548
rect 47516 20130 47572 20132
rect 47516 20078 47518 20130
rect 47518 20078 47570 20130
rect 47570 20078 47572 20130
rect 47516 20076 47572 20078
rect 48188 21084 48244 21140
rect 48076 20860 48132 20916
rect 46956 18396 47012 18452
rect 46844 16716 46900 16772
rect 46732 16268 46788 16324
rect 48188 18396 48244 18452
rect 47180 17612 47236 17668
rect 48188 17612 48244 17668
rect 47852 17164 47908 17220
rect 47404 16716 47460 16772
rect 47852 16156 47908 16212
rect 47628 15874 47684 15876
rect 47628 15822 47630 15874
rect 47630 15822 47682 15874
rect 47682 15822 47684 15874
rect 47628 15820 47684 15822
rect 48188 15820 48244 15876
rect 48188 15260 48244 15316
rect 45276 15092 45332 15148
rect 44268 13634 44324 13636
rect 44268 13582 44270 13634
rect 44270 13582 44322 13634
rect 44322 13582 44324 13634
rect 44268 13580 44324 13582
rect 44716 13132 44772 13188
rect 44940 13746 44996 13748
rect 44940 13694 44942 13746
rect 44942 13694 44994 13746
rect 44994 13694 44996 13746
rect 44940 13692 44996 13694
rect 41244 10108 41300 10164
rect 42364 9996 42420 10052
rect 40236 8146 40292 8148
rect 40236 8094 40238 8146
rect 40238 8094 40290 8146
rect 40290 8094 40292 8146
rect 40236 8092 40292 8094
rect 41244 8092 41300 8148
rect 40124 6748 40180 6804
rect 38780 6578 38836 6580
rect 38780 6526 38782 6578
rect 38782 6526 38834 6578
rect 38834 6526 38836 6578
rect 38780 6524 38836 6526
rect 39788 6524 39844 6580
rect 36988 6188 37044 6244
rect 36092 5068 36148 5124
rect 35196 3946 35252 3948
rect 35196 3894 35198 3946
rect 35198 3894 35250 3946
rect 35250 3894 35252 3946
rect 35196 3892 35252 3894
rect 35300 3946 35356 3948
rect 35300 3894 35302 3946
rect 35302 3894 35354 3946
rect 35354 3894 35356 3946
rect 35300 3892 35356 3894
rect 35404 3946 35460 3948
rect 35404 3894 35406 3946
rect 35406 3894 35458 3946
rect 35458 3894 35460 3946
rect 35404 3892 35460 3894
rect 36428 4898 36484 4900
rect 36428 4846 36430 4898
rect 36430 4846 36482 4898
rect 36482 4846 36484 4898
rect 36428 4844 36484 4846
rect 37772 6018 37828 6020
rect 37772 5966 37774 6018
rect 37774 5966 37826 6018
rect 37826 5966 37828 6018
rect 37772 5964 37828 5966
rect 38332 6300 38388 6356
rect 39676 6466 39732 6468
rect 39676 6414 39678 6466
rect 39678 6414 39730 6466
rect 39730 6414 39732 6466
rect 39676 6412 39732 6414
rect 38556 6076 38612 6132
rect 38444 5964 38500 6020
rect 39004 5906 39060 5908
rect 39004 5854 39006 5906
rect 39006 5854 39058 5906
rect 39058 5854 39060 5906
rect 39004 5852 39060 5854
rect 39452 5906 39508 5908
rect 39452 5854 39454 5906
rect 39454 5854 39506 5906
rect 39506 5854 39508 5906
rect 39452 5852 39508 5854
rect 40012 6466 40068 6468
rect 40012 6414 40014 6466
rect 40014 6414 40066 6466
rect 40066 6414 40068 6466
rect 40012 6412 40068 6414
rect 39900 6300 39956 6356
rect 41244 7250 41300 7252
rect 41244 7198 41246 7250
rect 41246 7198 41298 7250
rect 41298 7198 41300 7250
rect 41244 7196 41300 7198
rect 40684 6802 40740 6804
rect 40684 6750 40686 6802
rect 40686 6750 40738 6802
rect 40738 6750 40740 6802
rect 40684 6748 40740 6750
rect 41356 6636 41412 6692
rect 41580 9660 41636 9716
rect 41692 9154 41748 9156
rect 41692 9102 41694 9154
rect 41694 9102 41746 9154
rect 41746 9102 41748 9154
rect 41692 9100 41748 9102
rect 41804 8316 41860 8372
rect 41468 7644 41524 7700
rect 41580 7980 41636 8036
rect 42364 8428 42420 8484
rect 42700 9660 42756 9716
rect 42812 10780 42868 10836
rect 42476 8764 42532 8820
rect 42028 7980 42084 8036
rect 42140 8146 42196 8148
rect 42140 8094 42142 8146
rect 42142 8094 42194 8146
rect 42194 8094 42196 8146
rect 42140 8092 42196 8094
rect 42252 8034 42308 8036
rect 42252 7982 42254 8034
rect 42254 7982 42306 8034
rect 42306 7982 42308 8034
rect 42252 7980 42308 7982
rect 42140 7532 42196 7588
rect 41692 7196 41748 7252
rect 41804 6860 41860 6916
rect 41692 6636 41748 6692
rect 40460 6524 40516 6580
rect 40460 6300 40516 6356
rect 40908 6412 40964 6468
rect 40236 6188 40292 6244
rect 40012 6076 40068 6132
rect 39900 5964 39956 6020
rect 38668 5740 38724 5796
rect 38444 5628 38500 5684
rect 38332 5292 38388 5348
rect 37548 5122 37604 5124
rect 37548 5070 37550 5122
rect 37550 5070 37602 5122
rect 37602 5070 37604 5122
rect 37548 5068 37604 5070
rect 38444 4844 38500 4900
rect 41020 6076 41076 6132
rect 41244 6412 41300 6468
rect 41580 6018 41636 6020
rect 41580 5966 41582 6018
rect 41582 5966 41634 6018
rect 41634 5966 41636 6018
rect 41580 5964 41636 5966
rect 41244 5740 41300 5796
rect 40796 5180 40852 5236
rect 40012 5122 40068 5124
rect 40012 5070 40014 5122
rect 40014 5070 40066 5122
rect 40066 5070 40068 5122
rect 40012 5068 40068 5070
rect 42140 6748 42196 6804
rect 42700 8146 42756 8148
rect 42700 8094 42702 8146
rect 42702 8094 42754 8146
rect 42754 8094 42756 8146
rect 42700 8092 42756 8094
rect 43372 11394 43428 11396
rect 43372 11342 43374 11394
rect 43374 11342 43426 11394
rect 43426 11342 43428 11394
rect 43372 11340 43428 11342
rect 43484 11282 43540 11284
rect 43484 11230 43486 11282
rect 43486 11230 43538 11282
rect 43538 11230 43540 11282
rect 43484 11228 43540 11230
rect 43820 11004 43876 11060
rect 43484 8876 43540 8932
rect 43260 8316 43316 8372
rect 43148 8258 43204 8260
rect 43148 8206 43150 8258
rect 43150 8206 43202 8258
rect 43202 8206 43204 8258
rect 43148 8204 43204 8206
rect 43372 8092 43428 8148
rect 42476 6914 42532 6916
rect 42476 6862 42478 6914
rect 42478 6862 42530 6914
rect 42530 6862 42532 6914
rect 42476 6860 42532 6862
rect 42252 6524 42308 6580
rect 41804 6188 41860 6244
rect 42588 6748 42644 6804
rect 41916 5964 41972 6020
rect 42812 6466 42868 6468
rect 42812 6414 42814 6466
rect 42814 6414 42866 6466
rect 42866 6414 42868 6466
rect 42812 6412 42868 6414
rect 41692 5234 41748 5236
rect 41692 5182 41694 5234
rect 41694 5182 41746 5234
rect 41746 5182 41748 5234
rect 41692 5180 41748 5182
rect 43148 7474 43204 7476
rect 43148 7422 43150 7474
rect 43150 7422 43202 7474
rect 43202 7422 43204 7474
rect 43148 7420 43204 7422
rect 43484 7586 43540 7588
rect 43484 7534 43486 7586
rect 43486 7534 43538 7586
rect 43538 7534 43540 7586
rect 43484 7532 43540 7534
rect 43820 8764 43876 8820
rect 43820 8092 43876 8148
rect 45388 13746 45444 13748
rect 45388 13694 45390 13746
rect 45390 13694 45442 13746
rect 45442 13694 45444 13746
rect 45388 13692 45444 13694
rect 45052 13580 45108 13636
rect 44828 11170 44884 11172
rect 44828 11118 44830 11170
rect 44830 11118 44882 11170
rect 44882 11118 44884 11170
rect 44828 11116 44884 11118
rect 44268 10332 44324 10388
rect 44940 10332 44996 10388
rect 45388 10332 45444 10388
rect 46956 13916 47012 13972
rect 45612 13132 45668 13188
rect 45724 13020 45780 13076
rect 47740 13074 47796 13076
rect 47740 13022 47742 13074
rect 47742 13022 47794 13074
rect 47794 13022 47796 13074
rect 47740 13020 47796 13022
rect 45948 10668 46004 10724
rect 44828 9884 44884 9940
rect 44940 9660 44996 9716
rect 44492 8930 44548 8932
rect 44492 8878 44494 8930
rect 44494 8878 44546 8930
rect 44546 8878 44548 8930
rect 44492 8876 44548 8878
rect 44044 8652 44100 8708
rect 45388 9714 45444 9716
rect 45388 9662 45390 9714
rect 45390 9662 45442 9714
rect 45442 9662 45444 9714
rect 45388 9660 45444 9662
rect 45276 9602 45332 9604
rect 45276 9550 45278 9602
rect 45278 9550 45330 9602
rect 45330 9550 45332 9602
rect 45276 9548 45332 9550
rect 45052 8652 45108 8708
rect 44828 8316 44884 8372
rect 43932 7532 43988 7588
rect 45052 8316 45108 8372
rect 44044 7474 44100 7476
rect 44044 7422 44046 7474
rect 44046 7422 44098 7474
rect 44098 7422 44100 7474
rect 44044 7420 44100 7422
rect 43260 6860 43316 6916
rect 45836 9938 45892 9940
rect 45836 9886 45838 9938
rect 45838 9886 45890 9938
rect 45890 9886 45892 9938
rect 45836 9884 45892 9886
rect 45724 8876 45780 8932
rect 43596 6748 43652 6804
rect 44380 7420 44436 7476
rect 43372 6412 43428 6468
rect 43820 6690 43876 6692
rect 43820 6638 43822 6690
rect 43822 6638 43874 6690
rect 43874 6638 43876 6690
rect 43820 6636 43876 6638
rect 43708 5964 43764 6020
rect 40124 4956 40180 5012
rect 39228 4338 39284 4340
rect 39228 4286 39230 4338
rect 39230 4286 39282 4338
rect 39282 4286 39284 4338
rect 39228 4284 39284 4286
rect 40012 4284 40068 4340
rect 42924 4898 42980 4900
rect 42924 4846 42926 4898
rect 42926 4846 42978 4898
rect 42978 4846 42980 4898
rect 42924 4844 42980 4846
rect 40796 4284 40852 4340
rect 44268 6578 44324 6580
rect 44268 6526 44270 6578
rect 44270 6526 44322 6578
rect 44322 6526 44324 6578
rect 44268 6524 44324 6526
rect 44156 6412 44212 6468
rect 44044 5068 44100 5124
rect 44828 6860 44884 6916
rect 44492 6636 44548 6692
rect 46620 9548 46676 9604
rect 47628 9436 47684 9492
rect 48188 9436 48244 9492
rect 46060 8370 46116 8372
rect 46060 8318 46062 8370
rect 46062 8318 46114 8370
rect 46114 8318 46116 8370
rect 46060 8316 46116 8318
rect 46956 6578 47012 6580
rect 46956 6526 46958 6578
rect 46958 6526 47010 6578
rect 47010 6526 47012 6578
rect 46956 6524 47012 6526
rect 47068 5068 47124 5124
rect 46284 4844 46340 4900
rect 45948 4284 46004 4340
rect 47628 4338 47684 4340
rect 47628 4286 47630 4338
rect 47630 4286 47682 4338
rect 47682 4286 47684 4338
rect 47628 4284 47684 4286
rect 48300 3666 48356 3668
rect 48300 3614 48302 3666
rect 48302 3614 48354 3666
rect 48354 3614 48356 3666
rect 48300 3612 48356 3614
rect 19836 3162 19892 3164
rect 19836 3110 19838 3162
rect 19838 3110 19890 3162
rect 19890 3110 19892 3162
rect 19836 3108 19892 3110
rect 19940 3162 19996 3164
rect 19940 3110 19942 3162
rect 19942 3110 19994 3162
rect 19994 3110 19996 3162
rect 19940 3108 19996 3110
rect 20044 3162 20100 3164
rect 20044 3110 20046 3162
rect 20046 3110 20098 3162
rect 20098 3110 20100 3162
rect 20044 3108 20100 3110
<< metal3 >>
rect 38098 57036 38108 57092
rect 38164 57036 44604 57092
rect 44660 57036 44670 57092
rect 19826 56420 19836 56476
rect 19892 56420 19940 56476
rect 19996 56420 20044 56476
rect 20100 56420 20110 56476
rect 15362 56252 15372 56308
rect 15428 56252 16156 56308
rect 16212 56252 16222 56308
rect 20850 56252 20860 56308
rect 20916 56252 22092 56308
rect 22148 56252 22158 56308
rect 25554 56252 25564 56308
rect 25620 56252 27468 56308
rect 27524 56252 27534 56308
rect 36530 56252 36540 56308
rect 36596 56252 40796 56308
rect 40852 56252 40862 56308
rect 22418 56140 22428 56196
rect 22484 56140 25340 56196
rect 25396 56140 25406 56196
rect 49200 56084 50000 56112
rect 35074 56028 35084 56084
rect 35140 56028 35868 56084
rect 35924 56028 38780 56084
rect 38836 56028 38846 56084
rect 41122 56028 41132 56084
rect 41188 56028 47852 56084
rect 47908 56028 47918 56084
rect 48076 56028 50000 56084
rect 48076 55972 48132 56028
rect 49200 56000 50000 56028
rect 17714 55916 17724 55972
rect 17780 55916 18508 55972
rect 18564 55916 18574 55972
rect 38098 55916 38108 55972
rect 38164 55916 38668 55972
rect 42914 55916 42924 55972
rect 42980 55916 43708 55972
rect 44034 55916 44044 55972
rect 44100 55916 48132 55972
rect 38612 55748 38668 55916
rect 43652 55860 43708 55916
rect 43652 55804 47628 55860
rect 47684 55804 47694 55860
rect 38612 55692 39340 55748
rect 39396 55692 39406 55748
rect 4466 55636 4476 55692
rect 4532 55636 4580 55692
rect 4636 55636 4684 55692
rect 4740 55636 4750 55692
rect 35186 55636 35196 55692
rect 35252 55636 35300 55692
rect 35356 55636 35404 55692
rect 35460 55636 35470 55692
rect 32162 55468 32172 55524
rect 32228 55468 33628 55524
rect 33684 55468 33694 55524
rect 35970 55468 35980 55524
rect 36036 55468 37548 55524
rect 37604 55468 37996 55524
rect 38052 55468 38556 55524
rect 38612 55468 38622 55524
rect 43250 55468 43260 55524
rect 43316 55468 43596 55524
rect 43652 55468 43662 55524
rect 25778 55356 25788 55412
rect 25844 55356 27020 55412
rect 27076 55356 27086 55412
rect 31826 55356 31836 55412
rect 31892 55356 34188 55412
rect 34244 55356 34254 55412
rect 41458 55356 41468 55412
rect 41524 55356 43260 55412
rect 43316 55356 43326 55412
rect 43652 55356 45276 55412
rect 45332 55356 45342 55412
rect 43652 55300 43708 55356
rect 27122 55244 27132 55300
rect 27188 55244 43708 55300
rect 10882 55132 10892 55188
rect 10948 55132 13468 55188
rect 13524 55132 13534 55188
rect 21858 55132 21868 55188
rect 21924 55132 23772 55188
rect 23828 55132 25452 55188
rect 25508 55132 25518 55188
rect 30706 55132 30716 55188
rect 30772 55132 32508 55188
rect 32564 55132 32574 55188
rect 42354 55132 42364 55188
rect 42420 55132 43036 55188
rect 43092 55132 43102 55188
rect 43698 55132 43708 55188
rect 43764 55132 44940 55188
rect 44996 55132 45006 55188
rect 6850 55020 6860 55076
rect 6916 55020 11564 55076
rect 11620 55020 11630 55076
rect 22194 55020 22204 55076
rect 22260 55020 22540 55076
rect 22596 55020 22606 55076
rect 23650 55020 23660 55076
rect 23716 55020 24332 55076
rect 24388 55020 25788 55076
rect 25844 55020 25854 55076
rect 28242 55020 28252 55076
rect 28308 55020 30156 55076
rect 30212 55020 30222 55076
rect 40450 55020 40460 55076
rect 40516 55020 42588 55076
rect 42644 55020 42654 55076
rect 43586 55020 43596 55076
rect 43652 55020 44828 55076
rect 44884 55020 44894 55076
rect 11442 54908 11452 54964
rect 11508 54908 12236 54964
rect 12292 54908 12302 54964
rect 19826 54852 19836 54908
rect 19892 54852 19940 54908
rect 19996 54852 20044 54908
rect 20100 54852 20110 54908
rect 9314 54796 9324 54852
rect 9380 54796 10332 54852
rect 10388 54796 10398 54852
rect 42354 54796 42364 54852
rect 42420 54796 43372 54852
rect 43428 54796 43438 54852
rect 44258 54796 44268 54852
rect 44324 54796 45500 54852
rect 45556 54796 45566 54852
rect 27458 54684 27468 54740
rect 27524 54684 27916 54740
rect 27972 54684 27982 54740
rect 38434 54684 38444 54740
rect 38500 54684 38892 54740
rect 38948 54684 40068 54740
rect 43474 54684 43484 54740
rect 43540 54684 45724 54740
rect 45780 54684 45790 54740
rect 34962 54572 34972 54628
rect 35028 54572 37100 54628
rect 37156 54572 37166 54628
rect 37762 54572 37772 54628
rect 37828 54572 39452 54628
rect 39508 54572 39518 54628
rect 40012 54516 40068 54684
rect 41010 54572 41020 54628
rect 41076 54572 42812 54628
rect 42868 54572 42878 54628
rect 18050 54460 18060 54516
rect 18116 54460 19068 54516
rect 19124 54460 19134 54516
rect 23426 54460 23436 54516
rect 23492 54460 23884 54516
rect 23940 54460 23950 54516
rect 27122 54460 27132 54516
rect 27188 54460 27468 54516
rect 27524 54460 28028 54516
rect 28084 54460 28094 54516
rect 35830 54460 35868 54516
rect 35924 54460 35934 54516
rect 37874 54460 37884 54516
rect 37940 54460 39676 54516
rect 39732 54460 39742 54516
rect 40002 54460 40012 54516
rect 40068 54460 42476 54516
rect 42532 54460 44716 54516
rect 44772 54460 44782 54516
rect 13794 54348 13804 54404
rect 13860 54348 14588 54404
rect 14644 54348 16492 54404
rect 16548 54348 16940 54404
rect 16996 54348 17724 54404
rect 17780 54348 18284 54404
rect 18340 54348 18350 54404
rect 18722 54348 18732 54404
rect 18788 54348 21868 54404
rect 21924 54348 21934 54404
rect 30034 54348 30044 54404
rect 30100 54348 30940 54404
rect 30996 54348 31388 54404
rect 31444 54348 33292 54404
rect 33348 54348 33358 54404
rect 36530 54348 36540 54404
rect 36596 54348 38332 54404
rect 38388 54348 39228 54404
rect 39284 54348 39294 54404
rect 41458 54348 41468 54404
rect 41524 54348 42252 54404
rect 42308 54348 42318 54404
rect 10994 54236 11004 54292
rect 11060 54236 12460 54292
rect 12516 54236 12526 54292
rect 23314 54236 23324 54292
rect 23380 54236 24108 54292
rect 24164 54236 24174 54292
rect 4466 54068 4476 54124
rect 4532 54068 4580 54124
rect 4636 54068 4684 54124
rect 4740 54068 4750 54124
rect 35186 54068 35196 54124
rect 35252 54068 35300 54124
rect 35356 54068 35404 54124
rect 35460 54068 35470 54124
rect 22166 54012 22204 54068
rect 22260 54012 22270 54068
rect 27234 54012 27244 54068
rect 27300 54012 27310 54068
rect 44818 54012 44828 54068
rect 44884 54012 46508 54068
rect 46564 54012 46574 54068
rect 19842 53900 19852 53956
rect 19908 53900 22988 53956
rect 23044 53900 23054 53956
rect 12796 53788 13132 53844
rect 13188 53788 13692 53844
rect 13748 53788 13758 53844
rect 23090 53788 23100 53844
rect 23156 53788 24220 53844
rect 24276 53788 24286 53844
rect 12796 53732 12852 53788
rect 27244 53732 27300 54012
rect 31826 53900 31836 53956
rect 31892 53900 33740 53956
rect 33796 53900 33806 53956
rect 32498 53788 32508 53844
rect 32564 53788 33516 53844
rect 33572 53788 33582 53844
rect 37426 53788 37436 53844
rect 37492 53788 37996 53844
rect 38052 53788 38062 53844
rect 38630 53788 38668 53844
rect 38724 53788 38734 53844
rect 42802 53788 42812 53844
rect 42868 53788 45052 53844
rect 45108 53788 45276 53844
rect 45332 53788 45342 53844
rect 11218 53676 11228 53732
rect 11284 53676 12852 53732
rect 18274 53676 18284 53732
rect 18340 53676 18956 53732
rect 19012 53676 19022 53732
rect 24770 53676 24780 53732
rect 24836 53676 25340 53732
rect 25396 53676 26124 53732
rect 26180 53676 27300 53732
rect 27794 53676 27804 53732
rect 27860 53676 29148 53732
rect 29204 53676 29214 53732
rect 32946 53676 32956 53732
rect 33012 53676 38444 53732
rect 38500 53676 39116 53732
rect 39172 53676 40124 53732
rect 40180 53676 44268 53732
rect 44324 53676 44940 53732
rect 44996 53676 45006 53732
rect 10098 53564 10108 53620
rect 10164 53564 11116 53620
rect 11172 53564 11182 53620
rect 12450 53564 12460 53620
rect 12516 53564 14140 53620
rect 14196 53564 14924 53620
rect 14980 53564 14990 53620
rect 21634 53564 21644 53620
rect 21700 53564 22092 53620
rect 22148 53564 22158 53620
rect 27122 53564 27132 53620
rect 27188 53564 27692 53620
rect 27748 53564 27758 53620
rect 28578 53564 28588 53620
rect 28644 53564 30828 53620
rect 30884 53564 30894 53620
rect 37660 53564 40236 53620
rect 40292 53564 41692 53620
rect 41748 53564 41758 53620
rect 37660 53508 37716 53564
rect 12786 53452 12796 53508
rect 12852 53452 13580 53508
rect 13636 53452 13646 53508
rect 14354 53452 14364 53508
rect 14420 53452 15596 53508
rect 15652 53452 20972 53508
rect 21028 53452 21038 53508
rect 23090 53452 23100 53508
rect 23156 53452 24220 53508
rect 24276 53452 24286 53508
rect 24994 53452 25004 53508
rect 25060 53452 25900 53508
rect 25956 53452 25966 53508
rect 27010 53452 27020 53508
rect 27076 53452 29596 53508
rect 29652 53452 30268 53508
rect 30324 53452 30334 53508
rect 31266 53452 31276 53508
rect 31332 53452 32060 53508
rect 32116 53452 32956 53508
rect 33012 53452 33022 53508
rect 33394 53452 33404 53508
rect 33460 53452 34636 53508
rect 34692 53452 34702 53508
rect 37090 53452 37100 53508
rect 37156 53452 37716 53508
rect 41458 53452 41468 53508
rect 41524 53452 42700 53508
rect 42756 53452 42766 53508
rect 44034 53452 44044 53508
rect 44100 53452 48076 53508
rect 48132 53452 48142 53508
rect 12226 53340 12236 53396
rect 12292 53340 13916 53396
rect 13972 53340 15036 53396
rect 15092 53340 15102 53396
rect 40898 53340 40908 53396
rect 40964 53340 44156 53396
rect 44212 53340 44222 53396
rect 19826 53284 19836 53340
rect 19892 53284 19940 53340
rect 19996 53284 20044 53340
rect 20100 53284 20110 53340
rect 27346 53228 27356 53284
rect 27412 53228 28476 53284
rect 28532 53228 29260 53284
rect 29316 53228 29326 53284
rect 31714 53228 31724 53284
rect 31780 53228 37324 53284
rect 37380 53228 39452 53284
rect 39508 53228 39518 53284
rect 43138 53228 43148 53284
rect 43204 53228 44828 53284
rect 44884 53228 44894 53284
rect 19282 53116 19292 53172
rect 19348 53116 20524 53172
rect 20580 53116 20590 53172
rect 24210 53116 24220 53172
rect 24276 53116 25228 53172
rect 25284 53116 25788 53172
rect 25844 53116 25854 53172
rect 35074 53116 35084 53172
rect 35140 53116 37492 53172
rect 39778 53116 39788 53172
rect 39844 53116 41916 53172
rect 41972 53116 41982 53172
rect 33058 53004 33068 53060
rect 33124 53004 34300 53060
rect 34356 53004 37212 53060
rect 37268 53004 37278 53060
rect 37436 52948 37492 53116
rect 43810 53004 43820 53060
rect 43876 53004 44380 53060
rect 44436 53004 44446 53060
rect 4162 52892 4172 52948
rect 4228 52892 6188 52948
rect 6244 52892 7980 52948
rect 8036 52892 8988 52948
rect 9044 52892 11228 52948
rect 11284 52892 11294 52948
rect 15698 52892 15708 52948
rect 15764 52892 16492 52948
rect 16548 52892 16558 52948
rect 21746 52892 21756 52948
rect 21812 52892 22428 52948
rect 22484 52892 22494 52948
rect 24098 52892 24108 52948
rect 24164 52892 25340 52948
rect 25396 52892 25406 52948
rect 34962 52892 34972 52948
rect 35028 52892 36204 52948
rect 36260 52892 36270 52948
rect 37314 52892 37324 52948
rect 37380 52892 37492 52948
rect 37650 52892 37660 52948
rect 37716 52892 38332 52948
rect 38388 52892 38398 52948
rect 13794 52780 13804 52836
rect 13860 52780 14588 52836
rect 14644 52780 14654 52836
rect 29698 52780 29708 52836
rect 29764 52780 30828 52836
rect 30884 52780 31388 52836
rect 31444 52780 31454 52836
rect 35074 52780 35084 52836
rect 35140 52780 35868 52836
rect 35924 52780 37100 52836
rect 37156 52780 37166 52836
rect 43586 52780 43596 52836
rect 43652 52780 47516 52836
rect 47572 52780 47582 52836
rect 6962 52668 6972 52724
rect 7028 52668 8092 52724
rect 8148 52668 8158 52724
rect 34290 52668 34300 52724
rect 34356 52668 35196 52724
rect 35252 52668 35262 52724
rect 4844 52556 16828 52612
rect 16884 52556 17500 52612
rect 17556 52556 21644 52612
rect 21700 52556 21710 52612
rect 38994 52556 39004 52612
rect 39060 52556 47740 52612
rect 47796 52556 47964 52612
rect 48020 52556 48030 52612
rect 4466 52500 4476 52556
rect 4532 52500 4580 52556
rect 4636 52500 4684 52556
rect 4740 52500 4750 52556
rect 4844 52388 4900 52556
rect 35186 52500 35196 52556
rect 35252 52500 35300 52556
rect 35356 52500 35404 52556
rect 35460 52500 35470 52556
rect 15362 52444 15372 52500
rect 15428 52444 16044 52500
rect 16100 52444 16110 52500
rect 15372 52388 15428 52444
rect 1586 52332 1596 52388
rect 1652 52332 4900 52388
rect 7634 52332 7644 52388
rect 7700 52332 15428 52388
rect 25778 52332 25788 52388
rect 25844 52332 26348 52388
rect 26404 52332 26908 52388
rect 26964 52332 26974 52388
rect 4834 52220 4844 52276
rect 4900 52220 6076 52276
rect 6132 52220 6142 52276
rect 10434 52220 10444 52276
rect 10500 52220 11116 52276
rect 11172 52220 13580 52276
rect 13636 52220 13646 52276
rect 34710 52220 34748 52276
rect 34804 52220 34814 52276
rect 35522 52220 35532 52276
rect 35588 52220 36204 52276
rect 36260 52220 38220 52276
rect 38276 52220 38286 52276
rect 41682 52220 41692 52276
rect 41748 52220 42364 52276
rect 42420 52220 42430 52276
rect 44146 52220 44156 52276
rect 44212 52220 45164 52276
rect 45220 52220 45230 52276
rect 6860 52108 10332 52164
rect 10388 52108 10398 52164
rect 16594 52108 16604 52164
rect 16660 52108 17612 52164
rect 17668 52108 17678 52164
rect 22642 52108 22652 52164
rect 22708 52108 23548 52164
rect 23604 52108 23614 52164
rect 24210 52108 24220 52164
rect 24276 52108 29260 52164
rect 29316 52108 29326 52164
rect 30146 52108 30156 52164
rect 30212 52108 34300 52164
rect 34356 52108 34366 52164
rect 35970 52108 35980 52164
rect 36036 52108 37436 52164
rect 37492 52108 37502 52164
rect 38098 52108 38108 52164
rect 38164 52108 39116 52164
rect 39172 52108 39182 52164
rect 44818 52108 44828 52164
rect 44884 52108 45612 52164
rect 45668 52108 45678 52164
rect 6860 51940 6916 52108
rect 29586 51996 29596 52052
rect 29652 51996 30604 52052
rect 30660 51996 30670 52052
rect 30818 51996 30828 52052
rect 30884 51996 31612 52052
rect 31668 51996 31678 52052
rect 33618 51996 33628 52052
rect 33684 51996 36372 52052
rect 38546 51996 38556 52052
rect 38612 51996 38668 52052
rect 38724 51996 38734 52052
rect 43474 51996 43484 52052
rect 43540 51996 44604 52052
rect 44660 51996 44670 52052
rect 36316 51940 36372 51996
rect 6850 51884 6860 51940
rect 6916 51884 6926 51940
rect 7522 51884 7532 51940
rect 7588 51884 8092 51940
rect 8148 51884 8158 51940
rect 14354 51884 14364 51940
rect 14420 51884 15148 51940
rect 15204 51884 15214 51940
rect 19730 51884 19740 51940
rect 19796 51884 20412 51940
rect 20468 51884 21308 51940
rect 21364 51884 21374 51940
rect 21634 51884 21644 51940
rect 21700 51884 22092 51940
rect 22148 51884 22158 51940
rect 22866 51884 22876 51940
rect 22932 51884 23324 51940
rect 23380 51884 23390 51940
rect 35410 51884 35420 51940
rect 35476 51884 36092 51940
rect 36148 51884 36158 51940
rect 36316 51884 42924 51940
rect 42980 51884 44268 51940
rect 44324 51884 44334 51940
rect 14130 51772 14140 51828
rect 14196 51772 15372 51828
rect 15428 51772 16156 51828
rect 16212 51772 16222 51828
rect 19826 51716 19836 51772
rect 19892 51716 19940 51772
rect 19996 51716 20044 51772
rect 20100 51716 20110 51772
rect 39330 51660 39340 51716
rect 39396 51660 40460 51716
rect 40516 51660 41468 51716
rect 41524 51660 41534 51716
rect 5730 51548 5740 51604
rect 5796 51548 6188 51604
rect 6244 51548 6254 51604
rect 13570 51548 13580 51604
rect 13636 51548 21140 51604
rect 21298 51548 21308 51604
rect 21364 51548 21980 51604
rect 22036 51548 22046 51604
rect 26786 51548 26796 51604
rect 26852 51548 28028 51604
rect 28084 51548 28094 51604
rect 35522 51548 35532 51604
rect 35588 51548 35868 51604
rect 35924 51548 37660 51604
rect 37716 51548 37726 51604
rect 39218 51548 39228 51604
rect 39284 51548 41356 51604
rect 41412 51548 41422 51604
rect 10994 51436 11004 51492
rect 11060 51436 12124 51492
rect 12180 51436 12190 51492
rect 20066 51436 20076 51492
rect 20132 51436 20860 51492
rect 20916 51436 20926 51492
rect 21084 51380 21140 51548
rect 27010 51436 27020 51492
rect 27076 51436 28140 51492
rect 28196 51436 28206 51492
rect 36978 51436 36988 51492
rect 37044 51436 38108 51492
rect 38164 51436 38174 51492
rect 41234 51436 41244 51492
rect 41300 51436 42028 51492
rect 42084 51436 42094 51492
rect 44034 51436 44044 51492
rect 44100 51436 47404 51492
rect 47460 51436 47470 51492
rect 5506 51324 5516 51380
rect 5572 51324 5964 51380
rect 6020 51324 6412 51380
rect 6468 51324 6478 51380
rect 8306 51324 8316 51380
rect 8372 51324 9324 51380
rect 9380 51324 10332 51380
rect 10388 51324 10398 51380
rect 12898 51324 12908 51380
rect 12964 51324 21028 51380
rect 21084 51324 28308 51380
rect 30258 51324 30268 51380
rect 30324 51324 32508 51380
rect 32564 51324 32574 51380
rect 39778 51324 39788 51380
rect 39844 51324 40796 51380
rect 40852 51324 40862 51380
rect 20972 51268 21028 51324
rect 3714 51212 3724 51268
rect 3780 51212 4844 51268
rect 4900 51212 4910 51268
rect 8978 51212 8988 51268
rect 9044 51212 9772 51268
rect 9828 51212 9838 51268
rect 18722 51212 18732 51268
rect 18788 51212 20636 51268
rect 20692 51212 20702 51268
rect 20972 51212 22540 51268
rect 22596 51212 22606 51268
rect 22754 51212 22764 51268
rect 22820 51212 28028 51268
rect 28084 51212 28094 51268
rect 28252 51156 28308 51324
rect 38770 51212 38780 51268
rect 38836 51212 39676 51268
rect 39732 51212 39742 51268
rect 42354 51212 42364 51268
rect 42420 51212 43932 51268
rect 43988 51212 45276 51268
rect 45332 51212 45342 51268
rect 21410 51100 21420 51156
rect 21476 51100 21868 51156
rect 21924 51100 23660 51156
rect 23716 51100 23726 51156
rect 25666 51100 25676 51156
rect 25732 51100 26908 51156
rect 28252 51100 31388 51156
rect 31444 51100 31454 51156
rect 26852 51044 26908 51100
rect 19170 50988 19180 51044
rect 19236 50988 20300 51044
rect 20356 50988 22204 51044
rect 22260 50988 22270 51044
rect 26852 50988 31276 51044
rect 31332 50988 32732 51044
rect 32788 50988 32798 51044
rect 4466 50932 4476 50988
rect 4532 50932 4580 50988
rect 4636 50932 4684 50988
rect 4740 50932 4750 50988
rect 35186 50932 35196 50988
rect 35252 50932 35300 50988
rect 35356 50932 35404 50988
rect 35460 50932 35470 50988
rect 21970 50876 21980 50932
rect 22036 50876 23324 50932
rect 23380 50876 23390 50932
rect 26852 50876 30828 50932
rect 30884 50876 32620 50932
rect 32676 50876 33180 50932
rect 33236 50876 33246 50932
rect 21186 50764 21196 50820
rect 21252 50764 22092 50820
rect 22148 50764 22158 50820
rect 26852 50708 26908 50876
rect 29586 50764 29596 50820
rect 29652 50764 31164 50820
rect 31220 50764 31230 50820
rect 37090 50764 37100 50820
rect 37156 50764 39228 50820
rect 39284 50764 39294 50820
rect 14914 50652 14924 50708
rect 14980 50652 15876 50708
rect 16034 50652 16044 50708
rect 16100 50652 26908 50708
rect 28018 50652 28028 50708
rect 28084 50652 28700 50708
rect 28756 50652 28766 50708
rect 30146 50652 30156 50708
rect 30212 50652 33964 50708
rect 34020 50652 34030 50708
rect 35746 50652 35756 50708
rect 35812 50652 36876 50708
rect 36932 50652 37548 50708
rect 37604 50652 37614 50708
rect 38612 50652 39844 50708
rect 42018 50652 42028 50708
rect 42084 50652 43708 50708
rect 15820 50596 15876 50652
rect 38612 50596 38668 50652
rect 8866 50540 8876 50596
rect 8932 50540 9884 50596
rect 9940 50540 11116 50596
rect 11172 50540 11182 50596
rect 14354 50540 14364 50596
rect 14420 50540 15372 50596
rect 15428 50540 15438 50596
rect 15820 50540 23100 50596
rect 23156 50540 23166 50596
rect 23762 50540 23772 50596
rect 23828 50540 28252 50596
rect 28308 50540 28924 50596
rect 28980 50540 28990 50596
rect 29586 50540 29596 50596
rect 29652 50540 30268 50596
rect 30324 50540 30334 50596
rect 32498 50540 32508 50596
rect 32564 50540 33516 50596
rect 33572 50540 33582 50596
rect 33842 50540 33852 50596
rect 33908 50540 38668 50596
rect 23100 50484 23156 50540
rect 39788 50484 39844 50652
rect 43652 50484 43708 50652
rect 1810 50428 1820 50484
rect 1876 50428 4172 50484
rect 4228 50428 4844 50484
rect 4900 50428 6076 50484
rect 6132 50428 6142 50484
rect 23100 50428 23884 50484
rect 23940 50428 23950 50484
rect 26226 50428 26236 50484
rect 26292 50428 26796 50484
rect 26852 50428 26862 50484
rect 28466 50428 28476 50484
rect 28532 50428 29484 50484
rect 29540 50428 29550 50484
rect 29922 50428 29932 50484
rect 29988 50428 30380 50484
rect 30436 50428 31052 50484
rect 31108 50428 31118 50484
rect 34402 50428 34412 50484
rect 34468 50428 34478 50484
rect 36306 50428 36316 50484
rect 36372 50428 36988 50484
rect 37044 50428 37054 50484
rect 39788 50428 40460 50484
rect 40516 50428 40526 50484
rect 41804 50428 43036 50484
rect 43092 50428 43102 50484
rect 43652 50428 44604 50484
rect 44660 50428 45052 50484
rect 45108 50428 45118 50484
rect 46834 50428 46844 50484
rect 46900 50428 47852 50484
rect 47908 50428 47918 50484
rect 34412 50372 34468 50428
rect 6738 50316 6748 50372
rect 6804 50316 7980 50372
rect 8036 50316 10892 50372
rect 10948 50316 11564 50372
rect 11620 50316 11630 50372
rect 18722 50316 18732 50372
rect 18788 50316 20524 50372
rect 20580 50316 20590 50372
rect 34412 50316 35084 50372
rect 35140 50316 35150 50372
rect 40114 50316 40124 50372
rect 40180 50316 41580 50372
rect 41636 50316 41646 50372
rect 41804 50260 41860 50428
rect 49200 50260 50000 50288
rect 34290 50204 34300 50260
rect 34356 50204 34636 50260
rect 34692 50204 34972 50260
rect 35028 50204 35038 50260
rect 35970 50204 35980 50260
rect 36036 50204 36764 50260
rect 36820 50204 38108 50260
rect 38164 50204 38174 50260
rect 41458 50204 41468 50260
rect 41524 50204 41860 50260
rect 42140 50204 43708 50260
rect 43764 50204 43774 50260
rect 48290 50204 48300 50260
rect 48356 50204 50000 50260
rect 19826 50148 19836 50204
rect 19892 50148 19940 50204
rect 19996 50148 20044 50204
rect 20100 50148 20110 50204
rect 11778 50092 11788 50148
rect 11844 50092 13804 50148
rect 13860 50092 13870 50148
rect 2146 49980 2156 50036
rect 2212 49980 13020 50036
rect 13076 49980 13086 50036
rect 13906 49980 13916 50036
rect 13972 49980 15036 50036
rect 15092 49980 15102 50036
rect 35858 49980 35868 50036
rect 35924 49980 36652 50036
rect 36708 49980 36718 50036
rect 42140 49924 42196 50204
rect 49200 50176 50000 50204
rect 43652 50092 44716 50148
rect 44772 50092 44782 50148
rect 43652 50036 43708 50092
rect 42364 49980 43708 50036
rect 23762 49868 23772 49924
rect 23828 49868 23996 49924
rect 24052 49868 24220 49924
rect 24276 49868 24286 49924
rect 33506 49868 33516 49924
rect 33572 49868 42140 49924
rect 42196 49868 42206 49924
rect 0 49812 800 49840
rect 42364 49812 42420 49980
rect 42914 49868 42924 49924
rect 42980 49868 46396 49924
rect 46452 49868 46462 49924
rect 0 49756 1708 49812
rect 1764 49756 1774 49812
rect 26450 49756 26460 49812
rect 26516 49756 27580 49812
rect 27636 49756 27646 49812
rect 28690 49756 28700 49812
rect 28756 49756 29372 49812
rect 29428 49756 29438 49812
rect 35522 49756 35532 49812
rect 35588 49756 36316 49812
rect 36372 49756 36382 49812
rect 38994 49756 39004 49812
rect 39060 49756 42420 49812
rect 44482 49756 44492 49812
rect 44548 49756 46732 49812
rect 46788 49756 46798 49812
rect 0 49728 800 49756
rect 4610 49644 4620 49700
rect 4676 49644 4956 49700
rect 5012 49644 5628 49700
rect 5684 49644 5694 49700
rect 23426 49644 23436 49700
rect 23492 49644 25676 49700
rect 25732 49644 25742 49700
rect 35970 49644 35980 49700
rect 36036 49644 38220 49700
rect 38276 49644 38286 49700
rect 45042 49644 45052 49700
rect 45108 49644 46284 49700
rect 46340 49644 46350 49700
rect 13570 49532 13580 49588
rect 13636 49532 14252 49588
rect 14308 49532 14318 49588
rect 25890 49532 25900 49588
rect 25956 49532 27916 49588
rect 27972 49532 27982 49588
rect 37090 49532 37100 49588
rect 37156 49532 38668 49588
rect 38724 49532 39116 49588
rect 39172 49532 41244 49588
rect 41300 49532 44380 49588
rect 44436 49532 44446 49588
rect 37426 49420 37436 49476
rect 37492 49420 39452 49476
rect 39508 49420 39518 49476
rect 4466 49364 4476 49420
rect 4532 49364 4580 49420
rect 4636 49364 4684 49420
rect 4740 49364 4750 49420
rect 35186 49364 35196 49420
rect 35252 49364 35300 49420
rect 35356 49364 35404 49420
rect 35460 49364 35470 49420
rect 2482 49196 2492 49252
rect 2548 49196 3388 49252
rect 35410 49196 35420 49252
rect 35476 49196 35980 49252
rect 36036 49196 36046 49252
rect 45378 49196 45388 49252
rect 45444 49196 47404 49252
rect 47460 49196 47470 49252
rect 3332 49140 3388 49196
rect 3332 49084 7420 49140
rect 7476 49084 7486 49140
rect 15092 49084 25340 49140
rect 25396 49084 27356 49140
rect 27412 49084 29708 49140
rect 29764 49084 29774 49140
rect 32834 49084 32844 49140
rect 32900 49084 33740 49140
rect 33796 49084 36988 49140
rect 37044 49084 37054 49140
rect 37762 49084 37772 49140
rect 37828 49084 39004 49140
rect 39060 49084 39070 49140
rect 40226 49084 40236 49140
rect 40292 49084 41356 49140
rect 41412 49084 42028 49140
rect 42084 49084 42094 49140
rect 4722 48972 4732 49028
rect 4788 48972 5516 49028
rect 5572 48972 5582 49028
rect 5058 48860 5068 48916
rect 5124 48860 5740 48916
rect 5796 48860 9996 48916
rect 10052 48860 10062 48916
rect 11106 48860 11116 48916
rect 11172 48860 11564 48916
rect 11620 48860 12236 48916
rect 12292 48860 13244 48916
rect 13300 48860 13310 48916
rect 1474 48748 1484 48804
rect 1540 48748 2268 48804
rect 2324 48748 2334 48804
rect 9874 48748 9884 48804
rect 9940 48748 10444 48804
rect 10500 48748 10510 48804
rect 11666 48748 11676 48804
rect 11732 48748 13020 48804
rect 13076 48748 13086 48804
rect 15092 48692 15148 49084
rect 40236 49028 40292 49084
rect 17490 48972 17500 49028
rect 17556 48972 18732 49028
rect 18788 48972 18798 49028
rect 25554 48972 25564 49028
rect 25620 48972 26460 49028
rect 26516 48972 26526 49028
rect 28018 48972 28028 49028
rect 28084 48972 28588 49028
rect 28644 48972 29260 49028
rect 29316 48972 31500 49028
rect 31556 48972 31566 49028
rect 34178 48972 34188 49028
rect 34244 48972 36764 49028
rect 36820 48972 36830 49028
rect 38322 48972 38332 49028
rect 38388 48972 40292 49028
rect 46386 48972 46396 49028
rect 46452 48972 47628 49028
rect 47684 48972 47694 49028
rect 16706 48860 16716 48916
rect 16772 48860 18060 48916
rect 18116 48860 18126 48916
rect 20290 48860 20300 48916
rect 20356 48860 22820 48916
rect 36082 48860 36092 48916
rect 36148 48860 37100 48916
rect 37156 48860 37166 48916
rect 22764 48804 22820 48860
rect 15698 48748 15708 48804
rect 15764 48748 18284 48804
rect 18340 48748 18350 48804
rect 19730 48748 19740 48804
rect 19796 48748 20412 48804
rect 20468 48748 20478 48804
rect 22754 48748 22764 48804
rect 22820 48748 24332 48804
rect 24388 48748 26460 48804
rect 26516 48748 26526 48804
rect 33394 48748 33404 48804
rect 33460 48748 37212 48804
rect 37268 48748 40572 48804
rect 40628 48748 41916 48804
rect 41972 48748 41982 48804
rect 45826 48748 45836 48804
rect 45892 48748 46004 48804
rect 47394 48748 47404 48804
rect 47460 48748 48188 48804
rect 48244 48748 48254 48804
rect 45948 48692 46004 48748
rect 5058 48636 5068 48692
rect 5124 48636 5852 48692
rect 5908 48636 8428 48692
rect 8484 48636 8494 48692
rect 12786 48636 12796 48692
rect 12852 48636 15148 48692
rect 42466 48636 42476 48692
rect 42532 48636 44268 48692
rect 44324 48636 44334 48692
rect 44930 48636 44940 48692
rect 44996 48636 48076 48692
rect 48132 48636 48142 48692
rect 19826 48580 19836 48636
rect 19892 48580 19940 48636
rect 19996 48580 20044 48636
rect 20100 48580 20110 48636
rect 44268 48580 44324 48636
rect 44268 48524 45948 48580
rect 46004 48524 46014 48580
rect 15698 48412 15708 48468
rect 15764 48412 16380 48468
rect 16436 48412 16828 48468
rect 16884 48412 22092 48468
rect 22148 48412 22158 48468
rect 43362 48412 43372 48468
rect 43428 48412 44044 48468
rect 44100 48412 44110 48468
rect 8642 48300 8652 48356
rect 8708 48300 9100 48356
rect 9156 48300 9660 48356
rect 9716 48300 9726 48356
rect 10658 48300 10668 48356
rect 10724 48300 11228 48356
rect 11284 48300 11788 48356
rect 11844 48300 12908 48356
rect 12964 48300 12974 48356
rect 20290 48300 20300 48356
rect 20356 48300 22204 48356
rect 22260 48300 22270 48356
rect 27906 48300 27916 48356
rect 27972 48300 29484 48356
rect 29540 48300 29550 48356
rect 34738 48300 34748 48356
rect 34804 48300 40012 48356
rect 40068 48300 40078 48356
rect 41682 48300 41692 48356
rect 41748 48300 42364 48356
rect 42420 48300 42430 48356
rect 46610 48300 46620 48356
rect 46676 48300 47404 48356
rect 47460 48300 47470 48356
rect 2370 48188 2380 48244
rect 2436 48188 3164 48244
rect 3220 48188 3948 48244
rect 4004 48188 4014 48244
rect 4162 48188 4172 48244
rect 4228 48188 4844 48244
rect 4900 48188 4910 48244
rect 11890 48188 11900 48244
rect 11956 48188 12684 48244
rect 12740 48188 12750 48244
rect 24434 48188 24444 48244
rect 24500 48188 25564 48244
rect 25620 48188 25630 48244
rect 40338 48188 40348 48244
rect 40404 48188 41468 48244
rect 41524 48188 41534 48244
rect 18610 48076 18620 48132
rect 18676 48076 20636 48132
rect 20692 48076 20702 48132
rect 22418 48076 22428 48132
rect 22484 48076 23324 48132
rect 23380 48076 23390 48132
rect 24658 48076 24668 48132
rect 24724 48076 25340 48132
rect 25396 48076 25406 48132
rect 27010 48076 27020 48132
rect 27076 48076 28364 48132
rect 28420 48076 28430 48132
rect 40450 48076 40460 48132
rect 40516 48076 41244 48132
rect 41300 48076 41310 48132
rect 17602 47964 17612 48020
rect 17668 47964 21084 48020
rect 21140 47964 23996 48020
rect 24052 47964 24556 48020
rect 24612 47964 24622 48020
rect 26786 47964 26796 48020
rect 26852 47964 28700 48020
rect 28756 47964 28766 48020
rect 38882 47964 38892 48020
rect 38948 47964 39564 48020
rect 39620 47964 39630 48020
rect 4466 47796 4476 47852
rect 4532 47796 4580 47852
rect 4636 47796 4684 47852
rect 4740 47796 4750 47852
rect 35186 47796 35196 47852
rect 35252 47796 35300 47852
rect 35356 47796 35404 47852
rect 35460 47796 35470 47852
rect 11666 47740 11676 47796
rect 11732 47740 12124 47796
rect 12180 47740 12190 47796
rect 27122 47740 27132 47796
rect 27188 47740 27804 47796
rect 27860 47740 27870 47796
rect 29474 47628 29484 47684
rect 29540 47628 30268 47684
rect 30324 47628 30334 47684
rect 37538 47628 37548 47684
rect 37604 47628 38444 47684
rect 38500 47628 38510 47684
rect 1810 47516 1820 47572
rect 1876 47516 5068 47572
rect 5124 47516 5134 47572
rect 8530 47516 8540 47572
rect 8596 47516 9548 47572
rect 9604 47516 9614 47572
rect 16034 47516 16044 47572
rect 16100 47516 17388 47572
rect 17444 47516 17454 47572
rect 23986 47516 23996 47572
rect 24052 47516 27916 47572
rect 27972 47516 27982 47572
rect 39778 47516 39788 47572
rect 39844 47516 41020 47572
rect 41076 47516 41086 47572
rect 46834 47516 46844 47572
rect 46900 47516 47964 47572
rect 48020 47516 48030 47572
rect 3266 47404 3276 47460
rect 3332 47404 4172 47460
rect 4228 47404 4620 47460
rect 4676 47404 4686 47460
rect 7074 47404 7084 47460
rect 7140 47404 7532 47460
rect 7588 47404 8876 47460
rect 8932 47404 8942 47460
rect 11554 47404 11564 47460
rect 11620 47404 12124 47460
rect 12180 47404 12190 47460
rect 20066 47404 20076 47460
rect 20132 47404 20860 47460
rect 20916 47404 20926 47460
rect 21634 47404 21644 47460
rect 21700 47404 23548 47460
rect 23604 47404 23614 47460
rect 24098 47404 24108 47460
rect 24164 47404 24668 47460
rect 24724 47404 24734 47460
rect 24994 47404 25004 47460
rect 25060 47404 26908 47460
rect 26964 47404 28028 47460
rect 28084 47404 28094 47460
rect 29362 47404 29372 47460
rect 29428 47404 30716 47460
rect 30772 47404 31500 47460
rect 31556 47404 31566 47460
rect 32162 47404 32172 47460
rect 32228 47404 34972 47460
rect 35028 47404 35532 47460
rect 35588 47404 35598 47460
rect 39554 47404 39564 47460
rect 39620 47404 41692 47460
rect 41748 47404 41758 47460
rect 45042 47404 45052 47460
rect 45108 47404 47404 47460
rect 47460 47404 47470 47460
rect 7298 47292 7308 47348
rect 7364 47292 7644 47348
rect 7700 47292 7710 47348
rect 25330 47292 25340 47348
rect 25396 47292 27916 47348
rect 27972 47292 27982 47348
rect 33730 47292 33740 47348
rect 33796 47292 35756 47348
rect 35812 47292 35822 47348
rect 36418 47292 36428 47348
rect 36484 47292 37212 47348
rect 37268 47292 37278 47348
rect 41458 47292 41468 47348
rect 41524 47292 42588 47348
rect 42644 47292 42654 47348
rect 44818 47292 44828 47348
rect 44884 47292 46620 47348
rect 46676 47292 47628 47348
rect 47684 47292 47694 47348
rect 22866 47180 22876 47236
rect 22932 47180 24668 47236
rect 24724 47180 27132 47236
rect 27188 47180 27198 47236
rect 41346 47180 41356 47236
rect 41412 47180 42364 47236
rect 42420 47180 42430 47236
rect 42690 47180 42700 47236
rect 42756 47180 43596 47236
rect 43652 47180 43662 47236
rect 45378 47180 45388 47236
rect 45444 47180 46060 47236
rect 46116 47180 46126 47236
rect 9762 47068 9772 47124
rect 9828 47068 10332 47124
rect 10388 47068 10836 47124
rect 13682 47068 13692 47124
rect 13748 47068 17388 47124
rect 17444 47068 17454 47124
rect 22530 47068 22540 47124
rect 22596 47068 24444 47124
rect 24500 47068 24510 47124
rect 29810 47068 29820 47124
rect 29876 47068 29886 47124
rect 34524 47068 35196 47124
rect 35252 47068 36316 47124
rect 36372 47068 36382 47124
rect 41234 47068 41244 47124
rect 41300 47068 42476 47124
rect 42532 47068 43484 47124
rect 43540 47068 43550 47124
rect 6514 46956 6524 47012
rect 6580 46956 7756 47012
rect 7812 46956 7822 47012
rect 10780 46788 10836 47068
rect 19826 47012 19836 47068
rect 19892 47012 19940 47068
rect 19996 47012 20044 47068
rect 20100 47012 20110 47068
rect 29820 47012 29876 47068
rect 34524 47012 34580 47068
rect 29820 46956 30380 47012
rect 30436 46956 30446 47012
rect 34514 46956 34524 47012
rect 34580 46956 34590 47012
rect 37090 46956 37100 47012
rect 37156 46956 38220 47012
rect 38276 46956 38286 47012
rect 38612 46956 38780 47012
rect 38836 46956 38846 47012
rect 41010 46956 41020 47012
rect 41076 46956 42028 47012
rect 42084 46956 43708 47012
rect 14354 46844 14364 46900
rect 14420 46844 15932 46900
rect 15988 46844 15998 46900
rect 20962 46844 20972 46900
rect 21028 46844 25004 46900
rect 25060 46844 25340 46900
rect 25396 46844 25406 46900
rect 30930 46844 30940 46900
rect 30996 46844 33292 46900
rect 33348 46844 34748 46900
rect 34804 46844 34814 46900
rect 10770 46732 10780 46788
rect 10836 46732 10846 46788
rect 10994 46732 11004 46788
rect 11060 46732 11452 46788
rect 11508 46732 12236 46788
rect 12292 46732 12302 46788
rect 29250 46732 29260 46788
rect 29316 46732 29932 46788
rect 29988 46732 29998 46788
rect 34626 46732 34636 46788
rect 34692 46732 35308 46788
rect 35364 46732 35374 46788
rect 38612 46676 38668 46956
rect 3714 46620 3724 46676
rect 3780 46620 4844 46676
rect 4900 46620 10668 46676
rect 10724 46620 10734 46676
rect 15138 46620 15148 46676
rect 15204 46620 15596 46676
rect 15652 46620 15662 46676
rect 15810 46620 15820 46676
rect 15876 46620 16940 46676
rect 16996 46620 17006 46676
rect 21410 46620 21420 46676
rect 21476 46620 22540 46676
rect 22596 46620 23100 46676
rect 23156 46620 23166 46676
rect 29698 46620 29708 46676
rect 29764 46620 31276 46676
rect 31332 46620 31342 46676
rect 34402 46620 34412 46676
rect 34468 46620 38668 46676
rect 43652 46620 43708 46956
rect 43764 46620 44268 46676
rect 44324 46620 44334 46676
rect 9874 46508 9884 46564
rect 9940 46508 10220 46564
rect 10276 46508 10286 46564
rect 21298 46508 21308 46564
rect 21364 46508 23212 46564
rect 23268 46508 23278 46564
rect 23874 46508 23884 46564
rect 23940 46508 29596 46564
rect 29652 46508 29662 46564
rect 36978 46508 36988 46564
rect 37044 46508 38556 46564
rect 38612 46508 39116 46564
rect 39172 46508 39182 46564
rect 18610 46396 18620 46452
rect 18676 46396 20188 46452
rect 20244 46396 20254 46452
rect 35410 46396 35420 46452
rect 35476 46396 36092 46452
rect 36148 46396 36158 46452
rect 39218 46284 39228 46340
rect 39284 46284 39564 46340
rect 39620 46284 39630 46340
rect 4466 46228 4476 46284
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4740 46228 4750 46284
rect 35186 46228 35196 46284
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35460 46228 35470 46284
rect 34850 46060 34860 46116
rect 34916 46060 35868 46116
rect 35924 46060 37212 46116
rect 37268 46060 37278 46116
rect 15026 45948 15036 46004
rect 15092 45948 21308 46004
rect 21364 45948 21374 46004
rect 34738 45948 34748 46004
rect 34804 45948 35196 46004
rect 35252 45948 36876 46004
rect 36932 45948 36942 46004
rect 42802 45948 42812 46004
rect 42868 45948 44044 46004
rect 44100 45948 44828 46004
rect 44884 45948 44894 46004
rect 10658 45836 10668 45892
rect 10724 45836 11452 45892
rect 11508 45836 12684 45892
rect 12740 45836 13580 45892
rect 13636 45836 13646 45892
rect 15586 45836 15596 45892
rect 15652 45836 16492 45892
rect 16548 45836 16558 45892
rect 19282 45836 19292 45892
rect 19348 45836 20412 45892
rect 20468 45836 20478 45892
rect 22082 45836 22092 45892
rect 22148 45836 22988 45892
rect 23044 45836 23054 45892
rect 36306 45836 36316 45892
rect 36372 45836 36764 45892
rect 36820 45836 40348 45892
rect 40404 45836 40414 45892
rect 42466 45836 42476 45892
rect 42532 45836 43260 45892
rect 43316 45836 43326 45892
rect 43586 45836 43596 45892
rect 43652 45836 45836 45892
rect 45892 45836 45902 45892
rect 3602 45724 3612 45780
rect 3668 45724 4844 45780
rect 4900 45724 4910 45780
rect 6290 45724 6300 45780
rect 6356 45724 7084 45780
rect 7140 45724 7150 45780
rect 12898 45724 12908 45780
rect 12964 45724 13916 45780
rect 13972 45724 13982 45780
rect 18386 45724 18396 45780
rect 18452 45724 20300 45780
rect 20356 45724 20366 45780
rect 21858 45724 21868 45780
rect 21924 45724 23996 45780
rect 24052 45724 24062 45780
rect 43260 45668 43316 45836
rect 5954 45612 5964 45668
rect 6020 45612 6412 45668
rect 6468 45612 6860 45668
rect 6916 45612 6926 45668
rect 20178 45612 20188 45668
rect 20244 45612 22876 45668
rect 22932 45612 22942 45668
rect 24546 45612 24556 45668
rect 24612 45612 25340 45668
rect 25396 45612 25406 45668
rect 43260 45612 44156 45668
rect 44212 45612 44222 45668
rect 22204 45556 22260 45612
rect 21746 45500 21756 45556
rect 21812 45500 21980 45556
rect 22036 45500 22046 45556
rect 22194 45500 22204 45556
rect 22260 45500 22270 45556
rect 24994 45500 25004 45556
rect 25060 45500 25452 45556
rect 25508 45500 25518 45556
rect 28130 45500 28140 45556
rect 28196 45500 30380 45556
rect 30436 45500 30446 45556
rect 45042 45500 45052 45556
rect 45108 45500 47628 45556
rect 47684 45500 47694 45556
rect 19826 45444 19836 45500
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 20100 45444 20110 45500
rect 20402 45388 20412 45444
rect 20468 45388 21196 45444
rect 21252 45388 25788 45444
rect 25844 45388 25854 45444
rect 33852 45388 34300 45444
rect 34356 45388 34366 45444
rect 33852 45332 33908 45388
rect 2818 45276 2828 45332
rect 2884 45276 3836 45332
rect 3892 45276 3902 45332
rect 15138 45276 15148 45332
rect 15204 45276 16268 45332
rect 16324 45276 16716 45332
rect 16772 45276 26124 45332
rect 26180 45276 26190 45332
rect 33730 45276 33740 45332
rect 33796 45276 33964 45332
rect 34020 45276 34030 45332
rect 34402 45276 34412 45332
rect 34468 45276 35756 45332
rect 35812 45276 35822 45332
rect 38658 45276 38668 45332
rect 38724 45276 40236 45332
rect 40292 45276 40908 45332
rect 40964 45276 40974 45332
rect 44930 45276 44940 45332
rect 44996 45276 45388 45332
rect 45444 45276 46172 45332
rect 46228 45276 46238 45332
rect 2370 45164 2380 45220
rect 2436 45164 3724 45220
rect 3780 45164 3790 45220
rect 7074 45164 7084 45220
rect 7140 45164 8316 45220
rect 8372 45164 8382 45220
rect 10070 45164 10108 45220
rect 10164 45164 10174 45220
rect 23426 45164 23436 45220
rect 23492 45164 24332 45220
rect 24388 45164 25004 45220
rect 25060 45164 25070 45220
rect 32386 45164 32396 45220
rect 32452 45164 33404 45220
rect 33460 45164 38332 45220
rect 38388 45164 38556 45220
rect 38612 45164 38622 45220
rect 38770 45164 38780 45220
rect 38836 45164 40012 45220
rect 40068 45164 40078 45220
rect 43362 45164 43372 45220
rect 43428 45164 45612 45220
rect 45668 45164 46284 45220
rect 46340 45164 46350 45220
rect 2594 45052 2604 45108
rect 2660 45052 3276 45108
rect 3332 45052 3836 45108
rect 3892 45052 3902 45108
rect 4834 45052 4844 45108
rect 4900 45052 8988 45108
rect 9044 45052 12908 45108
rect 12964 45052 13580 45108
rect 13636 45052 14476 45108
rect 14532 45052 14542 45108
rect 15362 45052 15372 45108
rect 15428 45052 15932 45108
rect 15988 45052 15998 45108
rect 16818 45052 16828 45108
rect 16884 45052 19180 45108
rect 19236 45052 19246 45108
rect 21074 45052 21084 45108
rect 21140 45052 21756 45108
rect 21812 45052 21822 45108
rect 25442 45052 25452 45108
rect 25508 45052 26012 45108
rect 26068 45052 26078 45108
rect 29586 45052 29596 45108
rect 29652 45052 31948 45108
rect 32004 45052 32014 45108
rect 38098 45052 38108 45108
rect 38164 45052 39116 45108
rect 39172 45052 39182 45108
rect 40338 45052 40348 45108
rect 40404 45052 41580 45108
rect 41636 45052 42812 45108
rect 42868 45052 42878 45108
rect 45154 45052 45164 45108
rect 45220 45052 46508 45108
rect 46564 45052 46574 45108
rect 3042 44940 3052 44996
rect 3108 44940 3500 44996
rect 3556 44940 4172 44996
rect 4228 44940 4238 44996
rect 4386 44940 4396 44996
rect 4452 44940 5740 44996
rect 5796 44940 5806 44996
rect 22530 44940 22540 44996
rect 22596 44940 23548 44996
rect 23604 44940 23614 44996
rect 24658 44940 24668 44996
rect 24724 44940 25004 44996
rect 25060 44940 25070 44996
rect 38210 44940 38220 44996
rect 38276 44940 39564 44996
rect 39620 44940 39630 44996
rect 42354 44940 42364 44996
rect 42420 44940 43596 44996
rect 43652 44940 43662 44996
rect 46172 44940 46732 44996
rect 46788 44940 47516 44996
rect 47572 44940 47582 44996
rect 46172 44884 46228 44940
rect 3266 44828 3276 44884
rect 3332 44828 4060 44884
rect 4116 44828 8764 44884
rect 8820 44828 9772 44884
rect 9828 44828 9838 44884
rect 39218 44828 39228 44884
rect 39284 44828 42028 44884
rect 42084 44828 42094 44884
rect 42690 44828 42700 44884
rect 42756 44828 46228 44884
rect 47170 44828 47180 44884
rect 47236 44828 47740 44884
rect 47796 44828 47806 44884
rect 3378 44716 3388 44772
rect 3444 44716 4284 44772
rect 4340 44716 4350 44772
rect 4466 44660 4476 44716
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4740 44660 4750 44716
rect 35186 44660 35196 44716
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35460 44660 35470 44716
rect 24658 44492 24668 44548
rect 24724 44492 25452 44548
rect 25508 44492 25518 44548
rect 26226 44492 26236 44548
rect 26292 44492 27580 44548
rect 27636 44492 27646 44548
rect 42914 44492 42924 44548
rect 42980 44492 43932 44548
rect 43988 44492 43998 44548
rect 49200 44436 50000 44464
rect 17938 44380 17948 44436
rect 18004 44380 18620 44436
rect 18676 44380 19852 44436
rect 19908 44380 19918 44436
rect 31490 44380 31500 44436
rect 31556 44380 34748 44436
rect 34804 44380 34814 44436
rect 39666 44380 39676 44436
rect 39732 44380 40236 44436
rect 40292 44380 40302 44436
rect 41906 44380 41916 44436
rect 41972 44380 42364 44436
rect 42420 44380 42430 44436
rect 45266 44380 45276 44436
rect 45332 44380 46620 44436
rect 46676 44380 47292 44436
rect 47348 44380 47358 44436
rect 48178 44380 48188 44436
rect 48244 44380 50000 44436
rect 49200 44352 50000 44380
rect 6850 44268 6860 44324
rect 6916 44268 7644 44324
rect 7700 44268 7710 44324
rect 23650 44268 23660 44324
rect 23716 44268 24556 44324
rect 24612 44268 24622 44324
rect 24882 44268 24892 44324
rect 24948 44268 25452 44324
rect 25508 44268 25900 44324
rect 25956 44268 25966 44324
rect 27906 44268 27916 44324
rect 27972 44268 29372 44324
rect 29428 44268 29438 44324
rect 32946 44268 32956 44324
rect 33012 44268 33852 44324
rect 33908 44268 33918 44324
rect 41122 44268 41132 44324
rect 41188 44268 41580 44324
rect 41636 44268 44044 44324
rect 44100 44268 44110 44324
rect 44258 44268 44268 44324
rect 44324 44268 45164 44324
rect 45220 44268 45230 44324
rect 19282 44156 19292 44212
rect 19348 44156 20748 44212
rect 20804 44156 20814 44212
rect 43810 44156 43820 44212
rect 43876 44156 44940 44212
rect 44996 44156 45006 44212
rect 6738 44044 6748 44100
rect 6804 44044 7644 44100
rect 7700 44044 7980 44100
rect 8036 44044 9548 44100
rect 9604 44044 9614 44100
rect 11442 44044 11452 44100
rect 11508 44044 12236 44100
rect 12292 44044 12302 44100
rect 17490 44044 17500 44100
rect 17556 44044 19404 44100
rect 19460 44044 20300 44100
rect 20356 44044 20366 44100
rect 21970 44044 21980 44100
rect 22036 44044 22764 44100
rect 22820 44044 22830 44100
rect 31042 44044 31052 44100
rect 31108 44044 31836 44100
rect 31892 44044 31902 44100
rect 44034 44044 44044 44100
rect 44100 44044 46172 44100
rect 46228 44044 47180 44100
rect 47236 44044 47246 44100
rect 19826 43876 19836 43932
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 20100 43876 20110 43932
rect 26898 43820 26908 43876
rect 26964 43820 30604 43876
rect 30660 43820 30670 43876
rect 40226 43820 40236 43876
rect 40292 43820 40302 43876
rect 43362 43820 43372 43876
rect 43428 43820 44044 43876
rect 44100 43820 44110 43876
rect 40236 43764 40292 43820
rect 18274 43708 18284 43764
rect 18340 43708 20300 43764
rect 20356 43708 20366 43764
rect 29474 43708 29484 43764
rect 29540 43708 30828 43764
rect 30884 43708 30894 43764
rect 37538 43708 37548 43764
rect 37604 43708 41020 43764
rect 41076 43708 41468 43764
rect 41524 43708 41534 43764
rect 4274 43596 4284 43652
rect 4340 43596 5404 43652
rect 5460 43596 5470 43652
rect 9986 43596 9996 43652
rect 10052 43596 11228 43652
rect 11284 43596 11294 43652
rect 12674 43596 12684 43652
rect 12740 43596 15372 43652
rect 15428 43596 16716 43652
rect 16772 43596 16782 43652
rect 20178 43596 20188 43652
rect 20244 43596 21868 43652
rect 21924 43596 21934 43652
rect 23986 43596 23996 43652
rect 24052 43596 24892 43652
rect 24948 43596 24958 43652
rect 26674 43596 26684 43652
rect 26740 43596 27356 43652
rect 27412 43596 27422 43652
rect 36306 43596 36316 43652
rect 36372 43596 36988 43652
rect 37044 43596 37324 43652
rect 37380 43596 37772 43652
rect 37828 43596 37838 43652
rect 8194 43484 8204 43540
rect 8260 43484 8988 43540
rect 9044 43484 9054 43540
rect 9314 43484 9324 43540
rect 9380 43484 10444 43540
rect 10500 43484 10510 43540
rect 15026 43484 15036 43540
rect 15092 43484 15708 43540
rect 15764 43484 15774 43540
rect 16258 43484 16268 43540
rect 16324 43484 16334 43540
rect 26562 43484 26572 43540
rect 26628 43484 28028 43540
rect 28084 43484 28094 43540
rect 36866 43484 36876 43540
rect 36932 43484 38780 43540
rect 38836 43484 38846 43540
rect 38994 43484 39004 43540
rect 39060 43484 42028 43540
rect 42084 43484 42094 43540
rect 43586 43484 43596 43540
rect 43652 43484 45052 43540
rect 45108 43484 45118 43540
rect 16268 43428 16324 43484
rect 39004 43428 39060 43484
rect 3490 43372 3500 43428
rect 3556 43372 4396 43428
rect 4452 43372 5516 43428
rect 5572 43372 5582 43428
rect 14690 43372 14700 43428
rect 14756 43372 16324 43428
rect 38434 43372 38444 43428
rect 38500 43372 39060 43428
rect 13122 43260 13132 43316
rect 13188 43260 27692 43316
rect 27748 43260 27758 43316
rect 30482 43260 30492 43316
rect 30548 43260 33068 43316
rect 33124 43260 33134 43316
rect 38546 43260 38556 43316
rect 38612 43260 40124 43316
rect 40180 43260 40684 43316
rect 40740 43260 40750 43316
rect 5292 43148 14924 43204
rect 14980 43148 16828 43204
rect 16884 43148 16894 43204
rect 26450 43148 26460 43204
rect 26516 43148 29148 43204
rect 29204 43148 29596 43204
rect 29652 43148 29662 43204
rect 4466 43092 4476 43148
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4740 43092 4750 43148
rect 5292 42868 5348 43148
rect 35186 43092 35196 43148
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35460 43092 35470 43148
rect 5506 42924 5516 42980
rect 5572 42924 8540 42980
rect 8596 42924 10332 42980
rect 10388 42924 10398 42980
rect 11116 42924 11676 42980
rect 11732 42924 12236 42980
rect 12292 42924 12302 42980
rect 38770 42924 38780 42980
rect 38836 42924 39228 42980
rect 39284 42924 40236 42980
rect 40292 42924 40302 42980
rect 11116 42868 11172 42924
rect 4162 42812 4172 42868
rect 4228 42812 5348 42868
rect 11106 42812 11116 42868
rect 11172 42812 11182 42868
rect 21746 42812 21756 42868
rect 21812 42812 22652 42868
rect 22708 42812 22718 42868
rect 23986 42812 23996 42868
rect 24052 42812 24556 42868
rect 24612 42812 24622 42868
rect 4834 42700 4844 42756
rect 4900 42700 5180 42756
rect 5236 42700 5246 42756
rect 8642 42700 8652 42756
rect 8708 42700 9324 42756
rect 9380 42700 9884 42756
rect 9940 42700 9950 42756
rect 14690 42700 14700 42756
rect 14756 42700 16492 42756
rect 16548 42700 16558 42756
rect 20850 42700 20860 42756
rect 20916 42700 21980 42756
rect 22036 42700 22046 42756
rect 3154 42588 3164 42644
rect 3220 42588 4004 42644
rect 5730 42588 5740 42644
rect 5796 42588 6636 42644
rect 6692 42588 6702 42644
rect 10322 42588 10332 42644
rect 10388 42588 11788 42644
rect 11844 42588 11854 42644
rect 18498 42588 18508 42644
rect 18564 42588 19292 42644
rect 19348 42588 19358 42644
rect 20514 42588 20524 42644
rect 20580 42588 20748 42644
rect 20804 42588 21420 42644
rect 21476 42588 21486 42644
rect 3948 42532 4004 42588
rect 24556 42532 24612 42812
rect 26226 42700 26236 42756
rect 26292 42700 27356 42756
rect 27412 42700 27422 42756
rect 32050 42700 32060 42756
rect 32116 42700 33068 42756
rect 33124 42700 33134 42756
rect 33282 42700 33292 42756
rect 33348 42700 34076 42756
rect 34132 42700 34142 42756
rect 38210 42700 38220 42756
rect 38276 42700 39004 42756
rect 39060 42700 39070 42756
rect 33068 42644 33124 42700
rect 33068 42588 33628 42644
rect 33684 42588 33694 42644
rect 2818 42476 2828 42532
rect 2884 42476 3052 42532
rect 3108 42476 3724 42532
rect 3780 42476 3790 42532
rect 3938 42476 3948 42532
rect 4004 42476 4732 42532
rect 4788 42476 4798 42532
rect 14802 42476 14812 42532
rect 14868 42476 16268 42532
rect 16324 42476 16334 42532
rect 24556 42476 28364 42532
rect 28420 42476 28430 42532
rect 32946 42476 32956 42532
rect 33012 42476 34300 42532
rect 34356 42476 34366 42532
rect 36306 42476 36316 42532
rect 36372 42476 37100 42532
rect 37156 42476 37166 42532
rect 38098 42476 38108 42532
rect 38164 42476 38556 42532
rect 38612 42476 38622 42532
rect 47170 42476 47180 42532
rect 47236 42476 48412 42532
rect 48468 42476 48478 42532
rect 2594 42364 2604 42420
rect 2660 42364 4060 42420
rect 4116 42364 4126 42420
rect 19826 42308 19836 42364
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 20100 42308 20110 42364
rect 9090 42252 9100 42308
rect 9156 42252 9996 42308
rect 10052 42252 10444 42308
rect 10500 42252 10510 42308
rect 34514 42252 34524 42308
rect 34580 42252 38668 42308
rect 38612 42196 38668 42252
rect 8754 42140 8764 42196
rect 8820 42140 8988 42196
rect 9044 42140 10892 42196
rect 10948 42140 10958 42196
rect 31826 42140 31836 42196
rect 31892 42140 37212 42196
rect 37268 42140 37278 42196
rect 38612 42140 39340 42196
rect 39396 42140 39406 42196
rect 3490 42028 3500 42084
rect 3556 42028 4284 42084
rect 4340 42028 4350 42084
rect 5954 42028 5964 42084
rect 6020 42028 6748 42084
rect 6804 42028 8204 42084
rect 8260 42028 11116 42084
rect 11172 42028 11182 42084
rect 17826 42028 17836 42084
rect 17892 42028 19068 42084
rect 19124 42028 19134 42084
rect 20514 42028 20524 42084
rect 20580 42028 23884 42084
rect 23940 42028 23950 42084
rect 34738 42028 34748 42084
rect 34804 42028 41356 42084
rect 41412 42028 41422 42084
rect 46050 42028 46060 42084
rect 46116 42028 47068 42084
rect 47124 42028 47134 42084
rect 1810 41916 1820 41972
rect 1876 41916 5404 41972
rect 5460 41916 8652 41972
rect 8708 41916 12572 41972
rect 12628 41916 12638 41972
rect 20626 41916 20636 41972
rect 20692 41916 21644 41972
rect 21700 41916 22652 41972
rect 22708 41916 22718 41972
rect 24658 41916 24668 41972
rect 24724 41916 25340 41972
rect 25396 41916 25406 41972
rect 27682 41916 27692 41972
rect 27748 41916 29260 41972
rect 29316 41916 29326 41972
rect 33394 41916 33404 41972
rect 33460 41916 35196 41972
rect 35252 41916 35262 41972
rect 45714 41916 45724 41972
rect 45780 41916 48076 41972
rect 48132 41916 48142 41972
rect 8194 41804 8204 41860
rect 8260 41804 9660 41860
rect 9716 41804 9726 41860
rect 13346 41804 13356 41860
rect 13412 41804 15148 41860
rect 15204 41804 15214 41860
rect 16706 41804 16716 41860
rect 16772 41804 25228 41860
rect 25284 41804 25564 41860
rect 25620 41804 25630 41860
rect 28578 41804 28588 41860
rect 28644 41804 29820 41860
rect 29876 41804 30716 41860
rect 30772 41804 30782 41860
rect 33842 41804 33852 41860
rect 33908 41804 36764 41860
rect 36820 41804 39116 41860
rect 39172 41804 39182 41860
rect 8082 41692 8092 41748
rect 8148 41692 9212 41748
rect 9268 41692 9278 41748
rect 17602 41692 17612 41748
rect 17668 41692 19180 41748
rect 19236 41692 19246 41748
rect 33058 41692 33068 41748
rect 33124 41692 34524 41748
rect 34580 41692 36540 41748
rect 36596 41692 36606 41748
rect 40114 41692 40124 41748
rect 40180 41692 41468 41748
rect 41524 41692 41534 41748
rect 43474 41692 43484 41748
rect 43540 41692 45724 41748
rect 45780 41692 45790 41748
rect 15250 41580 15260 41636
rect 15316 41580 15820 41636
rect 15876 41580 15886 41636
rect 4466 41524 4476 41580
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4740 41524 4750 41580
rect 35186 41524 35196 41580
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35460 41524 35470 41580
rect 10770 41468 10780 41524
rect 10836 41468 16492 41524
rect 16548 41468 16558 41524
rect 38770 41468 38780 41524
rect 38836 41468 39340 41524
rect 39396 41468 39406 41524
rect 8194 41356 8204 41412
rect 8260 41356 11004 41412
rect 11060 41356 11070 41412
rect 14466 41356 14476 41412
rect 14532 41356 25676 41412
rect 25732 41356 25900 41412
rect 25956 41356 25966 41412
rect 31490 41356 31500 41412
rect 31556 41356 37212 41412
rect 37268 41356 42812 41412
rect 42868 41356 42878 41412
rect 7298 41244 7308 41300
rect 7364 41244 9884 41300
rect 9940 41244 9950 41300
rect 15026 41244 15036 41300
rect 15092 41244 15260 41300
rect 15316 41244 15326 41300
rect 25106 41244 25116 41300
rect 25172 41244 25452 41300
rect 25508 41244 25518 41300
rect 25778 41244 25788 41300
rect 25844 41244 28700 41300
rect 28756 41244 32508 41300
rect 32564 41244 33852 41300
rect 33908 41244 33918 41300
rect 10434 41132 10444 41188
rect 10500 41132 11228 41188
rect 11284 41132 11294 41188
rect 11554 41132 11564 41188
rect 11620 41132 13804 41188
rect 13860 41132 13870 41188
rect 27794 41132 27804 41188
rect 27860 41132 29036 41188
rect 29092 41132 29102 41188
rect 32834 41132 32844 41188
rect 32900 41132 33404 41188
rect 33460 41132 36988 41188
rect 37044 41132 37054 41188
rect 38770 41132 38780 41188
rect 38836 41132 39564 41188
rect 39620 41132 39630 41188
rect 17938 41020 17948 41076
rect 18004 41020 18396 41076
rect 18452 41020 18462 41076
rect 29922 41020 29932 41076
rect 29988 41020 33068 41076
rect 33124 41020 33134 41076
rect 35746 41020 35756 41076
rect 35812 41020 37100 41076
rect 37156 41020 37166 41076
rect 37650 41020 37660 41076
rect 37716 41020 38444 41076
rect 38500 41020 38510 41076
rect 8978 40908 8988 40964
rect 9044 40908 9660 40964
rect 9716 40908 9996 40964
rect 10052 40908 10780 40964
rect 10836 40908 10846 40964
rect 15250 40908 15260 40964
rect 15316 40908 15932 40964
rect 15988 40908 15998 40964
rect 19170 40908 19180 40964
rect 19236 40908 19628 40964
rect 19684 40908 20524 40964
rect 20580 40908 20590 40964
rect 33842 40908 33852 40964
rect 33908 40908 34972 40964
rect 35028 40908 35038 40964
rect 38322 40908 38332 40964
rect 38388 40908 38668 40964
rect 38724 40908 40348 40964
rect 40404 40908 40414 40964
rect 9884 40796 13132 40852
rect 13188 40796 14140 40852
rect 14196 40796 14206 40852
rect 9884 40628 9940 40796
rect 19826 40740 19836 40796
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 20100 40740 20110 40796
rect 10892 40684 14028 40740
rect 14084 40684 14094 40740
rect 31714 40684 31724 40740
rect 31780 40684 33180 40740
rect 33236 40684 34636 40740
rect 34692 40684 34702 40740
rect 4162 40572 4172 40628
rect 4228 40572 9884 40628
rect 9940 40572 9950 40628
rect 10892 40516 10948 40684
rect 11106 40572 11116 40628
rect 11172 40572 13580 40628
rect 13636 40572 13646 40628
rect 28466 40572 28476 40628
rect 28532 40572 28924 40628
rect 28980 40572 29820 40628
rect 29876 40572 29886 40628
rect 33506 40572 33516 40628
rect 33572 40572 34412 40628
rect 34468 40572 36428 40628
rect 36484 40572 36494 40628
rect 1698 40460 1708 40516
rect 1764 40460 3164 40516
rect 3220 40460 4508 40516
rect 4564 40460 4574 40516
rect 4722 40460 4732 40516
rect 4788 40460 7980 40516
rect 8036 40460 8046 40516
rect 8978 40460 8988 40516
rect 9044 40460 10780 40516
rect 10836 40460 10948 40516
rect 11778 40460 11788 40516
rect 11844 40460 13468 40516
rect 13524 40460 13534 40516
rect 15362 40460 15372 40516
rect 15428 40460 16156 40516
rect 16212 40460 17612 40516
rect 17668 40460 17678 40516
rect 23874 40460 23884 40516
rect 23940 40460 24668 40516
rect 24724 40460 24734 40516
rect 27906 40460 27916 40516
rect 27972 40460 29036 40516
rect 29092 40460 29708 40516
rect 29764 40460 29774 40516
rect 32050 40460 32060 40516
rect 32116 40460 33628 40516
rect 33684 40460 33964 40516
rect 34020 40460 34030 40516
rect 34738 40460 34748 40516
rect 34804 40460 35756 40516
rect 35812 40460 35822 40516
rect 40908 40460 41916 40516
rect 41972 40460 43820 40516
rect 43876 40460 43886 40516
rect 45602 40460 45612 40516
rect 45668 40460 46172 40516
rect 46228 40460 47516 40516
rect 47572 40460 47582 40516
rect 47954 40460 47964 40516
rect 48020 40460 48188 40516
rect 48244 40460 48254 40516
rect 4732 40404 4788 40460
rect 40908 40404 40964 40460
rect 2818 40348 2828 40404
rect 2884 40348 4788 40404
rect 7858 40348 7868 40404
rect 7924 40348 11396 40404
rect 7868 40292 7924 40348
rect 11340 40292 11396 40348
rect 11788 40348 15596 40404
rect 15652 40348 19404 40404
rect 19460 40348 19470 40404
rect 24434 40348 24444 40404
rect 24500 40348 25228 40404
rect 25284 40348 25294 40404
rect 28018 40348 28028 40404
rect 28084 40348 30044 40404
rect 30100 40348 30110 40404
rect 35298 40348 35308 40404
rect 35364 40348 36540 40404
rect 36596 40348 37436 40404
rect 37492 40348 38892 40404
rect 38948 40348 38958 40404
rect 39788 40348 40908 40404
rect 40964 40348 40974 40404
rect 41122 40348 41132 40404
rect 41188 40348 42252 40404
rect 42308 40348 42700 40404
rect 42756 40348 45388 40404
rect 45444 40348 45454 40404
rect 11788 40292 11844 40348
rect 35308 40292 35364 40348
rect 5730 40236 5740 40292
rect 5796 40236 7924 40292
rect 8418 40236 8428 40292
rect 8484 40236 8652 40292
rect 8708 40236 8718 40292
rect 11340 40236 11844 40292
rect 21186 40236 21196 40292
rect 21252 40236 27356 40292
rect 27412 40236 27422 40292
rect 32386 40236 32396 40292
rect 32452 40236 35364 40292
rect 35746 40236 35756 40292
rect 35812 40236 37100 40292
rect 37156 40236 37166 40292
rect 39788 40180 39844 40348
rect 45490 40236 45500 40292
rect 45556 40236 46396 40292
rect 46452 40236 47012 40292
rect 46956 40180 47012 40236
rect 8306 40124 8316 40180
rect 8372 40124 9436 40180
rect 9492 40124 9502 40180
rect 20738 40124 20748 40180
rect 20804 40124 21980 40180
rect 22036 40124 22428 40180
rect 22484 40124 22494 40180
rect 32162 40124 32172 40180
rect 32228 40124 39844 40180
rect 44146 40124 44156 40180
rect 44212 40124 45836 40180
rect 45892 40124 45902 40180
rect 46946 40124 46956 40180
rect 47012 40124 47404 40180
rect 47460 40124 47470 40180
rect 12562 40012 12572 40068
rect 12628 40012 12638 40068
rect 17938 40012 17948 40068
rect 18004 40012 19516 40068
rect 19572 40012 19582 40068
rect 28354 40012 28364 40068
rect 28420 40012 30940 40068
rect 30996 40012 31006 40068
rect 47058 40012 47068 40068
rect 47124 40012 47964 40068
rect 48020 40012 48030 40068
rect 4466 39956 4476 40012
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4740 39956 4750 40012
rect 12572 39620 12628 40012
rect 35186 39956 35196 40012
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35460 39956 35470 40012
rect 16594 39900 16604 39956
rect 16660 39900 28812 39956
rect 28868 39900 29260 39956
rect 29316 39900 30380 39956
rect 30436 39900 30446 39956
rect 38994 39900 39004 39956
rect 39060 39900 42476 39956
rect 42532 39900 42542 39956
rect 44156 39900 47180 39956
rect 47236 39900 47246 39956
rect 13010 39788 13020 39844
rect 13076 39788 14028 39844
rect 14084 39788 14094 39844
rect 20066 39788 20076 39844
rect 20132 39788 27468 39844
rect 27524 39788 27534 39844
rect 34178 39788 34188 39844
rect 34244 39788 35644 39844
rect 35700 39788 35710 39844
rect 44156 39732 44212 39900
rect 12898 39676 12908 39732
rect 12964 39676 15148 39732
rect 22194 39676 22204 39732
rect 22260 39676 27132 39732
rect 27188 39676 27198 39732
rect 33282 39676 33292 39732
rect 33348 39676 34076 39732
rect 34132 39676 35308 39732
rect 35364 39676 35374 39732
rect 43362 39676 43372 39732
rect 43428 39676 44156 39732
rect 44212 39676 44222 39732
rect 46722 39676 46732 39732
rect 46788 39676 47068 39732
rect 47124 39676 47134 39732
rect 4834 39564 4844 39620
rect 4900 39564 5740 39620
rect 5796 39564 5806 39620
rect 11778 39564 11788 39620
rect 11844 39564 12236 39620
rect 12292 39564 12302 39620
rect 12562 39564 12572 39620
rect 12628 39564 14028 39620
rect 14084 39564 14094 39620
rect 7410 39452 7420 39508
rect 7476 39452 8540 39508
rect 8596 39452 10444 39508
rect 10500 39452 10510 39508
rect 12786 39452 12796 39508
rect 12852 39452 13356 39508
rect 13412 39452 13422 39508
rect 6514 39340 6524 39396
rect 6580 39340 8988 39396
rect 9044 39340 9054 39396
rect 13122 39340 13132 39396
rect 13188 39340 13692 39396
rect 13748 39340 13758 39396
rect 15092 39284 15148 39676
rect 15362 39564 15372 39620
rect 15428 39564 15820 39620
rect 15876 39564 15886 39620
rect 24098 39564 24108 39620
rect 24164 39564 25004 39620
rect 25060 39564 25070 39620
rect 28578 39564 28588 39620
rect 28644 39564 28924 39620
rect 28980 39564 28990 39620
rect 43250 39564 43260 39620
rect 43316 39564 47628 39620
rect 47684 39564 47694 39620
rect 15474 39452 15484 39508
rect 15540 39452 22316 39508
rect 22372 39452 22382 39508
rect 23538 39452 23548 39508
rect 23604 39452 23996 39508
rect 24052 39452 24062 39508
rect 27906 39452 27916 39508
rect 27972 39452 29036 39508
rect 29092 39452 30716 39508
rect 30772 39452 30782 39508
rect 31266 39452 31276 39508
rect 31332 39452 37548 39508
rect 37604 39452 37996 39508
rect 38052 39452 38062 39508
rect 45490 39452 45500 39508
rect 45556 39452 46732 39508
rect 46788 39452 46798 39508
rect 15362 39340 15372 39396
rect 15428 39340 16044 39396
rect 16100 39340 16110 39396
rect 17602 39340 17612 39396
rect 17668 39340 18508 39396
rect 18564 39340 18574 39396
rect 23314 39340 23324 39396
rect 23380 39340 24556 39396
rect 24612 39340 24622 39396
rect 26338 39340 26348 39396
rect 26404 39340 27356 39396
rect 27412 39340 27422 39396
rect 32050 39340 32060 39396
rect 32116 39340 32396 39396
rect 32452 39340 32462 39396
rect 33730 39340 33740 39396
rect 33796 39340 36428 39396
rect 36484 39340 36494 39396
rect 7634 39228 7644 39284
rect 7700 39228 8204 39284
rect 8260 39228 8652 39284
rect 8708 39228 10892 39284
rect 10948 39228 10958 39284
rect 15092 39228 17948 39284
rect 18004 39228 18014 39284
rect 31714 39228 31724 39284
rect 31780 39228 33292 39284
rect 33348 39228 33358 39284
rect 33506 39228 33516 39284
rect 33572 39228 35980 39284
rect 36036 39228 36046 39284
rect 19826 39172 19836 39228
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 20100 39172 20110 39228
rect 5170 39116 5180 39172
rect 5236 39116 6300 39172
rect 6356 39116 6972 39172
rect 7028 39116 7308 39172
rect 7364 39116 15652 39172
rect 15810 39116 15820 39172
rect 15876 39116 19516 39172
rect 19572 39116 19582 39172
rect 22418 39116 22428 39172
rect 22484 39116 28028 39172
rect 28084 39116 28094 39172
rect 8306 39004 8316 39060
rect 8372 39004 9212 39060
rect 9268 39004 11788 39060
rect 11844 39004 11854 39060
rect 13346 39004 13356 39060
rect 13412 39004 14028 39060
rect 14084 39004 14094 39060
rect 15596 38948 15652 39116
rect 17154 39004 17164 39060
rect 17220 39004 17948 39060
rect 18004 39004 30380 39060
rect 30436 39004 31276 39060
rect 31332 39004 31342 39060
rect 31826 39004 31836 39060
rect 31892 39004 33180 39060
rect 33236 39004 33246 39060
rect 8978 38892 8988 38948
rect 9044 38892 11844 38948
rect 12674 38892 12684 38948
rect 12740 38892 15372 38948
rect 15428 38892 15438 38948
rect 15596 38892 17388 38948
rect 17444 38892 17454 38948
rect 18386 38892 18396 38948
rect 18452 38892 19628 38948
rect 19684 38892 21084 38948
rect 21140 38892 21150 38948
rect 24658 38892 24668 38948
rect 24724 38892 26124 38948
rect 26180 38892 26190 38948
rect 33954 38892 33964 38948
rect 34020 38892 38556 38948
rect 38612 38892 38622 38948
rect 11788 38836 11844 38892
rect 8082 38780 8092 38836
rect 8148 38780 9548 38836
rect 9604 38780 10220 38836
rect 10276 38780 10286 38836
rect 11778 38780 11788 38836
rect 11844 38780 12124 38836
rect 12180 38780 12190 38836
rect 12450 38780 12460 38836
rect 12516 38780 13692 38836
rect 13748 38780 13758 38836
rect 19170 38780 19180 38836
rect 19236 38780 22988 38836
rect 23044 38780 23054 38836
rect 23202 38780 23212 38836
rect 23268 38780 23772 38836
rect 23828 38780 24556 38836
rect 24612 38780 24622 38836
rect 31938 38780 31948 38836
rect 32004 38780 33068 38836
rect 33124 38780 33134 38836
rect 45938 38780 45948 38836
rect 46004 38780 46732 38836
rect 46788 38780 46798 38836
rect 47394 38780 47404 38836
rect 47460 38780 48076 38836
rect 48132 38780 48142 38836
rect 3826 38668 3836 38724
rect 3892 38668 5068 38724
rect 5124 38668 5134 38724
rect 7522 38668 7532 38724
rect 7588 38668 10108 38724
rect 10164 38668 10174 38724
rect 16370 38668 16380 38724
rect 16436 38668 21308 38724
rect 21364 38668 21374 38724
rect 24322 38668 24332 38724
rect 24388 38668 25228 38724
rect 25284 38668 25294 38724
rect 38882 38668 38892 38724
rect 38948 38668 40460 38724
rect 40516 38668 40526 38724
rect 42914 38668 42924 38724
rect 42980 38668 43932 38724
rect 43988 38668 43998 38724
rect 48178 38668 48188 38724
rect 48244 38668 48254 38724
rect 48188 38612 48244 38668
rect 49200 38612 50000 38640
rect 4162 38556 4172 38612
rect 4228 38556 4956 38612
rect 5012 38556 5022 38612
rect 5282 38556 5292 38612
rect 5348 38556 5740 38612
rect 5796 38556 5806 38612
rect 13794 38556 13804 38612
rect 13860 38556 14812 38612
rect 14868 38556 15148 38612
rect 15204 38556 15214 38612
rect 28354 38556 28364 38612
rect 28420 38556 31164 38612
rect 31220 38556 31836 38612
rect 31892 38556 31902 38612
rect 48188 38556 50000 38612
rect 49200 38528 50000 38556
rect 20066 38444 20076 38500
rect 20132 38444 21980 38500
rect 22036 38444 22046 38500
rect 4466 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4750 38444
rect 35186 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35470 38444
rect 15092 38332 24780 38388
rect 24836 38332 24846 38388
rect 15092 38276 15148 38332
rect 11778 38220 11788 38276
rect 11844 38220 15148 38276
rect 19282 38220 19292 38276
rect 19348 38220 21868 38276
rect 21924 38220 21934 38276
rect 39890 38220 39900 38276
rect 39956 38220 42028 38276
rect 42084 38220 42094 38276
rect 42354 38220 42364 38276
rect 42420 38220 43820 38276
rect 43876 38220 45276 38276
rect 45332 38220 45342 38276
rect 11218 38108 11228 38164
rect 11284 38108 13692 38164
rect 13748 38108 13758 38164
rect 19170 38108 19180 38164
rect 19236 38108 19628 38164
rect 19684 38108 19694 38164
rect 20178 38108 20188 38164
rect 20244 38108 28252 38164
rect 28308 38108 28318 38164
rect 38770 38108 38780 38164
rect 38836 38108 40124 38164
rect 40180 38108 40190 38164
rect 9986 37996 9996 38052
rect 10052 37996 10780 38052
rect 10836 37996 11900 38052
rect 11956 37996 11966 38052
rect 12674 37996 12684 38052
rect 12740 37996 13580 38052
rect 13636 37996 13646 38052
rect 14242 37996 14252 38052
rect 14308 37996 16156 38052
rect 16212 37996 16222 38052
rect 16594 37996 16604 38052
rect 16660 37996 23996 38052
rect 24052 37996 24062 38052
rect 24210 37996 24220 38052
rect 24276 37996 26572 38052
rect 26628 37996 26638 38052
rect 28018 37996 28028 38052
rect 28084 37996 29148 38052
rect 29204 37996 29214 38052
rect 30930 37996 30940 38052
rect 30996 37996 32396 38052
rect 32452 37996 32462 38052
rect 33618 37996 33628 38052
rect 33684 37996 34076 38052
rect 34132 37996 34142 38052
rect 41570 37996 41580 38052
rect 41636 37996 42476 38052
rect 42532 37996 42812 38052
rect 42868 37996 42878 38052
rect 46162 37996 46172 38052
rect 46228 37996 46844 38052
rect 46900 37996 46910 38052
rect 6514 37884 6524 37940
rect 6580 37884 7420 37940
rect 7476 37884 8204 37940
rect 8260 37884 8270 37940
rect 9314 37884 9324 37940
rect 9380 37884 9660 37940
rect 9716 37884 11004 37940
rect 11060 37884 11070 37940
rect 12338 37884 12348 37940
rect 12404 37884 13692 37940
rect 13748 37884 17612 37940
rect 17668 37884 17678 37940
rect 19170 37884 19180 37940
rect 19236 37884 20748 37940
rect 20804 37884 20814 37940
rect 21746 37884 21756 37940
rect 21812 37884 23100 37940
rect 23156 37884 26908 37940
rect 26964 37884 26974 37940
rect 45378 37884 45388 37940
rect 45444 37884 47292 37940
rect 47348 37884 47358 37940
rect 20748 37828 20804 37884
rect 6178 37772 6188 37828
rect 6244 37772 7196 37828
rect 7252 37772 7262 37828
rect 10210 37772 10220 37828
rect 10276 37772 13132 37828
rect 13188 37772 13198 37828
rect 18834 37772 18844 37828
rect 18900 37772 19404 37828
rect 19460 37772 20692 37828
rect 20748 37772 21644 37828
rect 21700 37772 22652 37828
rect 22708 37772 22718 37828
rect 25890 37772 25900 37828
rect 25956 37772 33068 37828
rect 33124 37772 33134 37828
rect 33394 37772 33404 37828
rect 33460 37772 33964 37828
rect 34020 37772 34030 37828
rect 38210 37772 38220 37828
rect 38276 37772 39676 37828
rect 39732 37772 40236 37828
rect 40292 37772 40302 37828
rect 7074 37660 7084 37716
rect 7140 37660 8652 37716
rect 8708 37660 8988 37716
rect 9044 37660 9054 37716
rect 19826 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20110 37660
rect 20636 37604 20692 37772
rect 21858 37660 21868 37716
rect 21924 37660 22316 37716
rect 22372 37660 22382 37716
rect 20636 37548 36988 37604
rect 37044 37548 37054 37604
rect 37538 37548 37548 37604
rect 37604 37548 38500 37604
rect 38444 37492 38500 37548
rect 18162 37436 18172 37492
rect 18228 37436 19852 37492
rect 19908 37436 19918 37492
rect 22754 37436 22764 37492
rect 22820 37436 23772 37492
rect 23828 37436 23838 37492
rect 24098 37436 24108 37492
rect 24164 37436 25452 37492
rect 25508 37436 26012 37492
rect 26068 37436 26078 37492
rect 37426 37436 37436 37492
rect 37492 37436 38220 37492
rect 38276 37436 38286 37492
rect 38444 37436 38556 37492
rect 38612 37436 39228 37492
rect 39284 37436 39294 37492
rect 41906 37436 41916 37492
rect 41972 37436 42700 37492
rect 42756 37436 42766 37492
rect 2930 37324 2940 37380
rect 2996 37324 4172 37380
rect 4228 37324 4238 37380
rect 12338 37324 12348 37380
rect 12404 37324 12684 37380
rect 12740 37324 15148 37380
rect 15204 37324 15214 37380
rect 16706 37324 16716 37380
rect 16772 37324 20860 37380
rect 20916 37324 20926 37380
rect 25330 37324 25340 37380
rect 25396 37324 27804 37380
rect 27860 37324 27870 37380
rect 39778 37324 39788 37380
rect 39844 37324 40348 37380
rect 40404 37324 43372 37380
rect 43428 37324 43438 37380
rect 43586 37324 43596 37380
rect 43652 37324 46284 37380
rect 46340 37324 47180 37380
rect 47236 37324 47246 37380
rect 2818 37212 2828 37268
rect 2884 37212 3724 37268
rect 3780 37212 3790 37268
rect 5170 37212 5180 37268
rect 5236 37212 8988 37268
rect 9044 37212 9660 37268
rect 9716 37212 9726 37268
rect 14690 37212 14700 37268
rect 14756 37212 15372 37268
rect 15428 37212 15438 37268
rect 18274 37212 18284 37268
rect 18340 37212 19740 37268
rect 19796 37212 19806 37268
rect 20962 37212 20972 37268
rect 21028 37212 21868 37268
rect 21924 37212 21934 37268
rect 22306 37212 22316 37268
rect 22372 37212 24556 37268
rect 24612 37212 24622 37268
rect 24770 37212 24780 37268
rect 24836 37212 25228 37268
rect 25284 37212 25564 37268
rect 25620 37212 26460 37268
rect 26516 37212 26526 37268
rect 26786 37212 26796 37268
rect 26852 37212 30044 37268
rect 30100 37212 32172 37268
rect 32228 37212 32238 37268
rect 32498 37212 32508 37268
rect 32564 37212 33852 37268
rect 33908 37212 33918 37268
rect 41570 37212 41580 37268
rect 41636 37212 42252 37268
rect 42308 37212 42318 37268
rect 46498 37212 46508 37268
rect 46564 37212 47068 37268
rect 47124 37212 47134 37268
rect 18162 37100 18172 37156
rect 18228 37100 18844 37156
rect 18900 37100 19964 37156
rect 20020 37100 20030 37156
rect 22194 37100 22204 37156
rect 22260 37100 23436 37156
rect 23492 37100 23502 37156
rect 27458 37100 27468 37156
rect 27524 37100 29484 37156
rect 29540 37100 29550 37156
rect 30706 37100 30716 37156
rect 30772 37100 34524 37156
rect 34580 37100 35084 37156
rect 35140 37100 35644 37156
rect 35700 37100 35710 37156
rect 42130 37100 42140 37156
rect 42196 37100 42924 37156
rect 42980 37100 42990 37156
rect 43148 37100 47180 37156
rect 47236 37100 47246 37156
rect 43148 37044 43204 37100
rect 4162 36988 4172 37044
rect 4228 36988 5068 37044
rect 5124 36988 5134 37044
rect 6626 36988 6636 37044
rect 6692 36988 7980 37044
rect 8036 36988 8652 37044
rect 8708 36988 8718 37044
rect 9874 36988 9884 37044
rect 9940 36988 9950 37044
rect 10658 36988 10668 37044
rect 10724 36988 11452 37044
rect 11508 36988 12012 37044
rect 12068 36988 12078 37044
rect 16034 36988 16044 37044
rect 16100 36988 16828 37044
rect 16884 36988 18060 37044
rect 18116 36988 18126 37044
rect 18386 36988 18396 37044
rect 18452 36988 19292 37044
rect 19348 36988 19358 37044
rect 20850 36988 20860 37044
rect 20916 36988 22540 37044
rect 22596 36988 22988 37044
rect 23044 36988 23054 37044
rect 28354 36988 28364 37044
rect 28420 36988 32956 37044
rect 33012 36988 33404 37044
rect 33460 36988 33470 37044
rect 40450 36988 40460 37044
rect 40516 36988 43204 37044
rect 46834 36988 46844 37044
rect 46900 36988 47852 37044
rect 47908 36988 47918 37044
rect 9884 36932 9940 36988
rect 9884 36876 11004 36932
rect 11060 36876 11070 36932
rect 11228 36876 16604 36932
rect 16660 36876 16670 36932
rect 16930 36876 16940 36932
rect 16996 36876 18844 36932
rect 18900 36876 18910 36932
rect 19170 36876 19180 36932
rect 19236 36876 20076 36932
rect 20132 36876 20142 36932
rect 21494 36876 21532 36932
rect 21588 36876 21598 36932
rect 4466 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4750 36876
rect 11228 36820 11284 36876
rect 16940 36820 16996 36876
rect 19180 36820 19236 36876
rect 35186 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35470 36876
rect 8978 36764 8988 36820
rect 9044 36764 11284 36820
rect 12002 36764 12012 36820
rect 12068 36764 16996 36820
rect 18274 36764 18284 36820
rect 18340 36764 19236 36820
rect 19366 36764 19404 36820
rect 19460 36764 19470 36820
rect 21410 36764 21420 36820
rect 21476 36764 21644 36820
rect 21700 36764 21710 36820
rect 1810 36652 1820 36708
rect 1876 36652 3948 36708
rect 4004 36652 5404 36708
rect 5460 36652 5740 36708
rect 5796 36652 8204 36708
rect 8260 36652 8270 36708
rect 10546 36652 10556 36708
rect 10612 36652 16492 36708
rect 16548 36652 16558 36708
rect 5506 36540 5516 36596
rect 5572 36540 5852 36596
rect 5908 36540 12012 36596
rect 12068 36540 12078 36596
rect 12562 36540 12572 36596
rect 12628 36540 17388 36596
rect 17444 36540 17454 36596
rect 18050 36540 18060 36596
rect 18116 36540 30940 36596
rect 30996 36540 31006 36596
rect 32162 36540 32172 36596
rect 32228 36540 33180 36596
rect 33236 36540 33246 36596
rect 41794 36540 41804 36596
rect 41860 36540 42812 36596
rect 42868 36540 42878 36596
rect 9986 36428 9996 36484
rect 10052 36428 10780 36484
rect 10836 36428 10846 36484
rect 11890 36428 11900 36484
rect 11956 36428 13580 36484
rect 13636 36428 13646 36484
rect 20402 36428 20412 36484
rect 20468 36428 21532 36484
rect 21588 36428 21598 36484
rect 30370 36428 30380 36484
rect 30436 36428 31164 36484
rect 31220 36428 33628 36484
rect 33684 36428 33694 36484
rect 10434 36316 10444 36372
rect 10500 36316 11676 36372
rect 11732 36316 12796 36372
rect 12852 36316 12862 36372
rect 20962 36316 20972 36372
rect 21028 36316 24668 36372
rect 24724 36316 24734 36372
rect 34738 36316 34748 36372
rect 34804 36316 35308 36372
rect 35364 36316 35374 36372
rect 35858 36316 35868 36372
rect 35924 36316 36316 36372
rect 36372 36316 36988 36372
rect 37044 36316 37054 36372
rect 40114 36316 40124 36372
rect 40180 36316 42140 36372
rect 42196 36316 42206 36372
rect 20188 36204 21308 36260
rect 21364 36204 21374 36260
rect 29474 36204 29484 36260
rect 29540 36204 30716 36260
rect 30772 36204 30782 36260
rect 36194 36204 36204 36260
rect 36260 36204 37772 36260
rect 37828 36204 37838 36260
rect 46946 36204 46956 36260
rect 47012 36204 47516 36260
rect 47572 36204 48188 36260
rect 48244 36204 48254 36260
rect 9874 36092 9884 36148
rect 9940 36092 11676 36148
rect 11732 36092 17276 36148
rect 17332 36092 17342 36148
rect 19826 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20110 36092
rect 16370 35980 16380 36036
rect 16436 35980 18956 36036
rect 19012 35980 19022 36036
rect 20188 35924 20244 36204
rect 20626 36092 20636 36148
rect 20692 36092 21868 36148
rect 21924 36092 22316 36148
rect 22372 36092 22382 36148
rect 27010 36092 27020 36148
rect 27076 36092 28364 36148
rect 28420 36092 29260 36148
rect 29316 36092 29326 36148
rect 4162 35868 4172 35924
rect 4228 35868 4732 35924
rect 4788 35868 4798 35924
rect 15698 35868 15708 35924
rect 15764 35868 19404 35924
rect 19460 35868 19470 35924
rect 19954 35868 19964 35924
rect 20020 35868 20244 35924
rect 10070 35756 10108 35812
rect 10164 35756 10174 35812
rect 16482 35756 16492 35812
rect 16548 35756 17500 35812
rect 17556 35756 17566 35812
rect 19506 35756 19516 35812
rect 19572 35756 21532 35812
rect 21588 35756 21598 35812
rect 28802 35756 28812 35812
rect 28868 35756 29596 35812
rect 29652 35756 29662 35812
rect 8754 35644 8764 35700
rect 8820 35644 9324 35700
rect 9380 35644 9390 35700
rect 11890 35644 11900 35700
rect 11956 35644 14252 35700
rect 14308 35644 14318 35700
rect 21074 35644 21084 35700
rect 21140 35644 22876 35700
rect 22932 35644 22942 35700
rect 26852 35644 28588 35700
rect 28644 35644 29372 35700
rect 29428 35644 29438 35700
rect 31154 35644 31164 35700
rect 31220 35644 36540 35700
rect 36596 35644 36606 35700
rect 4386 35532 4396 35588
rect 4452 35532 5516 35588
rect 5572 35532 5582 35588
rect 13794 35532 13804 35588
rect 13860 35532 15820 35588
rect 15876 35532 18172 35588
rect 18228 35532 18238 35588
rect 26852 35476 26908 35644
rect 33618 35532 33628 35588
rect 33684 35532 34412 35588
rect 34468 35532 34478 35588
rect 9650 35420 9660 35476
rect 9716 35420 9726 35476
rect 10434 35420 10444 35476
rect 10500 35420 15372 35476
rect 15428 35420 15438 35476
rect 24098 35420 24108 35476
rect 24164 35420 25340 35476
rect 25396 35420 26908 35476
rect 43250 35420 43260 35476
rect 43316 35420 45724 35476
rect 45780 35420 45948 35476
rect 46004 35420 46014 35476
rect 9660 35364 9716 35420
rect 9660 35308 10780 35364
rect 10836 35308 15260 35364
rect 15316 35308 15326 35364
rect 20626 35308 20636 35364
rect 20692 35308 21420 35364
rect 21476 35308 22204 35364
rect 22260 35308 22652 35364
rect 22708 35308 22718 35364
rect 42690 35308 42700 35364
rect 42756 35308 42766 35364
rect 4466 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4750 35308
rect 35186 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35470 35308
rect 42700 35252 42756 35308
rect 9398 35196 9436 35252
rect 9492 35196 9502 35252
rect 11442 35196 11452 35252
rect 11508 35196 12236 35252
rect 12292 35196 12302 35252
rect 16146 35196 16156 35252
rect 16212 35196 18620 35252
rect 18676 35196 18686 35252
rect 20066 35196 20076 35252
rect 20132 35196 20524 35252
rect 20580 35196 21924 35252
rect 22754 35196 22764 35252
rect 22820 35196 23548 35252
rect 23604 35196 23772 35252
rect 23828 35196 23838 35252
rect 38546 35196 38556 35252
rect 38612 35196 41356 35252
rect 41412 35196 43820 35252
rect 43876 35196 45388 35252
rect 45444 35196 45454 35252
rect 21868 35140 21924 35196
rect 10994 35084 11004 35140
rect 11060 35084 21700 35140
rect 21868 35084 23436 35140
rect 23492 35084 25340 35140
rect 25396 35084 25406 35140
rect 38612 35084 43260 35140
rect 43316 35084 43326 35140
rect 9538 34972 9548 35028
rect 9604 34972 9772 35028
rect 9828 34972 9838 35028
rect 13804 34972 15260 35028
rect 15316 34972 15326 35028
rect 19394 34972 19404 35028
rect 19460 34972 21420 35028
rect 21476 34972 21486 35028
rect 13804 34916 13860 34972
rect 21644 34916 21700 35084
rect 23986 34972 23996 35028
rect 24052 34972 25116 35028
rect 25172 34972 25564 35028
rect 25620 34972 27132 35028
rect 27188 34972 29148 35028
rect 29204 34972 29214 35028
rect 4946 34860 4956 34916
rect 5012 34860 5852 34916
rect 5908 34860 5918 34916
rect 7746 34860 7756 34916
rect 7812 34860 8764 34916
rect 8820 34860 10444 34916
rect 10500 34860 10510 34916
rect 12226 34860 12236 34916
rect 12292 34860 13580 34916
rect 13636 34860 13804 34916
rect 13860 34860 13870 34916
rect 15092 34860 17276 34916
rect 17332 34860 17342 34916
rect 19618 34860 19628 34916
rect 19684 34860 20300 34916
rect 20356 34860 20366 34916
rect 21644 34860 26908 34916
rect 27570 34860 27580 34916
rect 27636 34860 29708 34916
rect 29764 34860 30828 34916
rect 30884 34860 30894 34916
rect 38546 34860 38556 34916
rect 38612 34860 38668 35084
rect 15092 34804 15148 34860
rect 26852 34804 26908 34860
rect 3602 34748 3612 34804
rect 3668 34748 7420 34804
rect 7476 34748 7486 34804
rect 8306 34748 8316 34804
rect 8372 34748 11340 34804
rect 11396 34748 11406 34804
rect 11666 34748 11676 34804
rect 11732 34748 13916 34804
rect 13972 34748 15148 34804
rect 15362 34748 15372 34804
rect 15428 34748 19292 34804
rect 19348 34748 19358 34804
rect 21298 34748 21308 34804
rect 21364 34748 21374 34804
rect 23202 34748 23212 34804
rect 23268 34748 24780 34804
rect 24836 34748 24846 34804
rect 26852 34748 29484 34804
rect 29540 34748 29550 34804
rect 38612 34748 38780 34804
rect 38836 34748 38846 34804
rect 21308 34692 21364 34748
rect 28700 34692 28756 34748
rect 38612 34692 38668 34748
rect 2482 34636 2492 34692
rect 2548 34636 3500 34692
rect 3556 34636 3566 34692
rect 4834 34636 4844 34692
rect 4900 34636 6972 34692
rect 7028 34636 7038 34692
rect 8194 34636 8204 34692
rect 8260 34636 8876 34692
rect 8932 34636 11116 34692
rect 11172 34636 15596 34692
rect 15652 34636 15662 34692
rect 16258 34636 16268 34692
rect 16324 34636 21364 34692
rect 28690 34636 28700 34692
rect 28756 34636 28766 34692
rect 36082 34636 36092 34692
rect 36148 34636 37436 34692
rect 37492 34636 37884 34692
rect 37940 34636 38668 34692
rect 43474 34636 43484 34692
rect 43540 34636 44380 34692
rect 44436 34636 44446 34692
rect 2370 34524 2380 34580
rect 2436 34524 2940 34580
rect 2996 34524 3388 34580
rect 5058 34524 5068 34580
rect 5124 34524 7532 34580
rect 7588 34524 8540 34580
rect 8596 34524 8606 34580
rect 3332 34468 3388 34524
rect 19826 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20110 34524
rect 3332 34412 5740 34468
rect 5796 34412 5806 34468
rect 10546 34412 10556 34468
rect 10612 34412 12460 34468
rect 12516 34412 13468 34468
rect 13524 34412 13534 34468
rect 6962 34300 6972 34356
rect 7028 34300 7420 34356
rect 7476 34300 7486 34356
rect 14140 34300 15708 34356
rect 15764 34300 16156 34356
rect 16212 34300 16222 34356
rect 31266 34300 31276 34356
rect 31332 34300 31948 34356
rect 32004 34300 33180 34356
rect 33236 34300 33246 34356
rect 14140 34244 14196 34300
rect 7634 34188 7644 34244
rect 7700 34188 14140 34244
rect 14196 34188 14206 34244
rect 15092 34188 16716 34244
rect 16772 34188 16782 34244
rect 18498 34188 18508 34244
rect 18564 34188 23212 34244
rect 23268 34188 23278 34244
rect 26002 34188 26012 34244
rect 26068 34188 26572 34244
rect 26628 34188 26638 34244
rect 30818 34188 30828 34244
rect 30884 34188 31836 34244
rect 31892 34188 31902 34244
rect 33814 34188 33852 34244
rect 33908 34188 33918 34244
rect 37314 34188 37324 34244
rect 37380 34188 41468 34244
rect 41524 34188 41534 34244
rect 15092 34132 15148 34188
rect 2706 34076 2716 34132
rect 2772 34076 3612 34132
rect 3668 34076 3678 34132
rect 12114 34076 12124 34132
rect 12180 34076 14028 34132
rect 14084 34076 15148 34132
rect 15250 34076 15260 34132
rect 15316 34076 15932 34132
rect 15988 34076 15998 34132
rect 24294 34076 24332 34132
rect 24388 34076 24398 34132
rect 24658 34076 24668 34132
rect 24724 34076 25900 34132
rect 25956 34076 25966 34132
rect 33282 34076 33292 34132
rect 33348 34076 34524 34132
rect 34580 34076 35084 34132
rect 35140 34076 35150 34132
rect 43250 34076 43260 34132
rect 43316 34076 43820 34132
rect 43876 34076 43886 34132
rect 13122 33964 13132 34020
rect 13188 33964 13468 34020
rect 13524 33964 14140 34020
rect 14196 33964 14206 34020
rect 22502 33964 22540 34020
rect 22596 33964 22606 34020
rect 41682 33964 41692 34020
rect 41748 33964 44268 34020
rect 44324 33964 44334 34020
rect 46834 33964 46844 34020
rect 46900 33964 48188 34020
rect 48244 33964 48254 34020
rect 11442 33852 11452 33908
rect 11508 33852 14476 33908
rect 14532 33852 14542 33908
rect 16594 33852 16604 33908
rect 16660 33852 19068 33908
rect 19124 33852 19134 33908
rect 21522 33852 21532 33908
rect 21588 33852 22092 33908
rect 22148 33852 23996 33908
rect 24052 33852 24062 33908
rect 28242 33852 28252 33908
rect 28308 33852 30828 33908
rect 30884 33852 30894 33908
rect 31042 33852 31052 33908
rect 31108 33852 31948 33908
rect 32004 33852 32014 33908
rect 14018 33740 14028 33796
rect 14084 33740 15036 33796
rect 15092 33740 15102 33796
rect 19170 33740 19180 33796
rect 19236 33740 20524 33796
rect 20580 33740 20748 33796
rect 20804 33740 20814 33796
rect 22082 33740 22092 33796
rect 22148 33740 23212 33796
rect 23268 33740 23278 33796
rect 4466 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4750 33740
rect 35186 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35470 33740
rect 1698 33628 1708 33684
rect 1764 33628 2492 33684
rect 2548 33628 2558 33684
rect 5058 33628 5068 33684
rect 5124 33628 5740 33684
rect 5796 33628 5806 33684
rect 8978 33628 8988 33684
rect 9044 33628 10556 33684
rect 10612 33628 10622 33684
rect 15138 33628 15148 33684
rect 15204 33628 17724 33684
rect 17780 33628 19628 33684
rect 19684 33628 21308 33684
rect 21364 33628 21374 33684
rect 22652 33628 23548 33684
rect 23604 33628 23614 33684
rect 26898 33628 26908 33684
rect 26964 33628 27916 33684
rect 27972 33628 32508 33684
rect 32564 33628 32574 33684
rect 36950 33628 36988 33684
rect 37044 33628 37054 33684
rect 22652 33572 22708 33628
rect 6402 33516 6412 33572
rect 6468 33516 7196 33572
rect 7252 33516 7262 33572
rect 8642 33516 8652 33572
rect 8708 33516 9100 33572
rect 9156 33516 9166 33572
rect 10322 33516 10332 33572
rect 10388 33516 12012 33572
rect 12068 33516 12078 33572
rect 13906 33516 13916 33572
rect 13972 33516 18508 33572
rect 18564 33516 18574 33572
rect 20962 33516 20972 33572
rect 21028 33516 22316 33572
rect 22372 33516 22382 33572
rect 22642 33516 22652 33572
rect 22708 33516 22718 33572
rect 27794 33516 27804 33572
rect 27860 33516 29484 33572
rect 29540 33516 29820 33572
rect 29876 33516 29886 33572
rect 30146 33516 30156 33572
rect 30212 33516 30604 33572
rect 30660 33516 30670 33572
rect 33394 33516 33404 33572
rect 33460 33516 37436 33572
rect 37492 33516 37502 33572
rect 39106 33516 39116 33572
rect 39172 33516 40796 33572
rect 40852 33516 40862 33572
rect 2594 33404 2604 33460
rect 2660 33404 3612 33460
rect 3668 33404 3678 33460
rect 5618 33404 5628 33460
rect 5684 33404 6636 33460
rect 6692 33404 6702 33460
rect 8530 33404 8540 33460
rect 8596 33404 8606 33460
rect 9986 33404 9996 33460
rect 10052 33404 12124 33460
rect 12180 33404 12190 33460
rect 12450 33404 12460 33460
rect 12516 33404 17836 33460
rect 17892 33404 17902 33460
rect 25778 33404 25788 33460
rect 25844 33404 26684 33460
rect 26740 33404 26750 33460
rect 26852 33404 31164 33460
rect 31220 33404 31230 33460
rect 33170 33404 33180 33460
rect 33236 33404 33852 33460
rect 33908 33404 34748 33460
rect 34804 33404 34814 33460
rect 41234 33404 41244 33460
rect 41300 33404 41692 33460
rect 41748 33404 43148 33460
rect 43204 33404 43214 33460
rect 8540 33348 8596 33404
rect 15260 33348 15316 33404
rect 26852 33348 26908 33404
rect 8540 33292 8764 33348
rect 8820 33292 8830 33348
rect 10770 33292 10780 33348
rect 10836 33292 13804 33348
rect 13860 33292 13870 33348
rect 15250 33292 15260 33348
rect 15316 33292 15326 33348
rect 17042 33292 17052 33348
rect 17108 33292 18172 33348
rect 18228 33292 18238 33348
rect 21634 33292 21644 33348
rect 21700 33292 22092 33348
rect 22148 33292 22158 33348
rect 26562 33292 26572 33348
rect 26628 33292 26908 33348
rect 28466 33292 28476 33348
rect 28532 33292 32284 33348
rect 32340 33292 32350 33348
rect 32722 33292 32732 33348
rect 32788 33292 33740 33348
rect 33796 33292 33806 33348
rect 33954 33292 33964 33348
rect 34020 33292 34030 33348
rect 39890 33292 39900 33348
rect 39956 33292 40348 33348
rect 40404 33292 41356 33348
rect 41412 33292 41422 33348
rect 43250 33292 43260 33348
rect 43316 33292 44716 33348
rect 44772 33292 44782 33348
rect 32284 33236 32340 33292
rect 33964 33236 34020 33292
rect 3602 33180 3612 33236
rect 3668 33180 4732 33236
rect 4788 33180 4798 33236
rect 12898 33180 12908 33236
rect 12964 33180 14364 33236
rect 14420 33180 16044 33236
rect 16100 33180 16110 33236
rect 19618 33180 19628 33236
rect 19684 33180 22876 33236
rect 22932 33180 22942 33236
rect 23426 33180 23436 33236
rect 23492 33180 28364 33236
rect 28420 33180 29148 33236
rect 29204 33180 29214 33236
rect 32284 33180 34020 33236
rect 37538 33180 37548 33236
rect 37604 33180 39116 33236
rect 39172 33180 39182 33236
rect 40002 33180 40012 33236
rect 40068 33180 41020 33236
rect 41076 33180 41086 33236
rect 44930 33180 44940 33236
rect 44996 33180 45388 33236
rect 45444 33180 45612 33236
rect 45668 33180 45678 33236
rect 2594 33068 2604 33124
rect 2660 33068 3388 33124
rect 3444 33068 3454 33124
rect 6290 33068 6300 33124
rect 6356 33068 7084 33124
rect 7140 33068 7756 33124
rect 7812 33068 7822 33124
rect 9426 33068 9436 33124
rect 9492 33068 9660 33124
rect 9716 33068 9726 33124
rect 10770 33068 10780 33124
rect 10836 33068 11676 33124
rect 11732 33068 11742 33124
rect 14018 33068 14028 33124
rect 14084 33068 20524 33124
rect 20580 33068 20590 33124
rect 21298 33068 21308 33124
rect 21364 33068 23772 33124
rect 23828 33068 23838 33124
rect 44594 33068 44604 33124
rect 44660 33068 45276 33124
rect 45332 33068 46284 33124
rect 46340 33068 46350 33124
rect 19826 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20110 32956
rect 43148 32844 47852 32900
rect 47908 32844 47918 32900
rect 4050 32732 4060 32788
rect 4116 32732 4620 32788
rect 4676 32732 5068 32788
rect 5124 32732 5134 32788
rect 22306 32732 22316 32788
rect 22372 32732 22382 32788
rect 33730 32732 33740 32788
rect 33796 32732 35756 32788
rect 35812 32732 35822 32788
rect 10882 32620 10892 32676
rect 10948 32620 13132 32676
rect 13188 32620 13198 32676
rect 14690 32620 14700 32676
rect 14756 32620 17388 32676
rect 17444 32620 17454 32676
rect 3826 32508 3836 32564
rect 3892 32508 4732 32564
rect 4788 32508 4798 32564
rect 12002 32508 12012 32564
rect 12068 32508 15148 32564
rect 15204 32508 15214 32564
rect 22054 32508 22092 32564
rect 22148 32508 22158 32564
rect 22316 32452 22372 32732
rect 26786 32620 26796 32676
rect 26852 32620 29092 32676
rect 31826 32620 31836 32676
rect 31892 32620 31902 32676
rect 29036 32564 29092 32620
rect 31836 32564 31892 32620
rect 24546 32508 24556 32564
rect 24612 32508 26908 32564
rect 27682 32508 27692 32564
rect 27748 32508 28364 32564
rect 28420 32508 28430 32564
rect 29026 32508 29036 32564
rect 29092 32508 29102 32564
rect 31836 32508 32396 32564
rect 32452 32508 35532 32564
rect 35588 32508 35598 32564
rect 26852 32452 26908 32508
rect 4946 32396 4956 32452
rect 5012 32396 6412 32452
rect 6468 32396 6478 32452
rect 7746 32396 7756 32452
rect 7812 32396 9772 32452
rect 9828 32396 11004 32452
rect 11060 32396 11676 32452
rect 11732 32396 11742 32452
rect 13010 32396 13020 32452
rect 13076 32396 13916 32452
rect 13972 32396 13982 32452
rect 16482 32396 16492 32452
rect 16548 32396 17164 32452
rect 17220 32396 17230 32452
rect 20178 32396 20188 32452
rect 20244 32396 22988 32452
rect 23044 32396 23054 32452
rect 23986 32396 23996 32452
rect 24052 32396 24062 32452
rect 25330 32396 25340 32452
rect 25396 32396 26572 32452
rect 26628 32396 26638 32452
rect 26852 32396 29372 32452
rect 29428 32396 29438 32452
rect 33618 32396 33628 32452
rect 33684 32396 34076 32452
rect 34132 32396 34860 32452
rect 34916 32396 34926 32452
rect 23996 32340 24052 32396
rect 43148 32340 43204 32844
rect 49200 32788 50000 32816
rect 47618 32732 47628 32788
rect 47684 32732 48188 32788
rect 48244 32732 50000 32788
rect 49200 32704 50000 32732
rect 43474 32620 43484 32676
rect 43540 32620 44044 32676
rect 44100 32620 44940 32676
rect 44996 32620 45276 32676
rect 45332 32620 45342 32676
rect 46386 32620 46396 32676
rect 46452 32620 47404 32676
rect 47460 32620 47470 32676
rect 8418 32284 8428 32340
rect 8484 32284 13692 32340
rect 13748 32284 13758 32340
rect 18050 32284 18060 32340
rect 18116 32284 18620 32340
rect 18676 32284 18686 32340
rect 23996 32284 24220 32340
rect 24276 32284 25116 32340
rect 25172 32284 25182 32340
rect 33394 32284 33404 32340
rect 33460 32284 34524 32340
rect 34580 32284 34590 32340
rect 40002 32284 40012 32340
rect 40068 32284 43204 32340
rect 15474 32172 15484 32228
rect 15540 32172 15550 32228
rect 15698 32172 15708 32228
rect 15764 32172 16044 32228
rect 16100 32172 16110 32228
rect 36530 32172 36540 32228
rect 36596 32172 40124 32228
rect 40180 32172 40190 32228
rect 43586 32172 43596 32228
rect 43652 32172 44604 32228
rect 44660 32172 44670 32228
rect 4466 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4750 32172
rect 15484 32116 15540 32172
rect 35186 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35470 32172
rect 9426 32060 9436 32116
rect 9492 32060 9884 32116
rect 9940 32060 9950 32116
rect 15372 32060 15540 32116
rect 20738 32060 20748 32116
rect 20804 32060 21756 32116
rect 21812 32060 21822 32116
rect 44258 32060 44268 32116
rect 44324 32060 44334 32116
rect 15372 32004 15428 32060
rect 6402 31948 6412 32004
rect 6468 31948 7644 32004
rect 7700 31948 7710 32004
rect 8866 31948 8876 32004
rect 8932 31948 9436 32004
rect 9492 31948 9502 32004
rect 15362 31948 15372 32004
rect 15428 31948 15438 32004
rect 16034 31948 16044 32004
rect 16100 31948 18284 32004
rect 18340 31948 21196 32004
rect 21252 31948 21262 32004
rect 25442 31948 25452 32004
rect 25508 31948 26348 32004
rect 26404 31948 26414 32004
rect 32162 31948 32172 32004
rect 32228 31948 33180 32004
rect 33236 31948 33246 32004
rect 33506 31948 33516 32004
rect 33572 31948 35756 32004
rect 35812 31948 36652 32004
rect 36708 31948 36718 32004
rect 4274 31836 4284 31892
rect 4340 31836 4956 31892
rect 5012 31836 7308 31892
rect 7364 31836 7374 31892
rect 7970 31836 7980 31892
rect 8036 31836 9884 31892
rect 9940 31836 12068 31892
rect 12338 31836 12348 31892
rect 12404 31836 13580 31892
rect 13636 31836 13646 31892
rect 14354 31836 14364 31892
rect 14420 31836 15148 31892
rect 20402 31836 20412 31892
rect 20468 31836 21868 31892
rect 21924 31836 21934 31892
rect 23538 31836 23548 31892
rect 23604 31836 27468 31892
rect 27524 31836 29148 31892
rect 29204 31836 29214 31892
rect 39890 31836 39900 31892
rect 39956 31836 41468 31892
rect 41524 31836 41534 31892
rect 12012 31780 12068 31836
rect 13580 31780 13636 31836
rect 15092 31780 15148 31836
rect 44268 31780 44324 32060
rect 6178 31724 6188 31780
rect 6244 31724 7084 31780
rect 7140 31724 7532 31780
rect 7588 31724 7598 31780
rect 8306 31724 8316 31780
rect 8372 31724 11116 31780
rect 11172 31724 11182 31780
rect 12012 31724 13020 31780
rect 13076 31724 13356 31780
rect 13412 31724 13422 31780
rect 13580 31724 14588 31780
rect 14644 31724 14654 31780
rect 15092 31724 15932 31780
rect 15988 31724 16604 31780
rect 16660 31724 16670 31780
rect 17042 31724 17052 31780
rect 17108 31724 17500 31780
rect 17556 31724 17566 31780
rect 17938 31724 17948 31780
rect 18004 31724 18284 31780
rect 18340 31724 19068 31780
rect 19124 31724 19134 31780
rect 20626 31724 20636 31780
rect 20692 31724 21532 31780
rect 21588 31724 21598 31780
rect 21970 31724 21980 31780
rect 22036 31724 24332 31780
rect 24388 31724 24398 31780
rect 26786 31724 26796 31780
rect 26852 31724 27916 31780
rect 27972 31724 30940 31780
rect 30996 31724 31006 31780
rect 17948 31668 18004 31724
rect 8950 31612 8988 31668
rect 9044 31612 9054 31668
rect 9398 31612 9436 31668
rect 9492 31612 9502 31668
rect 14242 31612 14252 31668
rect 14308 31612 18004 31668
rect 20710 31612 20748 31668
rect 20804 31612 20814 31668
rect 20962 31612 20972 31668
rect 21028 31612 24444 31668
rect 24500 31612 24510 31668
rect 28018 31612 28028 31668
rect 28084 31612 28364 31668
rect 28420 31612 28430 31668
rect 35252 31556 35308 31780
rect 35364 31724 36092 31780
rect 36148 31724 39564 31780
rect 39620 31724 39630 31780
rect 41570 31724 41580 31780
rect 41636 31724 43372 31780
rect 43428 31724 44324 31780
rect 36978 31612 36988 31668
rect 37044 31612 37548 31668
rect 37604 31612 37614 31668
rect 42018 31612 42028 31668
rect 42084 31612 43820 31668
rect 43876 31612 43886 31668
rect 46050 31612 46060 31668
rect 46116 31612 46844 31668
rect 46900 31612 46910 31668
rect 11218 31500 11228 31556
rect 11284 31500 11900 31556
rect 11956 31500 11966 31556
rect 18722 31500 18732 31556
rect 18788 31500 21420 31556
rect 21476 31500 21486 31556
rect 29474 31500 29484 31556
rect 29540 31500 33964 31556
rect 34020 31500 34030 31556
rect 34962 31500 34972 31556
rect 35028 31500 35308 31556
rect 10658 31388 10668 31444
rect 10724 31388 13468 31444
rect 13524 31388 14924 31444
rect 14980 31388 14990 31444
rect 16594 31388 16604 31444
rect 16660 31388 17500 31444
rect 17556 31388 17566 31444
rect 31154 31388 31164 31444
rect 31220 31388 37436 31444
rect 37492 31388 37502 31444
rect 19826 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20110 31388
rect 4498 31276 4508 31332
rect 4564 31276 7980 31332
rect 8036 31276 8046 31332
rect 15026 31276 15036 31332
rect 15092 31276 17052 31332
rect 17108 31276 17118 31332
rect 30370 31276 30380 31332
rect 30436 31276 31388 31332
rect 31444 31276 34188 31332
rect 34244 31276 34254 31332
rect 4274 31164 4284 31220
rect 4340 31164 5180 31220
rect 5236 31164 8988 31220
rect 9044 31164 9054 31220
rect 11106 31164 11116 31220
rect 11172 31164 11788 31220
rect 11844 31164 11854 31220
rect 20626 31164 20636 31220
rect 20692 31164 21980 31220
rect 22036 31164 22764 31220
rect 22820 31164 22830 31220
rect 24658 31164 24668 31220
rect 24724 31164 29596 31220
rect 29652 31164 32508 31220
rect 32564 31164 32574 31220
rect 37202 31164 37212 31220
rect 37268 31164 38108 31220
rect 38164 31164 39004 31220
rect 39060 31164 39070 31220
rect 41794 31164 41804 31220
rect 41860 31164 42476 31220
rect 42532 31164 42542 31220
rect 44594 31164 44604 31220
rect 44660 31164 45164 31220
rect 45220 31164 45230 31220
rect 2706 31052 2716 31108
rect 2772 31052 3500 31108
rect 3556 31052 3566 31108
rect 4284 30996 4340 31164
rect 5730 31052 5740 31108
rect 5796 31052 24444 31108
rect 24500 31052 25228 31108
rect 25284 31052 25294 31108
rect 30594 31052 30604 31108
rect 30660 31052 32396 31108
rect 32452 31052 32462 31108
rect 33954 31052 33964 31108
rect 34020 31052 34636 31108
rect 34692 31052 34702 31108
rect 38322 31052 38332 31108
rect 38388 31052 39228 31108
rect 39284 31052 39294 31108
rect 42802 31052 42812 31108
rect 42868 31052 43260 31108
rect 43316 31052 43596 31108
rect 43652 31052 44828 31108
rect 44884 31052 44894 31108
rect 47170 31052 47180 31108
rect 47236 31052 47628 31108
rect 47684 31052 47694 31108
rect 1810 30940 1820 30996
rect 1876 30940 4340 30996
rect 10546 30940 10556 30996
rect 10612 30940 12796 30996
rect 12852 30940 12862 30996
rect 13682 30940 13692 30996
rect 13748 30940 17388 30996
rect 17444 30940 18060 30996
rect 18116 30940 18126 30996
rect 20514 30940 20524 30996
rect 20580 30940 23660 30996
rect 23716 30940 23726 30996
rect 38210 30940 38220 30996
rect 38276 30940 38668 30996
rect 38724 30940 38734 30996
rect 47058 30940 47068 30996
rect 47124 30940 47740 30996
rect 47796 30940 47806 30996
rect 2370 30828 2380 30884
rect 2436 30828 3276 30884
rect 3332 30772 3388 30884
rect 3490 30828 3500 30884
rect 3556 30828 4396 30884
rect 4452 30828 4462 30884
rect 12338 30828 12348 30884
rect 12404 30828 15148 30884
rect 15204 30828 16492 30884
rect 16548 30828 16558 30884
rect 18610 30828 18620 30884
rect 18676 30828 18732 30884
rect 18788 30828 18798 30884
rect 19618 30828 19628 30884
rect 19684 30828 25116 30884
rect 25172 30828 25182 30884
rect 33394 30828 33404 30884
rect 33460 30828 36540 30884
rect 36596 30828 36606 30884
rect 38612 30828 39564 30884
rect 39620 30828 39630 30884
rect 46386 30828 46396 30884
rect 46452 30828 47292 30884
rect 47348 30828 47358 30884
rect 38612 30772 38668 30828
rect 3332 30716 4508 30772
rect 4564 30716 4574 30772
rect 6962 30716 6972 30772
rect 7028 30716 8316 30772
rect 8372 30716 9212 30772
rect 9268 30716 9548 30772
rect 9604 30716 9614 30772
rect 28018 30716 28028 30772
rect 28084 30716 32396 30772
rect 32452 30716 32462 30772
rect 35410 30716 35420 30772
rect 35476 30716 35588 30772
rect 36082 30716 36092 30772
rect 36148 30716 38668 30772
rect 20850 30604 20860 30660
rect 20916 30604 27916 30660
rect 27972 30604 27982 30660
rect 4466 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4750 30604
rect 35186 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35470 30604
rect 35532 30548 35588 30716
rect 20066 30492 20076 30548
rect 20132 30492 24220 30548
rect 24276 30492 24286 30548
rect 35532 30492 44100 30548
rect 10770 30380 10780 30436
rect 10836 30380 12012 30436
rect 12068 30380 13580 30436
rect 13636 30380 13646 30436
rect 22978 30380 22988 30436
rect 23044 30380 23054 30436
rect 33506 30380 33516 30436
rect 33572 30380 35980 30436
rect 36036 30380 36046 30436
rect 37538 30380 37548 30436
rect 37604 30380 38108 30436
rect 38164 30380 38780 30436
rect 38836 30380 38846 30436
rect 4946 30268 4956 30324
rect 5012 30268 9212 30324
rect 9268 30268 9278 30324
rect 11106 30268 11116 30324
rect 11172 30268 12684 30324
rect 12740 30268 13804 30324
rect 13860 30268 13870 30324
rect 14690 30268 14700 30324
rect 14756 30268 16828 30324
rect 16884 30268 16894 30324
rect 22988 30212 23044 30380
rect 28242 30268 28252 30324
rect 28308 30268 29036 30324
rect 29092 30268 29102 30324
rect 31154 30268 31164 30324
rect 31220 30268 31500 30324
rect 31556 30268 31566 30324
rect 35746 30268 35756 30324
rect 35812 30268 37100 30324
rect 37156 30268 37166 30324
rect 8530 30156 8540 30212
rect 8596 30156 9436 30212
rect 9492 30156 9502 30212
rect 11442 30156 11452 30212
rect 11508 30156 12348 30212
rect 12404 30156 12414 30212
rect 13682 30156 13692 30212
rect 13748 30156 15484 30212
rect 15540 30156 15550 30212
rect 16034 30156 16044 30212
rect 16100 30156 17052 30212
rect 17108 30156 17118 30212
rect 19618 30156 19628 30212
rect 19684 30156 20412 30212
rect 20468 30156 20478 30212
rect 20738 30156 20748 30212
rect 20804 30156 21868 30212
rect 21924 30156 21934 30212
rect 22988 30156 24556 30212
rect 24612 30156 24622 30212
rect 28578 30156 28588 30212
rect 28644 30156 29820 30212
rect 29876 30156 29886 30212
rect 30482 30156 30492 30212
rect 30548 30156 31780 30212
rect 31938 30156 31948 30212
rect 32004 30156 32844 30212
rect 32900 30156 33964 30212
rect 34020 30156 34030 30212
rect 31724 30100 31780 30156
rect 44044 30100 44100 30492
rect 45378 30156 45388 30212
rect 45444 30156 46060 30212
rect 46116 30156 46126 30212
rect 8978 30044 8988 30100
rect 9044 30044 10108 30100
rect 10164 30044 10174 30100
rect 12450 30044 12460 30100
rect 12516 30044 14924 30100
rect 14980 30044 14990 30100
rect 19170 30044 19180 30100
rect 19236 30044 21420 30100
rect 21476 30044 21486 30100
rect 21746 30044 21756 30100
rect 21812 30044 22316 30100
rect 22372 30044 23884 30100
rect 23940 30044 23950 30100
rect 24210 30044 24220 30100
rect 24276 30044 25564 30100
rect 25620 30044 27076 30100
rect 27234 30044 27244 30100
rect 27300 30044 28476 30100
rect 28532 30044 31276 30100
rect 31332 30044 31342 30100
rect 31724 30044 32396 30100
rect 32452 30044 34524 30100
rect 34580 30044 34590 30100
rect 35074 30044 35084 30100
rect 35140 30044 35532 30100
rect 35588 30044 35598 30100
rect 44034 30044 44044 30100
rect 44100 30044 44110 30100
rect 27020 29988 27076 30044
rect 4834 29932 4844 29988
rect 4900 29932 7756 29988
rect 7812 29932 7822 29988
rect 9986 29932 9996 29988
rect 10052 29932 14588 29988
rect 14644 29932 15652 29988
rect 16818 29932 16828 29988
rect 16884 29932 26908 29988
rect 27020 29932 29708 29988
rect 29764 29932 29932 29988
rect 29988 29932 29998 29988
rect 31042 29932 31052 29988
rect 31108 29932 33628 29988
rect 33684 29932 33694 29988
rect 33954 29932 33964 29988
rect 34020 29932 36428 29988
rect 36484 29932 36494 29988
rect 41346 29932 41356 29988
rect 41412 29932 42252 29988
rect 42308 29932 45388 29988
rect 45444 29932 45454 29988
rect 45602 29932 45612 29988
rect 45668 29932 47180 29988
rect 47236 29932 47246 29988
rect 0 29876 800 29904
rect 0 29820 1708 29876
rect 1764 29820 1774 29876
rect 0 29792 800 29820
rect 15596 29764 15652 29932
rect 26852 29876 26908 29932
rect 26852 29820 33180 29876
rect 33236 29820 33246 29876
rect 19826 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20110 29820
rect 15586 29708 15596 29764
rect 15652 29708 15662 29764
rect 29138 29708 29148 29764
rect 29204 29708 29932 29764
rect 29988 29708 29998 29764
rect 32274 29708 32284 29764
rect 32340 29708 33516 29764
rect 33572 29708 33582 29764
rect 43026 29708 43036 29764
rect 43092 29708 43484 29764
rect 43540 29708 45724 29764
rect 45780 29708 45790 29764
rect 8726 29596 8764 29652
rect 8820 29596 8830 29652
rect 12562 29596 12572 29652
rect 12628 29596 14700 29652
rect 14756 29596 14766 29652
rect 16258 29596 16268 29652
rect 16324 29596 18396 29652
rect 18452 29596 19404 29652
rect 19460 29596 19740 29652
rect 19796 29596 19806 29652
rect 20738 29596 20748 29652
rect 20804 29596 22092 29652
rect 22148 29596 22158 29652
rect 28578 29596 28588 29652
rect 28644 29596 30380 29652
rect 30436 29596 30446 29652
rect 30716 29596 31052 29652
rect 31108 29596 31836 29652
rect 31892 29596 38668 29652
rect 30716 29540 30772 29596
rect 6850 29484 6860 29540
rect 6916 29484 7084 29540
rect 7140 29484 9660 29540
rect 9716 29484 10892 29540
rect 10948 29484 10958 29540
rect 23986 29484 23996 29540
rect 24052 29484 24780 29540
rect 24836 29484 29708 29540
rect 29764 29484 29774 29540
rect 30034 29484 30044 29540
rect 30100 29484 30772 29540
rect 31154 29484 31164 29540
rect 31220 29484 32956 29540
rect 33012 29484 33022 29540
rect 33842 29484 33852 29540
rect 33908 29484 34524 29540
rect 34580 29484 34590 29540
rect 38612 29428 38668 29596
rect 14130 29372 14140 29428
rect 14196 29372 16044 29428
rect 16100 29372 16110 29428
rect 17378 29372 17388 29428
rect 17444 29372 17454 29428
rect 26786 29372 26796 29428
rect 26852 29372 27580 29428
rect 27636 29372 29372 29428
rect 29428 29372 29438 29428
rect 30156 29372 30940 29428
rect 30996 29372 32508 29428
rect 32564 29372 33292 29428
rect 33348 29372 33740 29428
rect 33796 29372 33806 29428
rect 34066 29372 34076 29428
rect 34132 29372 34748 29428
rect 34804 29372 34814 29428
rect 38612 29372 39228 29428
rect 39284 29372 39294 29428
rect 17388 29316 17444 29372
rect 30156 29316 30212 29372
rect 5954 29260 5964 29316
rect 6020 29260 8428 29316
rect 8484 29260 11116 29316
rect 11172 29260 13916 29316
rect 13972 29260 13982 29316
rect 14914 29260 14924 29316
rect 14980 29260 17444 29316
rect 24546 29260 24556 29316
rect 24612 29260 26012 29316
rect 26068 29260 26078 29316
rect 26852 29260 30212 29316
rect 30370 29260 30380 29316
rect 30436 29260 31500 29316
rect 31556 29260 31566 29316
rect 42354 29260 42364 29316
rect 42420 29260 42924 29316
rect 42980 29260 42990 29316
rect 26852 29204 26908 29260
rect 5170 29148 5180 29204
rect 5236 29148 10332 29204
rect 10388 29148 11228 29204
rect 11284 29148 11294 29204
rect 20626 29148 20636 29204
rect 20692 29148 21420 29204
rect 21476 29148 26908 29204
rect 27906 29148 27916 29204
rect 27972 29148 29148 29204
rect 29204 29148 29214 29204
rect 30930 29148 30940 29204
rect 30996 29148 31948 29204
rect 32004 29148 32014 29204
rect 7746 29036 7756 29092
rect 7812 29036 11004 29092
rect 11060 29036 14476 29092
rect 14532 29036 14542 29092
rect 20290 29036 20300 29092
rect 20356 29036 21644 29092
rect 21700 29036 21710 29092
rect 32050 29036 32060 29092
rect 32116 29036 33404 29092
rect 33460 29036 33470 29092
rect 4466 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4750 29036
rect 35186 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35470 29036
rect 10098 28924 10108 28980
rect 10164 28924 12236 28980
rect 12292 28924 12302 28980
rect 30146 28924 30156 28980
rect 30212 28924 32956 28980
rect 33012 28924 33022 28980
rect 4498 28812 4508 28868
rect 4564 28812 8428 28868
rect 8484 28812 8494 28868
rect 9510 28812 9548 28868
rect 9604 28812 9614 28868
rect 10882 28812 10892 28868
rect 10948 28812 18172 28868
rect 18228 28812 18238 28868
rect 21746 28812 21756 28868
rect 21812 28812 23436 28868
rect 23492 28812 23502 28868
rect 33506 28812 33516 28868
rect 33572 28812 35644 28868
rect 35700 28812 35710 28868
rect 6748 28700 10108 28756
rect 10164 28700 10174 28756
rect 12562 28700 12572 28756
rect 12628 28700 12908 28756
rect 12964 28700 14140 28756
rect 14196 28700 14206 28756
rect 16370 28700 16380 28756
rect 16436 28700 17836 28756
rect 17892 28700 17902 28756
rect 19842 28700 19852 28756
rect 19908 28700 21756 28756
rect 21812 28700 21822 28756
rect 22978 28700 22988 28756
rect 23044 28700 23548 28756
rect 23604 28700 23614 28756
rect 24098 28700 24108 28756
rect 24164 28700 27132 28756
rect 27188 28700 30380 28756
rect 30436 28700 30446 28756
rect 34178 28700 34188 28756
rect 34244 28700 35420 28756
rect 35476 28700 35486 28756
rect 6748 28644 6804 28700
rect 4610 28588 4620 28644
rect 4676 28588 6748 28644
rect 6804 28588 6814 28644
rect 6962 28588 6972 28644
rect 7028 28588 7308 28644
rect 7364 28588 9772 28644
rect 9828 28588 10556 28644
rect 10612 28588 10622 28644
rect 16258 28588 16268 28644
rect 16324 28588 17052 28644
rect 17108 28588 18396 28644
rect 18452 28588 18462 28644
rect 23762 28588 23772 28644
rect 23828 28588 25564 28644
rect 25620 28588 27804 28644
rect 27860 28588 27870 28644
rect 29362 28588 29372 28644
rect 29428 28588 30604 28644
rect 30660 28588 30670 28644
rect 42578 28588 42588 28644
rect 42644 28588 43484 28644
rect 43540 28588 43550 28644
rect 7858 28476 7868 28532
rect 7924 28476 11340 28532
rect 11396 28476 12012 28532
rect 12068 28476 12078 28532
rect 12786 28476 12796 28532
rect 12852 28476 17388 28532
rect 17444 28476 17454 28532
rect 27906 28476 27916 28532
rect 27972 28476 30156 28532
rect 30212 28476 30222 28532
rect 39890 28476 39900 28532
rect 39956 28476 40908 28532
rect 40964 28476 40974 28532
rect 42914 28476 42924 28532
rect 42980 28476 43596 28532
rect 43652 28476 44604 28532
rect 44660 28476 44670 28532
rect 9650 28364 9660 28420
rect 9716 28364 10444 28420
rect 10500 28364 10510 28420
rect 11414 28364 11452 28420
rect 11508 28364 11518 28420
rect 12226 28364 12236 28420
rect 12292 28364 14700 28420
rect 14756 28364 18956 28420
rect 19012 28364 19022 28420
rect 22306 28364 22316 28420
rect 22372 28364 23660 28420
rect 23716 28364 23726 28420
rect 24658 28364 24668 28420
rect 24724 28364 27412 28420
rect 46386 28364 46396 28420
rect 46452 28364 47180 28420
rect 47236 28364 47246 28420
rect 27356 28308 27412 28364
rect 27346 28252 27356 28308
rect 27412 28252 28812 28308
rect 28868 28252 33068 28308
rect 33124 28252 33134 28308
rect 34934 28252 34972 28308
rect 35028 28252 35038 28308
rect 19826 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20110 28252
rect 23314 28140 23324 28196
rect 23380 28140 24332 28196
rect 24388 28140 31276 28196
rect 31332 28140 31342 28196
rect 34066 28140 34076 28196
rect 34132 28140 35644 28196
rect 35700 28140 35710 28196
rect 18610 28028 18620 28084
rect 18676 28028 19180 28084
rect 19236 28028 19246 28084
rect 22754 28028 22764 28084
rect 22820 28028 25900 28084
rect 25956 28028 25966 28084
rect 26852 28028 27468 28084
rect 27524 28028 27692 28084
rect 27748 28028 27758 28084
rect 30146 28028 30156 28084
rect 30212 28028 35532 28084
rect 35588 28028 35598 28084
rect 26852 27972 26908 28028
rect 4274 27916 4284 27972
rect 4340 27916 9436 27972
rect 9492 27916 9502 27972
rect 23314 27916 23324 27972
rect 23380 27916 26908 27972
rect 27794 27916 27804 27972
rect 27860 27916 31836 27972
rect 31892 27916 33628 27972
rect 33684 27916 34412 27972
rect 34468 27916 34478 27972
rect 42130 27916 42140 27972
rect 42196 27916 42476 27972
rect 42532 27916 42812 27972
rect 42868 27916 42878 27972
rect 5170 27804 5180 27860
rect 5236 27804 9772 27860
rect 9828 27804 9838 27860
rect 26114 27804 26124 27860
rect 26180 27804 27916 27860
rect 27972 27804 27982 27860
rect 28354 27804 28364 27860
rect 28420 27804 29708 27860
rect 29764 27804 30716 27860
rect 30772 27804 30782 27860
rect 32498 27804 32508 27860
rect 32564 27804 34468 27860
rect 34412 27748 34468 27804
rect 9874 27692 9884 27748
rect 9940 27692 11788 27748
rect 11844 27692 11854 27748
rect 16034 27692 16044 27748
rect 16100 27692 17724 27748
rect 17780 27692 17790 27748
rect 26226 27692 26236 27748
rect 26292 27692 28476 27748
rect 28532 27692 28542 27748
rect 29026 27692 29036 27748
rect 29092 27692 31164 27748
rect 31220 27692 33180 27748
rect 33236 27692 33246 27748
rect 34402 27692 34412 27748
rect 34468 27692 37996 27748
rect 38052 27692 38062 27748
rect 39554 27692 39564 27748
rect 39620 27692 41356 27748
rect 41412 27692 43596 27748
rect 43652 27692 44268 27748
rect 44324 27692 44334 27748
rect 45266 27692 45276 27748
rect 45332 27692 46508 27748
rect 46564 27692 46574 27748
rect 2258 27580 2268 27636
rect 2324 27580 10892 27636
rect 10948 27580 15148 27636
rect 18694 27580 18732 27636
rect 18788 27580 18798 27636
rect 26852 27580 32508 27636
rect 32564 27580 32574 27636
rect 33282 27580 33292 27636
rect 33348 27580 34748 27636
rect 34804 27580 34814 27636
rect 35074 27580 35084 27636
rect 35140 27580 35868 27636
rect 35924 27580 35934 27636
rect 15092 27524 15148 27580
rect 26852 27524 26908 27580
rect 15092 27468 16492 27524
rect 16548 27468 26908 27524
rect 4466 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4750 27468
rect 35186 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35470 27468
rect 19170 27356 19180 27412
rect 19236 27356 19516 27412
rect 19572 27356 19582 27412
rect 32162 27356 32172 27412
rect 32228 27356 32956 27412
rect 33012 27356 33022 27412
rect 12114 27244 12124 27300
rect 12180 27244 13804 27300
rect 13860 27244 13870 27300
rect 16146 27244 16156 27300
rect 16212 27244 16492 27300
rect 16548 27244 16558 27300
rect 16818 27244 16828 27300
rect 16884 27244 18620 27300
rect 18676 27244 29372 27300
rect 29428 27244 29438 27300
rect 34626 27244 34636 27300
rect 34692 27244 35196 27300
rect 35252 27244 35262 27300
rect 8642 27132 8652 27188
rect 8708 27132 15708 27188
rect 15764 27132 18172 27188
rect 18228 27132 18238 27188
rect 24322 27132 24332 27188
rect 24388 27132 25340 27188
rect 25396 27132 25406 27188
rect 26852 27132 31276 27188
rect 31332 27132 37492 27188
rect 40226 27132 40236 27188
rect 40292 27132 41020 27188
rect 41076 27132 41086 27188
rect 26852 27076 26908 27132
rect 16034 27020 16044 27076
rect 16100 27020 16110 27076
rect 18396 27020 18956 27076
rect 19012 27020 20188 27076
rect 20244 27020 20254 27076
rect 26114 27020 26124 27076
rect 26180 27020 26908 27076
rect 28466 27020 28476 27076
rect 28532 27020 29148 27076
rect 29204 27020 29214 27076
rect 35186 27020 35196 27076
rect 35252 27020 36988 27076
rect 37044 27020 37054 27076
rect 9426 26908 9436 26964
rect 9492 26908 9996 26964
rect 10052 26908 10062 26964
rect 13906 26908 13916 26964
rect 13972 26908 15820 26964
rect 15876 26908 15886 26964
rect 5506 26796 5516 26852
rect 5572 26796 6300 26852
rect 6356 26796 6366 26852
rect 6850 26796 6860 26852
rect 6916 26796 7084 26852
rect 7140 26796 7150 26852
rect 16044 26740 16100 27020
rect 18396 26908 18452 27020
rect 19030 26908 19068 26964
rect 19124 26908 19134 26964
rect 23874 26908 23884 26964
rect 23940 26908 25788 26964
rect 25844 26908 26796 26964
rect 26852 26908 26862 26964
rect 36082 26908 36092 26964
rect 36148 26908 36876 26964
rect 36932 26908 37268 26964
rect 18386 26852 18396 26908
rect 18452 26852 18462 26908
rect 37212 26852 37268 26908
rect 19506 26796 19516 26852
rect 19572 26796 20300 26852
rect 20356 26796 20366 26852
rect 21858 26796 21868 26852
rect 21924 26796 26684 26852
rect 26740 26796 26750 26852
rect 35522 26796 35532 26852
rect 35588 26796 35756 26852
rect 35812 26796 35822 26852
rect 36418 26796 36428 26852
rect 36484 26796 36988 26852
rect 37044 26796 37054 26852
rect 37202 26796 37212 26852
rect 37268 26796 37278 26852
rect 37436 26740 37492 27132
rect 44930 27020 44940 27076
rect 44996 27020 46284 27076
rect 46340 27020 47740 27076
rect 47796 27020 47806 27076
rect 49200 26964 50000 26992
rect 37986 26908 37996 26964
rect 38052 26908 40348 26964
rect 40404 26908 40414 26964
rect 45938 26908 45948 26964
rect 46004 26908 47852 26964
rect 47908 26908 47918 26964
rect 48290 26908 48300 26964
rect 48356 26908 50000 26964
rect 49200 26880 50000 26908
rect 41906 26796 41916 26852
rect 41972 26796 43148 26852
rect 43204 26796 43214 26852
rect 15586 26684 15596 26740
rect 15652 26684 16100 26740
rect 19030 26684 19068 26740
rect 19124 26684 19134 26740
rect 20178 26684 20188 26740
rect 20244 26684 25228 26740
rect 25284 26684 25294 26740
rect 28578 26684 28588 26740
rect 28644 26684 32228 26740
rect 37436 26684 41244 26740
rect 41300 26684 41310 26740
rect 19826 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20110 26684
rect 32172 26628 32228 26684
rect 7186 26572 7196 26628
rect 7252 26572 8652 26628
rect 8708 26572 8718 26628
rect 26562 26572 26572 26628
rect 26628 26572 27132 26628
rect 27188 26572 30492 26628
rect 30548 26572 30558 26628
rect 32162 26572 32172 26628
rect 32228 26572 38220 26628
rect 38276 26572 38286 26628
rect 10098 26460 10108 26516
rect 10164 26460 11676 26516
rect 11732 26460 14924 26516
rect 14980 26460 14990 26516
rect 15922 26460 15932 26516
rect 15988 26460 17388 26516
rect 17444 26460 17454 26516
rect 17910 26460 17948 26516
rect 18004 26460 18014 26516
rect 20290 26460 20300 26516
rect 20356 26460 21196 26516
rect 21252 26460 21262 26516
rect 21970 26460 21980 26516
rect 22036 26460 23548 26516
rect 23604 26460 23614 26516
rect 26002 26460 26012 26516
rect 26068 26460 33852 26516
rect 33908 26460 33918 26516
rect 37426 26460 37436 26516
rect 37492 26460 37996 26516
rect 38052 26460 38892 26516
rect 38948 26460 38958 26516
rect 41122 26460 41132 26516
rect 41188 26460 42364 26516
rect 42420 26460 42924 26516
rect 42980 26460 42990 26516
rect 12898 26348 12908 26404
rect 12964 26348 14252 26404
rect 14308 26348 14318 26404
rect 18582 26348 18620 26404
rect 18676 26348 18686 26404
rect 18946 26348 18956 26404
rect 19012 26348 20524 26404
rect 20580 26348 20860 26404
rect 20916 26348 20926 26404
rect 25554 26348 25564 26404
rect 25620 26348 28700 26404
rect 28756 26348 28766 26404
rect 32498 26348 32508 26404
rect 32564 26348 39340 26404
rect 39396 26348 39406 26404
rect 5954 26236 5964 26292
rect 6020 26236 8764 26292
rect 8820 26236 8830 26292
rect 13122 26236 13132 26292
rect 13188 26236 14700 26292
rect 14756 26236 15372 26292
rect 15428 26236 16268 26292
rect 16324 26236 16334 26292
rect 20300 26236 22204 26292
rect 22260 26236 22270 26292
rect 29250 26236 29260 26292
rect 29316 26236 30716 26292
rect 30772 26236 32620 26292
rect 32676 26236 33180 26292
rect 33236 26236 33246 26292
rect 20300 26180 20356 26236
rect 4834 26124 4844 26180
rect 4900 26124 6412 26180
rect 6468 26124 7420 26180
rect 7476 26124 7486 26180
rect 14354 26124 14364 26180
rect 14420 26124 16156 26180
rect 16212 26124 16222 26180
rect 20290 26124 20300 26180
rect 20356 26124 20366 26180
rect 21410 26124 21420 26180
rect 21476 26124 24668 26180
rect 24724 26124 24734 26180
rect 24882 26124 24892 26180
rect 24948 26124 27916 26180
rect 27972 26124 27982 26180
rect 32620 26124 45052 26180
rect 45108 26124 45118 26180
rect 14802 26012 14812 26068
rect 14868 26012 15820 26068
rect 15876 26012 15886 26068
rect 16258 26012 16268 26068
rect 16324 26012 16604 26068
rect 16660 26012 17388 26068
rect 17444 26012 17454 26068
rect 19730 26012 19740 26068
rect 19796 26012 20860 26068
rect 20916 26012 20926 26068
rect 30034 26012 30044 26068
rect 30100 26012 32396 26068
rect 32452 26012 32462 26068
rect 32620 25956 32676 26124
rect 34738 26012 34748 26068
rect 34804 26012 34972 26068
rect 35028 26012 35038 26068
rect 23202 25900 23212 25956
rect 23268 25900 32676 25956
rect 40338 25900 40348 25956
rect 40404 25900 41132 25956
rect 41188 25900 41198 25956
rect 4466 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4750 25900
rect 35186 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35470 25900
rect 15138 25788 15148 25844
rect 15204 25788 26012 25844
rect 26068 25788 26078 25844
rect 26786 25788 26796 25844
rect 26852 25620 26908 25844
rect 31602 25676 31612 25732
rect 31668 25676 33628 25732
rect 33684 25676 36764 25732
rect 36820 25676 36830 25732
rect 4722 25564 4732 25620
rect 4788 25564 4956 25620
rect 5012 25564 8428 25620
rect 8484 25564 8494 25620
rect 20188 25564 21980 25620
rect 22036 25564 22652 25620
rect 22708 25564 22718 25620
rect 25666 25564 25676 25620
rect 25732 25564 27468 25620
rect 27524 25564 27534 25620
rect 33170 25564 33180 25620
rect 33236 25564 34076 25620
rect 34132 25564 34142 25620
rect 35942 25564 35980 25620
rect 36036 25564 36046 25620
rect 20188 25508 20244 25564
rect 6738 25452 6748 25508
rect 6804 25452 8092 25508
rect 8148 25452 11788 25508
rect 11844 25452 11854 25508
rect 13682 25452 13692 25508
rect 13748 25452 18620 25508
rect 18676 25452 18686 25508
rect 19058 25452 19068 25508
rect 19124 25452 19134 25508
rect 19292 25452 20188 25508
rect 20244 25452 20254 25508
rect 21186 25452 21196 25508
rect 21252 25452 23212 25508
rect 23268 25452 24892 25508
rect 24948 25452 24958 25508
rect 35522 25452 35532 25508
rect 35588 25452 36988 25508
rect 37044 25452 37054 25508
rect 39442 25452 39452 25508
rect 39508 25452 41356 25508
rect 41412 25452 41916 25508
rect 41972 25452 43036 25508
rect 43092 25452 43102 25508
rect 43362 25452 43372 25508
rect 43428 25452 43708 25508
rect 43764 25452 43774 25508
rect 19068 25396 19124 25452
rect 19292 25396 19348 25452
rect 5058 25340 5068 25396
rect 5124 25340 6860 25396
rect 6916 25340 6926 25396
rect 18722 25340 18732 25396
rect 18788 25340 19124 25396
rect 19282 25340 19292 25396
rect 19348 25340 19358 25396
rect 19954 25340 19964 25396
rect 20020 25340 20412 25396
rect 20468 25340 20478 25396
rect 21858 25340 21868 25396
rect 21924 25340 23548 25396
rect 23604 25340 23614 25396
rect 24546 25340 24556 25396
rect 24612 25340 27020 25396
rect 27076 25340 27086 25396
rect 34514 25340 34524 25396
rect 34580 25340 36428 25396
rect 36484 25340 36494 25396
rect 5394 25228 5404 25284
rect 5460 25228 5964 25284
rect 6020 25228 6030 25284
rect 9762 25228 9772 25284
rect 9828 25228 10444 25284
rect 10500 25228 13804 25284
rect 13860 25228 13870 25284
rect 14326 25228 14364 25284
rect 14420 25228 14430 25284
rect 15138 25228 15148 25284
rect 15204 25228 15708 25284
rect 15764 25228 15774 25284
rect 18162 25228 18172 25284
rect 18228 25228 20076 25284
rect 20132 25228 20142 25284
rect 23090 25228 23100 25284
rect 23156 25228 24780 25284
rect 24836 25228 24846 25284
rect 35868 25228 37212 25284
rect 37268 25228 37278 25284
rect 35868 25172 35924 25228
rect 16146 25116 16156 25172
rect 16212 25116 19404 25172
rect 19460 25116 19470 25172
rect 21634 25116 21644 25172
rect 21700 25116 22652 25172
rect 22708 25116 22988 25172
rect 23044 25116 23054 25172
rect 23426 25116 23436 25172
rect 23492 25116 25788 25172
rect 25844 25116 26796 25172
rect 26852 25116 26862 25172
rect 35858 25116 35868 25172
rect 35924 25116 35934 25172
rect 36866 25116 36876 25172
rect 36932 25116 36942 25172
rect 45042 25116 45052 25172
rect 45108 25116 45388 25172
rect 45444 25116 45454 25172
rect 19826 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20110 25116
rect 36876 25060 36932 25116
rect 17714 25004 17724 25060
rect 17780 25004 19516 25060
rect 19572 25004 19582 25060
rect 34850 25004 34860 25060
rect 34916 25004 36932 25060
rect 18834 24892 18844 24948
rect 18900 24892 21420 24948
rect 21476 24892 21756 24948
rect 21812 24892 21822 24948
rect 27682 24892 27692 24948
rect 27748 24892 28588 24948
rect 28644 24892 28654 24948
rect 43922 24892 43932 24948
rect 43988 24892 44828 24948
rect 44884 24892 44894 24948
rect 45154 24892 45164 24948
rect 45220 24892 46284 24948
rect 46340 24892 47572 24948
rect 15922 24780 15932 24836
rect 15988 24780 16716 24836
rect 16772 24780 20524 24836
rect 20580 24780 20590 24836
rect 22754 24780 22764 24836
rect 22820 24780 23884 24836
rect 23940 24780 24444 24836
rect 24500 24780 24510 24836
rect 45042 24780 45052 24836
rect 45108 24780 45612 24836
rect 45668 24780 45678 24836
rect 47516 24724 47572 24892
rect 18610 24668 18620 24724
rect 18676 24668 18956 24724
rect 19012 24668 19022 24724
rect 20066 24668 20076 24724
rect 20132 24668 21308 24724
rect 21364 24668 21374 24724
rect 24546 24668 24556 24724
rect 24612 24668 26124 24724
rect 26180 24668 29036 24724
rect 29092 24668 29102 24724
rect 29586 24668 29596 24724
rect 29652 24668 30492 24724
rect 30548 24668 30558 24724
rect 44594 24668 44604 24724
rect 44660 24668 45276 24724
rect 45332 24668 45724 24724
rect 45780 24668 46732 24724
rect 46788 24668 46798 24724
rect 47506 24668 47516 24724
rect 47572 24668 47582 24724
rect 18956 24612 19012 24668
rect 3154 24556 3164 24612
rect 3220 24556 3388 24612
rect 13794 24556 13804 24612
rect 13860 24556 14700 24612
rect 14756 24556 14766 24612
rect 18956 24556 20972 24612
rect 21028 24556 21038 24612
rect 29250 24556 29260 24612
rect 29316 24556 29708 24612
rect 29764 24556 32396 24612
rect 32452 24556 32462 24612
rect 35970 24556 35980 24612
rect 36036 24556 36316 24612
rect 36372 24556 36382 24612
rect 39218 24556 39228 24612
rect 39284 24556 39676 24612
rect 39732 24556 41580 24612
rect 41636 24556 41646 24612
rect 45378 24556 45388 24612
rect 45444 24556 46172 24612
rect 46228 24556 48300 24612
rect 48356 24556 48366 24612
rect 3332 24500 3388 24556
rect 3332 24444 4508 24500
rect 4564 24444 5852 24500
rect 5908 24444 5918 24500
rect 19506 24332 19516 24388
rect 19572 24332 23996 24388
rect 24052 24332 24062 24388
rect 4466 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4750 24332
rect 35186 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35470 24332
rect 6850 24220 6860 24276
rect 6916 24220 7196 24276
rect 7252 24220 7262 24276
rect 13682 24220 13692 24276
rect 13748 24220 15148 24276
rect 18274 24220 18284 24276
rect 18340 24220 20860 24276
rect 20916 24220 20926 24276
rect 22306 24220 22316 24276
rect 22372 24220 23212 24276
rect 23268 24220 30940 24276
rect 30996 24220 31006 24276
rect 12786 24108 12796 24164
rect 12852 24108 14924 24164
rect 14980 24108 14990 24164
rect 15092 24108 15148 24220
rect 15204 24108 28476 24164
rect 28532 24108 29708 24164
rect 29764 24108 29774 24164
rect 10994 23996 11004 24052
rect 11060 23996 11340 24052
rect 11396 23996 12404 24052
rect 18946 23996 18956 24052
rect 19012 23996 19516 24052
rect 19572 23996 19582 24052
rect 20178 23996 20188 24052
rect 20244 23996 21644 24052
rect 21700 23996 28140 24052
rect 28196 23996 31276 24052
rect 31332 23996 31836 24052
rect 31892 23996 31902 24052
rect 12348 23940 12404 23996
rect 4274 23884 4284 23940
rect 4340 23884 8428 23940
rect 8484 23884 8494 23940
rect 8642 23884 8652 23940
rect 8708 23884 10220 23940
rect 10276 23884 12124 23940
rect 12180 23884 12190 23940
rect 12338 23884 12348 23940
rect 12404 23884 14028 23940
rect 14084 23884 14094 23940
rect 14914 23884 14924 23940
rect 14980 23884 15484 23940
rect 15540 23884 15550 23940
rect 17938 23884 17948 23940
rect 18004 23884 20300 23940
rect 20356 23884 20366 23940
rect 23314 23884 23324 23940
rect 23380 23884 23390 23940
rect 31602 23884 31612 23940
rect 31668 23884 32284 23940
rect 32340 23884 33068 23940
rect 33124 23884 33134 23940
rect 34626 23884 34636 23940
rect 34692 23884 36092 23940
rect 36148 23884 36158 23940
rect 23324 23828 23380 23884
rect 6514 23772 6524 23828
rect 6580 23772 9044 23828
rect 14130 23772 14140 23828
rect 14196 23772 18284 23828
rect 18340 23772 18350 23828
rect 19506 23772 19516 23828
rect 19572 23772 20636 23828
rect 20692 23772 20702 23828
rect 22866 23772 22876 23828
rect 22932 23772 23380 23828
rect 24546 23772 24556 23828
rect 24612 23772 25676 23828
rect 25732 23772 25742 23828
rect 30930 23772 30940 23828
rect 30996 23772 32060 23828
rect 32116 23772 32126 23828
rect 35186 23772 35196 23828
rect 35252 23772 38556 23828
rect 38612 23772 38622 23828
rect 45602 23772 45612 23828
rect 45668 23772 46956 23828
rect 47012 23772 47022 23828
rect 8988 23604 9044 23772
rect 9314 23660 9324 23716
rect 9380 23660 13580 23716
rect 13636 23660 13646 23716
rect 17602 23660 17612 23716
rect 17668 23660 19964 23716
rect 20020 23660 20030 23716
rect 21522 23660 21532 23716
rect 21588 23660 22204 23716
rect 22260 23660 23436 23716
rect 23492 23660 23502 23716
rect 25442 23660 25452 23716
rect 25508 23660 28140 23716
rect 28196 23660 30828 23716
rect 30884 23660 33516 23716
rect 33572 23660 33582 23716
rect 5282 23548 5292 23604
rect 5348 23548 8484 23604
rect 8978 23548 8988 23604
rect 9044 23548 11452 23604
rect 11508 23548 11518 23604
rect 12674 23548 12684 23604
rect 12740 23548 12750 23604
rect 16706 23548 16716 23604
rect 16772 23548 17836 23604
rect 17892 23548 17902 23604
rect 22306 23548 22316 23604
rect 22372 23548 22764 23604
rect 22820 23548 23100 23604
rect 23156 23548 23166 23604
rect 24210 23548 24220 23604
rect 24276 23548 25340 23604
rect 25396 23548 25406 23604
rect 34962 23548 34972 23604
rect 35028 23548 35532 23604
rect 35588 23548 35598 23604
rect 8428 23492 8484 23548
rect 12684 23492 12740 23548
rect 19826 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20110 23548
rect 8428 23436 11788 23492
rect 11844 23436 11854 23492
rect 12684 23436 14924 23492
rect 14980 23436 14990 23492
rect 23174 23436 23212 23492
rect 23268 23436 23278 23492
rect 36306 23436 36316 23492
rect 36372 23436 37436 23492
rect 37492 23436 37502 23492
rect 44930 23436 44940 23492
rect 44996 23436 47740 23492
rect 47796 23436 47806 23492
rect 5954 23324 5964 23380
rect 6020 23324 8316 23380
rect 8372 23324 12124 23380
rect 12180 23324 12796 23380
rect 12852 23324 15036 23380
rect 15092 23324 15102 23380
rect 18386 23324 18396 23380
rect 18452 23324 19068 23380
rect 19124 23324 19134 23380
rect 26226 23324 26236 23380
rect 26292 23324 27916 23380
rect 27972 23324 27982 23380
rect 38612 23324 39564 23380
rect 39620 23324 39630 23380
rect 43698 23324 43708 23380
rect 43764 23324 45164 23380
rect 45220 23324 46620 23380
rect 46676 23324 48076 23380
rect 48132 23324 48142 23380
rect 12226 23212 12236 23268
rect 12292 23212 17612 23268
rect 17668 23212 17678 23268
rect 17836 23212 38556 23268
rect 38612 23212 38668 23324
rect 44706 23212 44716 23268
rect 44772 23212 46172 23268
rect 46228 23212 46238 23268
rect 17836 23156 17892 23212
rect 11218 23100 11228 23156
rect 11284 23100 12572 23156
rect 12628 23100 12638 23156
rect 13234 23100 13244 23156
rect 13300 23100 13468 23156
rect 13524 23100 13534 23156
rect 16146 23100 16156 23156
rect 16212 23100 17892 23156
rect 19058 23100 19068 23156
rect 19124 23100 19740 23156
rect 19796 23100 19806 23156
rect 21298 23100 21308 23156
rect 21364 23100 21868 23156
rect 21924 23100 21934 23156
rect 46834 23100 46844 23156
rect 46900 23100 47404 23156
rect 47460 23100 47470 23156
rect 3490 22988 3500 23044
rect 3556 22988 4956 23044
rect 5012 22988 7532 23044
rect 7588 22988 8316 23044
rect 8372 22988 8382 23044
rect 9986 22988 9996 23044
rect 10052 22988 12684 23044
rect 12740 22988 12750 23044
rect 18050 22988 18060 23044
rect 18116 22988 21980 23044
rect 22036 22988 22046 23044
rect 25330 22988 25340 23044
rect 25396 22988 27804 23044
rect 27860 22988 28140 23044
rect 28196 22988 28206 23044
rect 29026 22988 29036 23044
rect 29092 22988 29484 23044
rect 29540 22988 29550 23044
rect 30146 22988 30156 23044
rect 30212 22988 30604 23044
rect 30660 22988 31164 23044
rect 31220 22988 31230 23044
rect 40898 22988 40908 23044
rect 40964 22988 41580 23044
rect 41636 22988 43148 23044
rect 43204 22988 44268 23044
rect 44324 22988 44940 23044
rect 44996 22988 45006 23044
rect 8866 22876 8876 22932
rect 8932 22876 11676 22932
rect 11732 22876 14364 22932
rect 14420 22876 14430 22932
rect 18162 22876 18172 22932
rect 18228 22876 20524 22932
rect 20580 22876 20590 22932
rect 25218 22876 25228 22932
rect 25284 22876 40012 22932
rect 40068 22876 40078 22932
rect 16818 22764 16828 22820
rect 16884 22764 17724 22820
rect 17780 22764 18508 22820
rect 18564 22764 18574 22820
rect 4466 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4750 22764
rect 35186 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35470 22764
rect 15922 22652 15932 22708
rect 15988 22652 25452 22708
rect 25508 22652 25518 22708
rect 34822 22652 34860 22708
rect 34916 22652 34926 22708
rect 35830 22652 35868 22708
rect 35924 22652 35934 22708
rect 40450 22652 40460 22708
rect 40516 22652 40526 22708
rect 11106 22540 11116 22596
rect 11172 22540 13916 22596
rect 13972 22540 13982 22596
rect 17602 22540 17612 22596
rect 17668 22540 18844 22596
rect 18900 22540 28028 22596
rect 28084 22540 28094 22596
rect 28578 22540 28588 22596
rect 28644 22540 29372 22596
rect 29428 22540 38668 22596
rect 28028 22484 28084 22540
rect 38612 22484 38668 22540
rect 40460 22484 40516 22652
rect 12898 22428 12908 22484
rect 12964 22428 20244 22484
rect 20850 22428 20860 22484
rect 20916 22428 25900 22484
rect 25956 22428 25966 22484
rect 28028 22428 29148 22484
rect 29204 22428 29214 22484
rect 34188 22428 36428 22484
rect 36484 22428 36494 22484
rect 38612 22428 40516 22484
rect 20188 22372 20244 22428
rect 34188 22372 34244 22428
rect 13122 22316 13132 22372
rect 13188 22316 13198 22372
rect 14018 22316 14028 22372
rect 14084 22316 14094 22372
rect 14802 22316 14812 22372
rect 14868 22316 17612 22372
rect 17668 22316 17678 22372
rect 20178 22316 20188 22372
rect 20244 22316 20254 22372
rect 31948 22316 34188 22372
rect 34244 22316 34254 22372
rect 35074 22316 35084 22372
rect 35140 22316 35756 22372
rect 35812 22316 36316 22372
rect 36372 22316 36382 22372
rect 13132 22260 13188 22316
rect 6850 22204 6860 22260
rect 6916 22204 10332 22260
rect 10388 22204 11228 22260
rect 11284 22204 11294 22260
rect 12338 22204 12348 22260
rect 12404 22204 13580 22260
rect 13636 22204 13646 22260
rect 14028 22148 14084 22316
rect 31948 22260 32004 22316
rect 40460 22260 40516 22428
rect 14578 22204 14588 22260
rect 14644 22204 15820 22260
rect 15876 22204 15886 22260
rect 24434 22204 24444 22260
rect 24500 22204 32004 22260
rect 32162 22204 32172 22260
rect 32228 22204 34748 22260
rect 34804 22204 34814 22260
rect 40460 22204 41020 22260
rect 41076 22204 41086 22260
rect 41580 22204 41916 22260
rect 41972 22204 42476 22260
rect 42532 22204 42542 22260
rect 41580 22148 41636 22204
rect 2146 22092 2156 22148
rect 2212 22092 9436 22148
rect 9492 22092 9502 22148
rect 10994 22092 11004 22148
rect 11060 22092 14084 22148
rect 19842 22092 19852 22148
rect 19908 22092 20412 22148
rect 20468 22092 21084 22148
rect 21140 22092 21150 22148
rect 22978 22092 22988 22148
rect 23044 22092 23884 22148
rect 23940 22092 26236 22148
rect 26292 22092 26302 22148
rect 29922 22092 29932 22148
rect 29988 22092 30492 22148
rect 30548 22092 30558 22148
rect 35858 22092 35868 22148
rect 35924 22092 37100 22148
rect 37156 22092 37166 22148
rect 41570 22092 41580 22148
rect 41636 22092 41646 22148
rect 41794 22092 41804 22148
rect 41860 22092 43708 22148
rect 43764 22092 43774 22148
rect 5618 21980 5628 22036
rect 5684 21980 10332 22036
rect 10388 21980 10398 22036
rect 11078 21980 11116 22036
rect 11172 21980 11182 22036
rect 14018 21980 14028 22036
rect 14084 21980 14252 22036
rect 14308 21980 14318 22036
rect 21970 21980 21980 22036
rect 22036 21980 22876 22036
rect 22932 21980 23436 22036
rect 23492 21980 42140 22036
rect 42196 21980 42206 22036
rect 42578 21980 42588 22036
rect 42644 21980 44156 22036
rect 44212 21980 44222 22036
rect 19826 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20110 21980
rect 13234 21868 13244 21924
rect 13300 21868 15148 21924
rect 15204 21868 15214 21924
rect 15372 21868 16548 21924
rect 16706 21868 16716 21924
rect 16772 21868 18060 21924
rect 18116 21868 18126 21924
rect 20962 21868 20972 21924
rect 21028 21868 23548 21924
rect 23604 21868 23614 21924
rect 26114 21868 26124 21924
rect 26180 21868 27020 21924
rect 27076 21868 27086 21924
rect 28466 21868 28476 21924
rect 28532 21868 30828 21924
rect 30884 21868 31388 21924
rect 31444 21868 31454 21924
rect 15372 21812 15428 21868
rect 16492 21812 16548 21868
rect 1474 21756 1484 21812
rect 1540 21756 15428 21812
rect 15558 21756 15596 21812
rect 15652 21756 15662 21812
rect 16492 21756 17948 21812
rect 18004 21756 18732 21812
rect 18788 21756 18798 21812
rect 20066 21756 20076 21812
rect 20132 21756 20524 21812
rect 20580 21756 20590 21812
rect 26852 21756 28028 21812
rect 28084 21756 31612 21812
rect 31668 21756 34636 21812
rect 34692 21756 34702 21812
rect 37538 21756 37548 21812
rect 37604 21756 37884 21812
rect 37940 21756 40348 21812
rect 40404 21756 40414 21812
rect 45266 21756 45276 21812
rect 45332 21756 46620 21812
rect 46676 21756 47180 21812
rect 47236 21756 47246 21812
rect 26852 21700 26908 21756
rect 8194 21644 8204 21700
rect 8260 21644 10444 21700
rect 10500 21644 10510 21700
rect 11666 21644 11676 21700
rect 11732 21644 13916 21700
rect 13972 21644 13982 21700
rect 14130 21644 14140 21700
rect 14196 21644 14476 21700
rect 14532 21644 14542 21700
rect 14924 21644 18956 21700
rect 19012 21644 19022 21700
rect 19170 21644 19180 21700
rect 19236 21644 19740 21700
rect 19796 21644 19806 21700
rect 21074 21644 21084 21700
rect 21140 21644 22652 21700
rect 22708 21644 22718 21700
rect 23090 21644 23100 21700
rect 23156 21644 26908 21700
rect 30258 21644 30268 21700
rect 30324 21644 31052 21700
rect 31108 21644 32060 21700
rect 32116 21644 32126 21700
rect 35084 21644 39060 21700
rect 40002 21644 40012 21700
rect 40068 21644 40796 21700
rect 40852 21644 40862 21700
rect 46050 21644 46060 21700
rect 46116 21644 46126 21700
rect 46722 21644 46732 21700
rect 46788 21644 47068 21700
rect 47124 21644 47134 21700
rect 13916 21588 13972 21644
rect 14924 21588 14980 21644
rect 4834 21532 4844 21588
rect 4900 21532 5180 21588
rect 5236 21532 6300 21588
rect 6356 21532 6366 21588
rect 11106 21532 11116 21588
rect 11172 21532 11452 21588
rect 11508 21532 12572 21588
rect 12628 21532 12638 21588
rect 13682 21532 13692 21588
rect 13748 21532 13758 21588
rect 13916 21532 14980 21588
rect 15474 21532 15484 21588
rect 15540 21532 16156 21588
rect 16212 21532 16222 21588
rect 16930 21532 16940 21588
rect 16996 21532 18284 21588
rect 18340 21532 22764 21588
rect 22820 21532 22830 21588
rect 24658 21532 24668 21588
rect 24724 21532 25340 21588
rect 25396 21532 25406 21588
rect 26674 21532 26684 21588
rect 26740 21532 26750 21588
rect 27682 21532 27692 21588
rect 27748 21532 31388 21588
rect 31444 21532 33964 21588
rect 34020 21532 34860 21588
rect 34916 21532 34926 21588
rect 13692 21476 13748 21532
rect 26684 21476 26740 21532
rect 35084 21476 35140 21644
rect 38322 21532 38332 21588
rect 38388 21532 38668 21588
rect 38724 21532 38734 21588
rect 9874 21420 9884 21476
rect 9940 21420 12908 21476
rect 12964 21420 12974 21476
rect 13692 21420 14588 21476
rect 14644 21420 14654 21476
rect 23986 21420 23996 21476
rect 24052 21420 26348 21476
rect 26404 21420 26414 21476
rect 26684 21420 28700 21476
rect 28756 21420 35140 21476
rect 39004 21476 39060 21644
rect 46060 21588 46116 21644
rect 39218 21532 39228 21588
rect 39284 21532 39788 21588
rect 39844 21532 39854 21588
rect 40012 21532 46116 21588
rect 40012 21476 40068 21532
rect 39004 21420 40068 21476
rect 43586 21420 43596 21476
rect 43652 21420 44716 21476
rect 44772 21420 44782 21476
rect 9090 21308 9100 21364
rect 9156 21308 13244 21364
rect 13300 21308 13310 21364
rect 13990 21308 14028 21364
rect 14084 21308 14094 21364
rect 14326 21308 14364 21364
rect 14420 21308 14430 21364
rect 14690 21308 14700 21364
rect 14756 21308 15372 21364
rect 15428 21308 15438 21364
rect 17714 21308 17724 21364
rect 17780 21308 18508 21364
rect 18564 21308 18574 21364
rect 20626 21308 20636 21364
rect 20692 21308 21308 21364
rect 21364 21308 23660 21364
rect 23716 21308 23726 21364
rect 28130 21308 28140 21364
rect 28196 21308 38220 21364
rect 38276 21308 38286 21364
rect 38546 21308 38556 21364
rect 38612 21308 45500 21364
rect 45556 21308 45566 21364
rect 11078 21196 11116 21252
rect 11172 21196 11182 21252
rect 38658 21196 38668 21252
rect 38724 21196 39228 21252
rect 39284 21196 39294 21252
rect 4466 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4750 21196
rect 35186 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35470 21196
rect 49200 21140 50000 21168
rect 10658 21084 10668 21140
rect 10724 21084 11452 21140
rect 11508 21084 13468 21140
rect 13524 21084 15596 21140
rect 15652 21084 15662 21140
rect 19170 21084 19180 21140
rect 19236 21084 20188 21140
rect 20244 21084 20254 21140
rect 20626 21084 20636 21140
rect 20692 21084 21644 21140
rect 21700 21084 21710 21140
rect 23874 21084 23884 21140
rect 23940 21084 23950 21140
rect 25666 21084 25676 21140
rect 25732 21084 29596 21140
rect 29652 21084 29662 21140
rect 46274 21084 46284 21140
rect 46340 21084 48188 21140
rect 48244 21084 50000 21140
rect 4722 20972 4732 21028
rect 4788 20972 6748 21028
rect 6804 20972 6814 21028
rect 10770 20972 10780 21028
rect 10836 20972 14252 21028
rect 14308 20972 14318 21028
rect 19394 20972 19404 21028
rect 19460 20972 20412 21028
rect 20468 20972 21420 21028
rect 21476 20972 21486 21028
rect 23884 20916 23940 21084
rect 49200 21056 50000 21084
rect 25330 20972 25340 21028
rect 25396 20972 26460 21028
rect 26516 20972 26526 21028
rect 35746 20972 35756 21028
rect 35812 20972 37660 21028
rect 37716 20972 37726 21028
rect 4834 20860 4844 20916
rect 4900 20860 9996 20916
rect 10052 20860 10062 20916
rect 14130 20860 14140 20916
rect 14196 20860 15148 20916
rect 17938 20860 17948 20916
rect 18004 20860 21532 20916
rect 21588 20860 21598 20916
rect 23884 20860 24892 20916
rect 24948 20860 27356 20916
rect 27412 20860 27422 20916
rect 44370 20860 44380 20916
rect 44436 20860 44940 20916
rect 44996 20860 45388 20916
rect 45444 20860 46844 20916
rect 46900 20860 48076 20916
rect 48132 20860 48142 20916
rect 15092 20804 15148 20860
rect 6738 20748 6748 20804
rect 6804 20748 7980 20804
rect 8036 20748 8764 20804
rect 8820 20748 10668 20804
rect 10724 20748 10734 20804
rect 15092 20748 17724 20804
rect 17780 20748 17790 20804
rect 19292 20692 19348 20860
rect 19506 20748 19516 20804
rect 19572 20748 20188 20804
rect 20244 20748 20254 20804
rect 20402 20748 20412 20804
rect 20468 20748 21308 20804
rect 21364 20748 21374 20804
rect 38994 20748 39004 20804
rect 39060 20748 39564 20804
rect 39620 20748 39630 20804
rect 9538 20636 9548 20692
rect 9604 20636 11564 20692
rect 11620 20636 11630 20692
rect 12450 20636 12460 20692
rect 12516 20636 13244 20692
rect 13300 20636 13310 20692
rect 13458 20636 13468 20692
rect 13524 20636 14700 20692
rect 14756 20636 14766 20692
rect 15810 20636 15820 20692
rect 15876 20636 16268 20692
rect 16324 20636 16334 20692
rect 19292 20636 19404 20692
rect 19460 20636 19470 20692
rect 19730 20636 19740 20692
rect 19796 20636 20748 20692
rect 20804 20636 20814 20692
rect 21410 20636 21420 20692
rect 21476 20636 22092 20692
rect 22148 20636 22158 20692
rect 23426 20636 23436 20692
rect 23492 20636 23884 20692
rect 23940 20636 24332 20692
rect 24388 20636 24398 20692
rect 26562 20636 26572 20692
rect 26628 20636 26908 20692
rect 29250 20636 29260 20692
rect 29316 20636 31500 20692
rect 31556 20636 32508 20692
rect 32564 20636 34860 20692
rect 34916 20636 34926 20692
rect 36194 20636 36204 20692
rect 36260 20636 36988 20692
rect 37044 20636 37054 20692
rect 38546 20636 38556 20692
rect 38612 20636 40796 20692
rect 40852 20636 42700 20692
rect 42756 20636 42766 20692
rect 43110 20636 43148 20692
rect 43204 20636 43932 20692
rect 43988 20636 43998 20692
rect 11564 20468 11620 20636
rect 26852 20580 26908 20636
rect 12898 20524 12908 20580
rect 12964 20524 14476 20580
rect 14532 20524 14542 20580
rect 19058 20524 19068 20580
rect 19124 20524 22820 20580
rect 26852 20524 28364 20580
rect 28420 20524 29036 20580
rect 29092 20524 29102 20580
rect 33842 20524 33852 20580
rect 33908 20524 34020 20580
rect 35942 20524 35980 20580
rect 36036 20524 36652 20580
rect 36708 20524 36718 20580
rect 39218 20524 39228 20580
rect 39284 20524 40236 20580
rect 40292 20524 41244 20580
rect 41300 20524 41310 20580
rect 22764 20468 22820 20524
rect 33964 20468 34020 20524
rect 11564 20412 14588 20468
rect 14644 20412 15036 20468
rect 15092 20412 15102 20468
rect 18274 20412 18284 20468
rect 18340 20412 19180 20468
rect 19236 20412 19246 20468
rect 22754 20412 22764 20468
rect 22820 20412 22830 20468
rect 33964 20412 36988 20468
rect 37044 20412 37054 20468
rect 19826 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20110 20412
rect 11666 20300 11676 20356
rect 11732 20300 14924 20356
rect 14980 20300 14990 20356
rect 21858 20300 21868 20356
rect 21924 20300 26908 20356
rect 26964 20300 26974 20356
rect 33618 20300 33628 20356
rect 33684 20300 34188 20356
rect 34244 20300 34254 20356
rect 35522 20300 35532 20356
rect 35588 20300 35868 20356
rect 35924 20300 35934 20356
rect 44258 20300 44268 20356
rect 44324 20300 45276 20356
rect 45332 20300 45342 20356
rect 5506 20188 5516 20244
rect 5572 20188 8372 20244
rect 9762 20188 9772 20244
rect 9828 20188 11004 20244
rect 11060 20188 11070 20244
rect 12674 20188 12684 20244
rect 12740 20188 15484 20244
rect 15540 20188 15550 20244
rect 19618 20188 19628 20244
rect 19684 20188 20972 20244
rect 21028 20188 23660 20244
rect 23716 20188 23726 20244
rect 8316 20132 8372 20188
rect 26852 20132 26908 20300
rect 34962 20188 34972 20244
rect 35028 20188 35756 20244
rect 35812 20188 35822 20244
rect 38854 20188 38892 20244
rect 38948 20188 38958 20244
rect 8316 20076 12012 20132
rect 12068 20076 12078 20132
rect 12562 20076 12572 20132
rect 12628 20076 12638 20132
rect 13206 20076 13244 20132
rect 13300 20076 13310 20132
rect 13794 20076 13804 20132
rect 13860 20076 14700 20132
rect 14756 20076 14766 20132
rect 14924 20076 15148 20132
rect 15204 20076 15214 20132
rect 16482 20076 16492 20132
rect 16548 20076 17388 20132
rect 17444 20076 17454 20132
rect 17826 20076 17836 20132
rect 17892 20076 21868 20132
rect 21924 20076 21934 20132
rect 22614 20076 22652 20132
rect 22708 20076 22718 20132
rect 26852 20076 33740 20132
rect 33796 20076 33806 20132
rect 35074 20076 35084 20132
rect 35140 20076 35644 20132
rect 35700 20076 36092 20132
rect 36148 20076 36316 20132
rect 36372 20076 36382 20132
rect 37090 20076 37100 20132
rect 37156 20076 37772 20132
rect 37828 20076 38108 20132
rect 38164 20076 38174 20132
rect 39666 20076 39676 20132
rect 39732 20076 42140 20132
rect 42196 20076 43260 20132
rect 43316 20076 44380 20132
rect 44436 20076 44446 20132
rect 45490 20076 45500 20132
rect 45556 20076 47516 20132
rect 47572 20076 47582 20132
rect 12572 20020 12628 20076
rect 14924 20020 14980 20076
rect 6290 19964 6300 20020
rect 6356 19964 8652 20020
rect 8708 19964 8718 20020
rect 10658 19964 10668 20020
rect 10724 19964 12348 20020
rect 12404 19964 12414 20020
rect 12572 19964 14980 20020
rect 15092 19964 15260 20020
rect 15316 19964 16268 20020
rect 16324 19964 16334 20020
rect 16930 19964 16940 20020
rect 16996 19964 17612 20020
rect 17668 19964 17678 20020
rect 18050 19964 18060 20020
rect 18116 19964 18396 20020
rect 18452 19964 18462 20020
rect 18946 19964 18956 20020
rect 19012 19964 20188 20020
rect 20244 19964 22204 20020
rect 22260 19964 22270 20020
rect 31714 19964 31724 20020
rect 31780 19964 32172 20020
rect 32228 19964 32238 20020
rect 35756 19964 38668 20020
rect 41346 19964 41356 20020
rect 41412 19964 41916 20020
rect 41972 19964 41982 20020
rect 43698 19964 43708 20020
rect 43764 19964 45052 20020
rect 45108 19964 45724 20020
rect 45780 19964 46172 20020
rect 46228 19964 46238 20020
rect 15092 19908 15148 19964
rect 35756 19908 35812 19964
rect 38612 19908 38668 19964
rect 5058 19852 5068 19908
rect 5124 19852 5740 19908
rect 5796 19852 5806 19908
rect 13010 19852 13020 19908
rect 13076 19852 14028 19908
rect 14084 19852 14094 19908
rect 14914 19852 14924 19908
rect 14980 19852 15148 19908
rect 15698 19852 15708 19908
rect 15764 19852 17500 19908
rect 17556 19852 17566 19908
rect 18834 19852 18844 19908
rect 18900 19852 19628 19908
rect 19684 19852 19694 19908
rect 26226 19852 26236 19908
rect 26292 19852 28924 19908
rect 28980 19852 34412 19908
rect 34468 19852 35756 19908
rect 35812 19852 35822 19908
rect 35970 19852 35980 19908
rect 36036 19852 37100 19908
rect 37156 19852 37166 19908
rect 38612 19852 38892 19908
rect 38948 19852 40012 19908
rect 40068 19852 40078 19908
rect 40226 19852 40236 19908
rect 40292 19852 41020 19908
rect 41076 19852 41086 19908
rect 44258 19852 44268 19908
rect 44324 19852 46620 19908
rect 46676 19852 46686 19908
rect 4946 19740 4956 19796
rect 5012 19740 6748 19796
rect 6804 19740 6814 19796
rect 9762 19740 9772 19796
rect 9828 19740 12012 19796
rect 12068 19740 12078 19796
rect 14690 19740 14700 19796
rect 14756 19740 22652 19796
rect 22708 19740 22718 19796
rect 27916 19740 29708 19796
rect 29764 19740 30156 19796
rect 30212 19740 30222 19796
rect 34748 19740 36316 19796
rect 36372 19740 36382 19796
rect 38612 19740 41132 19796
rect 41188 19740 42812 19796
rect 42868 19740 42878 19796
rect 27916 19684 27972 19740
rect 34748 19684 34804 19740
rect 38612 19684 38668 19740
rect 10882 19628 10892 19684
rect 10948 19628 11452 19684
rect 11508 19628 12908 19684
rect 12964 19628 12974 19684
rect 19170 19628 19180 19684
rect 19236 19628 19628 19684
rect 19684 19628 21980 19684
rect 22036 19628 22046 19684
rect 25890 19628 25900 19684
rect 25956 19628 26796 19684
rect 26852 19628 26862 19684
rect 27906 19628 27916 19684
rect 27972 19628 27982 19684
rect 33730 19628 33740 19684
rect 33796 19628 34748 19684
rect 34804 19628 34814 19684
rect 35532 19628 38668 19684
rect 39218 19628 39228 19684
rect 39284 19628 41804 19684
rect 41860 19628 41870 19684
rect 4466 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4750 19628
rect 35186 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35470 19628
rect 15092 19516 18396 19572
rect 18452 19516 20188 19572
rect 20244 19516 24220 19572
rect 24276 19516 24286 19572
rect 15092 19460 15148 19516
rect 35532 19460 35588 19628
rect 37538 19516 37548 19572
rect 37604 19516 39116 19572
rect 39172 19516 39182 19572
rect 40450 19516 40460 19572
rect 40516 19516 42252 19572
rect 42308 19516 42318 19572
rect 1586 19404 1596 19460
rect 1652 19404 15148 19460
rect 16706 19404 16716 19460
rect 16772 19404 25564 19460
rect 25620 19404 25788 19460
rect 25844 19404 25854 19460
rect 30370 19404 30380 19460
rect 30436 19404 35588 19460
rect 36082 19404 36092 19460
rect 36148 19404 43708 19460
rect 43764 19404 43774 19460
rect 7858 19292 7868 19348
rect 7924 19292 12124 19348
rect 12180 19292 12190 19348
rect 13570 19292 13580 19348
rect 13636 19292 16044 19348
rect 16100 19292 17164 19348
rect 17220 19292 20300 19348
rect 20356 19292 20366 19348
rect 21746 19292 21756 19348
rect 21812 19292 22652 19348
rect 22708 19292 25116 19348
rect 25172 19292 30492 19348
rect 30548 19292 31052 19348
rect 31108 19292 31118 19348
rect 31266 19292 31276 19348
rect 31332 19292 32060 19348
rect 32116 19292 32126 19348
rect 33282 19292 33292 19348
rect 33348 19292 34524 19348
rect 34580 19292 34916 19348
rect 35970 19292 35980 19348
rect 36036 19292 38668 19348
rect 34860 19236 34916 19292
rect 38612 19236 38668 19292
rect 7298 19180 7308 19236
rect 7364 19180 8316 19236
rect 8372 19180 10220 19236
rect 10276 19180 13580 19236
rect 13636 19180 13646 19236
rect 14130 19180 14140 19236
rect 14196 19180 15596 19236
rect 15652 19180 15662 19236
rect 18722 19180 18732 19236
rect 18788 19180 21420 19236
rect 21476 19180 22092 19236
rect 22148 19180 24220 19236
rect 24276 19180 26236 19236
rect 26292 19180 26302 19236
rect 34860 19180 37212 19236
rect 37268 19180 37278 19236
rect 38612 19180 44268 19236
rect 44324 19180 44334 19236
rect 5730 19068 5740 19124
rect 5796 19068 9548 19124
rect 9604 19068 9614 19124
rect 11778 19068 11788 19124
rect 11844 19068 15148 19124
rect 15204 19068 18844 19124
rect 18900 19068 18910 19124
rect 25330 19068 25340 19124
rect 25396 19068 27916 19124
rect 27972 19068 27982 19124
rect 34626 19068 34636 19124
rect 34692 19068 35084 19124
rect 35140 19068 35150 19124
rect 35410 19068 35420 19124
rect 35476 19068 37772 19124
rect 37828 19068 37838 19124
rect 43362 19068 43372 19124
rect 43428 19068 44828 19124
rect 44884 19068 44894 19124
rect 11106 18956 11116 19012
rect 11172 18956 13580 19012
rect 13636 18956 13646 19012
rect 14802 18956 14812 19012
rect 14868 18956 16492 19012
rect 16548 18956 16558 19012
rect 16930 18956 16940 19012
rect 16996 18956 17388 19012
rect 17444 18956 17454 19012
rect 37538 18956 37548 19012
rect 37604 18956 37996 19012
rect 38052 18956 38668 19012
rect 38724 18956 38734 19012
rect 42130 18956 42140 19012
rect 42196 18956 42700 19012
rect 42756 18956 42766 19012
rect 34402 18844 34412 18900
rect 34468 18844 35196 18900
rect 35252 18844 35262 18900
rect 36194 18844 36204 18900
rect 36260 18844 36876 18900
rect 36932 18844 36942 18900
rect 19826 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20110 18844
rect 29026 18732 29036 18788
rect 29092 18732 30268 18788
rect 30324 18732 30334 18788
rect 32050 18732 32060 18788
rect 32116 18732 41804 18788
rect 41860 18732 41870 18788
rect 8866 18620 8876 18676
rect 8932 18620 11452 18676
rect 11508 18620 11518 18676
rect 23650 18620 23660 18676
rect 23716 18620 24668 18676
rect 24724 18620 25228 18676
rect 25284 18620 26572 18676
rect 26628 18620 26638 18676
rect 26786 18620 26796 18676
rect 26852 18620 29148 18676
rect 29204 18620 29214 18676
rect 35186 18620 35196 18676
rect 35252 18620 35868 18676
rect 35924 18620 36092 18676
rect 36148 18620 36158 18676
rect 44930 18620 44940 18676
rect 44996 18620 46396 18676
rect 46452 18620 46462 18676
rect 11778 18508 11788 18564
rect 11844 18508 12460 18564
rect 12516 18508 12526 18564
rect 17490 18508 17500 18564
rect 17556 18508 18620 18564
rect 18676 18508 20244 18564
rect 25442 18508 25452 18564
rect 25508 18508 25900 18564
rect 25956 18508 25966 18564
rect 42466 18508 42476 18564
rect 42532 18508 45164 18564
rect 45220 18508 45230 18564
rect 20188 18452 20244 18508
rect 13122 18396 13132 18452
rect 13188 18396 15596 18452
rect 15652 18396 15662 18452
rect 16930 18396 16940 18452
rect 16996 18396 17724 18452
rect 17780 18396 17790 18452
rect 20188 18396 22204 18452
rect 22260 18396 22270 18452
rect 23202 18396 23212 18452
rect 23268 18396 23996 18452
rect 24052 18396 24062 18452
rect 24658 18396 24668 18452
rect 24724 18396 33292 18452
rect 33348 18396 33358 18452
rect 35074 18396 35084 18452
rect 35140 18396 35308 18452
rect 35364 18396 35374 18452
rect 35522 18396 35532 18452
rect 35588 18396 35868 18452
rect 35924 18396 37212 18452
rect 37268 18396 37278 18452
rect 38210 18396 38220 18452
rect 38276 18396 38780 18452
rect 38836 18396 40012 18452
rect 40068 18396 40908 18452
rect 40964 18396 41692 18452
rect 41748 18396 41758 18452
rect 42252 18396 42924 18452
rect 42980 18396 43372 18452
rect 43428 18396 43438 18452
rect 43586 18396 43596 18452
rect 43652 18396 44828 18452
rect 44884 18396 46956 18452
rect 47012 18396 48188 18452
rect 48244 18396 48254 18452
rect 24668 18340 24724 18396
rect 42252 18340 42308 18396
rect 14690 18284 14700 18340
rect 14756 18284 16380 18340
rect 16436 18284 16446 18340
rect 17490 18284 17500 18340
rect 17556 18284 18060 18340
rect 18116 18284 18126 18340
rect 21522 18284 21532 18340
rect 21588 18284 23548 18340
rect 23604 18284 23614 18340
rect 23874 18284 23884 18340
rect 23940 18284 24724 18340
rect 28354 18284 28364 18340
rect 28420 18284 30044 18340
rect 30100 18284 30110 18340
rect 33506 18284 33516 18340
rect 33572 18284 34636 18340
rect 34692 18284 34702 18340
rect 40338 18284 40348 18340
rect 40404 18284 42308 18340
rect 42578 18284 42588 18340
rect 42644 18284 43932 18340
rect 43988 18284 43998 18340
rect 44342 18284 44380 18340
rect 44436 18284 44446 18340
rect 23548 18228 23604 18284
rect 23548 18172 25004 18228
rect 25060 18172 25070 18228
rect 33394 18172 33404 18228
rect 33460 18172 34300 18228
rect 34356 18172 34366 18228
rect 44034 18172 44044 18228
rect 44100 18172 45052 18228
rect 45108 18172 45118 18228
rect 38612 18060 39452 18116
rect 39508 18060 44380 18116
rect 44436 18060 44446 18116
rect 4466 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4750 18060
rect 35186 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35470 18060
rect 38612 18004 38668 18060
rect 13682 17948 13692 18004
rect 13748 17948 31724 18004
rect 31780 17948 31790 18004
rect 36306 17948 36316 18004
rect 36372 17948 36876 18004
rect 36932 17948 38668 18004
rect 18274 17836 18284 17892
rect 18340 17836 18844 17892
rect 18900 17836 20580 17892
rect 21746 17836 21756 17892
rect 21812 17836 23548 17892
rect 23604 17836 23614 17892
rect 23772 17836 28476 17892
rect 28532 17836 28542 17892
rect 32274 17836 32284 17892
rect 32340 17836 33180 17892
rect 33236 17836 33964 17892
rect 34020 17836 36428 17892
rect 36484 17836 37884 17892
rect 37940 17836 37950 17892
rect 20524 17780 20580 17836
rect 23772 17780 23828 17836
rect 12786 17724 12796 17780
rect 12852 17724 13580 17780
rect 13636 17724 15148 17780
rect 15204 17724 15214 17780
rect 19394 17724 19404 17780
rect 19460 17724 19740 17780
rect 19796 17724 19806 17780
rect 20514 17724 20524 17780
rect 20580 17724 23828 17780
rect 26012 17724 28588 17780
rect 28644 17724 28654 17780
rect 28914 17724 28924 17780
rect 28980 17724 29820 17780
rect 29876 17724 32956 17780
rect 33012 17724 33022 17780
rect 34178 17724 34188 17780
rect 34244 17724 34636 17780
rect 34692 17724 34702 17780
rect 34962 17724 34972 17780
rect 35028 17724 37660 17780
rect 37716 17724 43708 17780
rect 43764 17724 44044 17780
rect 44100 17724 44110 17780
rect 26012 17668 26068 17724
rect 34636 17668 34692 17724
rect 10882 17612 10892 17668
rect 10948 17612 13020 17668
rect 13076 17612 13086 17668
rect 16930 17612 16940 17668
rect 16996 17612 19628 17668
rect 19684 17612 19694 17668
rect 22194 17612 22204 17668
rect 22260 17612 22764 17668
rect 22820 17612 22830 17668
rect 24098 17612 24108 17668
rect 24164 17612 26012 17668
rect 26068 17612 26078 17668
rect 26226 17612 26236 17668
rect 26292 17612 28140 17668
rect 28196 17612 34356 17668
rect 34636 17612 34860 17668
rect 34916 17612 34926 17668
rect 36082 17612 36092 17668
rect 36148 17612 39116 17668
rect 39172 17612 39182 17668
rect 43586 17612 43596 17668
rect 43652 17612 44156 17668
rect 44212 17612 47180 17668
rect 47236 17612 48188 17668
rect 48244 17612 48254 17668
rect 34300 17556 34356 17612
rect 36092 17556 36148 17612
rect 17826 17500 17836 17556
rect 17892 17500 18732 17556
rect 18788 17500 19404 17556
rect 19460 17500 21644 17556
rect 21700 17500 21710 17556
rect 28466 17500 28476 17556
rect 28532 17500 29148 17556
rect 29204 17500 29214 17556
rect 29372 17500 31388 17556
rect 31444 17500 31454 17556
rect 34290 17500 34300 17556
rect 34356 17500 34366 17556
rect 34514 17500 34524 17556
rect 34580 17500 36148 17556
rect 38882 17500 38892 17556
rect 38948 17500 41804 17556
rect 41860 17500 41870 17556
rect 44342 17500 44380 17556
rect 44436 17500 44446 17556
rect 44930 17500 44940 17556
rect 44996 17500 46060 17556
rect 46116 17500 46126 17556
rect 29372 17444 29428 17500
rect 17938 17388 17948 17444
rect 18004 17388 19180 17444
rect 19236 17388 19246 17444
rect 22530 17388 22540 17444
rect 22596 17388 26460 17444
rect 26516 17388 28140 17444
rect 28196 17388 29260 17444
rect 29316 17388 29428 17444
rect 31154 17388 31164 17444
rect 31220 17388 32284 17444
rect 32340 17388 32350 17444
rect 43474 17388 43484 17444
rect 43540 17388 45388 17444
rect 45444 17388 45454 17444
rect 29362 17276 29372 17332
rect 29428 17276 29708 17332
rect 29764 17276 29774 17332
rect 41010 17276 41020 17332
rect 41076 17276 42924 17332
rect 42980 17276 43596 17332
rect 43652 17276 43662 17332
rect 44706 17276 44716 17332
rect 44772 17276 45164 17332
rect 45220 17276 45230 17332
rect 19826 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20110 17276
rect 26870 17164 26908 17220
rect 26964 17164 26974 17220
rect 33506 17164 33516 17220
rect 33572 17164 34188 17220
rect 34244 17164 34254 17220
rect 35420 17164 36652 17220
rect 36708 17164 36718 17220
rect 38434 17164 38444 17220
rect 38500 17164 41356 17220
rect 41412 17164 42252 17220
rect 42308 17164 42318 17220
rect 45042 17164 45052 17220
rect 45108 17164 45612 17220
rect 45668 17164 45678 17220
rect 46050 17164 46060 17220
rect 46116 17164 47852 17220
rect 47908 17164 47918 17220
rect 26908 17108 26964 17164
rect 35420 17108 35476 17164
rect 10546 17052 10556 17108
rect 10612 17052 12012 17108
rect 12068 17052 13580 17108
rect 13636 17052 13646 17108
rect 17042 17052 17052 17108
rect 17108 17052 17500 17108
rect 17556 17052 20076 17108
rect 20132 17052 21868 17108
rect 21924 17052 23100 17108
rect 23156 17052 23660 17108
rect 23716 17052 23726 17108
rect 26908 17052 34412 17108
rect 34468 17052 35420 17108
rect 35476 17052 35486 17108
rect 36306 17052 36316 17108
rect 36372 17052 37100 17108
rect 37156 17052 37166 17108
rect 42690 17052 42700 17108
rect 42756 17052 43372 17108
rect 43428 17052 43820 17108
rect 43876 17052 46564 17108
rect 16818 16940 16828 16996
rect 16884 16940 18172 16996
rect 18228 16940 18620 16996
rect 18676 16940 18686 16996
rect 27234 16940 27244 16996
rect 27300 16940 28364 16996
rect 28420 16940 36428 16996
rect 36484 16940 36494 16996
rect 39778 16940 39788 16996
rect 39844 16940 41132 16996
rect 41188 16940 42252 16996
rect 42308 16940 42318 16996
rect 43026 16940 43036 16996
rect 43092 16940 46340 16996
rect 46284 16884 46340 16940
rect 46508 16884 46564 17052
rect 11554 16828 11564 16884
rect 11620 16828 14028 16884
rect 14084 16828 14094 16884
rect 18722 16828 18732 16884
rect 18788 16828 22316 16884
rect 22372 16828 22382 16884
rect 30146 16828 30156 16884
rect 30212 16828 31388 16884
rect 31444 16828 34860 16884
rect 34916 16828 34926 16884
rect 35942 16828 35980 16884
rect 36036 16828 36046 16884
rect 36642 16828 36652 16884
rect 36708 16828 37884 16884
rect 37940 16828 37950 16884
rect 38770 16828 38780 16884
rect 38836 16828 39564 16884
rect 39620 16828 40908 16884
rect 40964 16828 40974 16884
rect 43250 16828 43260 16884
rect 43316 16828 45500 16884
rect 45556 16828 45566 16884
rect 46274 16828 46284 16884
rect 46340 16828 46350 16884
rect 46498 16828 46508 16884
rect 46564 16828 46574 16884
rect 21634 16716 21644 16772
rect 21700 16716 22988 16772
rect 23044 16716 23054 16772
rect 30482 16716 30492 16772
rect 30548 16716 31164 16772
rect 31220 16716 31230 16772
rect 32274 16716 32284 16772
rect 32340 16716 38556 16772
rect 38612 16716 38622 16772
rect 43138 16716 43148 16772
rect 43204 16716 44716 16772
rect 44772 16716 44782 16772
rect 44940 16716 46844 16772
rect 46900 16716 47404 16772
rect 47460 16716 47470 16772
rect 44940 16660 44996 16716
rect 21970 16604 21980 16660
rect 22036 16604 25676 16660
rect 25732 16604 25742 16660
rect 26898 16604 26908 16660
rect 26964 16604 32508 16660
rect 32564 16604 32574 16660
rect 33618 16604 33628 16660
rect 33684 16604 35588 16660
rect 36418 16604 36428 16660
rect 36484 16604 37100 16660
rect 37156 16604 37166 16660
rect 41458 16604 41468 16660
rect 41524 16604 42924 16660
rect 42980 16604 44996 16660
rect 45378 16604 45388 16660
rect 45444 16604 45948 16660
rect 46004 16604 46014 16660
rect 35532 16548 35588 16604
rect 35532 16492 39116 16548
rect 39172 16492 39182 16548
rect 41682 16492 41692 16548
rect 41748 16492 43148 16548
rect 43204 16492 43932 16548
rect 43988 16492 43998 16548
rect 44146 16492 44156 16548
rect 44212 16492 46060 16548
rect 46116 16492 46126 16548
rect 4466 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4750 16492
rect 35186 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35470 16492
rect 35532 16380 38668 16436
rect 41570 16380 41580 16436
rect 41636 16380 42924 16436
rect 42980 16380 45388 16436
rect 45444 16380 45454 16436
rect 35532 16324 35588 16380
rect 38612 16324 38668 16380
rect 14018 16268 14028 16324
rect 14084 16268 14924 16324
rect 14980 16268 17164 16324
rect 17220 16268 17612 16324
rect 17668 16268 17678 16324
rect 31938 16268 31948 16324
rect 32004 16268 35588 16324
rect 35858 16268 35868 16324
rect 35924 16268 36988 16324
rect 37044 16268 37054 16324
rect 38612 16268 44996 16324
rect 45154 16268 45164 16324
rect 45220 16268 45724 16324
rect 45780 16268 46732 16324
rect 46788 16268 46798 16324
rect 44940 16212 44996 16268
rect 16594 16156 16604 16212
rect 16660 16156 17500 16212
rect 17556 16156 21644 16212
rect 21700 16156 21710 16212
rect 35410 16156 35420 16212
rect 35476 16156 35868 16212
rect 35924 16156 35934 16212
rect 36306 16156 36316 16212
rect 36372 16156 37212 16212
rect 37268 16156 39564 16212
rect 39620 16156 39630 16212
rect 43372 16156 44044 16212
rect 44100 16156 44110 16212
rect 44940 16156 47852 16212
rect 47908 16156 47918 16212
rect 43372 16100 43428 16156
rect 20402 16044 20412 16100
rect 20468 16044 21196 16100
rect 21252 16044 22204 16100
rect 22260 16044 22270 16100
rect 22428 16044 27132 16100
rect 27188 16044 27198 16100
rect 33506 16044 33516 16100
rect 33572 16044 34636 16100
rect 34692 16044 34702 16100
rect 36530 16044 36540 16100
rect 36596 16044 37548 16100
rect 37604 16044 39004 16100
rect 39060 16044 39900 16100
rect 39956 16044 39966 16100
rect 42102 16044 42140 16100
rect 42196 16044 43372 16100
rect 43428 16044 43438 16100
rect 43698 16044 43708 16100
rect 43764 16044 45052 16100
rect 45108 16044 45118 16100
rect 22428 15988 22484 16044
rect 42140 15988 42196 16044
rect 18498 15932 18508 15988
rect 18564 15932 20748 15988
rect 20804 15932 22484 15988
rect 25778 15932 25788 15988
rect 25844 15932 26572 15988
rect 26628 15932 32172 15988
rect 32228 15932 33292 15988
rect 33348 15932 34300 15988
rect 34356 15932 34366 15988
rect 38612 15932 42196 15988
rect 42354 15932 42364 15988
rect 42420 15932 44940 15988
rect 44996 15932 45006 15988
rect 38612 15876 38668 15932
rect 16034 15820 16044 15876
rect 16100 15820 17276 15876
rect 17332 15820 17342 15876
rect 18386 15820 18396 15876
rect 18452 15820 18844 15876
rect 18900 15820 18910 15876
rect 19170 15820 19180 15876
rect 19236 15820 20412 15876
rect 20468 15820 20478 15876
rect 33954 15820 33964 15876
rect 34020 15820 38668 15876
rect 39442 15820 39452 15876
rect 39508 15820 42028 15876
rect 42084 15820 43372 15876
rect 43428 15820 43438 15876
rect 44370 15820 44380 15876
rect 44436 15820 45220 15876
rect 47618 15820 47628 15876
rect 47684 15820 48188 15876
rect 48244 15820 48254 15876
rect 19180 15652 19236 15820
rect 19590 15708 19628 15764
rect 19684 15708 19694 15764
rect 35634 15708 35644 15764
rect 35700 15708 35868 15764
rect 35924 15708 35980 15764
rect 36036 15708 36046 15764
rect 37650 15708 37660 15764
rect 37716 15708 38556 15764
rect 38612 15708 38622 15764
rect 19826 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20110 15708
rect 39452 15652 39508 15820
rect 44818 15708 44828 15764
rect 44884 15708 44894 15764
rect 18834 15596 18844 15652
rect 18900 15596 19236 15652
rect 35858 15596 35868 15652
rect 35924 15596 36876 15652
rect 36932 15596 36942 15652
rect 39004 15596 39508 15652
rect 39778 15596 39788 15652
rect 39844 15596 41020 15652
rect 41076 15596 41086 15652
rect 43026 15596 43036 15652
rect 43092 15596 43596 15652
rect 43652 15596 43662 15652
rect 39004 15540 39060 15596
rect 20738 15484 20748 15540
rect 20804 15484 21868 15540
rect 21924 15484 21934 15540
rect 23538 15484 23548 15540
rect 23604 15484 25228 15540
rect 25284 15484 25294 15540
rect 32386 15484 32396 15540
rect 32452 15484 33292 15540
rect 33348 15484 33852 15540
rect 33908 15484 34860 15540
rect 34916 15484 34926 15540
rect 37426 15484 37436 15540
rect 37492 15484 39060 15540
rect 39218 15484 39228 15540
rect 39284 15484 40236 15540
rect 40292 15484 40302 15540
rect 41570 15484 41580 15540
rect 41636 15484 42588 15540
rect 42644 15484 42654 15540
rect 22978 15372 22988 15428
rect 23044 15372 30940 15428
rect 30996 15372 31006 15428
rect 38098 15372 38108 15428
rect 38164 15372 38668 15428
rect 38724 15372 38892 15428
rect 38948 15372 38958 15428
rect 39228 15316 39284 15484
rect 44828 15428 44884 15708
rect 45164 15428 45220 15820
rect 41906 15372 41916 15428
rect 41972 15372 43036 15428
rect 43092 15372 44884 15428
rect 45154 15372 45164 15428
rect 45220 15372 45230 15428
rect 49200 15316 50000 15344
rect 16258 15260 16268 15316
rect 16324 15260 17164 15316
rect 17220 15260 17230 15316
rect 19730 15260 19740 15316
rect 19796 15260 20188 15316
rect 20244 15260 21308 15316
rect 21364 15260 21374 15316
rect 24098 15260 24108 15316
rect 24164 15260 26236 15316
rect 26292 15260 26302 15316
rect 27244 15260 33964 15316
rect 34020 15260 34030 15316
rect 34178 15260 34188 15316
rect 34244 15260 35084 15316
rect 35140 15260 39284 15316
rect 42242 15260 42252 15316
rect 42308 15260 42700 15316
rect 42756 15260 42766 15316
rect 43698 15260 43708 15316
rect 43764 15260 44604 15316
rect 44660 15260 44670 15316
rect 48178 15260 48188 15316
rect 48244 15260 50000 15316
rect 27244 15204 27300 15260
rect 49200 15232 50000 15260
rect 14690 15148 14700 15204
rect 14756 15148 16380 15204
rect 16436 15148 16446 15204
rect 16706 15148 16716 15204
rect 16772 15148 19292 15204
rect 19348 15148 19358 15204
rect 23846 15148 23884 15204
rect 23940 15148 23950 15204
rect 24770 15148 24780 15204
rect 24836 15148 25564 15204
rect 25620 15148 25630 15204
rect 26562 15148 26572 15204
rect 26628 15148 27300 15204
rect 27458 15148 27468 15204
rect 27524 15148 27916 15204
rect 27972 15148 34020 15204
rect 35858 15148 35868 15204
rect 35924 15148 38332 15204
rect 38388 15148 38398 15204
rect 38546 15148 38556 15204
rect 38612 15148 39116 15204
rect 39172 15148 39182 15204
rect 41010 15148 41020 15204
rect 41076 15148 41916 15204
rect 41972 15148 44156 15204
rect 44212 15148 44940 15204
rect 44996 15148 45006 15204
rect 26226 15036 26236 15092
rect 26292 15036 27132 15092
rect 27188 15036 27198 15092
rect 26870 14924 26908 14980
rect 26964 14924 26974 14980
rect 4466 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4750 14924
rect 33964 14756 34020 15148
rect 45266 15092 45276 15148
rect 45332 15092 45342 15148
rect 34188 15036 35420 15092
rect 35476 15036 35486 15092
rect 36194 15036 36204 15092
rect 36260 15036 45332 15092
rect 34188 14980 34244 15036
rect 34178 14924 34188 14980
rect 34244 14924 34254 14980
rect 38854 14924 38892 14980
rect 38948 14924 38958 14980
rect 35186 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35470 14924
rect 42886 14812 42924 14868
rect 42980 14812 42990 14868
rect 33964 14700 34076 14756
rect 34132 14700 36204 14756
rect 36260 14700 36270 14756
rect 29586 14588 29596 14644
rect 29652 14588 30492 14644
rect 30548 14588 30558 14644
rect 31938 14588 31948 14644
rect 32004 14588 32732 14644
rect 32788 14588 33404 14644
rect 33460 14588 33470 14644
rect 18050 14476 18060 14532
rect 18116 14476 25004 14532
rect 25060 14476 25070 14532
rect 20514 14364 20524 14420
rect 20580 14364 22876 14420
rect 22932 14364 22942 14420
rect 30818 14364 30828 14420
rect 30884 14364 31948 14420
rect 32004 14364 32014 14420
rect 43026 14364 43036 14420
rect 43092 14364 44268 14420
rect 44324 14364 44334 14420
rect 24994 14252 25004 14308
rect 25060 14252 26012 14308
rect 26068 14252 26078 14308
rect 34738 14140 34748 14196
rect 34804 14140 39340 14196
rect 39396 14140 39406 14196
rect 19826 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20110 14140
rect 30034 14028 30044 14084
rect 30100 14028 30828 14084
rect 30884 14028 38668 14084
rect 38612 13972 38668 14028
rect 18162 13916 18172 13972
rect 18228 13916 23996 13972
rect 24052 13916 24062 13972
rect 25554 13916 25564 13972
rect 25620 13916 26572 13972
rect 26628 13916 26638 13972
rect 31826 13916 31836 13972
rect 31892 13916 35196 13972
rect 35252 13916 35532 13972
rect 35588 13916 35598 13972
rect 38612 13916 46956 13972
rect 47012 13916 47022 13972
rect 16930 13804 16940 13860
rect 16996 13804 17836 13860
rect 17892 13804 17902 13860
rect 23846 13804 23884 13860
rect 23940 13804 23950 13860
rect 24108 13804 33740 13860
rect 33796 13804 33806 13860
rect 35746 13804 35756 13860
rect 35812 13804 36204 13860
rect 36260 13804 36270 13860
rect 16818 13692 16828 13748
rect 16884 13692 17948 13748
rect 18004 13692 18014 13748
rect 19618 13692 19628 13748
rect 19684 13692 20636 13748
rect 20692 13692 20702 13748
rect 14018 13580 14028 13636
rect 14084 13580 15260 13636
rect 15316 13580 16716 13636
rect 16772 13580 18732 13636
rect 18788 13580 18798 13636
rect 18946 13580 18956 13636
rect 19012 13580 20188 13636
rect 20244 13580 20254 13636
rect 24108 13524 24164 13804
rect 24322 13692 24332 13748
rect 24388 13692 26460 13748
rect 26516 13692 27972 13748
rect 33618 13692 33628 13748
rect 33684 13692 34412 13748
rect 34468 13692 34478 13748
rect 44930 13692 44940 13748
rect 44996 13692 45388 13748
rect 45444 13692 45454 13748
rect 25442 13580 25452 13636
rect 25508 13580 25518 13636
rect 26002 13580 26012 13636
rect 26068 13580 27692 13636
rect 27748 13580 27758 13636
rect 19394 13468 19404 13524
rect 19460 13468 24220 13524
rect 24276 13468 24286 13524
rect 25452 13412 25508 13580
rect 27916 13524 27972 13692
rect 33730 13580 33740 13636
rect 33796 13580 34076 13636
rect 34132 13580 34142 13636
rect 38770 13580 38780 13636
rect 38836 13580 44268 13636
rect 44324 13580 45052 13636
rect 45108 13580 45118 13636
rect 25666 13468 25676 13524
rect 25732 13468 27020 13524
rect 27076 13468 27086 13524
rect 27570 13468 27580 13524
rect 27636 13468 27972 13524
rect 28242 13468 28252 13524
rect 28308 13468 34188 13524
rect 34244 13468 34748 13524
rect 34804 13468 34814 13524
rect 36754 13468 36764 13524
rect 36820 13468 38556 13524
rect 38612 13468 38622 13524
rect 20150 13356 20188 13412
rect 20244 13356 20254 13412
rect 25452 13356 25788 13412
rect 25844 13356 26124 13412
rect 26180 13356 26190 13412
rect 26562 13356 26572 13412
rect 26628 13356 27132 13412
rect 27188 13356 27804 13412
rect 27860 13356 27870 13412
rect 4466 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4750 13356
rect 35186 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35470 13356
rect 22866 13244 22876 13300
rect 22932 13244 30268 13300
rect 30324 13244 30334 13300
rect 24546 13132 24556 13188
rect 24612 13132 25116 13188
rect 25172 13132 27692 13188
rect 27748 13132 27758 13188
rect 44706 13132 44716 13188
rect 44772 13132 45612 13188
rect 45668 13132 45678 13188
rect 21298 13020 21308 13076
rect 21364 13020 22092 13076
rect 22148 13020 22158 13076
rect 25666 13020 25676 13076
rect 25732 13020 26908 13076
rect 34178 13020 34188 13076
rect 34244 13020 35084 13076
rect 35140 13020 35150 13076
rect 37762 13020 37772 13076
rect 37828 13020 41132 13076
rect 41188 13020 41198 13076
rect 45714 13020 45724 13076
rect 45780 13020 47740 13076
rect 47796 13020 47806 13076
rect 26852 12852 26908 13020
rect 33954 12908 33964 12964
rect 34020 12908 34412 12964
rect 34468 12908 37436 12964
rect 37492 12908 37502 12964
rect 18162 12796 18172 12852
rect 18228 12796 19068 12852
rect 19124 12796 19134 12852
rect 19730 12796 19740 12852
rect 19796 12796 22092 12852
rect 22148 12796 22158 12852
rect 26852 12796 29372 12852
rect 29428 12796 29932 12852
rect 29988 12796 29998 12852
rect 34066 12796 34076 12852
rect 34132 12796 35084 12852
rect 35140 12796 35644 12852
rect 35700 12796 35710 12852
rect 34290 12684 34300 12740
rect 34356 12684 34636 12740
rect 34692 12684 34702 12740
rect 42018 12684 42028 12740
rect 42084 12684 42364 12740
rect 42420 12684 42430 12740
rect 29586 12572 29596 12628
rect 29652 12572 29820 12628
rect 29876 12572 30156 12628
rect 30212 12572 41916 12628
rect 41972 12572 42700 12628
rect 42756 12572 43148 12628
rect 43204 12572 43214 12628
rect 19826 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20110 12572
rect 30034 12460 30044 12516
rect 30100 12460 31724 12516
rect 31780 12460 32172 12516
rect 32228 12460 32238 12516
rect 16594 12348 16604 12404
rect 16660 12348 17500 12404
rect 17556 12348 17566 12404
rect 17938 12348 17948 12404
rect 18004 12348 18732 12404
rect 18788 12348 18798 12404
rect 20514 12348 20524 12404
rect 20580 12348 21308 12404
rect 21364 12348 21374 12404
rect 26786 12348 26796 12404
rect 26852 12348 33852 12404
rect 33908 12348 33918 12404
rect 17500 12292 17556 12348
rect 17500 12236 19740 12292
rect 19796 12236 19806 12292
rect 24098 12236 24108 12292
rect 24164 12236 24556 12292
rect 24612 12236 25676 12292
rect 25732 12236 25900 12292
rect 25956 12236 25966 12292
rect 27906 12236 27916 12292
rect 27972 12236 28476 12292
rect 28532 12236 28542 12292
rect 30268 12236 30380 12292
rect 30436 12236 30446 12292
rect 30604 12236 31612 12292
rect 31668 12236 31678 12292
rect 32162 12236 32172 12292
rect 32228 12236 42028 12292
rect 42084 12236 42094 12292
rect 16930 12124 16940 12180
rect 16996 12124 17948 12180
rect 18004 12124 18014 12180
rect 18834 12124 18844 12180
rect 18900 12124 20300 12180
rect 20356 12124 20366 12180
rect 23762 12012 23772 12068
rect 23828 12012 25116 12068
rect 25172 12012 25340 12068
rect 25396 12012 25406 12068
rect 30268 11956 30324 12236
rect 30604 12180 30660 12236
rect 32172 12180 32228 12236
rect 30594 12124 30604 12180
rect 30660 12124 30670 12180
rect 31154 12124 31164 12180
rect 31220 12124 32228 12180
rect 33618 12124 33628 12180
rect 33684 12124 37772 12180
rect 37828 12124 37838 12180
rect 34066 12012 34076 12068
rect 34132 12012 34636 12068
rect 34692 12012 34702 12068
rect 19730 11900 19740 11956
rect 19796 11900 20300 11956
rect 20356 11900 20366 11956
rect 25666 11900 25676 11956
rect 25732 11900 26796 11956
rect 26852 11900 26862 11956
rect 30268 11900 30940 11956
rect 30996 11900 31006 11956
rect 21746 11788 21756 11844
rect 21812 11788 25116 11844
rect 25172 11788 25788 11844
rect 25844 11788 25854 11844
rect 29138 11788 29148 11844
rect 29204 11788 30044 11844
rect 30100 11788 31164 11844
rect 31220 11788 31230 11844
rect 4466 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4750 11788
rect 35186 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35470 11788
rect 31042 11676 31052 11732
rect 31108 11676 31948 11732
rect 32004 11676 32014 11732
rect 38770 11676 38780 11732
rect 38836 11676 40236 11732
rect 40292 11676 40302 11732
rect 23650 11564 23660 11620
rect 23716 11564 24892 11620
rect 24948 11564 24958 11620
rect 38098 11564 38108 11620
rect 38164 11564 38892 11620
rect 38948 11564 38958 11620
rect 39106 11564 39116 11620
rect 39172 11564 39182 11620
rect 17714 11452 17724 11508
rect 17780 11452 18060 11508
rect 18116 11452 23212 11508
rect 23268 11452 23278 11508
rect 24210 11452 24220 11508
rect 24276 11452 32396 11508
rect 32452 11452 32462 11508
rect 32620 11452 35924 11508
rect 37650 11452 37660 11508
rect 37716 11452 38780 11508
rect 38836 11452 38846 11508
rect 24220 11396 24276 11452
rect 32620 11396 32676 11452
rect 35868 11396 35924 11452
rect 18722 11340 18732 11396
rect 18788 11340 21868 11396
rect 21924 11340 21934 11396
rect 22978 11340 22988 11396
rect 23044 11340 24276 11396
rect 25778 11340 25788 11396
rect 25844 11340 25854 11396
rect 26002 11340 26012 11396
rect 26068 11340 26684 11396
rect 26740 11340 26750 11396
rect 27794 11340 27804 11396
rect 27860 11340 28364 11396
rect 28420 11340 32676 11396
rect 33058 11340 33068 11396
rect 33124 11340 34300 11396
rect 34356 11340 35644 11396
rect 35700 11340 35710 11396
rect 35868 11340 38892 11396
rect 38948 11340 38958 11396
rect 25788 11284 25844 11340
rect 20626 11228 20636 11284
rect 20692 11228 21420 11284
rect 21476 11228 21486 11284
rect 25788 11228 27132 11284
rect 27188 11228 27198 11284
rect 34738 11228 34748 11284
rect 34804 11228 34972 11284
rect 35028 11228 36092 11284
rect 36148 11228 36158 11284
rect 38546 11228 38556 11284
rect 38612 11172 38668 11284
rect 39116 11172 39172 11564
rect 41122 11452 41132 11508
rect 41188 11452 42252 11508
rect 42308 11452 42318 11508
rect 40002 11340 40012 11396
rect 40068 11340 41468 11396
rect 41524 11340 43372 11396
rect 43428 11340 43438 11396
rect 41122 11228 41132 11284
rect 41188 11228 41198 11284
rect 41682 11228 41692 11284
rect 41748 11228 43484 11284
rect 43540 11228 43550 11284
rect 41132 11172 41188 11228
rect 16482 11116 16492 11172
rect 16548 11116 18060 11172
rect 18116 11116 18126 11172
rect 18834 11116 18844 11172
rect 18900 11116 19404 11172
rect 19460 11116 19470 11172
rect 23874 11116 23884 11172
rect 23940 11116 25676 11172
rect 25732 11116 25742 11172
rect 29586 11116 29596 11172
rect 29652 11116 30716 11172
rect 30772 11116 30782 11172
rect 35522 11116 35532 11172
rect 35588 11116 36988 11172
rect 37044 11116 37054 11172
rect 38612 11116 39676 11172
rect 39732 11116 41188 11172
rect 42466 11116 42476 11172
rect 42532 11116 44828 11172
rect 44884 11116 44894 11172
rect 26674 11004 26684 11060
rect 26740 11004 26908 11060
rect 34626 11004 34636 11060
rect 34692 11004 35868 11060
rect 35924 11004 35934 11060
rect 38882 11004 38892 11060
rect 38948 11004 38958 11060
rect 39554 11004 39564 11060
rect 39620 11004 40236 11060
rect 40292 11004 43820 11060
rect 43876 11004 43886 11060
rect 19826 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20110 11004
rect 26852 10948 26908 11004
rect 38892 10948 38948 11004
rect 16034 10892 16044 10948
rect 16100 10892 16604 10948
rect 16660 10892 17164 10948
rect 17220 10892 18620 10948
rect 18676 10892 18686 10948
rect 26852 10892 36092 10948
rect 36148 10892 36158 10948
rect 38892 10892 42868 10948
rect 42812 10836 42868 10892
rect 15026 10780 15036 10836
rect 15092 10780 17052 10836
rect 17108 10780 17612 10836
rect 17668 10780 18284 10836
rect 18340 10780 19180 10836
rect 19236 10780 19246 10836
rect 25452 10780 26012 10836
rect 26068 10780 26078 10836
rect 29810 10780 29820 10836
rect 29876 10780 30156 10836
rect 30212 10780 30222 10836
rect 38882 10780 38892 10836
rect 38948 10780 40572 10836
rect 40628 10780 41132 10836
rect 41188 10780 41198 10836
rect 42802 10780 42812 10836
rect 42868 10780 42878 10836
rect 25452 10612 25508 10780
rect 26674 10668 26684 10724
rect 26740 10668 28140 10724
rect 28196 10668 28206 10724
rect 30706 10668 30716 10724
rect 30772 10668 37660 10724
rect 37716 10668 40796 10724
rect 40852 10668 40862 10724
rect 42018 10668 42028 10724
rect 42084 10668 45948 10724
rect 46004 10668 46014 10724
rect 16930 10556 16940 10612
rect 16996 10556 18060 10612
rect 18116 10556 18126 10612
rect 23874 10556 23884 10612
rect 23940 10556 25452 10612
rect 25508 10556 25518 10612
rect 28018 10556 28028 10612
rect 28084 10556 29148 10612
rect 29204 10556 30828 10612
rect 30884 10556 30894 10612
rect 31266 10556 31276 10612
rect 31332 10556 31948 10612
rect 32004 10556 39564 10612
rect 39620 10556 40012 10612
rect 40068 10556 40078 10612
rect 40226 10556 40236 10612
rect 40292 10556 41356 10612
rect 41412 10556 41422 10612
rect 27458 10444 27468 10500
rect 27524 10444 29260 10500
rect 29316 10444 29326 10500
rect 35858 10444 35868 10500
rect 35924 10444 36372 10500
rect 36316 10388 36372 10444
rect 34626 10332 34636 10388
rect 34692 10332 35756 10388
rect 35812 10332 35822 10388
rect 36306 10332 36316 10388
rect 36372 10332 37324 10388
rect 37380 10332 37390 10388
rect 44258 10332 44268 10388
rect 44324 10332 44940 10388
rect 44996 10332 45388 10388
rect 45444 10332 45454 10388
rect 21522 10220 21532 10276
rect 21588 10220 22092 10276
rect 22148 10220 32508 10276
rect 32564 10220 32574 10276
rect 4466 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4750 10220
rect 35186 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35470 10220
rect 19618 10108 19628 10164
rect 19684 10108 20972 10164
rect 21028 10108 23100 10164
rect 23156 10108 24556 10164
rect 24612 10108 24622 10164
rect 27122 10108 27132 10164
rect 27188 10108 27198 10164
rect 27794 10108 27804 10164
rect 27860 10108 28588 10164
rect 28644 10108 28654 10164
rect 35532 10108 36092 10164
rect 36148 10108 36158 10164
rect 37202 10108 37212 10164
rect 37268 10108 37548 10164
rect 37604 10108 37614 10164
rect 41234 10108 41244 10164
rect 41300 10108 41310 10164
rect 24434 9996 24444 10052
rect 24500 9996 25452 10052
rect 25508 9996 25518 10052
rect 0 9940 800 9968
rect 0 9884 5964 9940
rect 6020 9884 6030 9940
rect 22642 9884 22652 9940
rect 22708 9884 24668 9940
rect 24724 9884 24734 9940
rect 0 9856 800 9884
rect 27132 9828 27188 10108
rect 35532 10052 35588 10108
rect 31154 9996 31164 10052
rect 31220 9996 31948 10052
rect 32004 9996 32396 10052
rect 32452 9996 32462 10052
rect 33170 9996 33180 10052
rect 33236 9996 33852 10052
rect 33908 9996 34524 10052
rect 34580 9996 34590 10052
rect 35410 9996 35420 10052
rect 35476 9996 35588 10052
rect 41244 10052 41300 10108
rect 41244 9996 42364 10052
rect 42420 9996 42430 10052
rect 44818 9884 44828 9940
rect 44884 9884 45836 9940
rect 45892 9884 45902 9940
rect 27132 9772 35084 9828
rect 35140 9772 36540 9828
rect 36596 9772 36606 9828
rect 25442 9660 25452 9716
rect 25508 9660 26012 9716
rect 26068 9660 26572 9716
rect 26628 9660 26638 9716
rect 30258 9660 30268 9716
rect 30324 9660 31052 9716
rect 31108 9660 31118 9716
rect 41570 9660 41580 9716
rect 41636 9660 42700 9716
rect 42756 9660 42766 9716
rect 44930 9660 44940 9716
rect 44996 9660 45388 9716
rect 45444 9660 45454 9716
rect 19058 9548 19068 9604
rect 19124 9548 21980 9604
rect 22036 9548 22046 9604
rect 45266 9548 45276 9604
rect 45332 9548 46620 9604
rect 46676 9548 46686 9604
rect 49200 9492 50000 9520
rect 47618 9436 47628 9492
rect 47684 9436 48188 9492
rect 48244 9436 50000 9492
rect 19826 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20110 9436
rect 49200 9408 50000 9436
rect 33506 9324 33516 9380
rect 33572 9324 35868 9380
rect 35924 9324 37324 9380
rect 37380 9324 38108 9380
rect 38164 9324 38174 9380
rect 18610 9212 18620 9268
rect 18676 9212 19852 9268
rect 19908 9212 20412 9268
rect 20468 9212 20478 9268
rect 34178 9212 34188 9268
rect 34244 9212 35084 9268
rect 35140 9212 35150 9268
rect 16482 9100 16492 9156
rect 16548 9100 17948 9156
rect 18004 9100 18014 9156
rect 18386 9100 18396 9156
rect 18452 9100 19068 9156
rect 19124 9100 19134 9156
rect 21298 9100 21308 9156
rect 21364 9100 22092 9156
rect 22148 9100 22158 9156
rect 31490 9100 31500 9156
rect 31556 9100 34076 9156
rect 34132 9100 34142 9156
rect 39778 9100 39788 9156
rect 39844 9100 41692 9156
rect 41748 9100 41758 9156
rect 17826 8988 17836 9044
rect 17892 8988 23772 9044
rect 23828 8988 23838 9044
rect 33394 8988 33404 9044
rect 33460 8988 33852 9044
rect 33908 8988 33918 9044
rect 24882 8876 24892 8932
rect 24948 8876 25788 8932
rect 25844 8876 37772 8932
rect 37828 8876 38668 8932
rect 43474 8876 43484 8932
rect 43540 8876 44492 8932
rect 44548 8876 45724 8932
rect 45780 8876 45790 8932
rect 38612 8708 38668 8876
rect 42466 8764 42476 8820
rect 42532 8764 43820 8820
rect 43876 8764 43886 8820
rect 38612 8652 44044 8708
rect 44100 8652 45052 8708
rect 45108 8652 45118 8708
rect 4466 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4750 8652
rect 35186 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35470 8652
rect 19058 8540 19068 8596
rect 19124 8540 20300 8596
rect 20356 8540 20366 8596
rect 42354 8428 42364 8484
rect 42420 8428 42430 8484
rect 42364 8372 42420 8428
rect 22978 8316 22988 8372
rect 23044 8316 23772 8372
rect 23828 8316 26684 8372
rect 26740 8316 26750 8372
rect 31602 8316 31612 8372
rect 31668 8316 37660 8372
rect 37716 8316 37726 8372
rect 41794 8316 41804 8372
rect 41860 8316 43260 8372
rect 43316 8316 44828 8372
rect 44884 8316 44894 8372
rect 45042 8316 45052 8372
rect 45108 8316 46060 8372
rect 46116 8316 46126 8372
rect 17938 8204 17948 8260
rect 18004 8204 18732 8260
rect 18788 8204 18798 8260
rect 18946 8204 18956 8260
rect 19012 8204 23996 8260
rect 24052 8204 24062 8260
rect 24322 8204 24332 8260
rect 24388 8204 25452 8260
rect 25508 8204 25518 8260
rect 32722 8204 32732 8260
rect 32788 8204 34636 8260
rect 34692 8204 35644 8260
rect 35700 8204 35710 8260
rect 39666 8204 39676 8260
rect 39732 8204 43148 8260
rect 43204 8204 43214 8260
rect 25004 8036 25060 8204
rect 37548 8092 40236 8148
rect 40292 8092 40302 8148
rect 41234 8092 41244 8148
rect 41300 8092 42140 8148
rect 42196 8092 42206 8148
rect 42690 8092 42700 8148
rect 42756 8092 43372 8148
rect 43428 8092 43820 8148
rect 43876 8092 43886 8148
rect 37548 8036 37604 8092
rect 41244 8036 41300 8092
rect 22754 7980 22764 8036
rect 22820 7980 23884 8036
rect 23940 7980 23950 8036
rect 24994 7980 25004 8036
rect 25060 7980 25070 8036
rect 34402 7980 34412 8036
rect 34468 7980 36204 8036
rect 36260 7980 36428 8036
rect 36484 7980 37100 8036
rect 37156 7980 37166 8036
rect 37538 7980 37548 8036
rect 37604 7980 37614 8036
rect 38994 7980 39004 8036
rect 39060 7980 41300 8036
rect 41570 7980 41580 8036
rect 41636 7980 42028 8036
rect 42084 7980 42252 8036
rect 42308 7980 42318 8036
rect 19826 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20110 7868
rect 22082 7756 22092 7812
rect 22148 7756 35084 7812
rect 35140 7756 35150 7812
rect 35298 7756 35308 7812
rect 35364 7756 36540 7812
rect 36596 7756 36606 7812
rect 17042 7644 17052 7700
rect 17108 7644 18060 7700
rect 18116 7644 18126 7700
rect 27010 7644 27020 7700
rect 27076 7644 29036 7700
rect 29092 7644 30268 7700
rect 30324 7644 31612 7700
rect 31668 7644 31678 7700
rect 34860 7644 35756 7700
rect 35812 7644 35822 7700
rect 38882 7644 38892 7700
rect 38948 7644 41468 7700
rect 41524 7644 41534 7700
rect 34860 7588 34916 7644
rect 25890 7532 25900 7588
rect 25956 7532 28924 7588
rect 28980 7532 28990 7588
rect 33170 7532 33180 7588
rect 33236 7532 33740 7588
rect 33796 7532 34748 7588
rect 34804 7532 34916 7588
rect 35410 7532 35420 7588
rect 35476 7532 36092 7588
rect 36148 7532 37996 7588
rect 38052 7532 38668 7588
rect 38724 7532 39564 7588
rect 39620 7532 39630 7588
rect 42130 7532 42140 7588
rect 42196 7532 43484 7588
rect 43540 7532 43932 7588
rect 43988 7532 43998 7588
rect 18162 7420 18172 7476
rect 18228 7420 23884 7476
rect 23940 7420 23950 7476
rect 24210 7420 24220 7476
rect 24276 7420 25228 7476
rect 25284 7420 25294 7476
rect 30034 7420 30044 7476
rect 30100 7420 31500 7476
rect 31556 7420 31566 7476
rect 34402 7420 34412 7476
rect 34468 7420 34860 7476
rect 34916 7420 34926 7476
rect 35746 7420 35756 7476
rect 35812 7420 35822 7476
rect 43138 7420 43148 7476
rect 43204 7420 44044 7476
rect 44100 7420 44380 7476
rect 44436 7420 44446 7476
rect 35756 7364 35812 7420
rect 16594 7308 16604 7364
rect 16660 7308 17500 7364
rect 17556 7308 18396 7364
rect 18452 7308 22876 7364
rect 22932 7308 22942 7364
rect 24882 7308 24892 7364
rect 24948 7308 25340 7364
rect 25396 7308 25406 7364
rect 26852 7308 35812 7364
rect 26852 7252 26908 7308
rect 22194 7196 22204 7252
rect 22260 7196 26908 7252
rect 30818 7196 30828 7252
rect 30884 7196 32172 7252
rect 32228 7196 32238 7252
rect 41234 7196 41244 7252
rect 41300 7196 41692 7252
rect 41748 7196 41758 7252
rect 4466 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4750 7084
rect 35186 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35470 7084
rect 23762 6860 23772 6916
rect 23828 6860 25788 6916
rect 25844 6860 25854 6916
rect 41794 6860 41804 6916
rect 41860 6860 42476 6916
rect 42532 6860 42542 6916
rect 43250 6860 43260 6916
rect 43316 6860 44828 6916
rect 44884 6860 44894 6916
rect 21970 6748 21980 6804
rect 22036 6748 25116 6804
rect 25172 6748 25182 6804
rect 27346 6748 27356 6804
rect 27412 6748 27692 6804
rect 27748 6748 28476 6804
rect 28532 6748 30380 6804
rect 30436 6748 30446 6804
rect 31266 6748 31276 6804
rect 31332 6748 32172 6804
rect 32228 6748 33068 6804
rect 33124 6748 33134 6804
rect 34402 6748 34412 6804
rect 34468 6748 34748 6804
rect 34804 6748 34814 6804
rect 40114 6748 40124 6804
rect 40180 6748 40684 6804
rect 40740 6748 40750 6804
rect 42130 6748 42140 6804
rect 42196 6748 42588 6804
rect 42644 6748 43596 6804
rect 43652 6748 43662 6804
rect 15362 6636 15372 6692
rect 15428 6636 16492 6692
rect 16548 6636 16558 6692
rect 19394 6636 19404 6692
rect 19460 6636 19740 6692
rect 19796 6636 21308 6692
rect 21364 6636 22540 6692
rect 22596 6636 22606 6692
rect 22978 6636 22988 6692
rect 23044 6636 23324 6692
rect 23380 6636 23390 6692
rect 24322 6636 24332 6692
rect 24388 6636 26124 6692
rect 26180 6636 26190 6692
rect 28354 6636 28364 6692
rect 28420 6636 29260 6692
rect 29316 6636 30044 6692
rect 30100 6636 30110 6692
rect 34290 6636 34300 6692
rect 34356 6636 34860 6692
rect 34916 6636 35308 6692
rect 35364 6636 35374 6692
rect 35970 6636 35980 6692
rect 36036 6636 36876 6692
rect 36932 6636 36942 6692
rect 41346 6636 41356 6692
rect 41412 6636 41692 6692
rect 41748 6636 43820 6692
rect 43876 6636 44492 6692
rect 44548 6636 44558 6692
rect 35308 6580 35364 6636
rect 24658 6524 24668 6580
rect 24724 6524 26012 6580
rect 26068 6524 26684 6580
rect 26740 6524 26750 6580
rect 28578 6524 28588 6580
rect 28644 6524 30268 6580
rect 30324 6524 31052 6580
rect 31108 6524 31724 6580
rect 31780 6524 31790 6580
rect 35308 6524 36092 6580
rect 36148 6524 36158 6580
rect 36530 6524 36540 6580
rect 36596 6524 37548 6580
rect 37604 6524 37614 6580
rect 37762 6524 37772 6580
rect 37828 6524 38780 6580
rect 38836 6524 39788 6580
rect 39844 6524 39854 6580
rect 40450 6524 40460 6580
rect 40516 6524 42252 6580
rect 42308 6524 42318 6580
rect 44258 6524 44268 6580
rect 44324 6524 46956 6580
rect 47012 6524 47022 6580
rect 23426 6412 23436 6468
rect 23492 6412 28364 6468
rect 28420 6412 30492 6468
rect 30548 6412 32844 6468
rect 32900 6412 32910 6468
rect 39666 6412 39676 6468
rect 39732 6412 39742 6468
rect 40002 6412 40012 6468
rect 40068 6412 40908 6468
rect 40964 6412 40974 6468
rect 41234 6412 41244 6468
rect 41300 6412 42812 6468
rect 42868 6412 42878 6468
rect 43362 6412 43372 6468
rect 43428 6412 44156 6468
rect 44212 6412 44222 6468
rect 39676 6356 39732 6412
rect 22418 6300 22428 6356
rect 22484 6300 23660 6356
rect 23716 6300 25564 6356
rect 25620 6300 25630 6356
rect 26852 6300 36540 6356
rect 36596 6300 36606 6356
rect 38322 6300 38332 6356
rect 38388 6300 39732 6356
rect 39890 6300 39900 6356
rect 39956 6300 40460 6356
rect 40516 6300 40526 6356
rect 19826 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20110 6300
rect 26852 6244 26908 6300
rect 20626 6188 20636 6244
rect 20692 6188 21532 6244
rect 21588 6188 26908 6244
rect 27010 6188 27020 6244
rect 27076 6188 29260 6244
rect 29316 6188 31332 6244
rect 32610 6188 32620 6244
rect 32676 6188 34076 6244
rect 34132 6188 36988 6244
rect 37044 6188 37054 6244
rect 40226 6188 40236 6244
rect 40292 6188 41804 6244
rect 41860 6188 41870 6244
rect 31276 6132 31332 6188
rect 20962 6076 20972 6132
rect 21028 6076 21644 6132
rect 21700 6076 21710 6132
rect 22530 6076 22540 6132
rect 22596 6076 24668 6132
rect 24724 6076 25340 6132
rect 25396 6076 25406 6132
rect 26852 6076 27916 6132
rect 27972 6076 29820 6132
rect 29876 6076 29886 6132
rect 31266 6076 31276 6132
rect 31332 6076 33068 6132
rect 33124 6076 33134 6132
rect 35830 6076 35868 6132
rect 35924 6076 38052 6132
rect 38546 6076 38556 6132
rect 38612 6076 40012 6132
rect 40068 6076 41020 6132
rect 41076 6076 41086 6132
rect 26852 6020 26908 6076
rect 26012 5964 26908 6020
rect 29586 5964 29596 6020
rect 29652 5964 31500 6020
rect 31556 5964 33740 6020
rect 33796 5964 34972 6020
rect 35028 5964 36316 6020
rect 36372 5964 36382 6020
rect 37762 5964 37772 6020
rect 37828 5964 37838 6020
rect 26012 5908 26068 5964
rect 18386 5852 18396 5908
rect 18452 5852 18844 5908
rect 18900 5852 18910 5908
rect 19954 5852 19964 5908
rect 20020 5852 20524 5908
rect 20580 5852 20590 5908
rect 26002 5852 26012 5908
rect 26068 5852 26078 5908
rect 26226 5852 26236 5908
rect 26292 5852 27356 5908
rect 27412 5852 27692 5908
rect 27748 5852 27758 5908
rect 29026 5852 29036 5908
rect 29092 5852 29708 5908
rect 29764 5852 30268 5908
rect 30324 5852 30334 5908
rect 33506 5852 33516 5908
rect 33572 5852 35420 5908
rect 35476 5852 35486 5908
rect 37772 5796 37828 5964
rect 37996 5908 38052 6076
rect 38434 5964 38444 6020
rect 38500 5964 39900 6020
rect 39956 5964 41580 6020
rect 41636 5964 41646 6020
rect 41906 5964 41916 6020
rect 41972 5964 43708 6020
rect 43764 5964 43774 6020
rect 37996 5852 39004 5908
rect 39060 5852 39452 5908
rect 39508 5852 39518 5908
rect 23314 5740 23324 5796
rect 23380 5740 25452 5796
rect 25508 5740 25518 5796
rect 26338 5740 26348 5796
rect 26404 5740 27804 5796
rect 27860 5740 27870 5796
rect 35298 5740 35308 5796
rect 35364 5740 36652 5796
rect 36708 5740 36718 5796
rect 37772 5740 38668 5796
rect 38724 5740 41244 5796
rect 41300 5740 41310 5796
rect 36652 5684 36708 5740
rect 24770 5628 24780 5684
rect 24836 5628 27020 5684
rect 27076 5628 27086 5684
rect 35522 5628 35532 5684
rect 35588 5628 36092 5684
rect 36148 5628 36158 5684
rect 36652 5628 38444 5684
rect 38500 5628 38510 5684
rect 25442 5516 25452 5572
rect 25508 5516 26460 5572
rect 26516 5516 26526 5572
rect 4466 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4750 5516
rect 35186 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35470 5516
rect 18610 5404 18620 5460
rect 18676 5404 21420 5460
rect 21476 5404 21486 5460
rect 32386 5292 32396 5348
rect 32452 5292 35308 5348
rect 35364 5292 38332 5348
rect 38388 5292 38398 5348
rect 22866 5180 22876 5236
rect 22932 5180 25004 5236
rect 25060 5180 25070 5236
rect 31042 5180 31052 5236
rect 31108 5180 32732 5236
rect 32788 5180 32798 5236
rect 35830 5180 35868 5236
rect 35924 5180 35934 5236
rect 40786 5180 40796 5236
rect 40852 5180 41692 5236
rect 41748 5180 41758 5236
rect 16482 5068 16492 5124
rect 16548 5068 17948 5124
rect 18004 5068 18014 5124
rect 23314 5068 23324 5124
rect 23380 5068 24108 5124
rect 24164 5068 24174 5124
rect 28130 5068 28140 5124
rect 28196 5068 29036 5124
rect 29092 5068 29102 5124
rect 29922 5068 29932 5124
rect 29988 5068 33180 5124
rect 33236 5068 36092 5124
rect 36148 5068 36158 5124
rect 37538 5068 37548 5124
rect 37604 5068 40012 5124
rect 40068 5068 40078 5124
rect 44034 5068 44044 5124
rect 44100 5068 47068 5124
rect 47124 5068 47134 5124
rect 21522 4956 21532 5012
rect 21588 4956 22204 5012
rect 22260 4956 22270 5012
rect 25554 4956 25564 5012
rect 25620 4956 26572 5012
rect 26628 4956 27356 5012
rect 27412 4956 27422 5012
rect 33506 4956 33516 5012
rect 33572 4956 40124 5012
rect 40180 4956 40190 5012
rect 36418 4844 36428 4900
rect 36484 4844 38444 4900
rect 38500 4844 38510 4900
rect 42914 4844 42924 4900
rect 42980 4844 46284 4900
rect 46340 4844 46350 4900
rect 19826 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20110 4732
rect 39218 4284 39228 4340
rect 39284 4284 40012 4340
rect 40068 4284 40796 4340
rect 40852 4284 40862 4340
rect 45938 4284 45948 4340
rect 46004 4284 47628 4340
rect 47684 4284 47694 4340
rect 4466 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4750 3948
rect 35186 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35470 3948
rect 49200 3668 50000 3696
rect 48290 3612 48300 3668
rect 48356 3612 50000 3668
rect 49200 3584 50000 3612
rect 19826 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20110 3164
<< via3 >>
rect 19836 56420 19892 56476
rect 19940 56420 19996 56476
rect 20044 56420 20100 56476
rect 4476 55636 4532 55692
rect 4580 55636 4636 55692
rect 4684 55636 4740 55692
rect 35196 55636 35252 55692
rect 35300 55636 35356 55692
rect 35404 55636 35460 55692
rect 22204 55020 22260 55076
rect 19836 54852 19892 54908
rect 19940 54852 19996 54908
rect 20044 54852 20100 54908
rect 35868 54460 35924 54516
rect 4476 54068 4532 54124
rect 4580 54068 4636 54124
rect 4684 54068 4740 54124
rect 35196 54068 35252 54124
rect 35300 54068 35356 54124
rect 35404 54068 35460 54124
rect 22204 54012 22260 54068
rect 38668 53788 38724 53844
rect 19836 53284 19892 53340
rect 19940 53284 19996 53340
rect 20044 53284 20100 53340
rect 4476 52500 4532 52556
rect 4580 52500 4636 52556
rect 4684 52500 4740 52556
rect 35196 52500 35252 52556
rect 35300 52500 35356 52556
rect 35404 52500 35460 52556
rect 34748 52220 34804 52276
rect 38668 51996 38724 52052
rect 19836 51716 19892 51772
rect 19940 51716 19996 51772
rect 20044 51716 20100 51772
rect 35868 51548 35924 51604
rect 4476 50932 4532 50988
rect 4580 50932 4636 50988
rect 4684 50932 4740 50988
rect 35196 50932 35252 50988
rect 35300 50932 35356 50988
rect 35404 50932 35460 50988
rect 19836 50148 19892 50204
rect 19940 50148 19996 50204
rect 20044 50148 20100 50204
rect 4476 49364 4532 49420
rect 4580 49364 4636 49420
rect 4684 49364 4740 49420
rect 35196 49364 35252 49420
rect 35300 49364 35356 49420
rect 35404 49364 35460 49420
rect 19836 48580 19892 48636
rect 19940 48580 19996 48636
rect 20044 48580 20100 48636
rect 34748 48300 34804 48356
rect 4476 47796 4532 47852
rect 4580 47796 4636 47852
rect 4684 47796 4740 47852
rect 35196 47796 35252 47852
rect 35300 47796 35356 47852
rect 35404 47796 35460 47852
rect 22540 47068 22596 47124
rect 19836 47012 19892 47068
rect 19940 47012 19996 47068
rect 20044 47012 20100 47068
rect 4476 46228 4532 46284
rect 4580 46228 4636 46284
rect 4684 46228 4740 46284
rect 35196 46228 35252 46284
rect 35300 46228 35356 46284
rect 35404 46228 35460 46284
rect 21756 45500 21812 45556
rect 19836 45444 19892 45500
rect 19940 45444 19996 45500
rect 20044 45444 20100 45500
rect 10108 45164 10164 45220
rect 4476 44660 4532 44716
rect 4580 44660 4636 44716
rect 4684 44660 4740 44716
rect 35196 44660 35252 44716
rect 35300 44660 35356 44716
rect 35404 44660 35460 44716
rect 19836 43876 19892 43932
rect 19940 43876 19996 43932
rect 20044 43876 20100 43932
rect 4476 43092 4532 43148
rect 4580 43092 4636 43148
rect 4684 43092 4740 43148
rect 35196 43092 35252 43148
rect 35300 43092 35356 43148
rect 35404 43092 35460 43148
rect 19836 42308 19892 42364
rect 19940 42308 19996 42364
rect 20044 42308 20100 42364
rect 8764 42140 8820 42196
rect 4476 41524 4532 41580
rect 4580 41524 4636 41580
rect 4684 41524 4740 41580
rect 35196 41524 35252 41580
rect 35300 41524 35356 41580
rect 35404 41524 35460 41580
rect 19836 40740 19892 40796
rect 19940 40740 19996 40796
rect 20044 40740 20100 40796
rect 4476 39956 4532 40012
rect 4580 39956 4636 40012
rect 4684 39956 4740 40012
rect 35196 39956 35252 40012
rect 35300 39956 35356 40012
rect 35404 39956 35460 40012
rect 19836 39172 19892 39228
rect 19940 39172 19996 39228
rect 20044 39172 20100 39228
rect 4476 38388 4532 38444
rect 4580 38388 4636 38444
rect 4684 38388 4740 38444
rect 35196 38388 35252 38444
rect 35300 38388 35356 38444
rect 35404 38388 35460 38444
rect 19404 37772 19460 37828
rect 19836 37604 19892 37660
rect 19940 37604 19996 37660
rect 20044 37604 20100 37660
rect 8988 37212 9044 37268
rect 11452 36988 11508 37044
rect 21532 36876 21588 36932
rect 4476 36820 4532 36876
rect 4580 36820 4636 36876
rect 4684 36820 4740 36876
rect 35196 36820 35252 36876
rect 35300 36820 35356 36876
rect 35404 36820 35460 36876
rect 19404 36764 19460 36820
rect 21532 36428 21588 36484
rect 19836 36036 19892 36092
rect 19940 36036 19996 36092
rect 20044 36036 20100 36092
rect 10108 35756 10164 35812
rect 4476 35252 4532 35308
rect 4580 35252 4636 35308
rect 4684 35252 4740 35308
rect 35196 35252 35252 35308
rect 35300 35252 35356 35308
rect 35404 35252 35460 35308
rect 9436 35196 9492 35252
rect 9548 34972 9604 35028
rect 19836 34468 19892 34524
rect 19940 34468 19996 34524
rect 20044 34468 20100 34524
rect 33852 34188 33908 34244
rect 24332 34076 24388 34132
rect 22540 33964 22596 34020
rect 22092 33852 22148 33908
rect 20748 33740 20804 33796
rect 4476 33684 4532 33740
rect 4580 33684 4636 33740
rect 4684 33684 4740 33740
rect 35196 33684 35252 33740
rect 35300 33684 35356 33740
rect 35404 33684 35460 33740
rect 36988 33628 37044 33684
rect 9436 33068 9492 33124
rect 19836 32900 19892 32956
rect 19940 32900 19996 32956
rect 20044 32900 20100 32956
rect 22092 32508 22148 32564
rect 4476 32116 4532 32172
rect 4580 32116 4636 32172
rect 4684 32116 4740 32172
rect 35196 32116 35252 32172
rect 35300 32116 35356 32172
rect 35404 32116 35460 32172
rect 9436 32060 9492 32116
rect 17948 31724 18004 31780
rect 24332 31724 24388 31780
rect 8988 31612 9044 31668
rect 9436 31612 9492 31668
rect 20748 31612 20804 31668
rect 19836 31332 19892 31388
rect 19940 31332 19996 31388
rect 20044 31332 20100 31388
rect 18732 30828 18788 30884
rect 4476 30548 4532 30604
rect 4580 30548 4636 30604
rect 4684 30548 4740 30604
rect 35196 30548 35252 30604
rect 35300 30548 35356 30604
rect 35404 30548 35460 30604
rect 36428 29932 36484 29988
rect 19836 29764 19892 29820
rect 19940 29764 19996 29820
rect 20044 29764 20100 29820
rect 8764 29596 8820 29652
rect 33852 29484 33908 29540
rect 4476 28980 4532 29036
rect 4580 28980 4636 29036
rect 4684 28980 4740 29036
rect 35196 28980 35252 29036
rect 35300 28980 35356 29036
rect 35404 28980 35460 29036
rect 9548 28812 9604 28868
rect 21756 28812 21812 28868
rect 11452 28364 11508 28420
rect 34972 28252 35028 28308
rect 19836 28196 19892 28252
rect 19940 28196 19996 28252
rect 20044 28196 20100 28252
rect 18732 27580 18788 27636
rect 4476 27412 4532 27468
rect 4580 27412 4636 27468
rect 4684 27412 4740 27468
rect 35196 27412 35252 27468
rect 35300 27412 35356 27468
rect 35404 27412 35460 27468
rect 19068 26908 19124 26964
rect 36428 26796 36484 26852
rect 19068 26684 19124 26740
rect 19836 26628 19892 26684
rect 19940 26628 19996 26684
rect 20044 26628 20100 26684
rect 17948 26460 18004 26516
rect 33852 26460 33908 26516
rect 18620 26348 18676 26404
rect 34972 26012 35028 26068
rect 4476 25844 4532 25900
rect 4580 25844 4636 25900
rect 4684 25844 4740 25900
rect 35196 25844 35252 25900
rect 35300 25844 35356 25900
rect 35404 25844 35460 25900
rect 35980 25564 36036 25620
rect 18620 25452 18676 25508
rect 23212 25452 23268 25508
rect 14364 25228 14420 25284
rect 36876 25116 36932 25172
rect 19836 25060 19892 25116
rect 19940 25060 19996 25116
rect 20044 25060 20100 25116
rect 35980 24556 36036 24612
rect 4476 24276 4532 24332
rect 4580 24276 4636 24332
rect 4684 24276 4740 24332
rect 35196 24276 35252 24332
rect 35300 24276 35356 24332
rect 35404 24276 35460 24332
rect 14924 23884 14980 23940
rect 19836 23492 19892 23548
rect 19940 23492 19996 23548
rect 20044 23492 20100 23548
rect 14924 23436 14980 23492
rect 23212 23436 23268 23492
rect 13244 23100 13300 23156
rect 14364 22876 14420 22932
rect 4476 22708 4532 22764
rect 4580 22708 4636 22764
rect 4684 22708 4740 22764
rect 35196 22708 35252 22764
rect 35300 22708 35356 22764
rect 35404 22708 35460 22764
rect 34860 22652 34916 22708
rect 35868 22652 35924 22708
rect 13580 22204 13636 22260
rect 11116 21980 11172 22036
rect 14028 21980 14084 22036
rect 19836 21924 19892 21980
rect 19940 21924 19996 21980
rect 20044 21924 20100 21980
rect 13244 21868 13300 21924
rect 15596 21756 15652 21812
rect 22652 21644 22708 21700
rect 14028 21308 14084 21364
rect 14364 21308 14420 21364
rect 11116 21196 11172 21252
rect 4476 21140 4532 21196
rect 4580 21140 4636 21196
rect 4684 21140 4740 21196
rect 35196 21140 35252 21196
rect 35300 21140 35356 21196
rect 35404 21140 35460 21196
rect 15596 21084 15652 21140
rect 43148 20636 43204 20692
rect 35980 20524 36036 20580
rect 19836 20356 19892 20412
rect 19940 20356 19996 20412
rect 20044 20356 20100 20412
rect 38892 20188 38948 20244
rect 13244 20076 13300 20132
rect 22652 20076 22708 20132
rect 19628 19628 19684 19684
rect 4476 19572 4532 19628
rect 4580 19572 4636 19628
rect 4684 19572 4740 19628
rect 35196 19572 35252 19628
rect 35300 19572 35356 19628
rect 35404 19572 35460 19628
rect 13580 19292 13636 19348
rect 35980 19292 36036 19348
rect 19836 18788 19892 18844
rect 19940 18788 19996 18844
rect 20044 18788 20100 18844
rect 44380 18284 44436 18340
rect 44380 18060 44436 18116
rect 4476 18004 4532 18060
rect 4580 18004 4636 18060
rect 4684 18004 4740 18060
rect 35196 18004 35252 18060
rect 35300 18004 35356 18060
rect 35404 18004 35460 18060
rect 19628 17612 19684 17668
rect 44380 17500 44436 17556
rect 19836 17220 19892 17276
rect 19940 17220 19996 17276
rect 20044 17220 20100 17276
rect 26908 17164 26964 17220
rect 35980 16828 36036 16884
rect 4476 16436 4532 16492
rect 4580 16436 4636 16492
rect 4684 16436 4740 16492
rect 35196 16436 35252 16492
rect 35300 16436 35356 16492
rect 35404 16436 35460 16492
rect 42924 16380 42980 16436
rect 35868 16156 35924 16212
rect 19628 15708 19684 15764
rect 35868 15708 35924 15764
rect 19836 15652 19892 15708
rect 19940 15652 19996 15708
rect 20044 15652 20100 15708
rect 34860 15484 34916 15540
rect 20188 15260 20244 15316
rect 23884 15148 23940 15204
rect 26908 14924 26964 14980
rect 4476 14868 4532 14924
rect 4580 14868 4636 14924
rect 4684 14868 4740 14924
rect 38892 14924 38948 14980
rect 35196 14868 35252 14924
rect 35300 14868 35356 14924
rect 35404 14868 35460 14924
rect 42924 14812 42980 14868
rect 19836 14084 19892 14140
rect 19940 14084 19996 14140
rect 20044 14084 20100 14140
rect 23884 13804 23940 13860
rect 20188 13356 20244 13412
rect 4476 13300 4532 13356
rect 4580 13300 4636 13356
rect 4684 13300 4740 13356
rect 35196 13300 35252 13356
rect 35300 13300 35356 13356
rect 35404 13300 35460 13356
rect 43148 12572 43204 12628
rect 19836 12516 19892 12572
rect 19940 12516 19996 12572
rect 20044 12516 20100 12572
rect 4476 11732 4532 11788
rect 4580 11732 4636 11788
rect 4684 11732 4740 11788
rect 35196 11732 35252 11788
rect 35300 11732 35356 11788
rect 35404 11732 35460 11788
rect 38892 11564 38948 11620
rect 38892 11004 38948 11060
rect 19836 10948 19892 11004
rect 19940 10948 19996 11004
rect 20044 10948 20100 11004
rect 4476 10164 4532 10220
rect 4580 10164 4636 10220
rect 4684 10164 4740 10220
rect 35196 10164 35252 10220
rect 35300 10164 35356 10220
rect 35404 10164 35460 10220
rect 19836 9380 19892 9436
rect 19940 9380 19996 9436
rect 20044 9380 20100 9436
rect 4476 8596 4532 8652
rect 4580 8596 4636 8652
rect 4684 8596 4740 8652
rect 35196 8596 35252 8652
rect 35300 8596 35356 8652
rect 35404 8596 35460 8652
rect 19836 7812 19892 7868
rect 19940 7812 19996 7868
rect 20044 7812 20100 7868
rect 4476 7028 4532 7084
rect 4580 7028 4636 7084
rect 4684 7028 4740 7084
rect 35196 7028 35252 7084
rect 35300 7028 35356 7084
rect 35404 7028 35460 7084
rect 19836 6244 19892 6300
rect 19940 6244 19996 6300
rect 20044 6244 20100 6300
rect 35868 6076 35924 6132
rect 4476 5460 4532 5516
rect 4580 5460 4636 5516
rect 4684 5460 4740 5516
rect 35196 5460 35252 5516
rect 35300 5460 35356 5516
rect 35404 5460 35460 5516
rect 35868 5180 35924 5236
rect 19836 4676 19892 4732
rect 19940 4676 19996 4732
rect 20044 4676 20100 4732
rect 4476 3892 4532 3948
rect 4580 3892 4636 3948
rect 4684 3892 4740 3948
rect 35196 3892 35252 3948
rect 35300 3892 35356 3948
rect 35404 3892 35460 3948
rect 19836 3108 19892 3164
rect 19940 3108 19996 3164
rect 20044 3108 20100 3164
<< metal4 >>
rect 4448 55692 4768 56508
rect 4448 55636 4476 55692
rect 4532 55636 4580 55692
rect 4636 55636 4684 55692
rect 4740 55636 4768 55692
rect 4448 54124 4768 55636
rect 4448 54068 4476 54124
rect 4532 54068 4580 54124
rect 4636 54068 4684 54124
rect 4740 54068 4768 54124
rect 4448 52556 4768 54068
rect 4448 52500 4476 52556
rect 4532 52500 4580 52556
rect 4636 52500 4684 52556
rect 4740 52500 4768 52556
rect 4448 50988 4768 52500
rect 4448 50932 4476 50988
rect 4532 50932 4580 50988
rect 4636 50932 4684 50988
rect 4740 50932 4768 50988
rect 4448 49420 4768 50932
rect 4448 49364 4476 49420
rect 4532 49364 4580 49420
rect 4636 49364 4684 49420
rect 4740 49364 4768 49420
rect 4448 47852 4768 49364
rect 4448 47796 4476 47852
rect 4532 47796 4580 47852
rect 4636 47796 4684 47852
rect 4740 47796 4768 47852
rect 4448 46284 4768 47796
rect 4448 46228 4476 46284
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4740 46228 4768 46284
rect 4448 44716 4768 46228
rect 19808 56476 20128 56508
rect 19808 56420 19836 56476
rect 19892 56420 19940 56476
rect 19996 56420 20044 56476
rect 20100 56420 20128 56476
rect 19808 54908 20128 56420
rect 35168 55692 35488 56508
rect 35168 55636 35196 55692
rect 35252 55636 35300 55692
rect 35356 55636 35404 55692
rect 35460 55636 35488 55692
rect 19808 54852 19836 54908
rect 19892 54852 19940 54908
rect 19996 54852 20044 54908
rect 20100 54852 20128 54908
rect 19808 53340 20128 54852
rect 22204 55076 22260 55086
rect 22204 54068 22260 55020
rect 22204 54002 22260 54012
rect 35168 54124 35488 55636
rect 35168 54068 35196 54124
rect 35252 54068 35300 54124
rect 35356 54068 35404 54124
rect 35460 54068 35488 54124
rect 19808 53284 19836 53340
rect 19892 53284 19940 53340
rect 19996 53284 20044 53340
rect 20100 53284 20128 53340
rect 19808 51772 20128 53284
rect 35168 52556 35488 54068
rect 35168 52500 35196 52556
rect 35252 52500 35300 52556
rect 35356 52500 35404 52556
rect 35460 52500 35488 52556
rect 19808 51716 19836 51772
rect 19892 51716 19940 51772
rect 19996 51716 20044 51772
rect 20100 51716 20128 51772
rect 19808 50204 20128 51716
rect 19808 50148 19836 50204
rect 19892 50148 19940 50204
rect 19996 50148 20044 50204
rect 20100 50148 20128 50204
rect 19808 48636 20128 50148
rect 19808 48580 19836 48636
rect 19892 48580 19940 48636
rect 19996 48580 20044 48636
rect 20100 48580 20128 48636
rect 19808 47068 20128 48580
rect 34748 52276 34804 52286
rect 34748 48356 34804 52220
rect 34748 48290 34804 48300
rect 35168 50988 35488 52500
rect 35868 54516 35924 54526
rect 35868 51604 35924 54460
rect 38668 53844 38724 53854
rect 38668 52052 38724 53788
rect 38668 51986 38724 51996
rect 35868 51538 35924 51548
rect 35168 50932 35196 50988
rect 35252 50932 35300 50988
rect 35356 50932 35404 50988
rect 35460 50932 35488 50988
rect 35168 49420 35488 50932
rect 35168 49364 35196 49420
rect 35252 49364 35300 49420
rect 35356 49364 35404 49420
rect 35460 49364 35488 49420
rect 35168 47852 35488 49364
rect 35168 47796 35196 47852
rect 35252 47796 35300 47852
rect 35356 47796 35404 47852
rect 35460 47796 35488 47852
rect 19808 47012 19836 47068
rect 19892 47012 19940 47068
rect 19996 47012 20044 47068
rect 20100 47012 20128 47068
rect 19808 45500 20128 47012
rect 22540 47124 22596 47134
rect 19808 45444 19836 45500
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 20100 45444 20128 45500
rect 4448 44660 4476 44716
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4740 44660 4768 44716
rect 4448 43148 4768 44660
rect 4448 43092 4476 43148
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4740 43092 4768 43148
rect 4448 41580 4768 43092
rect 10108 45220 10164 45230
rect 4448 41524 4476 41580
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4740 41524 4768 41580
rect 4448 40012 4768 41524
rect 4448 39956 4476 40012
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4740 39956 4768 40012
rect 4448 38444 4768 39956
rect 4448 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4768 38444
rect 4448 36876 4768 38388
rect 4448 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4768 36876
rect 4448 35308 4768 36820
rect 4448 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4768 35308
rect 4448 33740 4768 35252
rect 4448 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4768 33740
rect 4448 32172 4768 33684
rect 4448 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4768 32172
rect 4448 30604 4768 32116
rect 4448 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4768 30604
rect 4448 29036 4768 30548
rect 8764 42196 8820 42206
rect 8764 29652 8820 42140
rect 8988 37268 9044 37278
rect 8988 31668 9044 37212
rect 10108 35812 10164 45164
rect 19808 43932 20128 45444
rect 19808 43876 19836 43932
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 20100 43876 20128 43932
rect 19808 42364 20128 43876
rect 19808 42308 19836 42364
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 20100 42308 20128 42364
rect 19808 40796 20128 42308
rect 19808 40740 19836 40796
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 20100 40740 20128 40796
rect 19808 39228 20128 40740
rect 19808 39172 19836 39228
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 20100 39172 20128 39228
rect 19404 37828 19460 37838
rect 10108 35746 10164 35756
rect 11452 37044 11508 37054
rect 9436 35252 9492 35262
rect 9436 33124 9492 35196
rect 9436 33058 9492 33068
rect 9548 35028 9604 35038
rect 8988 31602 9044 31612
rect 9436 32116 9492 32126
rect 9436 31668 9492 32060
rect 9436 31602 9492 31612
rect 8764 29586 8820 29596
rect 4448 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4768 29036
rect 4448 27468 4768 28980
rect 9548 28868 9604 34972
rect 9548 28802 9604 28812
rect 11452 28420 11508 36988
rect 19404 36820 19460 37772
rect 19404 36754 19460 36764
rect 19808 37660 20128 39172
rect 19808 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20128 37660
rect 19808 36092 20128 37604
rect 21756 45556 21812 45566
rect 21532 36932 21588 36942
rect 21532 36484 21588 36876
rect 21532 36418 21588 36428
rect 19808 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20128 36092
rect 19808 34524 20128 36036
rect 19808 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20128 34524
rect 19808 32956 20128 34468
rect 19808 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20128 32956
rect 11452 28354 11508 28364
rect 17948 31780 18004 31790
rect 4448 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4768 27468
rect 4448 25900 4768 27412
rect 17948 26516 18004 31724
rect 19808 31388 20128 32900
rect 20748 33796 20804 33806
rect 20748 31668 20804 33740
rect 20748 31602 20804 31612
rect 19808 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20128 31388
rect 18732 30884 18788 30894
rect 18732 27636 18788 30828
rect 18732 27570 18788 27580
rect 19808 29820 20128 31332
rect 19808 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20128 29820
rect 19808 28252 20128 29764
rect 21756 28868 21812 45500
rect 22540 34020 22596 47068
rect 35168 46284 35488 47796
rect 35168 46228 35196 46284
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35460 46228 35488 46284
rect 35168 44716 35488 46228
rect 35168 44660 35196 44716
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35460 44660 35488 44716
rect 35168 43148 35488 44660
rect 35168 43092 35196 43148
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35460 43092 35488 43148
rect 35168 41580 35488 43092
rect 35168 41524 35196 41580
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35460 41524 35488 41580
rect 35168 40012 35488 41524
rect 35168 39956 35196 40012
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35460 39956 35488 40012
rect 35168 38444 35488 39956
rect 35168 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35488 38444
rect 35168 36876 35488 38388
rect 35168 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35488 36876
rect 35168 35308 35488 36820
rect 35168 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35488 35308
rect 33852 34244 33908 34254
rect 22540 33954 22596 33964
rect 24332 34132 24388 34142
rect 22092 33908 22148 33918
rect 22092 32564 22148 33852
rect 22092 32498 22148 32508
rect 24332 31780 24388 34076
rect 24332 31714 24388 31724
rect 21756 28802 21812 28812
rect 33852 29540 33908 34188
rect 19808 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20128 28252
rect 19068 26964 19124 26974
rect 19068 26740 19124 26908
rect 19068 26674 19124 26684
rect 19808 26684 20128 28196
rect 17948 26450 18004 26460
rect 19808 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20128 26684
rect 4448 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4768 25900
rect 4448 24332 4768 25844
rect 18620 26404 18676 26414
rect 18620 25508 18676 26348
rect 18620 25442 18676 25452
rect 4448 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4768 24332
rect 4448 22764 4768 24276
rect 14364 25284 14420 25294
rect 4448 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4768 22764
rect 4448 21196 4768 22708
rect 13244 23156 13300 23166
rect 4448 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4768 21196
rect 11116 22036 11172 22046
rect 11116 21252 11172 21980
rect 11116 21186 11172 21196
rect 13244 21924 13300 23100
rect 14364 22932 14420 25228
rect 19808 25116 20128 26628
rect 33852 26516 33908 29484
rect 35168 33740 35488 35252
rect 35168 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35488 33740
rect 35168 32172 35488 33684
rect 35168 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35488 32172
rect 35168 30604 35488 32116
rect 35168 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35488 30604
rect 35168 29036 35488 30548
rect 36988 33684 37044 33694
rect 35168 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35488 29036
rect 33852 26450 33908 26460
rect 34972 28308 35028 28318
rect 34972 26068 35028 28252
rect 34972 26002 35028 26012
rect 35168 27468 35488 28980
rect 35168 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35488 27468
rect 35168 25900 35488 27412
rect 36428 29988 36484 29998
rect 36428 26852 36484 29932
rect 36988 26908 37044 33628
rect 36428 26786 36484 26796
rect 36876 26852 37044 26908
rect 35168 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35488 25900
rect 19808 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20128 25116
rect 14924 23940 14980 23950
rect 14924 23492 14980 23884
rect 14924 23426 14980 23436
rect 19808 23548 20128 25060
rect 19808 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20128 23548
rect 4448 19628 4768 21140
rect 13244 20132 13300 21868
rect 13244 20066 13300 20076
rect 13580 22260 13636 22270
rect 4448 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4768 19628
rect 4448 18060 4768 19572
rect 13580 19348 13636 22204
rect 14028 22036 14084 22046
rect 14028 21364 14084 21980
rect 14028 21298 14084 21308
rect 14364 21364 14420 22876
rect 19808 21980 20128 23492
rect 23212 25508 23268 25518
rect 23212 23492 23268 25452
rect 23212 23426 23268 23436
rect 35168 24332 35488 25844
rect 35980 25620 36036 25630
rect 35980 24612 36036 25564
rect 36876 25172 36932 26852
rect 36876 25106 36932 25116
rect 35980 24546 36036 24556
rect 35168 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35488 24332
rect 35168 22764 35488 24276
rect 19808 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20128 21980
rect 14364 21298 14420 21308
rect 15596 21812 15652 21822
rect 15596 21140 15652 21756
rect 15596 21074 15652 21084
rect 19808 20412 20128 21924
rect 34860 22708 34916 22718
rect 19808 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20128 20412
rect 13580 19282 13636 19292
rect 19628 19684 19684 19694
rect 4448 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4768 18060
rect 4448 16492 4768 18004
rect 4448 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4768 16492
rect 4448 14924 4768 16436
rect 19628 17668 19684 19628
rect 19628 15764 19684 17612
rect 19628 15698 19684 15708
rect 19808 18844 20128 20356
rect 22652 21700 22708 21710
rect 22652 20132 22708 21644
rect 22652 20066 22708 20076
rect 19808 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20128 18844
rect 19808 17276 20128 18788
rect 19808 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20128 17276
rect 19808 15708 20128 17220
rect 4448 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4768 14924
rect 4448 13356 4768 14868
rect 4448 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4768 13356
rect 4448 11788 4768 13300
rect 4448 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4768 11788
rect 4448 10220 4768 11732
rect 4448 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4768 10220
rect 4448 8652 4768 10164
rect 4448 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4768 8652
rect 4448 7084 4768 8596
rect 4448 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4768 7084
rect 4448 5516 4768 7028
rect 4448 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4768 5516
rect 4448 3948 4768 5460
rect 4448 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4768 3948
rect 4448 3076 4768 3892
rect 19808 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20128 15708
rect 19808 14140 20128 15652
rect 26908 17220 26964 17230
rect 19808 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20128 14140
rect 19808 12572 20128 14084
rect 20188 15316 20244 15326
rect 20188 13412 20244 15260
rect 23884 15204 23940 15214
rect 23884 13860 23940 15148
rect 26908 14980 26964 17164
rect 34860 15540 34916 22652
rect 34860 15474 34916 15484
rect 35168 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35488 22764
rect 35168 21196 35488 22708
rect 35168 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35488 21196
rect 35168 19628 35488 21140
rect 35168 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35488 19628
rect 35168 18060 35488 19572
rect 35168 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35488 18060
rect 35168 16492 35488 18004
rect 35168 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35488 16492
rect 26908 14914 26964 14924
rect 35168 14924 35488 16436
rect 35868 22708 35924 22718
rect 35868 16212 35924 22652
rect 43148 20692 43204 20702
rect 35980 20580 36036 20590
rect 35980 19348 36036 20524
rect 35980 16884 36036 19292
rect 35980 16818 36036 16828
rect 38892 20244 38948 20254
rect 35868 15764 35924 16156
rect 35868 15698 35924 15708
rect 23884 13794 23940 13804
rect 35168 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35488 14924
rect 38892 14980 38948 20188
rect 38892 14914 38948 14924
rect 42924 16436 42980 16446
rect 20188 13346 20244 13356
rect 35168 13356 35488 14868
rect 42924 14868 42980 16380
rect 42924 14802 42980 14812
rect 19808 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20128 12572
rect 19808 11004 20128 12516
rect 19808 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20128 11004
rect 19808 9436 20128 10948
rect 19808 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20128 9436
rect 19808 7868 20128 9380
rect 19808 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20128 7868
rect 19808 6300 20128 7812
rect 19808 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20128 6300
rect 19808 4732 20128 6244
rect 19808 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20128 4732
rect 19808 3164 20128 4676
rect 19808 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20128 3164
rect 19808 3076 20128 3108
rect 35168 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35488 13356
rect 35168 11788 35488 13300
rect 43148 12628 43204 20636
rect 44380 18340 44436 18350
rect 44380 18116 44436 18284
rect 44380 17556 44436 18060
rect 44380 17490 44436 17500
rect 43148 12562 43204 12572
rect 35168 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35488 11788
rect 35168 10220 35488 11732
rect 38892 11620 38948 11630
rect 38892 11060 38948 11564
rect 38892 10994 38948 11004
rect 35168 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35488 10220
rect 35168 8652 35488 10164
rect 35168 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35488 8652
rect 35168 7084 35488 8596
rect 35168 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35488 7084
rect 35168 5516 35488 7028
rect 35168 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35488 5516
rect 35168 3948 35488 5460
rect 35868 6132 35924 6142
rect 35868 5236 35924 6076
rect 35868 5170 35924 5180
rect 35168 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35488 3948
rect 35168 3076 35488 3892
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1259_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 18928 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1260_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 18256 0 -1 31360
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1261_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 21168 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1262_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 19376 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1263_
timestamp 1698431365
transform 1 0 20272 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1264_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 19152 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_4  _1265_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 21168 0 -1 31360
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1266_
timestamp 1698431365
transform -1 0 20944 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1267_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 19376 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1268_
timestamp 1698431365
transform 1 0 18480 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1269_
timestamp 1698431365
transform 1 0 19264 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _1270_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 24080 0 1 32928
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1271_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 18480 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1272_
timestamp 1698431365
transform 1 0 19824 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_4  _1273_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 22288 0 1 34496
box -86 -86 4006 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1274_
timestamp 1698431365
transform 1 0 20048 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1275_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 18816 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _1276_
timestamp 1698431365
transform 1 0 19040 0 -1 29792
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1277_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 16464 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1278_
timestamp 1698431365
transform 1 0 16128 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1279_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 22960 0 -1 36064
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1280_
timestamp 1698431365
transform -1 0 28784 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  _1281_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 29568 0 -1 28224
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1282_
timestamp 1698431365
transform -1 0 27776 0 -1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1283_
timestamp 1698431365
transform -1 0 24640 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1284_
timestamp 1698431365
transform 1 0 26656 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1285_
timestamp 1698431365
transform 1 0 30576 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _1286_
timestamp 1698431365
transform 1 0 24864 0 1 26656
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1287_
timestamp 1698431365
transform 1 0 25088 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_2  _1288_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 26656 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1289_
timestamp 1698431365
transform -1 0 32368 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1290_
timestamp 1698431365
transform -1 0 32032 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1291_
timestamp 1698431365
transform -1 0 29680 0 -1 29792
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1292_
timestamp 1698431365
transform 1 0 27776 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  _1293_
timestamp 1698431365
transform 1 0 29008 0 1 26656
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_4  _1294_
timestamp 1698431365
transform -1 0 29344 0 -1 32928
box -86 -86 4006 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1295_
timestamp 1698431365
transform -1 0 28000 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _1296_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 26656 0 1 25088
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1297_
timestamp 1698431365
transform 1 0 24192 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1298_
timestamp 1698431365
transform -1 0 29904 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1299_
timestamp 1698431365
transform -1 0 27552 0 1 32928
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _1300_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 25200 0 -1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _1301_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 17248 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _1302_
timestamp 1698431365
transform 1 0 17248 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  _1303_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 15904 0 -1 29792
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1304_
timestamp 1698431365
transform -1 0 15120 0 1 31360
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  _1305_
timestamp 1698431365
transform -1 0 16688 0 -1 23520
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _1306_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 13104 0 1 28224
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  _1307_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 13104 0 1 31360
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1308_
timestamp 1698431365
transform -1 0 12992 0 1 29792
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  _1309_
timestamp 1698431365
transform -1 0 17024 0 -1 31360
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _1310_
timestamp 1698431365
transform 1 0 13328 0 -1 28224
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__or2_4  _1311_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 11872 0 1 29792
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _1312_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 12768 0 -1 31360
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _1313_
timestamp 1698431365
transform 1 0 16576 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1314_
timestamp 1698431365
transform 1 0 14784 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _1315_
timestamp 1698431365
transform -1 0 17248 0 1 32928
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1316_
timestamp 1698431365
transform -1 0 12768 0 -1 31360
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1317_
timestamp 1698431365
transform 1 0 11312 0 -1 32928
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1318_
timestamp 1698431365
transform 1 0 5824 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _1319_
timestamp 1698431365
transform -1 0 7504 0 1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  _1320_
timestamp 1698431365
transform -1 0 8176 0 -1 23520
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1321_
timestamp 1698431365
transform -1 0 7280 0 1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  _1322_
timestamp 1698431365
transform -1 0 7840 0 1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _1323_
timestamp 1698431365
transform 1 0 6272 0 -1 25088
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _1324_
timestamp 1698431365
transform -1 0 11200 0 -1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1325_
timestamp 1698431365
transform -1 0 5264 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  _1326_
timestamp 1698431365
transform 1 0 9968 0 -1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_4  _1327_
timestamp 1698431365
transform 1 0 8064 0 1 23520
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1328_
timestamp 1698431365
transform 1 0 9408 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_4  _1329_
timestamp 1698431365
transform -1 0 11424 0 1 20384
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_4  _1330_
timestamp 1698431365
transform -1 0 7392 0 -1 28224
box -86 -86 4006 870
use gf180mcu_fd_sc_mcu7t5v0__inv_2  _1331_
timestamp 1698431365
transform 1 0 5600 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  _1332_
timestamp 1698431365
transform -1 0 9408 0 1 20384
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _1333_
timestamp 1698431365
transform -1 0 12432 0 -1 23520
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1334_
timestamp 1698431365
transform 1 0 4480 0 -1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1335_
timestamp 1698431365
transform 1 0 5936 0 1 28224
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__and4_2  _1336_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 10080 0 1 31360
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1337_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 9408 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1338_
timestamp 1698431365
transform 1 0 25088 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1339_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 29008 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1340_
timestamp 1698431365
transform 1 0 26208 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1341_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 26880 0 1 34496
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1342_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 27552 0 -1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _1343_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 20944 0 1 31360
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1344_
timestamp 1698431365
transform 1 0 21168 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_2  _1345_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 21504 0 -1 32928
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1346_
timestamp 1698431365
transform 1 0 28448 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _1347_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 30688 0 -1 31360
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1348_
timestamp 1698431365
transform -1 0 34496 0 1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1349_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 33712 0 -1 28224
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _1350_
timestamp 1698431365
transform 1 0 29008 0 1 29792
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1351_
timestamp 1698431365
transform -1 0 32704 0 -1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_4  _1352_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 28784 0 1 31360
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1353_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 27664 0 -1 34496
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1354_
timestamp 1698431365
transform -1 0 16912 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1355_
timestamp 1698431365
transform -1 0 10304 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1356_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 13328 0 1 29792
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_4  _1357_
timestamp 1698431365
transform 1 0 16464 0 1 31360
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _1358_
timestamp 1698431365
transform 1 0 17248 0 -1 34496
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _1359_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 13104 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1360_
timestamp 1698431365
transform -1 0 8624 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _1361_
timestamp 1698431365
transform 1 0 15568 0 -1 34496
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1362_
timestamp 1698431365
transform -1 0 9184 0 -1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1363_
timestamp 1698431365
transform 1 0 8176 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1364_
timestamp 1698431365
transform 1 0 6160 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _1365_
timestamp 1698431365
transform -1 0 8400 0 -1 26656
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  _1366_
timestamp 1698431365
transform 1 0 12320 0 -1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _1367_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 15120 0 -1 23520
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1368_
timestamp 1698431365
transform 1 0 4144 0 1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _1369_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 11536 0 -1 28224
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_2  _1370_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 7952 0 1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1371_
timestamp 1698431365
transform 1 0 29008 0 1 36064
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1372_
timestamp 1698431365
transform -1 0 30464 0 1 37632
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1373_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 29008 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1374_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 27552 0 1 32928
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1375_
timestamp 1698431365
transform 1 0 28784 0 -1 36064
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_4  _1376_
timestamp 1698431365
transform 1 0 9968 0 -1 25088
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_4  _1377_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 13104 0 1 25088
box -86 -86 4902 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1378_
timestamp 1698431365
transform 1 0 10640 0 1 36064
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1379_
timestamp 1698431365
transform -1 0 9184 0 -1 34496
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1380_
timestamp 1698431365
transform 1 0 8848 0 1 37632
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1381_
timestamp 1698431365
transform 1 0 10528 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1382_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 4368 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1383_
timestamp 1698431365
transform 1 0 4368 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1384_
timestamp 1698431365
transform 1 0 13440 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _1385_
timestamp 1698431365
transform -1 0 9184 0 1 21952
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _1386_
timestamp 1698431365
transform -1 0 12656 0 1 26656
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _1387_
timestamp 1698431365
transform -1 0 12544 0 1 23520
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1388_
timestamp 1698431365
transform -1 0 9968 0 -1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _1389_
timestamp 1698431365
transform 1 0 13776 0 1 25088
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1390_
timestamp 1698431365
transform 1 0 10192 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_4  _1391_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 11088 0 1 32928
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_4  _1392_
timestamp 1698431365
transform -1 0 17024 0 -1 32928
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1393_
timestamp 1698431365
transform 1 0 17248 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_4  _1394_
timestamp 1698431365
transform 1 0 17248 0 1 32928
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  _1395_
timestamp 1698431365
transform -1 0 10640 0 1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _1396_
timestamp 1698431365
transform 1 0 12992 0 -1 29792
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _1397_
timestamp 1698431365
transform -1 0 12544 0 -1 34496
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  _1398_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 17808 0 1 36064
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1399_
timestamp 1698431365
transform 1 0 11648 0 1 37632
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1400_
timestamp 1698431365
transform -1 0 32256 0 -1 29792
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1401_
timestamp 1698431365
transform -1 0 28224 0 -1 28224
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1402_
timestamp 1698431365
transform -1 0 20272 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _1403_
timestamp 1698431365
transform 1 0 29680 0 -1 29792
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _1404_
timestamp 1698431365
transform 1 0 25088 0 -1 25088
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _1405_
timestamp 1698431365
transform 1 0 25088 0 -1 29792
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  _1406_
timestamp 1698431365
transform 1 0 24304 0 1 29792
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1407_
timestamp 1698431365
transform -1 0 21840 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1408_
timestamp 1698431365
transform -1 0 22848 0 1 29792
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _1409_
timestamp 1698431365
transform -1 0 20944 0 -1 32928
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _1410_
timestamp 1698431365
transform -1 0 21168 0 -1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1411_
timestamp 1698431365
transform -1 0 20944 0 1 32928
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1412_
timestamp 1698431365
transform 1 0 19936 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _1413_
timestamp 1698431365
transform 1 0 21168 0 1 36064
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1414_
timestamp 1698431365
transform -1 0 22512 0 -1 39200
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _1415_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 14336 0 -1 39200
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1416_
timestamp 1698431365
transform -1 0 30576 0 -1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1417_
timestamp 1698431365
transform 1 0 28672 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1418_
timestamp 1698431365
transform -1 0 28784 0 1 39200
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1419_
timestamp 1698431365
transform 1 0 14336 0 1 39200
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1420_
timestamp 1698431365
transform 1 0 22848 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1421_
timestamp 1698431365
transform -1 0 20272 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1422_
timestamp 1698431365
transform -1 0 23408 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1423_
timestamp 1698431365
transform 1 0 21952 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1424_
timestamp 1698431365
transform -1 0 26544 0 -1 28224
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1425_
timestamp 1698431365
transform 1 0 23184 0 -1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _1426_
timestamp 1698431365
transform -1 0 24864 0 -1 29792
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  _1427_
timestamp 1698431365
transform 1 0 24192 0 1 28224
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1428_
timestamp 1698431365
transform -1 0 19040 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1429_
timestamp 1698431365
transform 1 0 21168 0 1 34496
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1430_
timestamp 1698431365
transform 1 0 13776 0 1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1431_
timestamp 1698431365
transform 1 0 14896 0 1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1432_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 19824 0 1 34496
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1433_
timestamp 1698431365
transform -1 0 20832 0 -1 39200
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1434_
timestamp 1698431365
transform 1 0 8400 0 -1 26656
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1435_
timestamp 1698431365
transform -1 0 9968 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and3_2  _1436_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 9968 0 1 26656
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1437_
timestamp 1698431365
transform -1 0 14336 0 -1 39200
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1438_
timestamp 1698431365
transform -1 0 11536 0 -1 31360
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _1439_
timestamp 1698431365
transform -1 0 15456 0 -1 34496
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_4  _1440_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 12320 0 -1 36064
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1441_
timestamp 1698431365
transform 1 0 11760 0 1 39200
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1442_
timestamp 1698431365
transform -1 0 10640 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1443_
timestamp 1698431365
transform -1 0 11312 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1444_
timestamp 1698431365
transform 1 0 13888 0 -1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1445_
timestamp 1698431365
transform 1 0 14336 0 1 37632
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1446_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 17696 0 1 39200
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1447_
timestamp 1698431365
transform 1 0 26768 0 -1 40768
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1448_
timestamp 1698431365
transform 1 0 27104 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1449_
timestamp 1698431365
transform 1 0 29008 0 1 40768
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1450_
timestamp 1698431365
transform 1 0 19152 0 -1 40768
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1451_
timestamp 1698431365
transform -1 0 22176 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1452_
timestamp 1698431365
transform -1 0 20160 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1453_
timestamp 1698431365
transform 1 0 20384 0 1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1454_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 21504 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1455_
timestamp 1698431365
transform 1 0 20272 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1456_
timestamp 1698431365
transform 1 0 23296 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1457_
timestamp 1698431365
transform -1 0 22960 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1458_
timestamp 1698431365
transform 1 0 23968 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1459_
timestamp 1698431365
transform 1 0 23856 0 1 40768
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1460_
timestamp 1698431365
transform 1 0 10640 0 -1 36064
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1461_
timestamp 1698431365
transform 1 0 8400 0 1 28224
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1462_
timestamp 1698431365
transform 1 0 10416 0 1 40768
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1463_
timestamp 1698431365
transform 1 0 11424 0 -1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1464_
timestamp 1698431365
transform -1 0 8512 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1465_
timestamp 1698431365
transform -1 0 9184 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1466_
timestamp 1698431365
transform 1 0 10640 0 -1 42336
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1467_
timestamp 1698431365
transform -1 0 14224 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1468_
timestamp 1698431365
transform 1 0 13328 0 1 40768
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1469_
timestamp 1698431365
transform 1 0 25088 0 1 42336
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _1470_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 26768 0 -1 42336
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1471_
timestamp 1698431365
transform 1 0 29904 0 -1 43904
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1472_
timestamp 1698431365
transform 1 0 31696 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1473_
timestamp 1698431365
transform 1 0 26992 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1474_
timestamp 1698431365
transform 1 0 29120 0 -1 42336
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1475_
timestamp 1698431365
transform 1 0 23744 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1476_
timestamp 1698431365
transform 1 0 23968 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1477_
timestamp 1698431365
transform 1 0 25312 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1478_
timestamp 1698431365
transform -1 0 26768 0 -1 42336
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1479_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 23296 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1480_
timestamp 1698431365
transform 1 0 23072 0 1 36064
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1481_
timestamp 1698431365
transform 1 0 20272 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1482_
timestamp 1698431365
transform 1 0 24528 0 1 32928
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1483_
timestamp 1698431365
transform 1 0 25648 0 -1 43904
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1484_
timestamp 1698431365
transform 1 0 9968 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _1485_
timestamp 1698431365
transform -1 0 13216 0 -1 40768
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _1486_
timestamp 1698431365
transform 1 0 13328 0 1 34496
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1487_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 9408 0 1 32928
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1488_
timestamp 1698431365
transform 1 0 5264 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1489_
timestamp 1698431365
transform -1 0 7504 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1490_
timestamp 1698431365
transform 1 0 7504 0 1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1491_
timestamp 1698431365
transform -1 0 9072 0 -1 29792
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1492_
timestamp 1698431365
transform 1 0 9968 0 1 42336
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1493_
timestamp 1698431365
transform -1 0 12432 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _1494_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 11648 0 1 42336
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1495_
timestamp 1698431365
transform 1 0 12432 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1496_
timestamp 1698431365
transform 1 0 26768 0 1 43904
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1497_
timestamp 1698431365
transform 1 0 29008 0 1 43904
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1498_
timestamp 1698431365
transform 1 0 30352 0 1 43904
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1499_
timestamp 1698431365
transform -1 0 34720 0 1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1500_
timestamp 1698431365
transform -1 0 24080 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1501_
timestamp 1698431365
transform 1 0 21728 0 -1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1502_
timestamp 1698431365
transform -1 0 23296 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _1503_
timestamp 1698431365
transform 1 0 21840 0 1 31360
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1504_
timestamp 1698431365
transform 1 0 22848 0 1 29792
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1505_
timestamp 1698431365
transform -1 0 22064 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1506_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 21168 0 -1 34496
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1507_
timestamp 1698431365
transform -1 0 24976 0 1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1508_
timestamp 1698431365
transform 1 0 21504 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1509_
timestamp 1698431365
transform 1 0 19040 0 1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1510_
timestamp 1698431365
transform 1 0 21168 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1511_
timestamp 1698431365
transform 1 0 21392 0 1 45472
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1512_
timestamp 1698431365
transform 1 0 13552 0 1 37632
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1513_
timestamp 1698431365
transform -1 0 17024 0 -1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _1514_
timestamp 1698431365
transform 1 0 17248 0 -1 36064
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1515_
timestamp 1698431365
transform -1 0 17472 0 1 37632
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1516_
timestamp 1698431365
transform 1 0 18256 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1517_
timestamp 1698431365
transform 1 0 12544 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _1518_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 13328 0 1 26656
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _1519_
timestamp 1698431365
transform -1 0 12096 0 -1 29792
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1520_
timestamp 1698431365
transform 1 0 10304 0 -1 45472
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1521_
timestamp 1698431365
transform 1 0 10976 0 -1 43904
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1522_
timestamp 1698431365
transform 1 0 11984 0 1 43904
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _1523_
timestamp 1698431365
transform 1 0 13328 0 1 45472
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1524_
timestamp 1698431365
transform 1 0 22736 0 -1 47040
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1525_
timestamp 1698431365
transform -1 0 27104 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1526_
timestamp 1698431365
transform 1 0 27104 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1527_
timestamp 1698431365
transform 1 0 25872 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1528_
timestamp 1698431365
transform -1 0 28448 0 -1 43904
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _1529_
timestamp 1698431365
transform 1 0 29008 0 1 47040
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1530_
timestamp 1698431365
transform 1 0 28784 0 -1 43904
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1531_
timestamp 1698431365
transform 1 0 29120 0 -1 45472
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_4  _1532_
timestamp 1698431365
transform 1 0 29680 0 -1 45472
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1533_
timestamp 1698431365
transform 1 0 31024 0 1 47040
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1534_
timestamp 1698431365
transform 1 0 35280 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1535_
timestamp 1698431365
transform -1 0 30912 0 -1 47040
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1536_
timestamp 1698431365
transform -1 0 29792 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1537_
timestamp 1698431365
transform 1 0 24192 0 -1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1538_
timestamp 1698431365
transform -1 0 23408 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1539_
timestamp 1698431365
transform 1 0 22624 0 1 47040
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1540_
timestamp 1698431365
transform 1 0 21168 0 1 47040
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1541_
timestamp 1698431365
transform 1 0 23184 0 1 47040
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1542_
timestamp 1698431365
transform -1 0 5264 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1543_
timestamp 1698431365
transform -1 0 9856 0 1 29792
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1544_
timestamp 1698431365
transform 1 0 14896 0 -1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _1545_
timestamp 1698431365
transform -1 0 10640 0 -1 36064
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1546_
timestamp 1698431365
transform 1 0 9968 0 -1 47040
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1547_
timestamp 1698431365
transform 1 0 9520 0 1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1548_
timestamp 1698431365
transform 1 0 10080 0 1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1549_
timestamp 1698431365
transform 1 0 9968 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1550_
timestamp 1698431365
transform 1 0 11088 0 1 47040
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1551_
timestamp 1698431365
transform -1 0 11088 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1552_
timestamp 1698431365
transform -1 0 11760 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1553_
timestamp 1698431365
transform 1 0 10528 0 -1 47040
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1554_
timestamp 1698431365
transform 1 0 12096 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1555_
timestamp 1698431365
transform -1 0 13104 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1556_
timestamp 1698431365
transform 1 0 11648 0 1 47040
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1557_
timestamp 1698431365
transform -1 0 21504 0 -1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1558_
timestamp 1698431365
transform 1 0 22288 0 -1 34496
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1559_
timestamp 1698431365
transform 1 0 20048 0 -1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _1560_
timestamp 1698431365
transform 1 0 23744 0 1 31360
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1561_
timestamp 1698431365
transform 1 0 25088 0 -1 48608
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1562_
timestamp 1698431365
transform 1 0 25648 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _1563_
timestamp 1698431365
transform 1 0 26768 0 1 48608
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_2  _1564_
timestamp 1698431365
transform 1 0 29792 0 1 48608
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1565_
timestamp 1698431365
transform 1 0 36848 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1566_
timestamp 1698431365
transform 1 0 29120 0 1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  _1567_
timestamp 1698431365
transform 1 0 27664 0 -1 48608
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1568_
timestamp 1698431365
transform 1 0 29792 0 1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1569_
timestamp 1698431365
transform -1 0 24864 0 1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1570_
timestamp 1698431365
transform 1 0 25536 0 1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1571_
timestamp 1698431365
transform 1 0 26208 0 1 48608
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1572_
timestamp 1698431365
transform 1 0 27552 0 -1 50176
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1573_
timestamp 1698431365
transform -1 0 24192 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1574_
timestamp 1698431365
transform -1 0 23968 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1575_
timestamp 1698431365
transform 1 0 20496 0 -1 37632
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1576_
timestamp 1698431365
transform 1 0 21728 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1577_
timestamp 1698431365
transform -1 0 21840 0 1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1578_
timestamp 1698431365
transform 1 0 21168 0 1 50176
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1579_
timestamp 1698431365
transform 1 0 22288 0 -1 53312
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1580_
timestamp 1698431365
transform -1 0 13104 0 1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1581_
timestamp 1698431365
transform -1 0 12656 0 -1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _1582_
timestamp 1698431365
transform -1 0 12992 0 -1 28224
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1583_
timestamp 1698431365
transform -1 0 10080 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1584_
timestamp 1698431365
transform -1 0 9296 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1585_
timestamp 1698431365
transform 1 0 9408 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1586_
timestamp 1698431365
transform -1 0 10416 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1587_
timestamp 1698431365
transform -1 0 9184 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1588_
timestamp 1698431365
transform 1 0 10080 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1589_
timestamp 1698431365
transform 1 0 10416 0 1 43904
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1590_
timestamp 1698431365
transform 1 0 11200 0 -1 47040
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1591_
timestamp 1698431365
transform 1 0 12320 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1592_
timestamp 1698431365
transform 1 0 10528 0 1 50176
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1593_
timestamp 1698431365
transform 1 0 23072 0 1 51744
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1594_
timestamp 1698431365
transform 1 0 29008 0 1 51744
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1595_
timestamp 1698431365
transform 1 0 33488 0 -1 51744
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1596_
timestamp 1698431365
transform 1 0 36064 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1597_
timestamp 1698431365
transform 1 0 29120 0 1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1598_
timestamp 1698431365
transform 1 0 29120 0 -1 53312
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _1599_
timestamp 1698431365
transform 1 0 30576 0 -1 51744
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1600_
timestamp 1698431365
transform -1 0 23072 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1601_
timestamp 1698431365
transform 1 0 24080 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1602_
timestamp 1698431365
transform 1 0 21952 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1603_
timestamp 1698431365
transform 1 0 23072 0 -1 48608
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _1604_
timestamp 1698431365
transform 1 0 9184 0 1 21952
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1605_
timestamp 1698431365
transform 1 0 9968 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1606_
timestamp 1698431365
transform 1 0 13216 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1607_
timestamp 1698431365
transform 1 0 13552 0 -1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1608_
timestamp 1698431365
transform 1 0 14112 0 -1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1609_
timestamp 1698431365
transform 1 0 13888 0 1 51744
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1610_
timestamp 1698431365
transform -1 0 15344 0 -1 50176
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1611_
timestamp 1698431365
transform -1 0 11424 0 -1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1612_
timestamp 1698431365
transform 1 0 11424 0 1 48608
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1613_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 12320 0 -1 48608
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1614_
timestamp 1698431365
transform 1 0 11424 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1615_
timestamp 1698431365
transform 1 0 13776 0 1 50176
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1616_
timestamp 1698431365
transform 1 0 22624 0 1 50176
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1617_
timestamp 1698431365
transform 1 0 28448 0 -1 51744
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1618_
timestamp 1698431365
transform 1 0 30576 0 -1 53312
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1619_
timestamp 1698431365
transform 1 0 39312 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1620_
timestamp 1698431365
transform -1 0 23072 0 1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1621_
timestamp 1698431365
transform -1 0 22624 0 1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1622_
timestamp 1698431365
transform 1 0 22400 0 -1 50176
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1623_
timestamp 1698431365
transform 1 0 23744 0 -1 50176
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1624_
timestamp 1698431365
transform -1 0 23744 0 -1 50176
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1625_
timestamp 1698431365
transform 1 0 13888 0 1 48608
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1626_
timestamp 1698431365
transform 1 0 15232 0 1 50176
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1627_
timestamp 1698431365
transform 1 0 31024 0 1 51744
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1628_
timestamp 1698431365
transform 1 0 27888 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1629_
timestamp 1698431365
transform -1 0 31584 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1630_
timestamp 1698431365
transform 1 0 32480 0 1 51744
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1631_
timestamp 1698431365
transform 1 0 42784 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1632_
timestamp 1698431365
transform 1 0 32032 0 -1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1633_
timestamp 1698431365
transform -1 0 33936 0 1 50176
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1634_
timestamp 1698431365
transform 1 0 43680 0 -1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1635_
timestamp 1698431365
transform -1 0 43232 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1636_
timestamp 1698431365
transform -1 0 45696 0 1 45472
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1637_
timestamp 1698431365
transform 1 0 41440 0 1 43904
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1638_
timestamp 1698431365
transform -1 0 44352 0 -1 45472
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1639_
timestamp 1698431365
transform -1 0 40544 0 -1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1640_
timestamp 1698431365
transform -1 0 31920 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1641_
timestamp 1698431365
transform -1 0 25424 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1642_
timestamp 1698431365
transform -1 0 26880 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1643_
timestamp 1698431365
transform -1 0 22848 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1644_
timestamp 1698431365
transform 1 0 16576 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1645_
timestamp 1698431365
transform -1 0 18592 0 -1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1646_
timestamp 1698431365
transform -1 0 22400 0 1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1647_
timestamp 1698431365
transform 1 0 26768 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1648_
timestamp 1698431365
transform 1 0 27664 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1649_
timestamp 1698431365
transform 1 0 28336 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1650_
timestamp 1698431365
transform -1 0 31472 0 -1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1651_
timestamp 1698431365
transform -1 0 32704 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1652_
timestamp 1698431365
transform -1 0 31808 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1653_
timestamp 1698431365
transform -1 0 28448 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1654_
timestamp 1698431365
transform -1 0 30912 0 -1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1655_
timestamp 1698431365
transform -1 0 47824 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1656_
timestamp 1698431365
transform -1 0 30240 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1657_
timestamp 1698431365
transform 1 0 29456 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1658_
timestamp 1698431365
transform 1 0 16352 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1659_
timestamp 1698431365
transform -1 0 27440 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1660_
timestamp 1698431365
transform -1 0 38192 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1661_
timestamp 1698431365
transform -1 0 31360 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1662_
timestamp 1698431365
transform 1 0 30800 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1663_
timestamp 1698431365
transform -1 0 29456 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1664_
timestamp 1698431365
transform 1 0 27888 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1665_
timestamp 1698431365
transform 1 0 29904 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1666_
timestamp 1698431365
transform 1 0 29008 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1667_
timestamp 1698431365
transform -1 0 48048 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1668_
timestamp 1698431365
transform 1 0 38304 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1669_
timestamp 1698431365
transform 1 0 29008 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1670_
timestamp 1698431365
transform 1 0 27888 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1671_
timestamp 1698431365
transform -1 0 45136 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1672_
timestamp 1698431365
transform -1 0 27888 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1673_
timestamp 1698431365
transform 1 0 26880 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1674_
timestamp 1698431365
transform -1 0 34160 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1675_
timestamp 1698431365
transform -1 0 39648 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1676_
timestamp 1698431365
transform 1 0 39648 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1677_
timestamp 1698431365
transform 1 0 41776 0 -1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1678_
timestamp 1698431365
transform 1 0 42112 0 1 10976
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1679_
timestamp 1698431365
transform -1 0 41664 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1680_
timestamp 1698431365
transform 1 0 39536 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1681_
timestamp 1698431365
transform 1 0 38304 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1682_
timestamp 1698431365
transform 1 0 43232 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1683_
timestamp 1698431365
transform 1 0 40992 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1684_
timestamp 1698431365
transform -1 0 40208 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1685_
timestamp 1698431365
transform 1 0 38416 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1686_
timestamp 1698431365
transform -1 0 43792 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1687_
timestamp 1698431365
transform 1 0 22624 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _1688_
timestamp 1698431365
transform -1 0 28448 0 -1 21952
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1689_
timestamp 1698431365
transform 1 0 38080 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1690_
timestamp 1698431365
transform 1 0 38640 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1691_
timestamp 1698431365
transform 1 0 42336 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1692_
timestamp 1698431365
transform 1 0 42560 0 1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1693_
timestamp 1698431365
transform 1 0 41664 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1694_
timestamp 1698431365
transform 1 0 40768 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1695_
timestamp 1698431365
transform 1 0 41440 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1696_
timestamp 1698431365
transform 1 0 40768 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1697_
timestamp 1698431365
transform -1 0 18816 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1698_
timestamp 1698431365
transform 1 0 17248 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1699_
timestamp 1698431365
transform -1 0 39648 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1700_
timestamp 1698431365
transform -1 0 40096 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1701_
timestamp 1698431365
transform -1 0 31920 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1702_
timestamp 1698431365
transform 1 0 30800 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1703_
timestamp 1698431365
transform -1 0 41216 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1704_
timestamp 1698431365
transform -1 0 39312 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1705_
timestamp 1698431365
transform -1 0 36288 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1706_
timestamp 1698431365
transform 1 0 31696 0 -1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1707_
timestamp 1698431365
transform 1 0 29344 0 -1 32928
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1708_
timestamp 1698431365
transform 1 0 31920 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1709_
timestamp 1698431365
transform 1 0 29680 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1710_
timestamp 1698431365
transform 1 0 29120 0 -1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1711_
timestamp 1698431365
transform 1 0 29904 0 1 32928
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1712_
timestamp 1698431365
transform 1 0 17248 0 -1 37632
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1713_
timestamp 1698431365
transform -1 0 18704 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1714_
timestamp 1698431365
transform 1 0 18704 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1715_
timestamp 1698431365
transform -1 0 39088 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1716_
timestamp 1698431365
transform -1 0 37744 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1717_
timestamp 1698431365
transform -1 0 18816 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1718_
timestamp 1698431365
transform -1 0 19376 0 -1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1719_
timestamp 1698431365
transform 1 0 19600 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1720_
timestamp 1698431365
transform -1 0 18592 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1721_
timestamp 1698431365
transform 1 0 16688 0 1 40768
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1722_
timestamp 1698431365
transform -1 0 18816 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1723_
timestamp 1698431365
transform 1 0 17472 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1724_
timestamp 1698431365
transform -1 0 19376 0 -1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1725_
timestamp 1698431365
transform -1 0 19152 0 -1 40768
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1726_
timestamp 1698431365
transform 1 0 16128 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1727_
timestamp 1698431365
transform -1 0 17024 0 -1 42336
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1728_
timestamp 1698431365
transform 1 0 15792 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1729_
timestamp 1698431365
transform 1 0 14896 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1730_
timestamp 1698431365
transform 1 0 14560 0 1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1731_
timestamp 1698431365
transform 1 0 15568 0 -1 43904
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1732_
timestamp 1698431365
transform 1 0 15120 0 1 42336
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1733_
timestamp 1698431365
transform -1 0 15904 0 1 43904
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1734_
timestamp 1698431365
transform 1 0 6608 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1735_
timestamp 1698431365
transform 1 0 16128 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1736_
timestamp 1698431365
transform 1 0 14672 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1737_
timestamp 1698431365
transform -1 0 17024 0 -1 47040
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1738_
timestamp 1698431365
transform -1 0 16464 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1739_
timestamp 1698431365
transform 1 0 16128 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1740_
timestamp 1698431365
transform -1 0 22736 0 -1 43904
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1741_
timestamp 1698431365
transform -1 0 18144 0 -1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1742_
timestamp 1698431365
transform -1 0 18816 0 -1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1743_
timestamp 1698431365
transform 1 0 18816 0 -1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1744_
timestamp 1698431365
transform 1 0 19488 0 1 45472
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1745_
timestamp 1698431365
transform -1 0 23072 0 -1 48608
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1746_
timestamp 1698431365
transform -1 0 18816 0 1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1747_
timestamp 1698431365
transform -1 0 20160 0 1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1748_
timestamp 1698431365
transform 1 0 20160 0 1 48608
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1749_
timestamp 1698431365
transform -1 0 20944 0 1 47040
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1750_
timestamp 1698431365
transform -1 0 23072 0 -1 51744
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1751_
timestamp 1698431365
transform -1 0 18928 0 1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1752_
timestamp 1698431365
transform -1 0 19600 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1753_
timestamp 1698431365
transform 1 0 19040 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1754_
timestamp 1698431365
transform -1 0 19936 0 1 51744
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1755_
timestamp 1698431365
transform -1 0 20608 0 1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1756_
timestamp 1698431365
transform -1 0 20944 0 1 50176
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1757_
timestamp 1698431365
transform 1 0 15344 0 1 48608
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1758_
timestamp 1698431365
transform -1 0 16240 0 -1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1759_
timestamp 1698431365
transform 1 0 15568 0 -1 48608
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1760_
timestamp 1698431365
transform -1 0 17024 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1761_
timestamp 1698431365
transform -1 0 18816 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1762_
timestamp 1698431365
transform -1 0 8736 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1763_
timestamp 1698431365
transform 1 0 3136 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1764_
timestamp 1698431365
transform 1 0 2240 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1765_
timestamp 1698431365
transform -1 0 4704 0 1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1766_
timestamp 1698431365
transform 1 0 1568 0 1 31360
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1767_
timestamp 1698431365
transform 1 0 4592 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1768_
timestamp 1698431365
transform -1 0 2912 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1769_
timestamp 1698431365
transform -1 0 3808 0 1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1770_
timestamp 1698431365
transform 1 0 2912 0 1 32928
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1771_
timestamp 1698431365
transform -1 0 4480 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1772_
timestamp 1698431365
transform -1 0 4704 0 1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1773_
timestamp 1698431365
transform -1 0 3136 0 -1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1774_
timestamp 1698431365
transform -1 0 3472 0 -1 36064
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1775_
timestamp 1698431365
transform 1 0 2464 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1776_
timestamp 1698431365
transform -1 0 5264 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1777_
timestamp 1698431365
transform -1 0 4592 0 -1 37632
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1778_
timestamp 1698431365
transform 1 0 1568 0 1 37632
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1779_
timestamp 1698431365
transform 1 0 4816 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1780_
timestamp 1698431365
transform 1 0 2688 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1781_
timestamp 1698431365
transform -1 0 4816 0 -1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1782_
timestamp 1698431365
transform -1 0 5040 0 1 39200
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1783_
timestamp 1698431365
transform -1 0 4704 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1784_
timestamp 1698431365
transform -1 0 4256 0 1 40768
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1785_
timestamp 1698431365
transform 1 0 3584 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1786_
timestamp 1698431365
transform 1 0 2688 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1787_
timestamp 1698431365
transform -1 0 5712 0 -1 43904
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1788_
timestamp 1698431365
transform -1 0 5040 0 1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1789_
timestamp 1698431365
transform -1 0 5152 0 -1 43904
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1790_
timestamp 1698431365
transform -1 0 3584 0 -1 45472
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1791_
timestamp 1698431365
transform -1 0 7280 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1792_
timestamp 1698431365
transform 1 0 3584 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1793_
timestamp 1698431365
transform 1 0 2128 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1794_
timestamp 1698431365
transform 1 0 3920 0 1 45472
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1795_
timestamp 1698431365
transform -1 0 3920 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1796_
timestamp 1698431365
transform -1 0 5040 0 1 45472
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1797_
timestamp 1698431365
transform -1 0 4032 0 -1 47040
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1798_
timestamp 1698431365
transform 1 0 2800 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1799_
timestamp 1698431365
transform -1 0 2800 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1800_
timestamp 1698431365
transform -1 0 38528 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1801_
timestamp 1698431365
transform -1 0 18144 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1802_
timestamp 1698431365
transform -1 0 5152 0 -1 48608
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1803_
timestamp 1698431365
transform -1 0 4592 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1804_
timestamp 1698431365
transform 1 0 4368 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1805_
timestamp 1698431365
transform 1 0 4816 0 -1 50176
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1806_
timestamp 1698431365
transform 1 0 7168 0 1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1807_
timestamp 1698431365
transform -1 0 6160 0 1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1808_
timestamp 1698431365
transform -1 0 5264 0 1 48608
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1809_
timestamp 1698431365
transform 1 0 5488 0 1 48608
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1810_
timestamp 1698431365
transform -1 0 8400 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1811_
timestamp 1698431365
transform -1 0 7504 0 1 50176
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1812_
timestamp 1698431365
transform -1 0 5936 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1813_
timestamp 1698431365
transform -1 0 6384 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1814_
timestamp 1698431365
transform -1 0 7728 0 -1 53312
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1815_
timestamp 1698431365
transform -1 0 7056 0 1 51744
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1816_
timestamp 1698431365
transform -1 0 7952 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _1817_
timestamp 1698431365
transform 1 0 14336 0 -1 51744
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1818_
timestamp 1698431365
transform 1 0 16352 0 1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1819_
timestamp 1698431365
transform -1 0 16128 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1820_
timestamp 1698431365
transform 1 0 32480 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1821_
timestamp 1698431365
transform 1 0 33600 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1822_
timestamp 1698431365
transform 1 0 16128 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1823_
timestamp 1698431365
transform -1 0 16576 0 1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1824_
timestamp 1698431365
transform -1 0 8176 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1825_
timestamp 1698431365
transform -1 0 6608 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1826_
timestamp 1698431365
transform -1 0 6720 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1827_
timestamp 1698431365
transform -1 0 7840 0 -1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1828_
timestamp 1698431365
transform -1 0 7952 0 -1 36064
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1829_
timestamp 1698431365
transform -1 0 4592 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1830_
timestamp 1698431365
transform -1 0 5264 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1831_
timestamp 1698431365
transform -1 0 7728 0 -1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1832_
timestamp 1698431365
transform -1 0 7280 0 1 34496
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1833_
timestamp 1698431365
transform -1 0 7392 0 1 36064
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1834_
timestamp 1698431365
transform -1 0 7952 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1835_
timestamp 1698431365
transform 1 0 7056 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1836_
timestamp 1698431365
transform 1 0 6160 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1837_
timestamp 1698431365
transform -1 0 9184 0 -1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1838_
timestamp 1698431365
transform -1 0 9072 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1839_
timestamp 1698431365
transform -1 0 8848 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1840_
timestamp 1698431365
transform -1 0 11312 0 1 39200
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1841_
timestamp 1698431365
transform -1 0 6720 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1842_
timestamp 1698431365
transform -1 0 7840 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1843_
timestamp 1698431365
transform 1 0 8064 0 -1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1844_
timestamp 1698431365
transform 1 0 9408 0 -1 39200
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1845_
timestamp 1698431365
transform -1 0 9856 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1846_
timestamp 1698431365
transform -1 0 8176 0 1 40768
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1847_
timestamp 1698431365
transform 1 0 6384 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1848_
timestamp 1698431365
transform -1 0 6384 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1849_
timestamp 1698431365
transform -1 0 9520 0 1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1850_
timestamp 1698431365
transform -1 0 8400 0 -1 43904
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1851_
timestamp 1698431365
transform 1 0 7280 0 1 42336
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1852_
timestamp 1698431365
transform -1 0 7504 0 1 43904
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1853_
timestamp 1698431365
transform 1 0 6720 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1854_
timestamp 1698431365
transform 1 0 5824 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1855_
timestamp 1698431365
transform 1 0 7504 0 1 43904
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1856_
timestamp 1698431365
transform 1 0 7840 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1857_
timestamp 1698431365
transform -1 0 8176 0 1 45472
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1858_
timestamp 1698431365
transform -1 0 8848 0 1 47040
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1859_
timestamp 1698431365
transform -1 0 7504 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1860_
timestamp 1698431365
transform -1 0 8064 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1861_
timestamp 1698431365
transform -1 0 37744 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1862_
timestamp 1698431365
transform -1 0 9968 0 -1 48608
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1863_
timestamp 1698431365
transform -1 0 9744 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1864_
timestamp 1698431365
transform -1 0 9520 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1865_
timestamp 1698431365
transform 1 0 9408 0 -1 51744
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1866_
timestamp 1698431365
transform -1 0 10864 0 1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1867_
timestamp 1698431365
transform 1 0 9184 0 1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1868_
timestamp 1698431365
transform 1 0 8176 0 1 50176
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1869_
timestamp 1698431365
transform 1 0 8736 0 1 50176
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1870_
timestamp 1698431365
transform 1 0 9408 0 -1 54880
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1871_
timestamp 1698431365
transform -1 0 11872 0 1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1872_
timestamp 1698431365
transform -1 0 9856 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1873_
timestamp 1698431365
transform 1 0 9184 0 1 54880
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1874_
timestamp 1698431365
transform -1 0 10528 0 1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1875_
timestamp 1698431365
transform -1 0 11200 0 1 54880
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1876_
timestamp 1698431365
transform -1 0 13104 0 1 53312
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1877_
timestamp 1698431365
transform 1 0 12320 0 -1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1878_
timestamp 1698431365
transform -1 0 15232 0 1 53312
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1879_
timestamp 1698431365
transform 1 0 30464 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1880_
timestamp 1698431365
transform -1 0 32256 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1881_
timestamp 1698431365
transform 1 0 13776 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1882_
timestamp 1698431365
transform 1 0 13328 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1883_
timestamp 1698431365
transform -1 0 47152 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1884_
timestamp 1698431365
transform 1 0 37744 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1885_
timestamp 1698431365
transform 1 0 45808 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1886_
timestamp 1698431365
transform -1 0 46928 0 -1 42336
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1887_
timestamp 1698431365
transform -1 0 43680 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1888_
timestamp 1698431365
transform 1 0 39088 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1889_
timestamp 1698431365
transform -1 0 47488 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1890_
timestamp 1698431365
transform 1 0 46592 0 -1 40768
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1891_
timestamp 1698431365
transform -1 0 47824 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1892_
timestamp 1698431365
transform -1 0 46368 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1893_
timestamp 1698431365
transform -1 0 46032 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1894_
timestamp 1698431365
transform 1 0 43568 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1895_
timestamp 1698431365
transform 1 0 37744 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1896_
timestamp 1698431365
transform -1 0 43232 0 1 37632
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1897_
timestamp 1698431365
transform -1 0 40096 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1898_
timestamp 1698431365
transform 1 0 42224 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1899_
timestamp 1698431365
transform 1 0 32928 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1900_
timestamp 1698431365
transform 1 0 40768 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1901_
timestamp 1698431365
transform -1 0 42560 0 -1 37632
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1902_
timestamp 1698431365
transform -1 0 41776 0 -1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1903_
timestamp 1698431365
transform 1 0 41552 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1904_
timestamp 1698431365
transform -1 0 43344 0 1 36064
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1905_
timestamp 1698431365
transform -1 0 40320 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1906_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 34944 0 -1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1907_
timestamp 1698431365
transform 1 0 39424 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1908_
timestamp 1698431365
transform 1 0 41104 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1909_
timestamp 1698431365
transform 1 0 42560 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1910_
timestamp 1698431365
transform -1 0 42896 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1911_
timestamp 1698431365
transform -1 0 42448 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1912_
timestamp 1698431365
transform 1 0 40656 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1913_
timestamp 1698431365
transform -1 0 42560 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1914_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 40880 0 -1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1915_
timestamp 1698431365
transform 1 0 42784 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1916_
timestamp 1698431365
transform 1 0 41216 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1917_
timestamp 1698431365
transform 1 0 44688 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1918_
timestamp 1698431365
transform -1 0 45360 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1919_
timestamp 1698431365
transform 1 0 43232 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1920_
timestamp 1698431365
transform -1 0 44016 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1921_
timestamp 1698431365
transform -1 0 45808 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1922_
timestamp 1698431365
transform -1 0 45920 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1923_
timestamp 1698431365
transform -1 0 46480 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1924_
timestamp 1698431365
transform -1 0 45920 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1925_
timestamp 1698431365
transform 1 0 44464 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1926_
timestamp 1698431365
transform 1 0 46368 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1927_
timestamp 1698431365
transform 1 0 47376 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1928_
timestamp 1698431365
transform 1 0 46928 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1929_
timestamp 1698431365
transform 1 0 47376 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1930_
timestamp 1698431365
transform -1 0 47376 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1931_
timestamp 1698431365
transform 1 0 46816 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1932_
timestamp 1698431365
transform 1 0 44464 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1933_
timestamp 1698431365
transform 1 0 46144 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1934_
timestamp 1698431365
transform 1 0 45920 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1935_
timestamp 1698431365
transform 1 0 46592 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1936_
timestamp 1698431365
transform 1 0 45472 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1937_
timestamp 1698431365
transform 1 0 46256 0 1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1938_
timestamp 1698431365
transform -1 0 47936 0 1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1939_
timestamp 1698431365
transform -1 0 47600 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1940_
timestamp 1698431365
transform -1 0 47376 0 1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1941_
timestamp 1698431365
transform 1 0 47600 0 -1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1942_
timestamp 1698431365
transform -1 0 47488 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1943_
timestamp 1698431365
transform 1 0 47264 0 -1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1944_
timestamp 1698431365
transform -1 0 47264 0 -1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1945_
timestamp 1698431365
transform 1 0 46704 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1946_
timestamp 1698431365
transform -1 0 47152 0 1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1947_
timestamp 1698431365
transform -1 0 44576 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1948_
timestamp 1698431365
transform 1 0 45136 0 -1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1949_
timestamp 1698431365
transform -1 0 45808 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1950_
timestamp 1698431365
transform 1 0 45696 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1951_
timestamp 1698431365
transform 1 0 42336 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1952_
timestamp 1698431365
transform 1 0 44688 0 1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1953_
timestamp 1698431365
transform 1 0 43344 0 -1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1954_
timestamp 1698431365
transform 1 0 43568 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1955_
timestamp 1698431365
transform 1 0 43008 0 1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1956_
timestamp 1698431365
transform 1 0 43456 0 1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1957_
timestamp 1698431365
transform 1 0 44016 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1958_
timestamp 1698431365
transform -1 0 45024 0 -1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1959_
timestamp 1698431365
transform -1 0 45136 0 -1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1960_
timestamp 1698431365
transform 1 0 43568 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1961_
timestamp 1698431365
transform -1 0 44016 0 1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1962_
timestamp 1698431365
transform -1 0 43120 0 -1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1963_
timestamp 1698431365
transform 1 0 42672 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1964_
timestamp 1698431365
transform -1 0 39648 0 -1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1965_
timestamp 1698431365
transform 1 0 38752 0 1 28224
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1966_
timestamp 1698431365
transform 1 0 41664 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1967_
timestamp 1698431365
transform 1 0 40768 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1968_
timestamp 1698431365
transform -1 0 48384 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _1969_
timestamp 1698431365
transform 1 0 42560 0 -1 37632
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1970_
timestamp 1698431365
transform -1 0 47824 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1971_
timestamp 1698431365
transform -1 0 46592 0 1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _1972_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 44240 0 -1 39200
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_4  _1973_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 44800 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1974_
timestamp 1698431365
transform -1 0 36064 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1975_
timestamp 1698431365
transform 1 0 33936 0 1 23520
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1976_
timestamp 1698431365
transform -1 0 35056 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1977_
timestamp 1698431365
transform 1 0 38304 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1978_
timestamp 1698431365
transform -1 0 48048 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1979_
timestamp 1698431365
transform -1 0 48384 0 -1 37632
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1980_
timestamp 1698431365
transform -1 0 33824 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1981_
timestamp 1698431365
transform 1 0 26432 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1982_
timestamp 1698431365
transform 1 0 33040 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1983_
timestamp 1698431365
transform -1 0 36176 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1984_
timestamp 1698431365
transform 1 0 35728 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1985_
timestamp 1698431365
transform -1 0 36624 0 1 25088
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1986_
timestamp 1698431365
transform -1 0 35840 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1987_
timestamp 1698431365
transform 1 0 36848 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1988_
timestamp 1698431365
transform -1 0 35952 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1989_
timestamp 1698431365
transform 1 0 35616 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1990_
timestamp 1698431365
transform -1 0 35280 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1991_
timestamp 1698431365
transform 1 0 36848 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1992_
timestamp 1698431365
transform 1 0 37744 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1993_
timestamp 1698431365
transform 1 0 34272 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1994_
timestamp 1698431365
transform 1 0 36848 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1995_
timestamp 1698431365
transform 1 0 37744 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1996_
timestamp 1698431365
transform 1 0 38528 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1997_
timestamp 1698431365
transform -1 0 38528 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1998_
timestamp 1698431365
transform -1 0 39424 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1999_
timestamp 1698431365
transform -1 0 38528 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2000_
timestamp 1698431365
transform -1 0 37632 0 -1 31360
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2001_
timestamp 1698431365
transform 1 0 37072 0 -1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2002_
timestamp 1698431365
transform 1 0 37296 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2003_
timestamp 1698431365
transform -1 0 36064 0 1 29792
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2004_
timestamp 1698431365
transform -1 0 35392 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2005_
timestamp 1698431365
transform 1 0 35280 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2006_
timestamp 1698431365
transform 1 0 33376 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2007_
timestamp 1698431365
transform -1 0 33936 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2008_
timestamp 1698431365
transform -1 0 36064 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2009_
timestamp 1698431365
transform 1 0 32032 0 1 32928
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2010_
timestamp 1698431365
transform 1 0 33712 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2011_
timestamp 1698431365
transform 1 0 34608 0 -1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2012_
timestamp 1698431365
transform 1 0 33152 0 -1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2013_
timestamp 1698431365
transform 1 0 34384 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2014_
timestamp 1698431365
transform -1 0 34608 0 -1 34496
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2015_
timestamp 1698431365
transform 1 0 23520 0 -1 39200
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2016_
timestamp 1698431365
transform -1 0 26320 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2017_
timestamp 1698431365
transform -1 0 26656 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2018_
timestamp 1698431365
transform 1 0 30240 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2019_
timestamp 1698431365
transform 1 0 23408 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2020_
timestamp 1698431365
transform 1 0 24192 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2021_
timestamp 1698431365
transform 1 0 24304 0 1 39200
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2022_
timestamp 1698431365
transform 1 0 21168 0 1 40768
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2023_
timestamp 1698431365
transform 1 0 23632 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2024_
timestamp 1698431365
transform 1 0 21280 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2025_
timestamp 1698431365
transform 1 0 20384 0 1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2026_
timestamp 1698431365
transform 1 0 21952 0 1 42336
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _2027_
timestamp 1698431365
transform 1 0 25088 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2028_
timestamp 1698431365
transform -1 0 26432 0 -1 45472
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2029_
timestamp 1698431365
transform 1 0 24192 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2030_
timestamp 1698431365
transform 1 0 23296 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2031_
timestamp 1698431365
transform -1 0 26208 0 1 45472
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2032_
timestamp 1698431365
transform -1 0 25648 0 1 45472
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2033_
timestamp 1698431365
transform -1 0 25872 0 1 43904
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2034_
timestamp 1698431365
transform 1 0 26656 0 -1 47040
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2035_
timestamp 1698431365
transform -1 0 33152 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2036_
timestamp 1698431365
transform -1 0 27328 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2037_
timestamp 1698431365
transform 1 0 27664 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2038_
timestamp 1698431365
transform 1 0 28000 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2039_
timestamp 1698431365
transform -1 0 28112 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2040_
timestamp 1698431365
transform -1 0 27552 0 -1 50176
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2041_
timestamp 1698431365
transform -1 0 27776 0 -1 51744
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2042_
timestamp 1698431365
transform -1 0 25760 0 1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2043_
timestamp 1698431365
transform 1 0 27776 0 -1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2044_
timestamp 1698431365
transform -1 0 27776 0 1 50176
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2045_
timestamp 1698431365
transform -1 0 27664 0 1 51744
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2046_
timestamp 1698431365
transform 1 0 26544 0 -1 54880
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2047_
timestamp 1698431365
transform 1 0 29008 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2048_
timestamp 1698431365
transform 1 0 27888 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2049_
timestamp 1698431365
transform -1 0 28560 0 1 53312
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2050_
timestamp 1698431365
transform -1 0 28000 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2051_
timestamp 1698431365
transform -1 0 27776 0 1 54880
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2052_
timestamp 1698431365
transform 1 0 25088 0 -1 54880
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2053_
timestamp 1698431365
transform 1 0 25760 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2054_
timestamp 1698431365
transform 1 0 24864 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2055_
timestamp 1698431365
transform -1 0 23968 0 1 54880
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2056_
timestamp 1698431365
transform 1 0 23968 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2057_
timestamp 1698431365
transform 1 0 22960 0 -1 53312
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _2058_
timestamp 1698431365
transform 1 0 22176 0 -1 54880
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2059_
timestamp 1698431365
transform -1 0 23520 0 1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2060_
timestamp 1698431365
transform -1 0 22512 0 1 54880
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2061_
timestamp 1698431365
transform -1 0 23296 0 1 54880
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2062_
timestamp 1698431365
transform -1 0 22848 0 1 53312
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2063_
timestamp 1698431365
transform -1 0 18928 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2064_
timestamp 1698431365
transform 1 0 43568 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2065_
timestamp 1698431365
transform -1 0 45920 0 -1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2066_
timestamp 1698431365
transform 1 0 37184 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or4_1  _2067_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 47600 0 -1 17248
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__or4_1  _2068_
timestamp 1698431365
transform 1 0 37632 0 1 17248
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _2069_
timestamp 1698431365
transform -1 0 43120 0 1 17248
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2070_
timestamp 1698431365
transform -1 0 46144 0 1 18816
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2071_
timestamp 1698431365
transform 1 0 43792 0 1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2072_
timestamp 1698431365
transform 1 0 44464 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2073_
timestamp 1698431365
transform 1 0 33264 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2074_
timestamp 1698431365
transform 1 0 40992 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2075_
timestamp 1698431365
transform 1 0 42896 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2076_
timestamp 1698431365
transform 1 0 44352 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2077_
timestamp 1698431365
transform 1 0 34160 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2078_
timestamp 1698431365
transform 1 0 33264 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2079_
timestamp 1698431365
transform -1 0 42896 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _2080_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 43792 0 -1 18816
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2081_
timestamp 1698431365
transform -1 0 46592 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2082_
timestamp 1698431365
transform 1 0 43232 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2083_
timestamp 1698431365
transform 1 0 45584 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2084_
timestamp 1698431365
transform 1 0 45248 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _2085_
timestamp 1698431365
transform 1 0 43120 0 1 17248
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2086_
timestamp 1698431365
transform 1 0 44688 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2087_
timestamp 1698431365
transform -1 0 40544 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2088_
timestamp 1698431365
transform 1 0 40768 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2089_
timestamp 1698431365
transform 1 0 42560 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2090_
timestamp 1698431365
transform 1 0 43456 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2091_
timestamp 1698431365
transform 1 0 37184 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _2092_
timestamp 1698431365
transform -1 0 44016 0 1 15680
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2093_
timestamp 1698431365
transform 1 0 43456 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2094_
timestamp 1698431365
transform 1 0 41664 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2095_
timestamp 1698431365
transform -1 0 43456 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2096_
timestamp 1698431365
transform 1 0 38416 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2097_
timestamp 1698431365
transform 1 0 44688 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _2098_
timestamp 1698431365
transform -1 0 42560 0 -1 15680
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2099_
timestamp 1698431365
transform 1 0 42224 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2100_
timestamp 1698431365
transform 1 0 37632 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2101_
timestamp 1698431365
transform -1 0 39088 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2102_
timestamp 1698431365
transform -1 0 39984 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2103_
timestamp 1698431365
transform 1 0 40768 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _2104_
timestamp 1698431365
transform -1 0 39984 0 -1 15680
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2105_
timestamp 1698431365
transform 1 0 38976 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2106_
timestamp 1698431365
transform -1 0 38416 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2107_
timestamp 1698431365
transform 1 0 35952 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2108_
timestamp 1698431365
transform 1 0 35952 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2109_
timestamp 1698431365
transform 1 0 36960 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2110_
timestamp 1698431365
transform 1 0 35392 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _2111_
timestamp 1698431365
transform 1 0 36848 0 -1 17248
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2112_
timestamp 1698431365
transform -1 0 38640 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2113_
timestamp 1698431365
transform -1 0 37296 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2114_
timestamp 1698431365
transform -1 0 35280 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2115_
timestamp 1698431365
transform 1 0 32816 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _2116_
timestamp 1698431365
transform -1 0 35952 0 -1 18816
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2117_
timestamp 1698431365
transform 1 0 35952 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2118_
timestamp 1698431365
transform 1 0 35056 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _2119_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 35168 0 1 20384
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2120_
timestamp 1698431365
transform 1 0 33824 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2121_
timestamp 1698431365
transform -1 0 34832 0 1 18816
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2122_
timestamp 1698431365
transform -1 0 45360 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2123_
timestamp 1698431365
transform 1 0 34720 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2124_
timestamp 1698431365
transform -1 0 36512 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2125_
timestamp 1698431365
transform 1 0 36848 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2126_
timestamp 1698431365
transform -1 0 32704 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2127_
timestamp 1698431365
transform 1 0 32928 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2128_
timestamp 1698431365
transform -1 0 33712 0 1 18816
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2129_
timestamp 1698431365
transform -1 0 32592 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2130_
timestamp 1698431365
transform -1 0 31360 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2131_
timestamp 1698431365
transform 1 0 32928 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2132_
timestamp 1698431365
transform -1 0 45808 0 1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or4_1  _2133_
timestamp 1698431365
transform -1 0 44464 0 1 7840
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__or4_1  _2134_
timestamp 1698431365
transform 1 0 36288 0 -1 7840
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _2135_
timestamp 1698431365
transform -1 0 41552 0 1 7840
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2136_
timestamp 1698431365
transform 1 0 43008 0 1 9408
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2137_
timestamp 1698431365
transform 1 0 44688 0 1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2138_
timestamp 1698431365
transform -1 0 45584 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2139_
timestamp 1698431365
transform 1 0 42000 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2140_
timestamp 1698431365
transform -1 0 42000 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2141_
timestamp 1698431365
transform 1 0 42000 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2142_
timestamp 1698431365
transform 1 0 37296 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _2143_
timestamp 1698431365
transform 1 0 42224 0 1 6272
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2144_
timestamp 1698431365
transform 1 0 44016 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2145_
timestamp 1698431365
transform 1 0 43344 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2146_
timestamp 1698431365
transform -1 0 43008 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2147_
timestamp 1698431365
transform -1 0 42224 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _2148_
timestamp 1698431365
transform 1 0 42000 0 -1 7840
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2149_
timestamp 1698431365
transform 1 0 42672 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2150_
timestamp 1698431365
transform -1 0 40432 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2151_
timestamp 1698431365
transform -1 0 39200 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2152_
timestamp 1698431365
transform 1 0 39536 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2153_
timestamp 1698431365
transform 1 0 40320 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2154_
timestamp 1698431365
transform -1 0 38416 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2155_
timestamp 1698431365
transform -1 0 40320 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _2156_
timestamp 1698431365
transform 1 0 40768 0 -1 6272
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2157_
timestamp 1698431365
transform 1 0 40992 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2158_
timestamp 1698431365
transform -1 0 38080 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2159_
timestamp 1698431365
transform -1 0 40208 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2160_
timestamp 1698431365
transform -1 0 38976 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _2161_
timestamp 1698431365
transform -1 0 39312 0 -1 6272
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2162_
timestamp 1698431365
transform 1 0 37296 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2163_
timestamp 1698431365
transform 1 0 35280 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2164_
timestamp 1698431365
transform -1 0 36064 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2165_
timestamp 1698431365
transform 1 0 35280 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2166_
timestamp 1698431365
transform -1 0 34272 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _2167_
timestamp 1698431365
transform 1 0 35840 0 -1 6272
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2168_
timestamp 1698431365
transform 1 0 36176 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2169_
timestamp 1698431365
transform -1 0 36176 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2170_
timestamp 1698431365
transform 1 0 34608 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2171_
timestamp 1698431365
transform 1 0 34496 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2172_
timestamp 1698431365
transform 1 0 33936 0 -1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2173_
timestamp 1698431365
transform -1 0 35056 0 -1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _2174_
timestamp 1698431365
transform 1 0 34496 0 -1 6272
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2175_
timestamp 1698431365
transform 1 0 33376 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2176_
timestamp 1698431365
transform -1 0 37296 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2177_
timestamp 1698431365
transform 1 0 32368 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _2178_
timestamp 1698431365
transform 1 0 33936 0 1 10976
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2179_
timestamp 1698431365
transform -1 0 34384 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2180_
timestamp 1698431365
transform 1 0 35504 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _2181_
timestamp 1698431365
transform 1 0 34496 0 1 9408
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2182_
timestamp 1698431365
transform 1 0 33264 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2183_
timestamp 1698431365
transform 1 0 34496 0 1 14112
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2184_
timestamp 1698431365
transform 1 0 34160 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2185_
timestamp 1698431365
transform 1 0 33936 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2186_
timestamp 1698431365
transform 1 0 35056 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2187_
timestamp 1698431365
transform -1 0 37744 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2188_
timestamp 1698431365
transform -1 0 32368 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2189_
timestamp 1698431365
transform 1 0 30576 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2190_
timestamp 1698431365
transform 1 0 31248 0 -1 14112
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2191_
timestamp 1698431365
transform 1 0 32928 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2192_
timestamp 1698431365
transform 1 0 33824 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2193_
timestamp 1698431365
transform 1 0 13328 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2194_
timestamp 1698431365
transform 1 0 10416 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2195_
timestamp 1698431365
transform -1 0 34384 0 -1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or4_1  _2196_
timestamp 1698431365
transform 1 0 30240 0 -1 7840
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__or4_1  _2197_
timestamp 1698431365
transform 1 0 24640 0 1 7840
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _2198_
timestamp 1698431365
transform -1 0 30240 0 -1 7840
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2199_
timestamp 1698431365
transform -1 0 31360 0 1 7840
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2200_
timestamp 1698431365
transform 1 0 32928 0 -1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2201_
timestamp 1698431365
transform -1 0 33824 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2202_
timestamp 1698431365
transform -1 0 33600 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2203_
timestamp 1698431365
transform 1 0 31584 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2204_
timestamp 1698431365
transform -1 0 31808 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2205_
timestamp 1698431365
transform 1 0 31808 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _2206_
timestamp 1698431365
transform -1 0 32144 0 -1 6272
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2207_
timestamp 1698431365
transform -1 0 31360 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2208_
timestamp 1698431365
transform 1 0 29008 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2209_
timestamp 1698431365
transform -1 0 28784 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2210_
timestamp 1698431365
transform -1 0 33376 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2211_
timestamp 1698431365
transform 1 0 29904 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _2212_
timestamp 1698431365
transform -1 0 30128 0 -1 6272
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2213_
timestamp 1698431365
transform -1 0 29456 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2214_
timestamp 1698431365
transform -1 0 27216 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2215_
timestamp 1698431365
transform 1 0 26992 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2216_
timestamp 1698431365
transform -1 0 26208 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2217_
timestamp 1698431365
transform 1 0 27552 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2218_
timestamp 1698431365
transform -1 0 27104 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _2219_
timestamp 1698431365
transform 1 0 26208 0 -1 6272
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2220_
timestamp 1698431365
transform -1 0 26880 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2221_
timestamp 1698431365
transform 1 0 23632 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2222_
timestamp 1698431365
transform -1 0 23184 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2223_
timestamp 1698431365
transform 1 0 23072 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _2224_
timestamp 1698431365
transform 1 0 23968 0 1 4704
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2225_
timestamp 1698431365
transform -1 0 23072 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2226_
timestamp 1698431365
transform 1 0 23520 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2227_
timestamp 1698431365
transform 1 0 25424 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2228_
timestamp 1698431365
transform -1 0 24080 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _2229_
timestamp 1698431365
transform 1 0 24080 0 1 6272
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2230_
timestamp 1698431365
transform 1 0 21840 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2231_
timestamp 1698431365
transform 1 0 22736 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2232_
timestamp 1698431365
transform 1 0 23408 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2233_
timestamp 1698431365
transform 1 0 23968 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2234_
timestamp 1698431365
transform 1 0 23408 0 -1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2235_
timestamp 1698431365
transform -1 0 25648 0 -1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _2236_
timestamp 1698431365
transform -1 0 25760 0 1 9408
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2237_
timestamp 1698431365
transform -1 0 22848 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2238_
timestamp 1698431365
transform 1 0 25984 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2239_
timestamp 1698431365
transform 1 0 23072 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _2240_
timestamp 1698431365
transform -1 0 26656 0 -1 12544
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2241_
timestamp 1698431365
transform -1 0 27328 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2242_
timestamp 1698431365
transform 1 0 25088 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _2243_
timestamp 1698431365
transform 1 0 25200 0 1 10976
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2244_
timestamp 1698431365
transform 1 0 24640 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2245_
timestamp 1698431365
transform 1 0 25984 0 -1 15680
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2246_
timestamp 1698431365
transform 1 0 27440 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2247_
timestamp 1698431365
transform 1 0 26544 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2248_
timestamp 1698431365
transform 1 0 26768 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2249_
timestamp 1698431365
transform -1 0 25984 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2250_
timestamp 1698431365
transform 1 0 23632 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2251_
timestamp 1698431365
transform 1 0 23408 0 -1 15680
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2252_
timestamp 1698431365
transform -1 0 24640 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2253_
timestamp 1698431365
transform -1 0 16016 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2254_
timestamp 1698431365
transform -1 0 18256 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2255_
timestamp 1698431365
transform 1 0 27216 0 1 36064
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2256_
timestamp 1698431365
transform 1 0 33264 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2257_
timestamp 1698431365
transform 1 0 32928 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2258_
timestamp 1698431365
transform 1 0 33824 0 -1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2259_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 26208 0 -1 34496
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _2260_
timestamp 1698431365
transform -1 0 27104 0 1 36064
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2261_
timestamp 1698431365
transform 1 0 28336 0 -1 37632
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2262_
timestamp 1698431365
transform 1 0 33936 0 -1 37632
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2263_
timestamp 1698431365
transform 1 0 35952 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2264_
timestamp 1698431365
transform 1 0 34384 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2265_
timestamp 1698431365
transform 1 0 35056 0 1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2266_
timestamp 1698431365
transform -1 0 35840 0 1 37632
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_2  _2267_
timestamp 1698431365
transform 1 0 29008 0 1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2268_
timestamp 1698431365
transform 1 0 31136 0 -1 39200
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2269_
timestamp 1698431365
transform 1 0 32928 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2270_
timestamp 1698431365
transform -1 0 32480 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2271_
timestamp 1698431365
transform 1 0 33040 0 -1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2272_
timestamp 1698431365
transform -1 0 34720 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2273_
timestamp 1698431365
transform -1 0 36400 0 1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2274_
timestamp 1698431365
transform 1 0 28560 0 -1 40768
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2275_
timestamp 1698431365
transform -1 0 36288 0 -1 40768
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2276_
timestamp 1698431365
transform 1 0 35504 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2277_
timestamp 1698431365
transform -1 0 37296 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2278_
timestamp 1698431365
transform 1 0 32928 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2279_
timestamp 1698431365
transform 1 0 29680 0 1 42336
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2280_
timestamp 1698431365
transform 1 0 32704 0 1 40768
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2281_
timestamp 1698431365
transform 1 0 32704 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2282_
timestamp 1698431365
transform -1 0 34496 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2283_
timestamp 1698431365
transform 1 0 34496 0 1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2284_
timestamp 1698431365
transform 1 0 34720 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2285_
timestamp 1698431365
transform 1 0 33264 0 -1 45472
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2286_
timestamp 1698431365
transform -1 0 34384 0 1 43904
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2287_
timestamp 1698431365
transform -1 0 34496 0 -1 47040
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2288_
timestamp 1698431365
transform 1 0 34384 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2289_
timestamp 1698431365
transform 1 0 32592 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2290_
timestamp 1698431365
transform 1 0 31808 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2291_
timestamp 1698431365
transform 1 0 38752 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2292_
timestamp 1698431365
transform 1 0 34384 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2293_
timestamp 1698431365
transform 1 0 34944 0 -1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2294_
timestamp 1698431365
transform 1 0 33936 0 -1 45472
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2295_
timestamp 1698431365
transform 1 0 35616 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2296_
timestamp 1698431365
transform 1 0 34048 0 1 45472
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2297_
timestamp 1698431365
transform 1 0 37072 0 1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2298_
timestamp 1698431365
transform -1 0 36288 0 1 48608
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _2299_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 35840 0 1 47040
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2300_
timestamp 1698431365
transform -1 0 35728 0 1 48608
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2301_
timestamp 1698431365
transform -1 0 38416 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2302_
timestamp 1698431365
transform 1 0 33488 0 1 48608
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2303_
timestamp 1698431365
transform 1 0 34832 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2304_
timestamp 1698431365
transform 1 0 33936 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2305_
timestamp 1698431365
transform -1 0 36512 0 1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2306_
timestamp 1698431365
transform 1 0 36176 0 -1 50176
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2307_
timestamp 1698431365
transform 1 0 35728 0 -1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2308_
timestamp 1698431365
transform 1 0 33488 0 -1 53312
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2309_
timestamp 1698431365
transform -1 0 38192 0 1 51744
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2310_
timestamp 1698431365
transform -1 0 37408 0 -1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2311_
timestamp 1698431365
transform -1 0 38752 0 1 54880
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2312_
timestamp 1698431365
transform -1 0 37408 0 1 54880
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2313_
timestamp 1698431365
transform -1 0 35840 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2314_
timestamp 1698431365
transform 1 0 36064 0 1 54880
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2315_
timestamp 1698431365
transform -1 0 37856 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2316_
timestamp 1698431365
transform 1 0 39088 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2317_
timestamp 1698431365
transform -1 0 37856 0 1 53312
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2318_
timestamp 1698431365
transform -1 0 38864 0 1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2319_
timestamp 1698431365
transform -1 0 39312 0 -1 53312
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _2320_
timestamp 1698431365
transform 1 0 41776 0 1 50176
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2321_
timestamp 1698431365
transform 1 0 43792 0 1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2322_
timestamp 1698431365
transform 1 0 44688 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2323_
timestamp 1698431365
transform 1 0 43792 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2324_
timestamp 1698431365
transform 1 0 46704 0 -1 50176
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2325_
timestamp 1698431365
transform 1 0 44688 0 1 50176
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2326_
timestamp 1698431365
transform 1 0 46368 0 -1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2327_
timestamp 1698431365
transform 1 0 40768 0 -1 54880
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2328_
timestamp 1698431365
transform -1 0 43232 0 -1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2329_
timestamp 1698431365
transform -1 0 48384 0 -1 56448
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2330_
timestamp 1698431365
transform 1 0 42112 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2331_
timestamp 1698431365
transform 1 0 42560 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2332_
timestamp 1698431365
transform -1 0 41888 0 1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2333_
timestamp 1698431365
transform -1 0 45920 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2334_
timestamp 1698431365
transform -1 0 44464 0 1 43904
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2335_
timestamp 1698431365
transform -1 0 45248 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2336_
timestamp 1698431365
transform 1 0 46704 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2337_
timestamp 1698431365
transform 1 0 46144 0 -1 45472
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2338_
timestamp 1698431365
transform -1 0 48160 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2339_
timestamp 1698431365
transform 1 0 45808 0 1 47040
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2340_
timestamp 1698431365
transform -1 0 46928 0 1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2341_
timestamp 1698431365
transform -1 0 48160 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2342_
timestamp 1698431365
transform -1 0 47264 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _2343_
timestamp 1698431365
transform 1 0 40320 0 1 43904
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _2344_
timestamp 1698431365
transform -1 0 41216 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2345_
timestamp 1698431365
transform -1 0 43232 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2346_
timestamp 1698431365
transform 1 0 44688 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2347_
timestamp 1698431365
transform -1 0 46592 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2348_
timestamp 1698431365
transform -1 0 43904 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2349_
timestamp 1698431365
transform -1 0 41440 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2350_
timestamp 1698431365
transform -1 0 38976 0 1 40768
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2351_
timestamp 1698431365
transform 1 0 37520 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2352_
timestamp 1698431365
transform 1 0 31920 0 1 37632
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2353_
timestamp 1698431365
transform -1 0 38864 0 1 42336
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2354_
timestamp 1698431365
transform 1 0 36848 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2355_
timestamp 1698431365
transform 1 0 41216 0 -1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2356_
timestamp 1698431365
transform 1 0 41440 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_1  _2357_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 38864 0 1 42336
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2358_
timestamp 1698431365
transform 1 0 39872 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2359_
timestamp 1698431365
transform -1 0 39424 0 -1 43904
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2360_
timestamp 1698431365
transform 1 0 36176 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2361_
timestamp 1698431365
transform -1 0 40544 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_1  _2362_
timestamp 1698431365
transform 1 0 38304 0 -1 45472
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2363_
timestamp 1698431365
transform -1 0 38416 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_1  _2364_
timestamp 1698431365
transform 1 0 38528 0 -1 47040
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2365_
timestamp 1698431365
transform -1 0 39872 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2366_
timestamp 1698431365
transform 1 0 41104 0 -1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2367_
timestamp 1698431365
transform 1 0 40992 0 1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_1  _2368_
timestamp 1698431365
transform 1 0 38864 0 -1 50176
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2369_
timestamp 1698431365
transform -1 0 38976 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_1  _2370_
timestamp 1698431365
transform 1 0 38976 0 -1 51744
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2371_
timestamp 1698431365
transform -1 0 39984 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_2  _2372_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 39984 0 1 51744
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2373_
timestamp 1698431365
transform -1 0 40544 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_1  _2374_
timestamp 1698431365
transform 1 0 42224 0 1 54880
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2375_
timestamp 1698431365
transform -1 0 45136 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_2  _2376_
timestamp 1698431365
transform 1 0 40992 0 -1 51744
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2377_
timestamp 1698431365
transform -1 0 46592 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2378_
timestamp 1698431365
transform -1 0 43120 0 -1 48608
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2379_
timestamp 1698431365
transform 1 0 41776 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2380_
timestamp 1698431365
transform 1 0 39760 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2381_
timestamp 1698431365
transform -1 0 26768 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2382_
timestamp 1698431365
transform 1 0 25088 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2383_
timestamp 1698431365
transform 1 0 18032 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2384_
timestamp 1698431365
transform -1 0 19376 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2385_
timestamp 1698431365
transform 1 0 18592 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _2386_
timestamp 1698431365
transform 1 0 18368 0 1 21952
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _2387_
timestamp 1698431365
transform 1 0 18928 0 -1 17248
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2388_
timestamp 1698431365
transform 1 0 24864 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2389_
timestamp 1698431365
transform 1 0 21280 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2390_
timestamp 1698431365
transform 1 0 30912 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2391_
timestamp 1698431365
transform 1 0 30016 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2392_
timestamp 1698431365
transform -1 0 20944 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2393_
timestamp 1698431365
transform 1 0 22064 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2394_
timestamp 1698431365
transform 1 0 30800 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2395_
timestamp 1698431365
transform 1 0 29904 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2396_
timestamp 1698431365
transform 1 0 23408 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2397_
timestamp 1698431365
transform -1 0 28784 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2398_
timestamp 1698431365
transform -1 0 29904 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2399_
timestamp 1698431365
transform 1 0 28560 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2400_
timestamp 1698431365
transform 1 0 27888 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2401_
timestamp 1698431365
transform -1 0 26320 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2402_
timestamp 1698431365
transform 1 0 25872 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2403_
timestamp 1698431365
transform 1 0 25088 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2404_
timestamp 1698431365
transform -1 0 24640 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2405_
timestamp 1698431365
transform -1 0 23632 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2406_
timestamp 1698431365
transform -1 0 21840 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2407_
timestamp 1698431365
transform -1 0 24304 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2408_
timestamp 1698431365
transform 1 0 22512 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _2409_
timestamp 1698431365
transform 1 0 18480 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__or2_2  _2410_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 17584 0 1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _2411_
timestamp 1698431365
transform 1 0 18928 0 -1 15680
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2412_
timestamp 1698431365
transform 1 0 18592 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2413_
timestamp 1698431365
transform 1 0 19264 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2414_
timestamp 1698431365
transform 1 0 20272 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2415_
timestamp 1698431365
transform 1 0 19376 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2416_
timestamp 1698431365
transform 1 0 29680 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2417_
timestamp 1698431365
transform 1 0 21168 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2418_
timestamp 1698431365
transform -1 0 19376 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2419_
timestamp 1698431365
transform 1 0 17472 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2420_
timestamp 1698431365
transform 1 0 20048 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2421_
timestamp 1698431365
transform 1 0 20944 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2422_
timestamp 1698431365
transform 1 0 19936 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2423_
timestamp 1698431365
transform 1 0 16128 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2424_
timestamp 1698431365
transform 1 0 18480 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2425_
timestamp 1698431365
transform 1 0 21168 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2426_
timestamp 1698431365
transform 1 0 19936 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2427_
timestamp 1698431365
transform -1 0 19824 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2428_
timestamp 1698431365
transform -1 0 19824 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2429_
timestamp 1698431365
transform -1 0 20944 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2430_
timestamp 1698431365
transform 1 0 21168 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _2431_
timestamp 1698431365
transform 1 0 18368 0 -1 18816
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2432_
timestamp 1698431365
transform -1 0 18592 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2433_
timestamp 1698431365
transform -1 0 18368 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2434_
timestamp 1698431365
transform 1 0 18592 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2435_
timestamp 1698431365
transform 1 0 17920 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2436_
timestamp 1698431365
transform -1 0 19376 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2437_
timestamp 1698431365
transform 1 0 17808 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2438_
timestamp 1698431365
transform 1 0 16128 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2439_
timestamp 1698431365
transform -1 0 19264 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2440_
timestamp 1698431365
transform 1 0 17808 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2441_
timestamp 1698431365
transform 1 0 16128 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2442_
timestamp 1698431365
transform 1 0 17696 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2443_
timestamp 1698431365
transform 1 0 16128 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2444_
timestamp 1698431365
transform 1 0 17584 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2445_
timestamp 1698431365
transform 1 0 16128 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2446_
timestamp 1698431365
transform -1 0 32480 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2447_
timestamp 1698431365
transform 1 0 17808 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2448_
timestamp 1698431365
transform 1 0 17024 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2449_
timestamp 1698431365
transform -1 0 24864 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _2450_
timestamp 1698431365
transform 1 0 19600 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2451_
timestamp 1698431365
transform -1 0 24192 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2452_
timestamp 1698431365
transform -1 0 21952 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2453_
timestamp 1698431365
transform 1 0 19488 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _2454_
timestamp 1698431365
transform 1 0 19824 0 1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2455_
timestamp 1698431365
transform 1 0 20832 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2456_
timestamp 1698431365
transform 1 0 21056 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2457_
timestamp 1698431365
transform 1 0 21728 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2458_
timestamp 1698431365
transform 1 0 24304 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2459_
timestamp 1698431365
transform 1 0 23632 0 1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2460_
timestamp 1698431365
transform 1 0 24304 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2461_
timestamp 1698431365
transform -1 0 21840 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2462_
timestamp 1698431365
transform -1 0 23632 0 1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2463_
timestamp 1698431365
transform -1 0 24080 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2464_
timestamp 1698431365
transform -1 0 22400 0 1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2465_
timestamp 1698431365
transform -1 0 23520 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2466_
timestamp 1698431365
transform 1 0 22400 0 1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2467_
timestamp 1698431365
transform -1 0 24192 0 1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2468_
timestamp 1698431365
transform 1 0 21840 0 -1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _2469_
timestamp 1698431365
transform 1 0 19824 0 -1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2470_
timestamp 1698431365
transform -1 0 20160 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2471_
timestamp 1698431365
transform -1 0 19600 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2472_
timestamp 1698431365
transform 1 0 19040 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2473_
timestamp 1698431365
transform -1 0 21168 0 -1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2474_
timestamp 1698431365
transform 1 0 19152 0 -1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2475_
timestamp 1698431365
transform -1 0 20608 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2476_
timestamp 1698431365
transform -1 0 20496 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2477_
timestamp 1698431365
transform -1 0 18704 0 -1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2478_
timestamp 1698431365
transform -1 0 19824 0 -1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2479_
timestamp 1698431365
transform 1 0 18928 0 1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2480_
timestamp 1698431365
transform -1 0 20832 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2481_
timestamp 1698431365
transform -1 0 18592 0 -1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2482_
timestamp 1698431365
transform -1 0 21728 0 1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _2483_
timestamp 1698431365
transform -1 0 20832 0 -1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2484_
timestamp 1698431365
transform -1 0 20720 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2485_
timestamp 1698431365
transform -1 0 13104 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2486_
timestamp 1698431365
transform -1 0 10080 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2487_
timestamp 1698431365
transform 1 0 11424 0 1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2488_
timestamp 1698431365
transform 1 0 11312 0 -1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2489_
timestamp 1698431365
transform -1 0 14784 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2490_
timestamp 1698431365
transform -1 0 16128 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2491_
timestamp 1698431365
transform -1 0 11312 0 -1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2492_
timestamp 1698431365
transform -1 0 15456 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2493_
timestamp 1698431365
transform -1 0 12320 0 -1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2494_
timestamp 1698431365
transform 1 0 9520 0 -1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2495_
timestamp 1698431365
transform -1 0 12656 0 1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _2496_
timestamp 1698431365
transform -1 0 19824 0 1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2497_
timestamp 1698431365
transform -1 0 22960 0 -1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2498_
timestamp 1698431365
transform -1 0 15008 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2499_
timestamp 1698431365
transform -1 0 14000 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2500_
timestamp 1698431365
transform -1 0 14896 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2501_
timestamp 1698431365
transform -1 0 14336 0 -1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2502_
timestamp 1698431365
transform 1 0 15344 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2503_
timestamp 1698431365
transform 1 0 28000 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2504_
timestamp 1698431365
transform -1 0 14448 0 1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2505_
timestamp 1698431365
transform 1 0 12544 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2506_
timestamp 1698431365
transform 1 0 14448 0 1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2507_
timestamp 1698431365
transform -1 0 15568 0 -1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2508_
timestamp 1698431365
transform -1 0 13104 0 1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2509_
timestamp 1698431365
transform -1 0 17024 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2510_
timestamp 1698431365
transform 1 0 17136 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2511_
timestamp 1698431365
transform 1 0 16240 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2512_
timestamp 1698431365
transform 1 0 17472 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2513_
timestamp 1698431365
transform 1 0 16128 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2514_
timestamp 1698431365
transform 1 0 17248 0 -1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2515_
timestamp 1698431365
transform 1 0 15568 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2516_
timestamp 1698431365
transform 1 0 34496 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2517_
timestamp 1698431365
transform -1 0 31808 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2518_
timestamp 1698431365
transform -1 0 30576 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2519_
timestamp 1698431365
transform 1 0 30240 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2520_
timestamp 1698431365
transform 1 0 29232 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2521_
timestamp 1698431365
transform 1 0 31248 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2522_
timestamp 1698431365
transform 1 0 30352 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2523_
timestamp 1698431365
transform -1 0 32704 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2524_
timestamp 1698431365
transform 1 0 29456 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2525_
timestamp 1698431365
transform -1 0 30464 0 1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2526_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 35280 0 -1 56448
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2527_
timestamp 1698431365
transform 1 0 29120 0 1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2528_
timestamp 1698431365
transform 1 0 29344 0 1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2529_
timestamp 1698431365
transform 1 0 26544 0 -1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2530_
timestamp 1698431365
transform 1 0 25760 0 -1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2531_
timestamp 1698431365
transform 1 0 42336 0 -1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2532_
timestamp 1698431365
transform 1 0 40768 0 -1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2533_
timestamp 1698431365
transform 1 0 40768 0 -1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2534_
timestamp 1698431365
transform 1 0 37072 0 1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2535_
timestamp 1698431365
transform 1 0 41664 0 -1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2536_
timestamp 1698431365
transform 1 0 39312 0 1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2537_
timestamp 1698431365
transform 1 0 40768 0 -1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2538_
timestamp 1698431365
transform 1 0 37408 0 1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2539_
timestamp 1698431365
transform 1 0 30128 0 1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2540_
timestamp 1698431365
transform -1 0 33264 0 1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2541_
timestamp 1698431365
transform 1 0 15456 0 1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2542_
timestamp 1698431365
transform -1 0 20272 0 1 42336
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2543_
timestamp 1698431365
transform 1 0 12432 0 -1 42336
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2544_
timestamp 1698431365
transform 1 0 12768 0 -1 45472
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2545_
timestamp 1698431365
transform 1 0 17248 0 -1 45472
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2546_
timestamp 1698431365
transform 1 0 17248 0 -1 48608
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2547_
timestamp 1698431365
transform 1 0 17248 0 -1 51744
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2548_
timestamp 1698431365
transform 1 0 13440 0 1 47040
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2549_
timestamp 1698431365
transform 1 0 16800 0 -1 56448
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2550_
timestamp 1698431365
transform 1 0 1568 0 1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2551_
timestamp 1698431365
transform -1 0 4816 0 -1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2552_
timestamp 1698431365
transform 1 0 1568 0 1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2553_
timestamp 1698431365
transform -1 0 4816 0 -1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2554_
timestamp 1698431365
transform 1 0 1568 0 -1 42336
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2555_
timestamp 1698431365
transform 1 0 1568 0 1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2556_
timestamp 1698431365
transform 1 0 1568 0 1 47040
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2557_
timestamp 1698431365
transform 1 0 1568 0 -1 50176
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2558_
timestamp 1698431365
transform 1 0 3920 0 -1 53312
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2559_
timestamp 1698431365
transform -1 0 18592 0 1 51744
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2560_
timestamp 1698431365
transform 1 0 14448 0 1 54880
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2561_
timestamp 1698431365
transform 1 0 4032 0 -1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2562_
timestamp 1698431365
transform 1 0 3920 0 -1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2563_
timestamp 1698431365
transform 1 0 4928 0 -1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2564_
timestamp 1698431365
transform 1 0 5488 0 1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2565_
timestamp 1698431365
transform 1 0 5152 0 -1 42336
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2566_
timestamp 1698431365
transform 1 0 4592 0 -1 45472
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2567_
timestamp 1698431365
transform 1 0 5600 0 -1 48608
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2568_
timestamp 1698431365
transform 1 0 5936 0 -1 51744
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2569_
timestamp 1698431365
transform 1 0 5936 0 -1 54880
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2570_
timestamp 1698431365
transform 1 0 11088 0 -1 53312
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2571_
timestamp 1698431365
transform 1 0 12992 0 -1 54880
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2572_
timestamp 1698431365
transform 1 0 45136 0 1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2573_
timestamp 1698431365
transform 1 0 42448 0 -1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2574_
timestamp 1698431365
transform 1 0 45136 0 1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2575_
timestamp 1698431365
transform 1 0 43680 0 -1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2576_
timestamp 1698431365
transform 1 0 38528 0 1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2577_
timestamp 1698431365
transform 1 0 40880 0 -1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2578_
timestamp 1698431365
transform 1 0 38752 0 1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2579_
timestamp 1698431365
transform -1 0 41328 0 1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2580_
timestamp 1698431365
transform -1 0 44464 0 -1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2581_
timestamp 1698431365
transform -1 0 47936 0 1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2582_
timestamp 1698431365
transform -1 0 48384 0 1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2583_
timestamp 1698431365
transform -1 0 48384 0 1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2584_
timestamp 1698431365
transform 1 0 45136 0 1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2585_
timestamp 1698431365
transform -1 0 48384 0 -1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2586_
timestamp 1698431365
transform 1 0 44688 0 -1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2587_
timestamp 1698431365
transform 1 0 45136 0 1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2588_
timestamp 1698431365
transform 1 0 45136 0 -1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2589_
timestamp 1698431365
transform 1 0 42448 0 -1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2590_
timestamp 1698431365
transform 1 0 40768 0 -1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2591_
timestamp 1698431365
transform 1 0 41104 0 1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2592_
timestamp 1698431365
transform 1 0 41216 0 1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2593_
timestamp 1698431365
transform 1 0 39312 0 1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2594_
timestamp 1698431365
transform 1 0 32928 0 -1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2595_
timestamp 1698431365
transform -1 0 39424 0 -1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2596_
timestamp 1698431365
transform 1 0 32368 0 1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2597_
timestamp 1698431365
transform -1 0 39312 0 -1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2598_
timestamp 1698431365
transform -1 0 40656 0 1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2599_
timestamp 1698431365
transform -1 0 40096 0 1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2600_
timestamp 1698431365
transform 1 0 32928 0 -1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2601_
timestamp 1698431365
transform 1 0 31136 0 1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2602_
timestamp 1698431365
transform 1 0 33376 0 1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2603_
timestamp 1698431365
transform -1 0 28336 0 -1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2604_
timestamp 1698431365
transform 1 0 19600 0 -1 42336
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2605_
timestamp 1698431365
transform 1 0 21616 0 -1 45472
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2606_
timestamp 1698431365
transform 1 0 24416 0 1 47040
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2607_
timestamp 1698431365
transform 1 0 23968 0 1 50176
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2608_
timestamp 1698431365
transform -1 0 31136 0 -1 54880
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2609_
timestamp 1698431365
transform 1 0 23968 0 1 54880
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2610_
timestamp 1698431365
transform 1 0 18928 0 -1 54880
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2611_
timestamp 1698431365
transform 1 0 17696 0 1 54880
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2612_
timestamp 1698431365
transform 1 0 44688 0 1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2613_
timestamp 1698431365
transform 1 0 45136 0 -1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2614_
timestamp 1698431365
transform 1 0 45136 0 1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2615_
timestamp 1698431365
transform 1 0 43904 0 -1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2616_
timestamp 1698431365
transform -1 0 44464 0 1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2617_
timestamp 1698431365
transform -1 0 41216 0 1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2618_
timestamp 1698431365
transform 1 0 34944 0 -1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2619_
timestamp 1698431365
transform 1 0 35056 0 -1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2620_
timestamp 1698431365
transform 1 0 35952 0 -1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2621_
timestamp 1698431365
transform 1 0 31360 0 1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2622_
timestamp 1698431365
transform 1 0 15904 0 1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2623_
timestamp 1698431365
transform -1 0 47600 0 -1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2624_
timestamp 1698431365
transform -1 0 47936 0 1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2625_
timestamp 1698431365
transform -1 0 47264 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2626_
timestamp 1698431365
transform 1 0 40768 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2627_
timestamp 1698431365
transform -1 0 40992 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2628_
timestamp 1698431365
transform -1 0 39424 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2629_
timestamp 1698431365
transform 1 0 32928 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2630_
timestamp 1698431365
transform 1 0 34272 0 -1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2631_
timestamp 1698431365
transform 1 0 34384 0 -1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2632_
timestamp 1698431365
transform -1 0 34496 0 1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_4  _2633_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 11536 0 1 18816
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2634_
timestamp 1698431365
transform -1 0 34608 0 1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2635_
timestamp 1698431365
transform 1 0 29680 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2636_
timestamp 1698431365
transform 1 0 27216 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2637_
timestamp 1698431365
transform 1 0 25312 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2638_
timestamp 1698431365
transform 1 0 21392 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2639_
timestamp 1698431365
transform 1 0 21168 0 -1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2640_
timestamp 1698431365
transform 1 0 21168 0 1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2641_
timestamp 1698431365
transform -1 0 24864 0 -1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2642_
timestamp 1698431365
transform -1 0 28784 0 1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2643_
timestamp 1698431365
transform 1 0 23408 0 1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_4  _2644_
timestamp 1698431365
transform -1 0 17360 0 1 28224
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2645_
timestamp 1698431365
transform 1 0 31136 0 1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2646_
timestamp 1698431365
transform -1 0 38752 0 -1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2647_
timestamp 1698431365
transform 1 0 32256 0 1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2648_
timestamp 1698431365
transform -1 0 37856 0 -1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2649_
timestamp 1698431365
transform -1 0 36176 0 -1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2650_
timestamp 1698431365
transform 1 0 30688 0 1 45472
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2651_
timestamp 1698431365
transform -1 0 39424 0 -1 48608
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2652_
timestamp 1698431365
transform 1 0 32928 0 -1 50176
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2653_
timestamp 1698431365
transform -1 0 36176 0 -1 54880
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2654_
timestamp 1698431365
transform -1 0 39088 0 -1 56448
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2655_
timestamp 1698431365
transform -1 0 48384 0 -1 51744
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2656_
timestamp 1698431365
transform -1 0 48384 0 1 53312
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2657_
timestamp 1698431365
transform -1 0 48384 0 1 54880
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2658_
timestamp 1698431365
transform 1 0 41104 0 1 42336
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2659_
timestamp 1698431365
transform 1 0 43456 0 -1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2660_
timestamp 1698431365
transform -1 0 48384 0 1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2661_
timestamp 1698431365
transform -1 0 48384 0 -1 48608
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2662_
timestamp 1698431365
transform -1 0 48384 0 -1 47040
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2663_
timestamp 1698431365
transform 1 0 29792 0 1 54880
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2664_
timestamp 1698431365
transform -1 0 44464 0 -1 47040
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2665_
timestamp 1698431365
transform 1 0 37296 0 -1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2666_
timestamp 1698431365
transform 1 0 35392 0 -1 42336
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2667_
timestamp 1698431365
transform -1 0 42448 0 1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2668_
timestamp 1698431365
transform 1 0 35056 0 -1 45472
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2669_
timestamp 1698431365
transform 1 0 36848 0 1 45472
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2670_
timestamp 1698431365
transform 1 0 37968 0 1 47040
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2671_
timestamp 1698431365
transform 1 0 37744 0 1 50176
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2672_
timestamp 1698431365
transform 1 0 38304 0 1 53312
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2673_
timestamp 1698431365
transform 1 0 38976 0 1 54880
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2674_
timestamp 1698431365
transform -1 0 44576 0 -1 54880
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2675_
timestamp 1698431365
transform -1 0 46032 0 -1 50176
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2676_
timestamp 1698431365
transform 1 0 41216 0 1 48608
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2677_
timestamp 1698431365
transform 1 0 40096 0 1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2678_
timestamp 1698431365
transform 1 0 29008 0 1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2679_
timestamp 1698431365
transform 1 0 29232 0 1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2680_
timestamp 1698431365
transform -1 0 30352 0 -1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2681_
timestamp 1698431365
transform 1 0 26768 0 -1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2682_
timestamp 1698431365
transform 1 0 25088 0 -1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2683_
timestamp 1698431365
transform 1 0 21616 0 1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2684_
timestamp 1698431365
transform 1 0 17696 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2685_
timestamp 1698431365
transform 1 0 18144 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2686_
timestamp 1698431365
transform 1 0 19040 0 -1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2687_
timestamp 1698431365
transform 1 0 19040 0 -1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2688_
timestamp 1698431365
transform 1 0 21168 0 1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2689_
timestamp 1698431365
transform 1 0 19824 0 -1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2690_
timestamp 1698431365
transform 1 0 16240 0 1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2691_
timestamp 1698431365
transform 1 0 15120 0 1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2692_
timestamp 1698431365
transform 1 0 14784 0 1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2693_
timestamp 1698431365
transform 1 0 14672 0 1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2694_
timestamp 1698431365
transform 1 0 13776 0 -1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2695_
timestamp 1698431365
transform 1 0 15120 0 1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2696_
timestamp 1698431365
transform 1 0 24752 0 1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2697_
timestamp 1698431365
transform 1 0 22736 0 1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _2698_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 21168 0 1 26656
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2699_
timestamp 1698431365
transform -1 0 24304 0 -1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2700_
timestamp 1698431365
transform 1 0 15232 0 1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2701_
timestamp 1698431365
transform 1 0 16128 0 1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2702_
timestamp 1698431365
transform 1 0 18480 0 -1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2703_
timestamp 1698431365
transform -1 0 19040 0 1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2704_
timestamp 1698431365
transform -1 0 6272 0 -1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2705_
timestamp 1698431365
transform -1 0 6608 0 -1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_4  _2706_
timestamp 1698431365
transform 1 0 4592 0 -1 21952
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2707_
timestamp 1698431365
transform -1 0 8848 0 -1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2708_
timestamp 1698431365
transform 1 0 13328 0 1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_4  _2709_
timestamp 1698431365
transform -1 0 15008 0 -1 26656
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _2710_
timestamp 1698431365
transform 1 0 12880 0 -1 25088
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _2711_
timestamp 1698431365
transform 1 0 11424 0 -1 18816
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2712_
timestamp 1698431365
transform 1 0 13888 0 1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2713_
timestamp 1698431365
transform 1 0 13776 0 -1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2714_
timestamp 1698431365
transform -1 0 17248 0 1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2715_
timestamp 1698431365
transform 1 0 37632 0 1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2716_
timestamp 1698431365
transform 1 0 28112 0 -1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2717_
timestamp 1698431365
transform 1 0 30576 0 1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2718_
timestamp 1698431365
transform 1 0 29008 0 -1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1338__A1 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 24192 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1338__A2
timestamp 1698431365
transform 1 0 26432 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1371__A2
timestamp 1698431365
transform 1 0 30688 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1375__A2
timestamp 1698431365
transform -1 0 28784 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1433__A1
timestamp 1698431365
transform 1 0 20720 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1451__I
timestamp 1698431365
transform 1 0 22400 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1506__A2
timestamp 1698431365
transform -1 0 19264 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1511__A1
timestamp 1698431365
transform 1 0 22736 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1537__I
timestamp 1698431365
transform 1 0 23968 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1546__A1
timestamp 1698431365
transform 1 0 9744 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1547__I
timestamp 1698431365
transform 1 0 10416 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1561__A2
timestamp 1698431365
transform 1 0 24640 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1563__A1
timestamp 1698431365
transform 1 0 25312 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1570__I
timestamp 1698431365
transform -1 0 25536 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1574__I
timestamp 1698431365
transform 1 0 23296 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1592__A2
timestamp 1698431365
transform 1 0 13552 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1603__A1
timestamp 1698431365
transform -1 0 24192 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1606__A1
timestamp 1698431365
transform 1 0 12992 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1607__I
timestamp 1698431365
transform 1 0 13328 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1611__I
timestamp 1698431365
transform -1 0 10752 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1612__A2
timestamp 1698431365
transform 1 0 12208 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1620__I
timestamp 1698431365
transform -1 0 23520 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1627__A2
timestamp 1698431365
transform 1 0 30800 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1633__A2
timestamp 1698431365
transform 1 0 33152 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1637__A1
timestamp 1698431365
transform -1 0 40320 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1641__I
timestamp 1698431365
transform -1 0 25648 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1642__I
timestamp 1698431365
transform -1 0 28112 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1643__I
timestamp 1698431365
transform -1 0 23408 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1644__I
timestamp 1698431365
transform 1 0 22624 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1645__A1
timestamp 1698431365
transform -1 0 18032 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1650__A1
timestamp 1698431365
transform 1 0 32144 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1651__I
timestamp 1698431365
transform 1 0 34384 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1654__C
timestamp 1698431365
transform 1 0 29568 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1656__I
timestamp 1698431365
transform -1 0 31136 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1657__I
timestamp 1698431365
transform 1 0 30464 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1658__I
timestamp 1698431365
transform -1 0 10976 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1659__I
timestamp 1698431365
transform 1 0 27664 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1660__I
timestamp 1698431365
transform 1 0 38416 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1662__A1
timestamp 1698431365
transform 1 0 31920 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1663__I
timestamp 1698431365
transform 1 0 31584 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1664__I
timestamp 1698431365
transform 1 0 29120 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1666__A1
timestamp 1698431365
transform -1 0 28784 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1668__I
timestamp 1698431365
transform -1 0 39648 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1670__A1
timestamp 1698431365
transform -1 0 27888 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1672__I
timestamp 1698431365
transform 1 0 28672 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1677__A1
timestamp 1698431365
transform 1 0 42336 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1678__C
timestamp 1698431365
transform 1 0 41888 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1680__A1
timestamp 1698431365
transform -1 0 39648 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1681__I
timestamp 1698431365
transform 1 0 38080 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1683__A1
timestamp 1698431365
transform -1 0 40992 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1685__A1
timestamp 1698431365
transform -1 0 39536 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1687__A1
timestamp 1698431365
transform 1 0 23408 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1691__A1
timestamp 1698431365
transform -1 0 44240 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1692__C
timestamp 1698431365
transform 1 0 43904 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1694__A1
timestamp 1698431365
transform 1 0 42784 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1696__A1
timestamp 1698431365
transform -1 0 40544 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1697__I
timestamp 1698431365
transform -1 0 13776 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1698__I
timestamp 1698431365
transform -1 0 13776 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1699__B
timestamp 1698431365
transform 1 0 39536 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1700__A1
timestamp 1698431365
transform -1 0 39200 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1701__B
timestamp 1698431365
transform 1 0 30800 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1703__I
timestamp 1698431365
transform 1 0 41440 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1708__A1
timestamp 1698431365
transform 1 0 31808 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1713__B
timestamp 1698431365
transform -1 0 16128 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1717__I
timestamp 1698431365
transform -1 0 17696 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1728__B
timestamp 1698431365
transform 1 0 16800 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1734__I
timestamp 1698431365
transform 1 0 8400 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1735__B
timestamp 1698431365
transform 1 0 14896 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1752__I
timestamp 1698431365
transform 1 0 18816 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1758__A1
timestamp 1698431365
transform -1 0 17136 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1760__B
timestamp 1698431365
transform 1 0 15344 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1763__B
timestamp 1698431365
transform 1 0 4928 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1767__A1
timestamp 1698431365
transform 1 0 5712 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1775__A1
timestamp 1698431365
transform -1 0 2464 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1779__A1
timestamp 1698431365
transform 1 0 5712 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1785__B
timestamp 1698431365
transform -1 0 2688 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1791__I
timestamp 1698431365
transform -1 0 6384 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1792__B
timestamp 1698431365
transform 1 0 5712 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1798__B
timestamp 1698431365
transform 1 0 3696 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1801__I
timestamp 1698431365
transform -1 0 17248 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1806__A1
timestamp 1698431365
transform 1 0 7840 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1812__B
timestamp 1698431365
transform 1 0 4816 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1818__A1
timestamp 1698431365
transform -1 0 17472 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1821__I
timestamp 1698431365
transform 1 0 33376 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1822__B
timestamp 1698431365
transform 1 0 17472 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1825__B
timestamp 1698431365
transform 1 0 6944 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1829__A1
timestamp 1698431365
transform 1 0 4704 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1834__I
timestamp 1698431365
transform -1 0 8400 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1841__A1
timestamp 1698431365
transform 1 0 6944 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1861__I
timestamp 1698431365
transform -1 0 37968 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1866__A1
timestamp 1698431365
transform 1 0 11088 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1871__A1
timestamp 1698431365
transform -1 0 12320 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1877__A1
timestamp 1698431365
transform 1 0 13552 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1879__I
timestamp 1698431365
transform 1 0 29344 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1881__B
timestamp 1698431365
transform -1 0 15680 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1885__A2
timestamp 1698431365
transform -1 0 45808 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1887__A1
timestamp 1698431365
transform 1 0 42784 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1891__A1
timestamp 1698431365
transform 1 0 46704 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1894__A1
timestamp 1698431365
transform 1 0 43344 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1895__I
timestamp 1698431365
transform 1 0 38080 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1897__A1
timestamp 1698431365
transform 1 0 40208 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1900__I
timestamp 1698431365
transform 1 0 41888 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1905__A1
timestamp 1698431365
transform 1 0 39536 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1906__I3
timestamp 1698431365
transform -1 0 35728 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1968__I
timestamp 1698431365
transform 1 0 48048 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1974__I
timestamp 1698431365
transform 1 0 37072 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1976__A1
timestamp 1698431365
transform 1 0 34832 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1980__I
timestamp 1698431365
transform -1 0 34272 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1984__A2
timestamp 1698431365
transform -1 0 35728 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1985__A3
timestamp 1698431365
transform 1 0 37520 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1987__A1
timestamp 1698431365
transform 1 0 37968 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1989__B
timestamp 1698431365
transform 1 0 36176 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1993__I
timestamp 1698431365
transform 1 0 35392 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1994__B
timestamp 1698431365
transform 1 0 37072 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1997__B
timestamp 1698431365
transform 1 0 37408 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2004__A1
timestamp 1698431365
transform 1 0 36064 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2006__B
timestamp 1698431365
transform -1 0 36512 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2016__B
timestamp 1698431365
transform 1 0 26544 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2018__I
timestamp 1698431365
transform 1 0 31360 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2023__A1
timestamp 1698431365
transform 1 0 24528 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2029__B
timestamp 1698431365
transform 1 0 25312 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2036__B
timestamp 1698431365
transform 1 0 26432 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2042__A1
timestamp 1698431365
transform 1 0 25760 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2047__B
timestamp 1698431365
transform -1 0 30352 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2052__A2
timestamp 1698431365
transform 1 0 25312 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2053__B
timestamp 1698431365
transform -1 0 27104 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2055__A2
timestamp 1698431365
transform -1 0 21952 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2056__A2
timestamp 1698431365
transform 1 0 23744 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2059__A1
timestamp 1698431365
transform 1 0 24192 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2062__C
timestamp 1698431365
transform -1 0 21728 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2064__I
timestamp 1698431365
transform -1 0 45808 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2065__A2
timestamp 1698431365
transform 1 0 46144 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2071__A1
timestamp 1698431365
transform -1 0 43792 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2072__B
timestamp 1698431365
transform 1 0 44240 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2079__B
timestamp 1698431365
transform -1 0 43008 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2080__C
timestamp 1698431365
transform 1 0 44240 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2084__B
timestamp 1698431365
transform 1 0 47824 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2085__C
timestamp 1698431365
transform -1 0 43120 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2090__B
timestamp 1698431365
transform 1 0 43344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2091__I
timestamp 1698431365
transform 1 0 36960 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2110__A1
timestamp 1698431365
transform 1 0 35168 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2114__I
timestamp 1698431365
transform -1 0 35728 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2119__A2
timestamp 1698431365
transform -1 0 36848 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2119__C
timestamp 1698431365
transform -1 0 37744 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2122__I
timestamp 1698431365
transform -1 0 46256 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2124__A2
timestamp 1698431365
transform 1 0 39424 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2125__B
timestamp 1698431365
transform 1 0 38640 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2129__A1
timestamp 1698431365
transform -1 0 31136 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2130__A1
timestamp 1698431365
transform 1 0 32480 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2130__B
timestamp 1698431365
transform 1 0 34496 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2131__A1
timestamp 1698431365
transform -1 0 34160 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2132__A2
timestamp 1698431365
transform 1 0 45360 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2137__A1
timestamp 1698431365
transform 1 0 46032 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2138__B
timestamp 1698431365
transform 1 0 45808 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2142__I
timestamp 1698431365
transform -1 0 37296 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2158__A1
timestamp 1698431365
transform -1 0 36624 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2166__I
timestamp 1698431365
transform -1 0 32704 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2173__A1
timestamp 1698431365
transform -1 0 34496 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2181__A2
timestamp 1698431365
transform -1 0 36176 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2181__C
timestamp 1698431365
transform -1 0 36624 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2185__A2
timestamp 1698431365
transform 1 0 35056 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2186__B
timestamp 1698431365
transform 1 0 36176 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2189__A2
timestamp 1698431365
transform 1 0 31696 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2191__A1
timestamp 1698431365
transform 1 0 33824 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2193__A2
timestamp 1698431365
transform 1 0 13552 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2193__B
timestamp 1698431365
transform -1 0 14672 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2194__A2
timestamp 1698431365
transform 1 0 11984 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2195__A2
timestamp 1698431365
transform 1 0 35056 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2200__A1
timestamp 1698431365
transform 1 0 33712 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2201__B
timestamp 1698431365
transform -1 0 34832 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2218__I
timestamp 1698431365
transform 1 0 27328 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2229__A2
timestamp 1698431365
transform 1 0 25424 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2235__A1
timestamp 1698431365
transform -1 0 26208 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2236__A2
timestamp 1698431365
transform 1 0 25760 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2243__A2
timestamp 1698431365
transform 1 0 26656 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2243__C
timestamp 1698431365
transform 1 0 27104 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2248__B
timestamp 1698431365
transform 1 0 27888 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2250__A2
timestamp 1698431365
transform -1 0 23632 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2252__A1
timestamp 1698431365
transform -1 0 23072 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2253__A2
timestamp 1698431365
transform -1 0 8736 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2253__B
timestamp 1698431365
transform 1 0 25984 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2254__A2
timestamp 1698431365
transform 1 0 18928 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2256__B
timestamp 1698431365
transform 1 0 32480 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2260__A1
timestamp 1698431365
transform 1 0 25984 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2260__A2
timestamp 1698431365
transform -1 0 24864 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2261__A2
timestamp 1698431365
transform -1 0 27552 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2263__A1
timestamp 1698431365
transform 1 0 37072 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2269__B
timestamp 1698431365
transform 1 0 36400 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2276__A1
timestamp 1698431365
transform -1 0 37184 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2289__B
timestamp 1698431365
transform 1 0 33712 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2296__A2
timestamp 1698431365
transform -1 0 37296 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2297__A1
timestamp 1698431365
transform 1 0 37744 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2298__A2
timestamp 1698431365
transform 1 0 37072 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2303__B
timestamp 1698431365
transform 1 0 37520 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2310__A1
timestamp 1698431365
transform 1 0 38080 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2315__B
timestamp 1698431365
transform 1 0 36400 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2321__A1
timestamp 1698431365
transform 1 0 44912 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2326__A2
timestamp 1698431365
transform 1 0 38976 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2329__C
timestamp 1698431365
transform 1 0 47152 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2334__C
timestamp 1698431365
transform 1 0 44912 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2345__B
timestamp 1698431365
transform 1 0 43456 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2348__A1
timestamp 1698431365
transform 1 0 44128 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2350__A2
timestamp 1698431365
transform 1 0 40992 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2353__A2
timestamp 1698431365
transform 1 0 40656 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2354__A2
timestamp 1698431365
transform 1 0 37744 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2359__A2
timestamp 1698431365
transform 1 0 40096 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2360__A2
timestamp 1698431365
transform 1 0 37296 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2368__C2
timestamp 1698431365
transform 1 0 38640 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2379__A2
timestamp 1698431365
transform 1 0 40544 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2380__A1
timestamp 1698431365
transform -1 0 39760 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2381__I
timestamp 1698431365
transform 1 0 28336 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2385__I
timestamp 1698431365
transform 1 0 19152 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2390__B
timestamp 1698431365
transform -1 0 32256 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2391__A1
timestamp 1698431365
transform 1 0 29792 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2392__I
timestamp 1698431365
transform 1 0 18480 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2395__A1
timestamp 1698431365
transform 1 0 30800 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2398__A1
timestamp 1698431365
transform 1 0 29680 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2400__A1
timestamp 1698431365
transform -1 0 27888 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2404__I
timestamp 1698431365
transform -1 0 24864 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2410__A2
timestamp 1698431365
transform -1 0 19824 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2414__A1
timestamp 1698431365
transform -1 0 21616 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2415__A1
timestamp 1698431365
transform 1 0 20272 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2416__I
timestamp 1698431365
transform 1 0 30800 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2418__A1
timestamp 1698431365
transform -1 0 18480 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2419__I
timestamp 1698431365
transform 1 0 19600 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2422__A1
timestamp 1698431365
transform -1 0 19936 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2423__I
timestamp 1698431365
transform 1 0 15120 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2426__A1
timestamp 1698431365
transform 1 0 19712 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2435__A1
timestamp 1698431365
transform 1 0 19040 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2438__A1
timestamp 1698431365
transform 1 0 17472 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2441__A1
timestamp 1698431365
transform -1 0 16128 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2443__A1
timestamp 1698431365
transform 1 0 17472 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2447__B
timestamp 1698431365
transform -1 0 18928 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2452__A1
timestamp 1698431365
transform 1 0 21952 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2452__A2
timestamp 1698431365
transform 1 0 22176 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2459__C
timestamp 1698431365
transform 1 0 25312 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2462__A1
timestamp 1698431365
transform 1 0 22288 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2464__A1
timestamp 1698431365
transform 1 0 22624 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2466__A1
timestamp 1698431365
transform -1 0 22400 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2477__A1
timestamp 1698431365
transform 1 0 20720 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2479__A1
timestamp 1698431365
transform 1 0 20720 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2481__A1
timestamp 1698431365
transform -1 0 15792 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2482__A2
timestamp 1698431365
transform 1 0 22400 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2490__I
timestamp 1698431365
transform -1 0 16352 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2491__A1
timestamp 1698431365
transform 1 0 11536 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2493__A1
timestamp 1698431365
transform -1 0 12544 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2495__A1
timestamp 1698431365
transform -1 0 12880 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2503__I
timestamp 1698431365
transform 1 0 30800 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2504__A1
timestamp 1698431365
transform 1 0 12880 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2504__C
timestamp 1698431365
transform -1 0 9184 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2506__A1
timestamp 1698431365
transform 1 0 15120 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2506__C
timestamp 1698431365
transform 1 0 15568 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2508__A1
timestamp 1698431365
transform 1 0 13552 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2508__C
timestamp 1698431365
transform -1 0 13104 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2510__B
timestamp 1698431365
transform 1 0 18032 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2512__B
timestamp 1698431365
transform 1 0 20496 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2514__C
timestamp 1698431365
transform -1 0 20272 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2516__A1
timestamp 1698431365
transform 1 0 36288 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2519__B
timestamp 1698431365
transform 1 0 31360 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2520__A1
timestamp 1698431365
transform 1 0 29568 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2522__A1
timestamp 1698431365
transform 1 0 32032 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2524__A1
timestamp 1698431365
transform 1 0 32368 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2525__C
timestamp 1698431365
transform 1 0 29680 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2526__CLK
timestamp 1698431365
transform 1 0 35504 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2526__D
timestamp 1698431365
transform 1 0 34720 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2531__CLK
timestamp 1698431365
transform 1 0 41776 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2532__CLK
timestamp 1698431365
transform 1 0 44464 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2533__CLK
timestamp 1698431365
transform 1 0 40544 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2534__CLK
timestamp 1698431365
transform 1 0 41216 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2535__CLK
timestamp 1698431365
transform 1 0 43120 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2536__CLK
timestamp 1698431365
transform 1 0 43232 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2537__CLK
timestamp 1698431365
transform 1 0 44240 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2538__CLK
timestamp 1698431365
transform 1 0 40880 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2539__CLK
timestamp 1698431365
transform 1 0 33600 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2540__CLK
timestamp 1698431365
transform -1 0 35840 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2541__CLK
timestamp 1698431365
transform 1 0 19376 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2542__CLK
timestamp 1698431365
transform 1 0 20272 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2543__CLK
timestamp 1698431365
transform 1 0 15344 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2544__CLK
timestamp 1698431365
transform -1 0 14560 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2545__CLK
timestamp 1698431365
transform 1 0 20720 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2548__CLK
timestamp 1698431365
transform 1 0 17360 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2549__CLK
timestamp 1698431365
transform 1 0 18256 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2550__CLK
timestamp 1698431365
transform -1 0 5264 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2551__CLK
timestamp 1698431365
transform 1 0 5040 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2552__CLK
timestamp 1698431365
transform 1 0 5712 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2553__CLK
timestamp 1698431365
transform 1 0 4928 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2554__CLK
timestamp 1698431365
transform 1 0 4928 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2555__CLK
timestamp 1698431365
transform 1 0 5040 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2556__CLK
timestamp 1698431365
transform 1 0 5040 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2557__CLK
timestamp 1698431365
transform 1 0 4816 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2558__CLK
timestamp 1698431365
transform 1 0 7952 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2560__CLK
timestamp 1698431365
transform 1 0 17696 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2561__CLK
timestamp 1698431365
transform 1 0 8960 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2562__CLK
timestamp 1698431365
transform 1 0 8176 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2563__CLK
timestamp 1698431365
transform 1 0 9632 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2564__CLK
timestamp 1698431365
transform 1 0 7840 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2565__CLK
timestamp 1698431365
transform 1 0 8624 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2566__CLK
timestamp 1698431365
transform 1 0 8960 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2567__CLK
timestamp 1698431365
transform 1 0 8400 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2568__CLK
timestamp 1698431365
transform 1 0 8960 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2569__CLK
timestamp 1698431365
transform 1 0 9184 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2570__CLK
timestamp 1698431365
transform 1 0 14560 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2571__CLK
timestamp 1698431365
transform 1 0 16464 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2576__CLK
timestamp 1698431365
transform 1 0 38192 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2578__CLK
timestamp 1698431365
transform 1 0 38528 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2579__CLK
timestamp 1698431365
transform 1 0 41552 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2580__CLK
timestamp 1698431365
transform 1 0 46144 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2581__CLK
timestamp 1698431365
transform 1 0 44240 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2582__CLK
timestamp 1698431365
transform 1 0 44912 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2583__CLK
timestamp 1698431365
transform 1 0 44912 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2584__CLK
timestamp 1698431365
transform 1 0 44912 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2585__CLK
timestamp 1698431365
transform 1 0 44240 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2586__CLK
timestamp 1698431365
transform 1 0 44464 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2592__CLK
timestamp 1698431365
transform 1 0 44912 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2593__CLK
timestamp 1698431365
transform 1 0 43568 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2594__CLK
timestamp 1698431365
transform 1 0 37072 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2595__CLK
timestamp 1698431365
transform 1 0 39648 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2596__CLK
timestamp 1698431365
transform 1 0 36624 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2597__CLK
timestamp 1698431365
transform 1 0 39536 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2598__CLK
timestamp 1698431365
transform 1 0 40992 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2600__CLK
timestamp 1698431365
transform -1 0 36624 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2601__CLK
timestamp 1698431365
transform 1 0 36400 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2602__CLK
timestamp 1698431365
transform 1 0 36624 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2603__CLK
timestamp 1698431365
transform 1 0 28336 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2604__CLK
timestamp 1698431365
transform 1 0 19376 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2608__CLK
timestamp 1698431365
transform 1 0 31360 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2612__CLK
timestamp 1698431365
transform 1 0 44464 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2613__CLK
timestamp 1698431365
transform 1 0 46816 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2614__CLK
timestamp 1698431365
transform 1 0 46704 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2615__CLK
timestamp 1698431365
transform 1 0 43792 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2616__CLK
timestamp 1698431365
transform 1 0 44912 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2617__CLK
timestamp 1698431365
transform 1 0 41888 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2618__CLK
timestamp 1698431365
transform 1 0 40208 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2619__CLK
timestamp 1698431365
transform 1 0 40320 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2620__CLK
timestamp 1698431365
transform 1 0 39088 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2621__CLK
timestamp 1698431365
transform 1 0 34832 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2622__CLK
timestamp 1698431365
transform -1 0 15792 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2623__CLK
timestamp 1698431365
transform 1 0 44912 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2624__CLK
timestamp 1698431365
transform 1 0 43792 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2625__CLK
timestamp 1698431365
transform -1 0 44016 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2626__CLK
timestamp 1698431365
transform 1 0 44016 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2627__CLK
timestamp 1698431365
transform 1 0 41664 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2628__CLK
timestamp 1698431365
transform -1 0 40096 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2629__CLK
timestamp 1698431365
transform -1 0 36400 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2630__CLK
timestamp 1698431365
transform 1 0 38864 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2631__CLK
timestamp 1698431365
transform 1 0 37632 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2632__CLK
timestamp 1698431365
transform 1 0 35504 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2633__CLK
timestamp 1698431365
transform 1 0 11536 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2634__CLK
timestamp 1698431365
transform 1 0 36400 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2635__CLK
timestamp 1698431365
transform 1 0 33152 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2638__CLK
timestamp 1698431365
transform 1 0 25312 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2639__CLK
timestamp 1698431365
transform 1 0 24640 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2640__CLK
timestamp 1698431365
transform 1 0 24528 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2644__CLK
timestamp 1698431365
transform 1 0 12880 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2645__CLK
timestamp 1698431365
transform 1 0 34384 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2647__CLK
timestamp 1698431365
transform 1 0 36512 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2648__CLK
timestamp 1698431365
transform 1 0 40320 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2649__CLK
timestamp 1698431365
transform -1 0 36400 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2650__CLK
timestamp 1698431365
transform 1 0 34720 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2651__CLK
timestamp 1698431365
transform 1 0 39424 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2652__CLK
timestamp 1698431365
transform 1 0 37408 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2653__CLK
timestamp 1698431365
transform 1 0 38080 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2654__CLK
timestamp 1698431365
transform 1 0 39088 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2655__CLK
timestamp 1698431365
transform 1 0 45808 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2656__CLK
timestamp 1698431365
transform 1 0 47488 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2657__CLK
timestamp 1698431365
transform -1 0 33040 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2659__CLK
timestamp 1698431365
transform 1 0 43232 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2660__CLK
timestamp 1698431365
transform -1 0 45136 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2661__CLK
timestamp 1698431365
transform 1 0 44912 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2662__CLK
timestamp 1698431365
transform 1 0 44240 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2663__CLK
timestamp 1698431365
transform 1 0 33264 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2663__D
timestamp 1698431365
transform 1 0 32480 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2664__CLK
timestamp 1698431365
transform 1 0 44688 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2665__CLK
timestamp 1698431365
transform 1 0 38864 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2666__CLK
timestamp 1698431365
transform -1 0 39872 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2668__CLK
timestamp 1698431365
transform 1 0 38640 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2669__CLK
timestamp 1698431365
transform 1 0 40992 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2670__CLK
timestamp 1698431365
transform 1 0 42112 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2671__CLK
timestamp 1698431365
transform 1 0 37632 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2672__CLK
timestamp 1698431365
transform 1 0 44912 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2673__CLK
timestamp 1698431365
transform 1 0 40096 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2674__CLK
timestamp 1698431365
transform 1 0 44016 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2675__CLK
timestamp 1698431365
transform 1 0 43344 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2676__CLK
timestamp 1698431365
transform 1 0 44464 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2678__CLK
timestamp 1698431365
transform 1 0 32480 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2680__CLK
timestamp 1698431365
transform -1 0 31472 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2681__CLK
timestamp 1698431365
transform 1 0 26544 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2682__CLK
timestamp 1698431365
transform 1 0 24640 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2683__CLK
timestamp 1698431365
transform 1 0 25312 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2684__CLK
timestamp 1698431365
transform 1 0 22288 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2685__CLK
timestamp 1698431365
transform -1 0 21616 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2686__CLK
timestamp 1698431365
transform 1 0 22512 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2687__CLK
timestamp 1698431365
transform 1 0 23072 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2688__CLK
timestamp 1698431365
transform 1 0 24864 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2689__CLK
timestamp 1698431365
transform 1 0 23072 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2690__CLK
timestamp 1698431365
transform 1 0 19712 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2691__CLK
timestamp 1698431365
transform 1 0 19712 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2692__CLK
timestamp 1698431365
transform 1 0 18256 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2693__CLK
timestamp 1698431365
transform 1 0 17584 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2694__CLK
timestamp 1698431365
transform 1 0 17024 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2695__CLK
timestamp 1698431365
transform 1 0 18704 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2696__CLK
timestamp 1698431365
transform 1 0 23856 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2697__CLK
timestamp 1698431365
transform 1 0 26208 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2698__CLK
timestamp 1698431365
transform 1 0 24640 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2699__CLK
timestamp 1698431365
transform 1 0 24304 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2700__CLK
timestamp 1698431365
transform 1 0 20272 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2701__CLK
timestamp 1698431365
transform 1 0 23072 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2702__CLK
timestamp 1698431365
transform 1 0 21728 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2703__CLK
timestamp 1698431365
transform 1 0 21392 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2704__CLK
timestamp 1698431365
transform 1 0 6272 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2705__CLK
timestamp 1698431365
transform 1 0 5040 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2706__CLK
timestamp 1698431365
transform 1 0 6272 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2707__CLK
timestamp 1698431365
transform 1 0 8848 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2708__CLK
timestamp 1698431365
transform 1 0 17360 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2709__CLK
timestamp 1698431365
transform 1 0 12320 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2710__CLK
timestamp 1698431365
transform 1 0 16016 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2711__CLK
timestamp 1698431365
transform 1 0 14896 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2712__CLK
timestamp 1698431365
transform 1 0 16800 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2713__CLK
timestamp 1698431365
transform -1 0 17696 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2714__CLK
timestamp 1698431365
transform 1 0 17472 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2715__CLK
timestamp 1698431365
transform 1 0 41104 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2716__CLK
timestamp 1698431365
transform 1 0 27888 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2717__CLK
timestamp 1698431365
transform 1 0 34048 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2718__CLK
timestamp 1698431365
transform 1 0 34048 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_0_wb_clk_i_I
timestamp 1698431365
transform -1 0 24528 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_0_0_wb_clk_i_I
timestamp 1698431365
transform 1 0 24304 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_1_0_wb_clk_i_I
timestamp 1698431365
transform -1 0 27776 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_2_0_wb_clk_i_I
timestamp 1698431365
transform 1 0 21392 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_3_0_wb_clk_i_I
timestamp 1698431365
transform 1 0 26208 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_4_0_wb_clk_i_I
timestamp 1698431365
transform 1 0 36400 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_5_0_wb_clk_i_I
timestamp 1698431365
transform 1 0 40208 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_6_0_wb_clk_i_I
timestamp 1698431365
transform 1 0 34384 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_7_0_wb_clk_i_I
timestamp 1698431365
transform 1 0 39984 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_8_0_wb_clk_i_I
timestamp 1698431365
transform 1 0 19824 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_9_0_wb_clk_i_I
timestamp 1698431365
transform 1 0 20720 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_10_0_wb_clk_i_I
timestamp 1698431365
transform 1 0 21168 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_11_0_wb_clk_i_I
timestamp 1698431365
transform 1 0 25760 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_12_0_wb_clk_i_I
timestamp 1698431365
transform 1 0 32480 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_13_0_wb_clk_i_I
timestamp 1698431365
transform 1 0 39312 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_14_0_wb_clk_i_I
timestamp 1698431365
transform -1 0 36288 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_15_0_wb_clk_i_I
timestamp 1698431365
transform 1 0 40320 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input1_I
timestamp 1698431365
transform -1 0 47488 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input2_I
timestamp 1698431365
transform -1 0 48160 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input3_I
timestamp 1698431365
transform -1 0 48384 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input4_I
timestamp 1698431365
transform -1 0 47712 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input5_I
timestamp 1698431365
transform -1 0 47712 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input6_I
timestamp 1698431365
transform -1 0 46368 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input7_I
timestamp 1698431365
transform -1 0 48384 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input8_I
timestamp 1698431365
transform -1 0 47712 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input9_I
timestamp 1698431365
transform -1 0 48384 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input10_I
timestamp 1698431365
transform -1 0 48384 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input11_I
timestamp 1698431365
transform 1 0 1792 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input12_I
timestamp 1698431365
transform 1 0 1792 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output15_I
timestamp 1698431365
transform -1 0 27552 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output16_I
timestamp 1698431365
transform 1 0 31808 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output21_I
timestamp 1698431365
transform 1 0 40992 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_rebuffer22_I
timestamp 1698431365
transform 1 0 30128 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_wb_clk_i $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 25088 0 -1 31360
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_0_0_wb_clk_i $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 24080 0 1 14112
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_1_0_wb_clk_i
timestamp 1698431365
transform 1 0 24416 0 1 12544
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_2_0_wb_clk_i
timestamp 1698431365
transform 1 0 18032 0 1 18816
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_3_0_wb_clk_i
timestamp 1698431365
transform 1 0 21952 0 1 18816
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_4_0_wb_clk_i
timestamp 1698431365
transform 1 0 36848 0 1 15680
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_5_0_wb_clk_i
timestamp 1698431365
transform 1 0 39760 0 1 15680
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_6_0_wb_clk_i
timestamp 1698431365
transform 1 0 35728 0 -1 20384
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_7_0_wb_clk_i
timestamp 1698431365
transform 1 0 39648 0 1 20384
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_8_0_wb_clk_i
timestamp 1698431365
transform -1 0 18816 0 1 43904
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_9_0_wb_clk_i
timestamp 1698431365
transform 1 0 17248 0 -1 43904
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_10_0_wb_clk_i
timestamp 1698431365
transform -1 0 19488 0 1 45472
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_11_0_wb_clk_i
timestamp 1698431365
transform 1 0 19824 0 -1 47040
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_12_0_wb_clk_i
timestamp 1698431365
transform 1 0 33712 0 1 40768
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_13_0_wb_clk_i
timestamp 1698431365
transform 1 0 38640 0 1 39200
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_14_0_wb_clk_i
timestamp 1698431365
transform 1 0 35616 0 -1 47040
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_15_0_wb_clk_i
timestamp 1698431365
transform 1 0 40096 0 1 45472
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_2 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1568 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_36
timestamp 1698431365
transform 1 0 5376 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_70
timestamp 1698431365
transform 1 0 9184 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_104
timestamp 1698431365
transform 1 0 12992 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_138
timestamp 1698431365
transform 1 0 16800 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_172 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 20608 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_176 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 21056 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_178 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 21280 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_181 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 21616 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_189
timestamp 1698431365
transform 1 0 22512 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_194
timestamp 1698431365
transform 1 0 23072 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_202
timestamp 1698431365
transform 1 0 23968 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_206
timestamp 1698431365
transform 1 0 24416 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_240
timestamp 1698431365
transform 1 0 28224 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_274
timestamp 1698431365
transform 1 0 32032 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_308
timestamp 1698431365
transform 1 0 35840 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_310
timestamp 1698431365
transform 1 0 36064 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_313 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 36400 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_329
timestamp 1698431365
transform 1 0 38192 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_337
timestamp 1698431365
transform 1 0 39088 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_339
timestamp 1698431365
transform 1 0 39312 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_342
timestamp 1698431365
transform 1 0 39648 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_346
timestamp 1698431365
transform 1 0 40096 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_362
timestamp 1698431365
transform 1 0 41888 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_370
timestamp 1698431365
transform 1 0 42784 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_376
timestamp 1698431365
transform 1 0 43456 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_378
timestamp 1698431365
transform 1 0 43680 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_381
timestamp 1698431365
transform 1 0 44016 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_397
timestamp 1698431365
transform 1 0 45808 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_405
timestamp 1698431365
transform 1 0 46704 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_407
timestamp 1698431365
transform 1 0 46928 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_410
timestamp 1698431365
transform 1 0 47264 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_2 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1568 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_66
timestamp 1698431365
transform 1 0 8736 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_72
timestamp 1698431365
transform 1 0 9408 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_136
timestamp 1698431365
transform 1 0 16576 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_142
timestamp 1698431365
transform 1 0 17248 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_208
timestamp 1698431365
transform 1 0 24640 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_212
timestamp 1698431365
transform 1 0 25088 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_216
timestamp 1698431365
transform 1 0 25536 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_228
timestamp 1698431365
transform 1 0 26880 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_230
timestamp 1698431365
transform 1 0 27104 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_260
timestamp 1698431365
transform 1 0 30464 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_268
timestamp 1698431365
transform 1 0 31360 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_276
timestamp 1698431365
transform 1 0 32256 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_340
timestamp 1698431365
transform 1 0 39424 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_342
timestamp 1698431365
transform 1 0 39648 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_349
timestamp 1698431365
transform 1 0 40432 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_410
timestamp 1698431365
transform 1 0 47264 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_2
timestamp 1698431365
transform 1 0 1568 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_34
timestamp 1698431365
transform 1 0 5152 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_37
timestamp 1698431365
transform 1 0 5488 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_101
timestamp 1698431365
transform 1 0 12656 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_107
timestamp 1698431365
transform 1 0 13328 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_139
timestamp 1698431365
transform 1 0 16912 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_143
timestamp 1698431365
transform 1 0 17360 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_145
timestamp 1698431365
transform 1 0 17584 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_185
timestamp 1698431365
transform 1 0 22064 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_189
timestamp 1698431365
transform 1 0 22512 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_193
timestamp 1698431365
transform 1 0 22960 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_243
timestamp 1698431365
transform 1 0 28560 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_251
timestamp 1698431365
transform 1 0 29456 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_282
timestamp 1698431365
transform 1 0 32928 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_290
timestamp 1698431365
transform 1 0 33824 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_298
timestamp 1698431365
transform 1 0 34720 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_302
timestamp 1698431365
transform 1 0 35168 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_317
timestamp 1698431365
transform 1 0 36848 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_358
timestamp 1698431365
transform 1 0 41440 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_362
timestamp 1698431365
transform 1 0 41888 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_366
timestamp 1698431365
transform 1 0 42336 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_368
timestamp 1698431365
transform 1 0 42560 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_373
timestamp 1698431365
transform 1 0 43120 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_383
timestamp 1698431365
transform 1 0 44240 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_387
timestamp 1698431365
transform 1 0 44688 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_419
timestamp 1698431365
transform 1 0 48272 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_2
timestamp 1698431365
transform 1 0 1568 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_66
timestamp 1698431365
transform 1 0 8736 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_72
timestamp 1698431365
transform 1 0 9408 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_136
timestamp 1698431365
transform 1 0 16576 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_3_142
timestamp 1698431365
transform 1 0 17248 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_150
timestamp 1698431365
transform 1 0 18144 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_206
timestamp 1698431365
transform 1 0 24416 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_212
timestamp 1698431365
transform 1 0 25088 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_242
timestamp 1698431365
transform 1 0 28448 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_244
timestamp 1698431365
transform 1 0 28672 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_257
timestamp 1698431365
transform 1 0 30128 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_261
timestamp 1698431365
transform 1 0 30576 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_275
timestamp 1698431365
transform 1 0 32144 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_277
timestamp 1698431365
transform 1 0 32368 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_294
timestamp 1698431365
transform 1 0 34272 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_320
timestamp 1698431365
transform 1 0 37184 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_347
timestamp 1698431365
transform 1 0 40208 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_349
timestamp 1698431365
transform 1 0 40432 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_3_372
timestamp 1698431365
transform 1 0 43008 0 -1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_3_404
timestamp 1698431365
transform 1 0 46592 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_2
timestamp 1698431365
transform 1 0 1568 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_34
timestamp 1698431365
transform 1 0 5152 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_37
timestamp 1698431365
transform 1 0 5488 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_101
timestamp 1698431365
transform 1 0 12656 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_4_107
timestamp 1698431365
transform 1 0 13328 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_123
timestamp 1698431365
transform 1 0 15120 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_131
timestamp 1698431365
transform 1 0 16016 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_162
timestamp 1698431365
transform 1 0 19488 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_166
timestamp 1698431365
transform 1 0 19936 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_168
timestamp 1698431365
transform 1 0 20160 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_171
timestamp 1698431365
transform 1 0 20496 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_177
timestamp 1698431365
transform 1 0 21168 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_181
timestamp 1698431365
transform 1 0 21616 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_223
timestamp 1698431365
transform 1 0 26320 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_227
timestamp 1698431365
transform 1 0 26768 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_263
timestamp 1698431365
transform 1 0 30800 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_286
timestamp 1698431365
transform 1 0 33376 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_310
timestamp 1698431365
transform 1 0 36064 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_312
timestamp 1698431365
transform 1 0 36288 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_317
timestamp 1698431365
transform 1 0 36848 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_319
timestamp 1698431365
transform 1 0 37072 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_336
timestamp 1698431365
transform 1 0 38976 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_356
timestamp 1698431365
transform 1 0 41216 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_377
timestamp 1698431365
transform 1 0 43568 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_416
timestamp 1698431365
transform 1 0 47936 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_2
timestamp 1698431365
transform 1 0 1568 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_66
timestamp 1698431365
transform 1 0 8736 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_5_72
timestamp 1698431365
transform 1 0 9408 0 -1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_5_104
timestamp 1698431365
transform 1 0 12992 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_120
timestamp 1698431365
transform 1 0 14784 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_128
timestamp 1698431365
transform 1 0 15680 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_142
timestamp 1698431365
transform 1 0 17248 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_146
timestamp 1698431365
transform 1 0 17696 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_155
timestamp 1698431365
transform 1 0 18704 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_157
timestamp 1698431365
transform 1 0 18928 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_187
timestamp 1698431365
transform 1 0 22288 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_191
timestamp 1698431365
transform 1 0 22736 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_195
timestamp 1698431365
transform 1 0 23184 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_197
timestamp 1698431365
transform 1 0 23408 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_206
timestamp 1698431365
transform 1 0 24416 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_212
timestamp 1698431365
transform 1 0 25088 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_214
timestamp 1698431365
transform 1 0 25312 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_217
timestamp 1698431365
transform 1 0 25648 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_278
timestamp 1698431365
transform 1 0 32480 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_287
timestamp 1698431365
transform 1 0 33488 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_301
timestamp 1698431365
transform 1 0 35056 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_311
timestamp 1698431365
transform 1 0 36176 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_324
timestamp 1698431365
transform 1 0 37632 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_337
timestamp 1698431365
transform 1 0 39088 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_349
timestamp 1698431365
transform 1 0 40432 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_352
timestamp 1698431365
transform 1 0 40768 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_354
timestamp 1698431365
transform 1 0 40992 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_383
timestamp 1698431365
transform 1 0 44240 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_387
timestamp 1698431365
transform 1 0 44688 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_391
timestamp 1698431365
transform 1 0 45136 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_5_395
timestamp 1698431365
transform 1 0 45584 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_411
timestamp 1698431365
transform 1 0 47376 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_419
timestamp 1698431365
transform 1 0 48272 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_2
timestamp 1698431365
transform 1 0 1568 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_34
timestamp 1698431365
transform 1 0 5152 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_37
timestamp 1698431365
transform 1 0 5488 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_101
timestamp 1698431365
transform 1 0 12656 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_6_107
timestamp 1698431365
transform 1 0 13328 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_152
timestamp 1698431365
transform 1 0 18368 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_162
timestamp 1698431365
transform 1 0 19488 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_166
timestamp 1698431365
transform 1 0 19936 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_174
timestamp 1698431365
transform 1 0 20832 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_6_177
timestamp 1698431365
transform 1 0 21168 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_193
timestamp 1698431365
transform 1 0 22960 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_197
timestamp 1698431365
transform 1 0 23408 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_207
timestamp 1698431365
transform 1 0 24528 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_220
timestamp 1698431365
transform 1 0 25984 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_224
timestamp 1698431365
transform 1 0 26432 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_231
timestamp 1698431365
transform 1 0 27216 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_239
timestamp 1698431365
transform 1 0 28112 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_243
timestamp 1698431365
transform 1 0 28560 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_247
timestamp 1698431365
transform 1 0 29008 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_311
timestamp 1698431365
transform 1 0 36176 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_317
timestamp 1698431365
transform 1 0 36848 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_321
timestamp 1698431365
transform 1 0 37296 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_359
timestamp 1698431365
transform 1 0 41552 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_371
timestamp 1698431365
transform 1 0 42896 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_397
timestamp 1698431365
transform 1 0 45808 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_6_401
timestamp 1698431365
transform 1 0 46256 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_417
timestamp 1698431365
transform 1 0 48048 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_419
timestamp 1698431365
transform 1 0 48272 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_2
timestamp 1698431365
transform 1 0 1568 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_66
timestamp 1698431365
transform 1 0 8736 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_72
timestamp 1698431365
transform 1 0 9408 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_136
timestamp 1698431365
transform 1 0 16576 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_142
timestamp 1698431365
transform 1 0 17248 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_146
timestamp 1698431365
transform 1 0 17696 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_156
timestamp 1698431365
transform 1 0 18816 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_160
timestamp 1698431365
transform 1 0 19264 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_174
timestamp 1698431365
transform 1 0 20832 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_183
timestamp 1698431365
transform 1 0 21840 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_205
timestamp 1698431365
transform 1 0 24304 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_209
timestamp 1698431365
transform 1 0 24752 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_212
timestamp 1698431365
transform 1 0 25088 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_216
timestamp 1698431365
transform 1 0 25536 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_220
timestamp 1698431365
transform 1 0 25984 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_224
timestamp 1698431365
transform 1 0 26432 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_254
timestamp 1698431365
transform 1 0 29792 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_270
timestamp 1698431365
transform 1 0 31584 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_278
timestamp 1698431365
transform 1 0 32480 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_295
timestamp 1698431365
transform 1 0 34384 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_299
timestamp 1698431365
transform 1 0 34832 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_303
timestamp 1698431365
transform 1 0 35280 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_311
timestamp 1698431365
transform 1 0 36176 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_319
timestamp 1698431365
transform 1 0 37072 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_328
timestamp 1698431365
transform 1 0 38080 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_338
timestamp 1698431365
transform 1 0 39200 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_342
timestamp 1698431365
transform 1 0 39648 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_381
timestamp 1698431365
transform 1 0 44016 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_383
timestamp 1698431365
transform 1 0 44240 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_413
timestamp 1698431365
transform 1 0 47600 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_417
timestamp 1698431365
transform 1 0 48048 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_419
timestamp 1698431365
transform 1 0 48272 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_2
timestamp 1698431365
transform 1 0 1568 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_34
timestamp 1698431365
transform 1 0 5152 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_37
timestamp 1698431365
transform 1 0 5488 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_101
timestamp 1698431365
transform 1 0 12656 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_107
timestamp 1698431365
transform 1 0 13328 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_115
timestamp 1698431365
transform 1 0 14224 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_119
timestamp 1698431365
transform 1 0 14672 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_149
timestamp 1698431365
transform 1 0 18032 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_8_153
timestamp 1698431365
transform 1 0 18480 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_169
timestamp 1698431365
transform 1 0 20272 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_173
timestamp 1698431365
transform 1 0 20720 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_218
timestamp 1698431365
transform 1 0 25760 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_222
timestamp 1698431365
transform 1 0 26208 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_230
timestamp 1698431365
transform 1 0 27104 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_234
timestamp 1698431365
transform 1 0 27552 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_242
timestamp 1698431365
transform 1 0 28448 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_247
timestamp 1698431365
transform 1 0 29008 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_249
timestamp 1698431365
transform 1 0 29232 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_8_279
timestamp 1698431365
transform 1 0 32592 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_295
timestamp 1698431365
transform 1 0 34384 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_307
timestamp 1698431365
transform 1 0 35728 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_311
timestamp 1698431365
transform 1 0 36176 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_317
timestamp 1698431365
transform 1 0 36848 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_348
timestamp 1698431365
transform 1 0 40320 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_354
timestamp 1698431365
transform 1 0 40992 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_358
timestamp 1698431365
transform 1 0 41440 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_360
timestamp 1698431365
transform 1 0 41664 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_371
timestamp 1698431365
transform 1 0 42896 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_395
timestamp 1698431365
transform 1 0 45584 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_399
timestamp 1698431365
transform 1 0 46032 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_407
timestamp 1698431365
transform 1 0 46928 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_411
timestamp 1698431365
transform 1 0 47376 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_2
timestamp 1698431365
transform 1 0 1568 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_66
timestamp 1698431365
transform 1 0 8736 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_9_72
timestamp 1698431365
transform 1 0 9408 0 -1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_9_104
timestamp 1698431365
transform 1 0 12992 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_120
timestamp 1698431365
transform 1 0 14784 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_128
timestamp 1698431365
transform 1 0 15680 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_142
timestamp 1698431365
transform 1 0 17248 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_144
timestamp 1698431365
transform 1 0 17472 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_155
timestamp 1698431365
transform 1 0 18704 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_157
timestamp 1698431365
transform 1 0 18928 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_187
timestamp 1698431365
transform 1 0 22288 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_192
timestamp 1698431365
transform 1 0 22848 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_196
timestamp 1698431365
transform 1 0 23296 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_208
timestamp 1698431365
transform 1 0 24640 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_217
timestamp 1698431365
transform 1 0 25648 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_271
timestamp 1698431365
transform 1 0 31696 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_275
timestamp 1698431365
transform 1 0 32144 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_279
timestamp 1698431365
transform 1 0 32592 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_282
timestamp 1698431365
transform 1 0 32928 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_289
timestamp 1698431365
transform 1 0 33712 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_293
timestamp 1698431365
transform 1 0 34160 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_329
timestamp 1698431365
transform 1 0 38192 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_333
timestamp 1698431365
transform 1 0 38640 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_337
timestamp 1698431365
transform 1 0 39088 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_349
timestamp 1698431365
transform 1 0 40432 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_360
timestamp 1698431365
transform 1 0 41664 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_9_395
timestamp 1698431365
transform 1 0 45584 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_415
timestamp 1698431365
transform 1 0 47824 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_419
timestamp 1698431365
transform 1 0 48272 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_2
timestamp 1698431365
transform 1 0 1568 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_34
timestamp 1698431365
transform 1 0 5152 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_37
timestamp 1698431365
transform 1 0 5488 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_101
timestamp 1698431365
transform 1 0 12656 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_107
timestamp 1698431365
transform 1 0 13328 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_115
timestamp 1698431365
transform 1 0 14224 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_174
timestamp 1698431365
transform 1 0 20832 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_185
timestamp 1698431365
transform 1 0 22064 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_189
timestamp 1698431365
transform 1 0 22512 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_191
timestamp 1698431365
transform 1 0 22736 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_208
timestamp 1698431365
transform 1 0 24640 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_212
timestamp 1698431365
transform 1 0 25088 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_224
timestamp 1698431365
transform 1 0 26432 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_228
timestamp 1698431365
transform 1 0 26880 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_232
timestamp 1698431365
transform 1 0 27328 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_234
timestamp 1698431365
transform 1 0 27552 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_255
timestamp 1698431365
transform 1 0 29904 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_259
timestamp 1698431365
transform 1 0 30352 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_268
timestamp 1698431365
transform 1 0 31360 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_276
timestamp 1698431365
transform 1 0 32256 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_313
timestamp 1698431365
transform 1 0 36400 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_321
timestamp 1698431365
transform 1 0 37296 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_323
timestamp 1698431365
transform 1 0 37520 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_326
timestamp 1698431365
transform 1 0 37856 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_330
timestamp 1698431365
transform 1 0 38304 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_347
timestamp 1698431365
transform 1 0 40208 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_349
timestamp 1698431365
transform 1 0 40432 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_352
timestamp 1698431365
transform 1 0 40768 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_362
timestamp 1698431365
transform 1 0 41888 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_382
timestamp 1698431365
transform 1 0 44128 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_384
timestamp 1698431365
transform 1 0 44352 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_391
timestamp 1698431365
transform 1 0 45136 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_407
timestamp 1698431365
transform 1 0 46928 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_415
timestamp 1698431365
transform 1 0 47824 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_419
timestamp 1698431365
transform 1 0 48272 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_2
timestamp 1698431365
transform 1 0 1568 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_66
timestamp 1698431365
transform 1 0 8736 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_11_72
timestamp 1698431365
transform 1 0 9408 0 -1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_104
timestamp 1698431365
transform 1 0 12992 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_120
timestamp 1698431365
transform 1 0 14784 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_128
timestamp 1698431365
transform 1 0 15680 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_142
timestamp 1698431365
transform 1 0 17248 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_160
timestamp 1698431365
transform 1 0 19264 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_166
timestamp 1698431365
transform 1 0 19936 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_173
timestamp 1698431365
transform 1 0 20720 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_232
timestamp 1698431365
transform 1 0 27328 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_234
timestamp 1698431365
transform 1 0 27552 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_247
timestamp 1698431365
transform 1 0 29008 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_251
timestamp 1698431365
transform 1 0 29456 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_273
timestamp 1698431365
transform 1 0 31920 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_277
timestamp 1698431365
transform 1 0 32368 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_279
timestamp 1698431365
transform 1 0 32592 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_282
timestamp 1698431365
transform 1 0 32928 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_286
timestamp 1698431365
transform 1 0 33376 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_288
timestamp 1698431365
transform 1 0 33600 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_348
timestamp 1698431365
transform 1 0 40320 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_381
timestamp 1698431365
transform 1 0 44016 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_11_387
timestamp 1698431365
transform 1 0 44688 0 -1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_419
timestamp 1698431365
transform 1 0 48272 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_2
timestamp 1698431365
transform 1 0 1568 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_34
timestamp 1698431365
transform 1 0 5152 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_37
timestamp 1698431365
transform 1 0 5488 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_101
timestamp 1698431365
transform 1 0 12656 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_107
timestamp 1698431365
transform 1 0 13328 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_139
timestamp 1698431365
transform 1 0 16912 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_142
timestamp 1698431365
transform 1 0 17248 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_152
timestamp 1698431365
transform 1 0 18368 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_159
timestamp 1698431365
transform 1 0 19152 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_232
timestamp 1698431365
transform 1 0 27328 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_236
timestamp 1698431365
transform 1 0 27776 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_244
timestamp 1698431365
transform 1 0 28672 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_247
timestamp 1698431365
transform 1 0 29008 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_277
timestamp 1698431365
transform 1 0 32368 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_285
timestamp 1698431365
transform 1 0 33264 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_289
timestamp 1698431365
transform 1 0 33712 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_299
timestamp 1698431365
transform 1 0 34832 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_303
timestamp 1698431365
transform 1 0 35280 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_311
timestamp 1698431365
transform 1 0 36176 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_317
timestamp 1698431365
transform 1 0 36848 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_349
timestamp 1698431365
transform 1 0 40432 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_357
timestamp 1698431365
transform 1 0 41328 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_361
timestamp 1698431365
transform 1 0 41776 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_364
timestamp 1698431365
transform 1 0 42112 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_368
timestamp 1698431365
transform 1 0 42560 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_376
timestamp 1698431365
transform 1 0 43456 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_384
timestamp 1698431365
transform 1 0 44352 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_416
timestamp 1698431365
transform 1 0 47936 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_2
timestamp 1698431365
transform 1 0 1568 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_66
timestamp 1698431365
transform 1 0 8736 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_13_72
timestamp 1698431365
transform 1 0 9408 0 -1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_104
timestamp 1698431365
transform 1 0 12992 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_108
timestamp 1698431365
transform 1 0 13440 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_110
timestamp 1698431365
transform 1 0 13664 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_142
timestamp 1698431365
transform 1 0 17248 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_144
timestamp 1698431365
transform 1 0 17472 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_153
timestamp 1698431365
transform 1 0 18480 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_194
timestamp 1698431365
transform 1 0 23072 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_196
timestamp 1698431365
transform 1 0 23296 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_207
timestamp 1698431365
transform 1 0 24528 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_209
timestamp 1698431365
transform 1 0 24752 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_224
timestamp 1698431365
transform 1 0 26432 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_241
timestamp 1698431365
transform 1 0 28336 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_249
timestamp 1698431365
transform 1 0 29232 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_261
timestamp 1698431365
transform 1 0 30576 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_265
timestamp 1698431365
transform 1 0 31024 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_282
timestamp 1698431365
transform 1 0 32928 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_284
timestamp 1698431365
transform 1 0 33152 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_309
timestamp 1698431365
transform 1 0 35952 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_313
timestamp 1698431365
transform 1 0 36400 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_317
timestamp 1698431365
transform 1 0 36848 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_320
timestamp 1698431365
transform 1 0 37184 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_340
timestamp 1698431365
transform 1 0 39424 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_348
timestamp 1698431365
transform 1 0 40320 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_352
timestamp 1698431365
transform 1 0 40768 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_360
timestamp 1698431365
transform 1 0 41664 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_364
timestamp 1698431365
transform 1 0 42112 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_369
timestamp 1698431365
transform 1 0 42672 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_373
timestamp 1698431365
transform 1 0 43120 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_377
timestamp 1698431365
transform 1 0 43568 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_381
timestamp 1698431365
transform 1 0 44016 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_398
timestamp 1698431365
transform 1 0 45920 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_402
timestamp 1698431365
transform 1 0 46368 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_418
timestamp 1698431365
transform 1 0 48160 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_2
timestamp 1698431365
transform 1 0 1568 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_34
timestamp 1698431365
transform 1 0 5152 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_37
timestamp 1698431365
transform 1 0 5488 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_101
timestamp 1698431365
transform 1 0 12656 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_107
timestamp 1698431365
transform 1 0 13328 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_152
timestamp 1698431365
transform 1 0 18368 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_154
timestamp 1698431365
transform 1 0 18592 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_165
timestamp 1698431365
transform 1 0 19824 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_203
timestamp 1698431365
transform 1 0 24080 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_207
timestamp 1698431365
transform 1 0 24528 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_247
timestamp 1698431365
transform 1 0 29008 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_249
timestamp 1698431365
transform 1 0 29232 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_258
timestamp 1698431365
transform 1 0 30240 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_262
timestamp 1698431365
transform 1 0 30688 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_266
timestamp 1698431365
transform 1 0 31136 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_303
timestamp 1698431365
transform 1 0 35280 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_307
timestamp 1698431365
transform 1 0 35728 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_311
timestamp 1698431365
transform 1 0 36176 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_317
timestamp 1698431365
transform 1 0 36848 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_319
timestamp 1698431365
transform 1 0 37072 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_326
timestamp 1698431365
transform 1 0 37856 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_387
timestamp 1698431365
transform 1 0 44688 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_391
timestamp 1698431365
transform 1 0 45136 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_407
timestamp 1698431365
transform 1 0 46928 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_415
timestamp 1698431365
transform 1 0 47824 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_419
timestamp 1698431365
transform 1 0 48272 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_2
timestamp 1698431365
transform 1 0 1568 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_66
timestamp 1698431365
transform 1 0 8736 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_15_72
timestamp 1698431365
transform 1 0 9408 0 -1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_104
timestamp 1698431365
transform 1 0 12992 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_120
timestamp 1698431365
transform 1 0 14784 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_128
timestamp 1698431365
transform 1 0 15680 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_142
timestamp 1698431365
transform 1 0 17248 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_146
timestamp 1698431365
transform 1 0 17696 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_155
timestamp 1698431365
transform 1 0 18704 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_194
timestamp 1698431365
transform 1 0 23072 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_196
timestamp 1698431365
transform 1 0 23296 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_235
timestamp 1698431365
transform 1 0 27664 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_239
timestamp 1698431365
transform 1 0 28112 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_247
timestamp 1698431365
transform 1 0 29008 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_259
timestamp 1698431365
transform 1 0 30352 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_277
timestamp 1698431365
transform 1 0 32368 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_279
timestamp 1698431365
transform 1 0 32592 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_288
timestamp 1698431365
transform 1 0 33600 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_292
timestamp 1698431365
transform 1 0 34048 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_345
timestamp 1698431365
transform 1 0 39984 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_349
timestamp 1698431365
transform 1 0 40432 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_352
timestamp 1698431365
transform 1 0 40768 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_409
timestamp 1698431365
transform 1 0 47152 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_417
timestamp 1698431365
transform 1 0 48048 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_419
timestamp 1698431365
transform 1 0 48272 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_2
timestamp 1698431365
transform 1 0 1568 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_34
timestamp 1698431365
transform 1 0 5152 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_37
timestamp 1698431365
transform 1 0 5488 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_101
timestamp 1698431365
transform 1 0 12656 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_107
timestamp 1698431365
transform 1 0 13328 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_115
timestamp 1698431365
transform 1 0 14224 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_119
timestamp 1698431365
transform 1 0 14672 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_123
timestamp 1698431365
transform 1 0 15120 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_131
timestamp 1698431365
transform 1 0 16016 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_134
timestamp 1698431365
transform 1 0 16352 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_148
timestamp 1698431365
transform 1 0 17920 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_152
timestamp 1698431365
transform 1 0 18368 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_161
timestamp 1698431365
transform 1 0 19376 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_167
timestamp 1698431365
transform 1 0 20048 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_191
timestamp 1698431365
transform 1 0 22736 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_193
timestamp 1698431365
transform 1 0 22960 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_196
timestamp 1698431365
transform 1 0 23296 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_226
timestamp 1698431365
transform 1 0 26656 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_242
timestamp 1698431365
transform 1 0 28448 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_244
timestamp 1698431365
transform 1 0 28672 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_247
timestamp 1698431365
transform 1 0 29008 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_278
timestamp 1698431365
transform 1 0 32480 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_282
timestamp 1698431365
transform 1 0 32928 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_284
timestamp 1698431365
transform 1 0 33152 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_299
timestamp 1698431365
transform 1 0 34832 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_301
timestamp 1698431365
transform 1 0 35056 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_381
timestamp 1698431365
transform 1 0 44016 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_403
timestamp 1698431365
transform 1 0 46480 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_407
timestamp 1698431365
transform 1 0 46928 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_411
timestamp 1698431365
transform 1 0 47376 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_2
timestamp 1698431365
transform 1 0 1568 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_66
timestamp 1698431365
transform 1 0 8736 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_72
timestamp 1698431365
transform 1 0 9408 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_88
timestamp 1698431365
transform 1 0 11200 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_90
timestamp 1698431365
transform 1 0 11424 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_93
timestamp 1698431365
transform 1 0 11760 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_97
timestamp 1698431365
transform 1 0 12208 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_103
timestamp 1698431365
transform 1 0 12880 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_107
timestamp 1698431365
transform 1 0 13328 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_142
timestamp 1698431365
transform 1 0 17248 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_146
timestamp 1698431365
transform 1 0 17696 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_148
timestamp 1698431365
transform 1 0 17920 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_151
timestamp 1698431365
transform 1 0 18256 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_194
timestamp 1698431365
transform 1 0 23072 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_212
timestamp 1698431365
transform 1 0 25088 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_216
timestamp 1698431365
transform 1 0 25536 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_259
timestamp 1698431365
transform 1 0 30352 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_265
timestamp 1698431365
transform 1 0 31024 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_269
timestamp 1698431365
transform 1 0 31472 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_273
timestamp 1698431365
transform 1 0 31920 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_277
timestamp 1698431365
transform 1 0 32368 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_279
timestamp 1698431365
transform 1 0 32592 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_282
timestamp 1698431365
transform 1 0 32928 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_290
timestamp 1698431365
transform 1 0 33824 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_302
timestamp 1698431365
transform 1 0 35168 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_306
timestamp 1698431365
transform 1 0 35616 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_308
timestamp 1698431365
transform 1 0 35840 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_345
timestamp 1698431365
transform 1 0 39984 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_349
timestamp 1698431365
transform 1 0 40432 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_400
timestamp 1698431365
transform 1 0 46144 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_413
timestamp 1698431365
transform 1 0 47600 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_417
timestamp 1698431365
transform 1 0 48048 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_419
timestamp 1698431365
transform 1 0 48272 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_2
timestamp 1698431365
transform 1 0 1568 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_34
timestamp 1698431365
transform 1 0 5152 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_37
timestamp 1698431365
transform 1 0 5488 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_69
timestamp 1698431365
transform 1 0 9072 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_71
timestamp 1698431365
transform 1 0 9296 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_80
timestamp 1698431365
transform 1 0 10304 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_89
timestamp 1698431365
transform 1 0 11312 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_93
timestamp 1698431365
transform 1 0 11760 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_97
timestamp 1698431365
transform 1 0 12208 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_100
timestamp 1698431365
transform 1 0 12544 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_102
timestamp 1698431365
transform 1 0 12768 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_107
timestamp 1698431365
transform 1 0 13328 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_111
timestamp 1698431365
transform 1 0 13776 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_141
timestamp 1698431365
transform 1 0 17136 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_145
timestamp 1698431365
transform 1 0 17584 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_157
timestamp 1698431365
transform 1 0 18928 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_161
timestamp 1698431365
transform 1 0 19376 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_165
timestamp 1698431365
transform 1 0 19824 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_169
timestamp 1698431365
transform 1 0 20272 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_173
timestamp 1698431365
transform 1 0 20720 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_177
timestamp 1698431365
transform 1 0 21168 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_216
timestamp 1698431365
transform 1 0 25536 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_218
timestamp 1698431365
transform 1 0 25760 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_233
timestamp 1698431365
transform 1 0 27440 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_271
timestamp 1698431365
transform 1 0 31696 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_279
timestamp 1698431365
transform 1 0 32592 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_289
timestamp 1698431365
transform 1 0 33712 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_314
timestamp 1698431365
transform 1 0 36512 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_317
timestamp 1698431365
transform 1 0 36848 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_323
timestamp 1698431365
transform 1 0 37520 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_2
timestamp 1698431365
transform 1 0 1568 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_66
timestamp 1698431365
transform 1 0 8736 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_69
timestamp 1698431365
transform 1 0 9072 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_72
timestamp 1698431365
transform 1 0 9408 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_76
timestamp 1698431365
transform 1 0 9856 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_87
timestamp 1698431365
transform 1 0 11088 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_89
timestamp 1698431365
transform 1 0 11312 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_121
timestamp 1698431365
transform 1 0 14896 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_125
timestamp 1698431365
transform 1 0 15344 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_129
timestamp 1698431365
transform 1 0 15792 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_131
timestamp 1698431365
transform 1 0 16016 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_142
timestamp 1698431365
transform 1 0 17248 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_205
timestamp 1698431365
transform 1 0 24304 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_207
timestamp 1698431365
transform 1 0 24528 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_241
timestamp 1698431365
transform 1 0 28336 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_251
timestamp 1698431365
transform 1 0 29456 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_255
timestamp 1698431365
transform 1 0 29904 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_271
timestamp 1698431365
transform 1 0 31696 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_290
timestamp 1698431365
transform 1 0 33824 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_294
timestamp 1698431365
transform 1 0 34272 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_338
timestamp 1698431365
transform 1 0 39200 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_342
timestamp 1698431365
transform 1 0 39648 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_360
timestamp 1698431365
transform 1 0 41664 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_362
timestamp 1698431365
transform 1 0 41888 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_2
timestamp 1698431365
transform 1 0 1568 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_34
timestamp 1698431365
transform 1 0 5152 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_37
timestamp 1698431365
transform 1 0 5488 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_101
timestamp 1698431365
transform 1 0 12656 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_120
timestamp 1698431365
transform 1 0 14784 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_122
timestamp 1698431365
transform 1 0 15008 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_125
timestamp 1698431365
transform 1 0 15344 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_129
timestamp 1698431365
transform 1 0 15792 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_177
timestamp 1698431365
transform 1 0 21168 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_210
timestamp 1698431365
transform 1 0 24864 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_220
timestamp 1698431365
transform 1 0 25984 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_224
timestamp 1698431365
transform 1 0 26432 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_232
timestamp 1698431365
transform 1 0 27328 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_234
timestamp 1698431365
transform 1 0 27552 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_289
timestamp 1698431365
transform 1 0 33712 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_291
timestamp 1698431365
transform 1 0 33936 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_299
timestamp 1698431365
transform 1 0 34832 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_331
timestamp 1698431365
transform 1 0 38416 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_335
timestamp 1698431365
transform 1 0 38864 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_368
timestamp 1698431365
transform 1 0 42560 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_372
timestamp 1698431365
transform 1 0 43008 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_382
timestamp 1698431365
transform 1 0 44128 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_384
timestamp 1698431365
transform 1 0 44352 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_404
timestamp 1698431365
transform 1 0 46592 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_408
timestamp 1698431365
transform 1 0 47040 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_416
timestamp 1698431365
transform 1 0 47936 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_2
timestamp 1698431365
transform 1 0 1568 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_18
timestamp 1698431365
transform 1 0 3360 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_26
timestamp 1698431365
transform 1 0 4256 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_67
timestamp 1698431365
transform 1 0 8848 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_69
timestamp 1698431365
transform 1 0 9072 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_72
timestamp 1698431365
transform 1 0 9408 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_131
timestamp 1698431365
transform 1 0 16016 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_133
timestamp 1698431365
transform 1 0 16240 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_152
timestamp 1698431365
transform 1 0 18368 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_161
timestamp 1698431365
transform 1 0 19376 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_175
timestamp 1698431365
transform 1 0 20944 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_193
timestamp 1698431365
transform 1 0 22960 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_203
timestamp 1698431365
transform 1 0 24080 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_207
timestamp 1698431365
transform 1 0 24528 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_212
timestamp 1698431365
transform 1 0 25088 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_214
timestamp 1698431365
transform 1 0 25312 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_217
timestamp 1698431365
transform 1 0 25648 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_272
timestamp 1698431365
transform 1 0 31808 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_276
timestamp 1698431365
transform 1 0 32256 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_282
timestamp 1698431365
transform 1 0 32928 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_286
timestamp 1698431365
transform 1 0 33376 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_293
timestamp 1698431365
transform 1 0 34160 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_303
timestamp 1698431365
transform 1 0 35280 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_339
timestamp 1698431365
transform 1 0 39312 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_343
timestamp 1698431365
transform 1 0 39760 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_347
timestamp 1698431365
transform 1 0 40208 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_349
timestamp 1698431365
transform 1 0 40432 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_368
timestamp 1698431365
transform 1 0 42560 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_372
timestamp 1698431365
transform 1 0 43008 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_376
timestamp 1698431365
transform 1 0 43456 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_393
timestamp 1698431365
transform 1 0 45360 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_397
timestamp 1698431365
transform 1 0 45808 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_401
timestamp 1698431365
transform 1 0 46256 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_409
timestamp 1698431365
transform 1 0 47152 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_417
timestamp 1698431365
transform 1 0 48048 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_419
timestamp 1698431365
transform 1 0 48272 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_2
timestamp 1698431365
transform 1 0 1568 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_18
timestamp 1698431365
transform 1 0 3360 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_22
timestamp 1698431365
transform 1 0 3808 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_24
timestamp 1698431365
transform 1 0 4032 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_37
timestamp 1698431365
transform 1 0 5488 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_41
timestamp 1698431365
transform 1 0 5936 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_43
timestamp 1698431365
transform 1 0 6160 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_142
timestamp 1698431365
transform 1 0 17248 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_144
timestamp 1698431365
transform 1 0 17472 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_182
timestamp 1698431365
transform 1 0 21728 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_192
timestamp 1698431365
transform 1 0 22848 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_208
timestamp 1698431365
transform 1 0 24640 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_215
timestamp 1698431365
transform 1 0 25424 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_235
timestamp 1698431365
transform 1 0 27664 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_239
timestamp 1698431365
transform 1 0 28112 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_243
timestamp 1698431365
transform 1 0 28560 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_247
timestamp 1698431365
transform 1 0 29008 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_251
timestamp 1698431365
transform 1 0 29456 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_253
timestamp 1698431365
transform 1 0 29680 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_256
timestamp 1698431365
transform 1 0 30016 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_264
timestamp 1698431365
transform 1 0 30912 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_297
timestamp 1698431365
transform 1 0 34608 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_301
timestamp 1698431365
transform 1 0 35056 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_313
timestamp 1698431365
transform 1 0 36400 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_321
timestamp 1698431365
transform 1 0 37296 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_325
timestamp 1698431365
transform 1 0 37744 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_327
timestamp 1698431365
transform 1 0 37968 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_378
timestamp 1698431365
transform 1 0 43680 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_382
timestamp 1698431365
transform 1 0 44128 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_384
timestamp 1698431365
transform 1 0 44352 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_387
timestamp 1698431365
transform 1 0 44688 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_2
timestamp 1698431365
transform 1 0 1568 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_18
timestamp 1698431365
transform 1 0 3360 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_26
timestamp 1698431365
transform 1 0 4256 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_28
timestamp 1698431365
transform 1 0 4480 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_65
timestamp 1698431365
transform 1 0 8624 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_67
timestamp 1698431365
transform 1 0 8848 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_78
timestamp 1698431365
transform 1 0 10080 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_105
timestamp 1698431365
transform 1 0 13104 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_142
timestamp 1698431365
transform 1 0 17248 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_162
timestamp 1698431365
transform 1 0 19488 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_184
timestamp 1698431365
transform 1 0 21952 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_188
timestamp 1698431365
transform 1 0 22400 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_195
timestamp 1698431365
transform 1 0 23184 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_220
timestamp 1698431365
transform 1 0 25984 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_242
timestamp 1698431365
transform 1 0 28448 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_246
timestamp 1698431365
transform 1 0 28896 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_250
timestamp 1698431365
transform 1 0 29344 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_254
timestamp 1698431365
transform 1 0 29792 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_262
timestamp 1698431365
transform 1 0 30688 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_272
timestamp 1698431365
transform 1 0 31808 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_279
timestamp 1698431365
transform 1 0 32592 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_282
timestamp 1698431365
transform 1 0 32928 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_298
timestamp 1698431365
transform 1 0 34720 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_300
timestamp 1698431365
transform 1 0 34944 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_346
timestamp 1698431365
transform 1 0 40096 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_389
timestamp 1698431365
transform 1 0 44912 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_397
timestamp 1698431365
transform 1 0 45808 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_399
timestamp 1698431365
transform 1 0 46032 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_412
timestamp 1698431365
transform 1 0 47488 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_2
timestamp 1698431365
transform 1 0 1568 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_18
timestamp 1698431365
transform 1 0 3360 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_26
timestamp 1698431365
transform 1 0 4256 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_28
timestamp 1698431365
transform 1 0 4480 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_37
timestamp 1698431365
transform 1 0 5488 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_96
timestamp 1698431365
transform 1 0 12096 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_161
timestamp 1698431365
transform 1 0 19376 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_173
timestamp 1698431365
transform 1 0 20720 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_177
timestamp 1698431365
transform 1 0 21168 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_181
timestamp 1698431365
transform 1 0 21616 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_183
timestamp 1698431365
transform 1 0 21840 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_186
timestamp 1698431365
transform 1 0 22176 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_190
timestamp 1698431365
transform 1 0 22624 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_220
timestamp 1698431365
transform 1 0 25984 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_224
timestamp 1698431365
transform 1 0 26432 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_247
timestamp 1698431365
transform 1 0 29008 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_257
timestamp 1698431365
transform 1 0 30128 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_266
timestamp 1698431365
transform 1 0 31136 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_284
timestamp 1698431365
transform 1 0 33152 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_310
timestamp 1698431365
transform 1 0 36064 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_314
timestamp 1698431365
transform 1 0 36512 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_317
timestamp 1698431365
transform 1 0 36848 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_321
timestamp 1698431365
transform 1 0 37296 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_351
timestamp 1698431365
transform 1 0 40656 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_355
timestamp 1698431365
transform 1 0 41104 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_357
timestamp 1698431365
transform 1 0 41328 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_371
timestamp 1698431365
transform 1 0 42896 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_379
timestamp 1698431365
transform 1 0 43792 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_383
timestamp 1698431365
transform 1 0 44240 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_387
timestamp 1698431365
transform 1 0 44688 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_2
timestamp 1698431365
transform 1 0 1568 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_69
timestamp 1698431365
transform 1 0 9072 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_72
timestamp 1698431365
transform 1 0 9408 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_137
timestamp 1698431365
transform 1 0 16688 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_139
timestamp 1698431365
transform 1 0 16912 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_142
timestamp 1698431365
transform 1 0 17248 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_154
timestamp 1698431365
transform 1 0 18592 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_156
timestamp 1698431365
transform 1 0 18816 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_167
timestamp 1698431365
transform 1 0 20048 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_171
timestamp 1698431365
transform 1 0 20496 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_175
timestamp 1698431365
transform 1 0 20944 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_188
timestamp 1698431365
transform 1 0 22400 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_192
timestamp 1698431365
transform 1 0 22848 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_198
timestamp 1698431365
transform 1 0 23520 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_200
timestamp 1698431365
transform 1 0 23744 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_203
timestamp 1698431365
transform 1 0 24080 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_207
timestamp 1698431365
transform 1 0 24528 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_209
timestamp 1698431365
transform 1 0 24752 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_212
timestamp 1698431365
transform 1 0 25088 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_216
timestamp 1698431365
transform 1 0 25536 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_232
timestamp 1698431365
transform 1 0 27328 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_236
timestamp 1698431365
transform 1 0 27776 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_268
timestamp 1698431365
transform 1 0 31360 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_272
timestamp 1698431365
transform 1 0 31808 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_282
timestamp 1698431365
transform 1 0 32928 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_314
timestamp 1698431365
transform 1 0 36512 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_317
timestamp 1698431365
transform 1 0 36848 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_333
timestamp 1698431365
transform 1 0 38640 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_335
timestamp 1698431365
transform 1 0 38864 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_338
timestamp 1698431365
transform 1 0 39200 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_342
timestamp 1698431365
transform 1 0 39648 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_346
timestamp 1698431365
transform 1 0 40096 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_381
timestamp 1698431365
transform 1 0 44016 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_419
timestamp 1698431365
transform 1 0 48272 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_2
timestamp 1698431365
transform 1 0 1568 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_18
timestamp 1698431365
transform 1 0 3360 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_26
timestamp 1698431365
transform 1 0 4256 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_30
timestamp 1698431365
transform 1 0 4704 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_32
timestamp 1698431365
transform 1 0 4928 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_37
timestamp 1698431365
transform 1 0 5488 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_39
timestamp 1698431365
transform 1 0 5712 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_58
timestamp 1698431365
transform 1 0 7840 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_127
timestamp 1698431365
transform 1 0 15568 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_164
timestamp 1698431365
transform 1 0 19712 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_171
timestamp 1698431365
transform 1 0 20496 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_183
timestamp 1698431365
transform 1 0 21840 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_244
timestamp 1698431365
transform 1 0 28672 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_251
timestamp 1698431365
transform 1 0 29456 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_261
timestamp 1698431365
transform 1 0 30576 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_265
timestamp 1698431365
transform 1 0 31024 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_272
timestamp 1698431365
transform 1 0 31808 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_276
timestamp 1698431365
transform 1 0 32256 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_284
timestamp 1698431365
transform 1 0 33152 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_288
timestamp 1698431365
transform 1 0 33600 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_290
timestamp 1698431365
transform 1 0 33824 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_303
timestamp 1698431365
transform 1 0 35280 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_317
timestamp 1698431365
transform 1 0 36848 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_321
timestamp 1698431365
transform 1 0 37296 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_323
timestamp 1698431365
transform 1 0 37520 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_353
timestamp 1698431365
transform 1 0 40880 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_357
timestamp 1698431365
transform 1 0 41328 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_373
timestamp 1698431365
transform 1 0 43120 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_381
timestamp 1698431365
transform 1 0 44016 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_416
timestamp 1698431365
transform 1 0 47936 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_2
timestamp 1698431365
transform 1 0 1568 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_10
timestamp 1698431365
transform 1 0 2464 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_14
timestamp 1698431365
transform 1 0 2912 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_134
timestamp 1698431365
transform 1 0 16352 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_142
timestamp 1698431365
transform 1 0 17248 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_144
timestamp 1698431365
transform 1 0 17472 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_155
timestamp 1698431365
transform 1 0 18704 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_174
timestamp 1698431365
transform 1 0 20832 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_250
timestamp 1698431365
transform 1 0 29344 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_256
timestamp 1698431365
transform 1 0 30016 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_258
timestamp 1698431365
transform 1 0 30240 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_275
timestamp 1698431365
transform 1 0 32144 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_279
timestamp 1698431365
transform 1 0 32592 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_340
timestamp 1698431365
transform 1 0 39424 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_344
timestamp 1698431365
transform 1 0 39872 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_348
timestamp 1698431365
transform 1 0 40320 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_352
timestamp 1698431365
transform 1 0 40768 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_385
timestamp 1698431365
transform 1 0 44464 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_387
timestamp 1698431365
transform 1 0 44688 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_398
timestamp 1698431365
transform 1 0 45920 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_402
timestamp 1698431365
transform 1 0 46368 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_416
timestamp 1698431365
transform 1 0 47936 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_2
timestamp 1698431365
transform 1 0 1568 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_18
timestamp 1698431365
transform 1 0 3360 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_26
timestamp 1698431365
transform 1 0 4256 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_37
timestamp 1698431365
transform 1 0 5488 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_41
timestamp 1698431365
transform 1 0 5936 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_43
timestamp 1698431365
transform 1 0 6160 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_46
timestamp 1698431365
transform 1 0 6496 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_107
timestamp 1698431365
transform 1 0 13328 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_172
timestamp 1698431365
transform 1 0 20608 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_174
timestamp 1698431365
transform 1 0 20832 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_177
timestamp 1698431365
transform 1 0 21168 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_203
timestamp 1698431365
transform 1 0 24080 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_210
timestamp 1698431365
transform 1 0 24864 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_238
timestamp 1698431365
transform 1 0 28000 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_247
timestamp 1698431365
transform 1 0 29008 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_249
timestamp 1698431365
transform 1 0 29232 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_260
timestamp 1698431365
transform 1 0 30464 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_290
timestamp 1698431365
transform 1 0 33824 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_294
timestamp 1698431365
transform 1 0 34272 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_301
timestamp 1698431365
transform 1 0 35056 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_303
timestamp 1698431365
transform 1 0 35280 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_325
timestamp 1698431365
transform 1 0 37744 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_327
timestamp 1698431365
transform 1 0 37968 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_357
timestamp 1698431365
transform 1 0 41328 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_367
timestamp 1698431365
transform 1 0 42448 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_371
timestamp 1698431365
transform 1 0 42896 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_381
timestamp 1698431365
transform 1 0 44016 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_387
timestamp 1698431365
transform 1 0 44688 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_2
timestamp 1698431365
transform 1 0 1568 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_34
timestamp 1698431365
transform 1 0 5152 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_36
timestamp 1698431365
transform 1 0 5376 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_80
timestamp 1698431365
transform 1 0 10304 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_122
timestamp 1698431365
transform 1 0 15008 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_139
timestamp 1698431365
transform 1 0 16912 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_165
timestamp 1698431365
transform 1 0 19824 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_177
timestamp 1698431365
transform 1 0 21168 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_181
timestamp 1698431365
transform 1 0 21616 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_184
timestamp 1698431365
transform 1 0 21952 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_188
timestamp 1698431365
transform 1 0 22400 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_192
timestamp 1698431365
transform 1 0 22848 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_196
timestamp 1698431365
transform 1 0 23296 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_203
timestamp 1698431365
transform 1 0 24080 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_207
timestamp 1698431365
transform 1 0 24528 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_218
timestamp 1698431365
transform 1 0 25760 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_222
timestamp 1698431365
transform 1 0 26208 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_244
timestamp 1698431365
transform 1 0 28672 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_246
timestamp 1698431365
transform 1 0 28896 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_290
timestamp 1698431365
transform 1 0 33824 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_294
timestamp 1698431365
transform 1 0 34272 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_298
timestamp 1698431365
transform 1 0 34720 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_309
timestamp 1698431365
transform 1 0 35952 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_313
timestamp 1698431365
transform 1 0 36400 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_317
timestamp 1698431365
transform 1 0 36848 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_321
timestamp 1698431365
transform 1 0 37296 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_325
timestamp 1698431365
transform 1 0 37744 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_329
timestamp 1698431365
transform 1 0 38192 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_342
timestamp 1698431365
transform 1 0 39648 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_352
timestamp 1698431365
transform 1 0 40768 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_363
timestamp 1698431365
transform 1 0 42000 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_371
timestamp 1698431365
transform 1 0 42896 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_373
timestamp 1698431365
transform 1 0 43120 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_380
timestamp 1698431365
transform 1 0 43904 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_388
timestamp 1698431365
transform 1 0 44800 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_390
timestamp 1698431365
transform 1 0 45024 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_397
timestamp 1698431365
transform 1 0 45808 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_401
timestamp 1698431365
transform 1 0 46256 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_403
timestamp 1698431365
transform 1 0 46480 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_412
timestamp 1698431365
transform 1 0 47488 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_416
timestamp 1698431365
transform 1 0 47936 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_2
timestamp 1698431365
transform 1 0 1568 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_18
timestamp 1698431365
transform 1 0 3360 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_26
timestamp 1698431365
transform 1 0 4256 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_37
timestamp 1698431365
transform 1 0 5488 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_41
timestamp 1698431365
transform 1 0 5936 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_53
timestamp 1698431365
transform 1 0 7280 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_61
timestamp 1698431365
transform 1 0 8176 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_63
timestamp 1698431365
transform 1 0 8400 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_101
timestamp 1698431365
transform 1 0 12656 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_130
timestamp 1698431365
transform 1 0 15904 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_173
timestamp 1698431365
transform 1 0 20720 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_208
timestamp 1698431365
transform 1 0 24640 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_242
timestamp 1698431365
transform 1 0 28448 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_244
timestamp 1698431365
transform 1 0 28672 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_314
timestamp 1698431365
transform 1 0 36512 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_331
timestamp 1698431365
transform 1 0 38416 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_368
timestamp 1698431365
transform 1 0 42560 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_375
timestamp 1698431365
transform 1 0 43344 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_379
timestamp 1698431365
transform 1 0 43792 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_383
timestamp 1698431365
transform 1 0 44240 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_393
timestamp 1698431365
transform 1 0 45360 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_397
timestamp 1698431365
transform 1 0 45808 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_399
timestamp 1698431365
transform 1 0 46032 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_413
timestamp 1698431365
transform 1 0 47600 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_2
timestamp 1698431365
transform 1 0 1568 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_18
timestamp 1698431365
transform 1 0 3360 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_54
timestamp 1698431365
transform 1 0 7392 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_72
timestamp 1698431365
transform 1 0 9408 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_104
timestamp 1698431365
transform 1 0 12992 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_106
timestamp 1698431365
transform 1 0 13216 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_133
timestamp 1698431365
transform 1 0 16240 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_150
timestamp 1698431365
transform 1 0 18144 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_152
timestamp 1698431365
transform 1 0 18368 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_193
timestamp 1698431365
transform 1 0 22960 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_208
timestamp 1698431365
transform 1 0 24640 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_212
timestamp 1698431365
transform 1 0 25088 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_214
timestamp 1698431365
transform 1 0 25312 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_240
timestamp 1698431365
transform 1 0 28224 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_248
timestamp 1698431365
transform 1 0 29120 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_289
timestamp 1698431365
transform 1 0 33712 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_293
timestamp 1698431365
transform 1 0 34160 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_303
timestamp 1698431365
transform 1 0 35280 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_307
timestamp 1698431365
transform 1 0 35728 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_309
timestamp 1698431365
transform 1 0 35952 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_339
timestamp 1698431365
transform 1 0 39312 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_343
timestamp 1698431365
transform 1 0 39760 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_347
timestamp 1698431365
transform 1 0 40208 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_349
timestamp 1698431365
transform 1 0 40432 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_373
timestamp 1698431365
transform 1 0 43120 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_381
timestamp 1698431365
transform 1 0 44016 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_2
timestamp 1698431365
transform 1 0 1568 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_6
timestamp 1698431365
transform 1 0 2016 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_22
timestamp 1698431365
transform 1 0 3808 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_26
timestamp 1698431365
transform 1 0 4256 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_37
timestamp 1698431365
transform 1 0 5488 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_56
timestamp 1698431365
transform 1 0 7616 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_60
timestamp 1698431365
transform 1 0 8064 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_62
timestamp 1698431365
transform 1 0 8288 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_78
timestamp 1698431365
transform 1 0 10080 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_185
timestamp 1698431365
transform 1 0 22064 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_187
timestamp 1698431365
transform 1 0 22288 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_244
timestamp 1698431365
transform 1 0 28672 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_259
timestamp 1698431365
transform 1 0 30352 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_311
timestamp 1698431365
transform 1 0 36176 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_331
timestamp 1698431365
transform 1 0 38416 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_333
timestamp 1698431365
transform 1 0 38640 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_346
timestamp 1698431365
transform 1 0 40096 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_354
timestamp 1698431365
transform 1 0 40992 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_387
timestamp 1698431365
transform 1 0 44688 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_391
timestamp 1698431365
transform 1 0 45136 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_393
timestamp 1698431365
transform 1 0 45360 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_400
timestamp 1698431365
transform 1 0 46144 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_416
timestamp 1698431365
transform 1 0 47936 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_33_10
timestamp 1698431365
transform 1 0 2464 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_26
timestamp 1698431365
transform 1 0 4256 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_34
timestamp 1698431365
transform 1 0 5152 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_51
timestamp 1698431365
transform 1 0 7056 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_53
timestamp 1698431365
transform 1 0 7280 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_69
timestamp 1698431365
transform 1 0 9072 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_96
timestamp 1698431365
transform 1 0 12096 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_276
timestamp 1698431365
transform 1 0 32256 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_298
timestamp 1698431365
transform 1 0 34720 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_33_332
timestamp 1698431365
transform 1 0 38528 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_348
timestamp 1698431365
transform 1 0 40320 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_352
timestamp 1698431365
transform 1 0 40768 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_356
timestamp 1698431365
transform 1 0 41216 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_364
timestamp 1698431365
transform 1 0 42112 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_368
timestamp 1698431365
transform 1 0 42560 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_377
timestamp 1698431365
transform 1 0 43568 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_416
timestamp 1698431365
transform 1 0 47936 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_31
timestamp 1698431365
transform 1 0 4816 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_37
timestamp 1698431365
transform 1 0 5488 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_45
timestamp 1698431365
transform 1 0 6384 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_60
timestamp 1698431365
transform 1 0 8064 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_104
timestamp 1698431365
transform 1 0 12992 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_128
timestamp 1698431365
transform 1 0 15680 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_159
timestamp 1698431365
transform 1 0 19152 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_284
timestamp 1698431365
transform 1 0 33152 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_294
timestamp 1698431365
transform 1 0 34272 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_310
timestamp 1698431365
transform 1 0 36064 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_314
timestamp 1698431365
transform 1 0 36512 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_317
timestamp 1698431365
transform 1 0 36848 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_321
timestamp 1698431365
transform 1 0 37296 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_359
timestamp 1698431365
transform 1 0 41552 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_361
timestamp 1698431365
transform 1 0 41776 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_374
timestamp 1698431365
transform 1 0 43232 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_381
timestamp 1698431365
transform 1 0 44016 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_34_387
timestamp 1698431365
transform 1 0 44688 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_403
timestamp 1698431365
transform 1 0 46480 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_412
timestamp 1698431365
transform 1 0 47488 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_2
timestamp 1698431365
transform 1 0 1568 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_6
timestamp 1698431365
transform 1 0 2016 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_66
timestamp 1698431365
transform 1 0 8736 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_91
timestamp 1698431365
transform 1 0 11536 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_150
timestamp 1698431365
transform 1 0 18144 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_311
timestamp 1698431365
transform 1 0 36176 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_315
timestamp 1698431365
transform 1 0 36624 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_344
timestamp 1698431365
transform 1 0 39872 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_348
timestamp 1698431365
transform 1 0 40320 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_352
timestamp 1698431365
transform 1 0 40768 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_362
timestamp 1698431365
transform 1 0 41888 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_372
timestamp 1698431365
transform 1 0 43008 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_376
timestamp 1698431365
transform 1 0 43456 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_390
timestamp 1698431365
transform 1 0 45024 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_397
timestamp 1698431365
transform 1 0 45808 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_404
timestamp 1698431365
transform 1 0 46592 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_418
timestamp 1698431365
transform 1 0 48160 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_30
timestamp 1698431365
transform 1 0 4704 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_34
timestamp 1698431365
transform 1 0 5152 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_37
timestamp 1698431365
transform 1 0 5488 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_55
timestamp 1698431365
transform 1 0 7504 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_78
timestamp 1698431365
transform 1 0 10080 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_107
timestamp 1698431365
transform 1 0 13328 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_123
timestamp 1698431365
transform 1 0 15120 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_161
timestamp 1698431365
transform 1 0 19376 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_163
timestamp 1698431365
transform 1 0 19600 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_255
timestamp 1698431365
transform 1 0 29904 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_296
timestamp 1698431365
transform 1 0 34496 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_304
timestamp 1698431365
transform 1 0 35392 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_308
timestamp 1698431365
transform 1 0 35840 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_312
timestamp 1698431365
transform 1 0 36288 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_314
timestamp 1698431365
transform 1 0 36512 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_317
timestamp 1698431365
transform 1 0 36848 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_321
timestamp 1698431365
transform 1 0 37296 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_36_338
timestamp 1698431365
transform 1 0 39200 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_354
timestamp 1698431365
transform 1 0 40992 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_384
timestamp 1698431365
transform 1 0 44352 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_387
timestamp 1698431365
transform 1 0 44688 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_31
timestamp 1698431365
transform 1 0 4816 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_35
timestamp 1698431365
transform 1 0 5264 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_39
timestamp 1698431365
transform 1 0 5712 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_48
timestamp 1698431365
transform 1 0 6720 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_52
timestamp 1698431365
transform 1 0 7168 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_61
timestamp 1698431365
transform 1 0 8176 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_88
timestamp 1698431365
transform 1 0 11200 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_112
timestamp 1698431365
transform 1 0 13888 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_142
timestamp 1698431365
transform 1 0 17248 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_144
timestamp 1698431365
transform 1 0 17472 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_209
timestamp 1698431365
transform 1 0 24752 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_212
timestamp 1698431365
transform 1 0 25088 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_214
timestamp 1698431365
transform 1 0 25312 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_279
timestamp 1698431365
transform 1 0 32592 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_282
timestamp 1698431365
transform 1 0 32928 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_301
timestamp 1698431365
transform 1 0 35056 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_305
timestamp 1698431365
transform 1 0 35504 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_310
timestamp 1698431365
transform 1 0 36064 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_314
timestamp 1698431365
transform 1 0 36512 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_317
timestamp 1698431365
transform 1 0 36848 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_327
timestamp 1698431365
transform 1 0 37968 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_335
timestamp 1698431365
transform 1 0 38864 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_339
timestamp 1698431365
transform 1 0 39312 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_349
timestamp 1698431365
transform 1 0 40432 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_352
timestamp 1698431365
transform 1 0 40768 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_354
timestamp 1698431365
transform 1 0 40992 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_363
timestamp 1698431365
transform 1 0 42000 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_371
timestamp 1698431365
transform 1 0 42896 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_396
timestamp 1698431365
transform 1 0 45696 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_404
timestamp 1698431365
transform 1 0 46592 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_415
timestamp 1698431365
transform 1 0 47824 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_419
timestamp 1698431365
transform 1 0 48272 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_2
timestamp 1698431365
transform 1 0 1568 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_6
timestamp 1698431365
transform 1 0 2016 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_37
timestamp 1698431365
transform 1 0 5488 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_41
timestamp 1698431365
transform 1 0 5936 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_59
timestamp 1698431365
transform 1 0 7952 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_63
timestamp 1698431365
transform 1 0 8400 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_65
timestamp 1698431365
transform 1 0 8624 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_107
timestamp 1698431365
transform 1 0 13328 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_203
timestamp 1698431365
transform 1 0 24080 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_253
timestamp 1698431365
transform 1 0 29680 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_270
timestamp 1698431365
transform 1 0 31584 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_375
timestamp 1698431365
transform 1 0 43344 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_381
timestamp 1698431365
transform 1 0 44016 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_392
timestamp 1698431365
transform 1 0 45248 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_409
timestamp 1698431365
transform 1 0 47152 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_411
timestamp 1698431365
transform 1 0 47376 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_2
timestamp 1698431365
transform 1 0 1568 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_10
timestamp 1698431365
transform 1 0 2464 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_14
timestamp 1698431365
transform 1 0 2912 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_16
timestamp 1698431365
transform 1 0 3136 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_72
timestamp 1698431365
transform 1 0 9408 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_126
timestamp 1698431365
transform 1 0 15456 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_155
timestamp 1698431365
transform 1 0 18704 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_157
timestamp 1698431365
transform 1 0 18928 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_185
timestamp 1698431365
transform 1 0 22064 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_212
timestamp 1698431365
transform 1 0 25088 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_230
timestamp 1698431365
transform 1 0 27104 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_234
timestamp 1698431365
transform 1 0 27552 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_259
timestamp 1698431365
transform 1 0 30352 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_276
timestamp 1698431365
transform 1 0 32256 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_302
timestamp 1698431365
transform 1 0 35168 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_312
timestamp 1698431365
transform 1 0 36288 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_316
timestamp 1698431365
transform 1 0 36736 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_318
timestamp 1698431365
transform 1 0 36960 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_39_324
timestamp 1698431365
transform 1 0 37632 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_340
timestamp 1698431365
transform 1 0 39424 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_348
timestamp 1698431365
transform 1 0 40320 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_389
timestamp 1698431365
transform 1 0 44912 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_2
timestamp 1698431365
transform 1 0 1568 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_6
timestamp 1698431365
transform 1 0 2016 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_16
timestamp 1698431365
transform 1 0 3136 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_22
timestamp 1698431365
transform 1 0 3808 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_37
timestamp 1698431365
transform 1 0 5488 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_88
timestamp 1698431365
transform 1 0 11200 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_173
timestamp 1698431365
transform 1 0 20720 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_184
timestamp 1698431365
transform 1 0 21952 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_186
timestamp 1698431365
transform 1 0 22176 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_222
timestamp 1698431365
transform 1 0 26208 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_226
timestamp 1698431365
transform 1 0 26656 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_240
timestamp 1698431365
transform 1 0 28224 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_242
timestamp 1698431365
transform 1 0 28448 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_255
timestamp 1698431365
transform 1 0 29904 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_286
timestamp 1698431365
transform 1 0 33376 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_40_290
timestamp 1698431365
transform 1 0 33824 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_306
timestamp 1698431365
transform 1 0 35616 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_314
timestamp 1698431365
transform 1 0 36512 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_339
timestamp 1698431365
transform 1 0 39312 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_40_343
timestamp 1698431365
transform 1 0 39760 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_359
timestamp 1698431365
transform 1 0 41552 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_367
timestamp 1698431365
transform 1 0 42448 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_371
timestamp 1698431365
transform 1 0 42896 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_387
timestamp 1698431365
transform 1 0 44688 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_2
timestamp 1698431365
transform 1 0 1568 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_6
timestamp 1698431365
transform 1 0 2016 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_19
timestamp 1698431365
transform 1 0 3472 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_28
timestamp 1698431365
transform 1 0 4480 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_32
timestamp 1698431365
transform 1 0 4928 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_59
timestamp 1698431365
transform 1 0 7952 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_63
timestamp 1698431365
transform 1 0 8400 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_134
timestamp 1698431365
transform 1 0 16352 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_159
timestamp 1698431365
transform 1 0 19152 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_208
timestamp 1698431365
transform 1 0 24640 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_212
timestamp 1698431365
transform 1 0 25088 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_258
timestamp 1698431365
transform 1 0 30240 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_262
timestamp 1698431365
transform 1 0 30688 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_273
timestamp 1698431365
transform 1 0 31920 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_277
timestamp 1698431365
transform 1 0 32368 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_279
timestamp 1698431365
transform 1 0 32592 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_282
timestamp 1698431365
transform 1 0 32928 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_290
timestamp 1698431365
transform 1 0 33824 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_294
timestamp 1698431365
transform 1 0 34272 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_297
timestamp 1698431365
transform 1 0 34608 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_348
timestamp 1698431365
transform 1 0 40320 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_352
timestamp 1698431365
transform 1 0 40768 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_360
timestamp 1698431365
transform 1 0 41664 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_364
timestamp 1698431365
transform 1 0 42112 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_366
timestamp 1698431365
transform 1 0 42336 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_396
timestamp 1698431365
transform 1 0 45696 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_403
timestamp 1698431365
transform 1 0 46480 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_407
timestamp 1698431365
transform 1 0 46928 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_415
timestamp 1698431365
transform 1 0 47824 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_419
timestamp 1698431365
transform 1 0 48272 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_37
timestamp 1698431365
transform 1 0 5488 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_41
timestamp 1698431365
transform 1 0 5936 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_54
timestamp 1698431365
transform 1 0 7392 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_58
timestamp 1698431365
transform 1 0 7840 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_60
timestamp 1698431365
transform 1 0 8064 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_67
timestamp 1698431365
transform 1 0 8848 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_90
timestamp 1698431365
transform 1 0 11424 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_163
timestamp 1698431365
transform 1 0 19600 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_165
timestamp 1698431365
transform 1 0 19824 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_174
timestamp 1698431365
transform 1 0 20832 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_230
timestamp 1698431365
transform 1 0 27104 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_243
timestamp 1698431365
transform 1 0 28560 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_260
timestamp 1698431365
transform 1 0 30464 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_264
timestamp 1698431365
transform 1 0 30912 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_306
timestamp 1698431365
transform 1 0 35616 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_308
timestamp 1698431365
transform 1 0 35840 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_317
timestamp 1698431365
transform 1 0 36848 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_321
timestamp 1698431365
transform 1 0 37296 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_329
timestamp 1698431365
transform 1 0 38192 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_331
timestamp 1698431365
transform 1 0 38416 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_375
timestamp 1698431365
transform 1 0 43344 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_383
timestamp 1698431365
transform 1 0 44240 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_387
timestamp 1698431365
transform 1 0 44688 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_397
timestamp 1698431365
transform 1 0 45808 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_401
timestamp 1698431365
transform 1 0 46256 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_417
timestamp 1698431365
transform 1 0 48048 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_419
timestamp 1698431365
transform 1 0 48272 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_2
timestamp 1698431365
transform 1 0 1568 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_10
timestamp 1698431365
transform 1 0 2464 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_29
timestamp 1698431365
transform 1 0 4592 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_31
timestamp 1698431365
transform 1 0 4816 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_69
timestamp 1698431365
transform 1 0 9072 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_72
timestamp 1698431365
transform 1 0 9408 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_76
timestamp 1698431365
transform 1 0 9856 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_89
timestamp 1698431365
transform 1 0 11312 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_102
timestamp 1698431365
transform 1 0 12768 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_110
timestamp 1698431365
transform 1 0 13664 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_114
timestamp 1698431365
transform 1 0 14112 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_128
timestamp 1698431365
transform 1 0 15680 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_154
timestamp 1698431365
transform 1 0 18592 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_178
timestamp 1698431365
transform 1 0 21280 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_204
timestamp 1698431365
transform 1 0 24192 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_218
timestamp 1698431365
transform 1 0 25760 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_222
timestamp 1698431365
transform 1 0 26208 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_226
timestamp 1698431365
transform 1 0 26656 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_230
timestamp 1698431365
transform 1 0 27104 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_239
timestamp 1698431365
transform 1 0 28112 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_264
timestamp 1698431365
transform 1 0 30912 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_272
timestamp 1698431365
transform 1 0 31808 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_276
timestamp 1698431365
transform 1 0 32256 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_290
timestamp 1698431365
transform 1 0 33824 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_314
timestamp 1698431365
transform 1 0 36512 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_322
timestamp 1698431365
transform 1 0 37408 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_324
timestamp 1698431365
transform 1 0 37632 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_327
timestamp 1698431365
transform 1 0 37968 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_345
timestamp 1698431365
transform 1 0 39984 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_349
timestamp 1698431365
transform 1 0 40432 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_352
timestamp 1698431365
transform 1 0 40768 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_30
timestamp 1698431365
transform 1 0 4704 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_34
timestamp 1698431365
transform 1 0 5152 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_37
timestamp 1698431365
transform 1 0 5488 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_41
timestamp 1698431365
transform 1 0 5936 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_80
timestamp 1698431365
transform 1 0 10304 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_90
timestamp 1698431365
transform 1 0 11424 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_107
timestamp 1698431365
transform 1 0 13328 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_144
timestamp 1698431365
transform 1 0 17472 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_154
timestamp 1698431365
transform 1 0 18592 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_183
timestamp 1698431365
transform 1 0 21840 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_190
timestamp 1698431365
transform 1 0 22624 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_198
timestamp 1698431365
transform 1 0 23520 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_212
timestamp 1698431365
transform 1 0 25088 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_214
timestamp 1698431365
transform 1 0 25312 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_223
timestamp 1698431365
transform 1 0 26320 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_227
timestamp 1698431365
transform 1 0 26768 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_235
timestamp 1698431365
transform 1 0 27664 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_239
timestamp 1698431365
transform 1 0 28112 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_243
timestamp 1698431365
transform 1 0 28560 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_266
timestamp 1698431365
transform 1 0 31136 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_270
timestamp 1698431365
transform 1 0 31584 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_272
timestamp 1698431365
transform 1 0 31808 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_313
timestamp 1698431365
transform 1 0 36400 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_331
timestamp 1698431365
transform 1 0 38416 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_374
timestamp 1698431365
transform 1 0 43232 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_376
timestamp 1698431365
transform 1 0 43456 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_387
timestamp 1698431365
transform 1 0 44688 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_37
timestamp 1698431365
transform 1 0 5488 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_41
timestamp 1698431365
transform 1 0 5936 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_48
timestamp 1698431365
transform 1 0 6720 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_87
timestamp 1698431365
transform 1 0 11088 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_89
timestamp 1698431365
transform 1 0 11312 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_174
timestamp 1698431365
transform 1 0 20832 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_176
timestamp 1698431365
transform 1 0 21056 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_197
timestamp 1698431365
transform 1 0 23408 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_241
timestamp 1698431365
transform 1 0 28336 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_243
timestamp 1698431365
transform 1 0 28560 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_45_250
timestamp 1698431365
transform 1 0 29344 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_278
timestamp 1698431365
transform 1 0 32480 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_295
timestamp 1698431365
transform 1 0 34384 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_326
timestamp 1698431365
transform 1 0 37856 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_338
timestamp 1698431365
transform 1 0 39200 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_346
timestamp 1698431365
transform 1 0 40096 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_352
timestamp 1698431365
transform 1 0 40768 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_382
timestamp 1698431365
transform 1 0 44128 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_2
timestamp 1698431365
transform 1 0 1568 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_10
timestamp 1698431365
transform 1 0 2464 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_33
timestamp 1698431365
transform 1 0 5040 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_89
timestamp 1698431365
transform 1 0 11312 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_115
timestamp 1698431365
transform 1 0 14224 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_134
timestamp 1698431365
transform 1 0 16352 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_138
timestamp 1698431365
transform 1 0 16800 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_142
timestamp 1698431365
transform 1 0 17248 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_169
timestamp 1698431365
transform 1 0 20272 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_177
timestamp 1698431365
transform 1 0 21168 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_192
timestamp 1698431365
transform 1 0 22848 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_196
timestamp 1698431365
transform 1 0 23296 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_226
timestamp 1698431365
transform 1 0 26656 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_230
timestamp 1698431365
transform 1 0 27104 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_311
timestamp 1698431365
transform 1 0 36176 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_325
timestamp 1698431365
transform 1 0 37744 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_332
timestamp 1698431365
transform 1 0 38528 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_373
timestamp 1698431365
transform 1 0 43120 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_377
timestamp 1698431365
transform 1 0 43568 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_387
timestamp 1698431365
transform 1 0 44688 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_47_2
timestamp 1698431365
transform 1 0 1568 0 -1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_47_18
timestamp 1698431365
transform 1 0 3360 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_47_31
timestamp 1698431365
transform 1 0 4816 0 -1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_47_47
timestamp 1698431365
transform 1 0 6608 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_55
timestamp 1698431365
transform 1 0 7504 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_57
timestamp 1698431365
transform 1 0 7728 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_72
timestamp 1698431365
transform 1 0 9408 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_74
timestamp 1698431365
transform 1 0 9632 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_117
timestamp 1698431365
transform 1 0 14448 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_121
timestamp 1698431365
transform 1 0 14896 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_123
timestamp 1698431365
transform 1 0 15120 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_136
timestamp 1698431365
transform 1 0 16576 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_142
timestamp 1698431365
transform 1 0 17248 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_186
timestamp 1698431365
transform 1 0 22176 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_47_190
timestamp 1698431365
transform 1 0 22624 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_198
timestamp 1698431365
transform 1 0 23520 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_208
timestamp 1698431365
transform 1 0 24640 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_47_212
timestamp 1698431365
transform 1 0 25088 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_220
timestamp 1698431365
transform 1 0 25984 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_224
timestamp 1698431365
transform 1 0 26432 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_226
timestamp 1698431365
transform 1 0 26656 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_240
timestamp 1698431365
transform 1 0 28224 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_242
timestamp 1698431365
transform 1 0 28448 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_47_261
timestamp 1698431365
transform 1 0 30576 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_269
timestamp 1698431365
transform 1 0 31472 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_278
timestamp 1698431365
transform 1 0 32480 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_282
timestamp 1698431365
transform 1 0 32928 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_288
timestamp 1698431365
transform 1 0 33600 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_312
timestamp 1698431365
transform 1 0 36288 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_316
timestamp 1698431365
transform 1 0 36736 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_320
timestamp 1698431365
transform 1 0 37184 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_360
timestamp 1698431365
transform 1 0 41664 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_364
timestamp 1698431365
transform 1 0 42112 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_366
timestamp 1698431365
transform 1 0 42336 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_402
timestamp 1698431365
transform 1 0 46368 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_48_2
timestamp 1698431365
transform 1 0 1568 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_10
timestamp 1698431365
transform 1 0 2464 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_30
timestamp 1698431365
transform 1 0 4704 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_34
timestamp 1698431365
transform 1 0 5152 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_48_37
timestamp 1698431365
transform 1 0 5488 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_45
timestamp 1698431365
transform 1 0 6384 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_61
timestamp 1698431365
transform 1 0 8176 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_70
timestamp 1698431365
transform 1 0 9184 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_74
timestamp 1698431365
transform 1 0 9632 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_119
timestamp 1698431365
transform 1 0 14672 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_160
timestamp 1698431365
transform 1 0 19264 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_168
timestamp 1698431365
transform 1 0 20160 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_200
timestamp 1698431365
transform 1 0 23744 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_48_222
timestamp 1698431365
transform 1 0 26208 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_238
timestamp 1698431365
transform 1 0 28000 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_242
timestamp 1698431365
transform 1 0 28448 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_244
timestamp 1698431365
transform 1 0 28672 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_48_262
timestamp 1698431365
transform 1 0 30688 0 1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_321
timestamp 1698431365
transform 1 0 37296 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_336
timestamp 1698431365
transform 1 0 38976 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_367
timestamp 1698431365
transform 1 0 42448 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_369
timestamp 1698431365
transform 1 0 42672 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_378
timestamp 1698431365
transform 1 0 43680 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_382
timestamp 1698431365
transform 1 0 44128 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_384
timestamp 1698431365
transform 1 0 44352 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_387
timestamp 1698431365
transform 1 0 44688 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_31
timestamp 1698431365
transform 1 0 4816 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_33
timestamp 1698431365
transform 1 0 5040 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_63
timestamp 1698431365
transform 1 0 8400 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_67
timestamp 1698431365
transform 1 0 8848 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_69
timestamp 1698431365
transform 1 0 9072 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_76
timestamp 1698431365
transform 1 0 9856 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_142
timestamp 1698431365
transform 1 0 17248 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_161
timestamp 1698431365
transform 1 0 19376 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_49_192
timestamp 1698431365
transform 1 0 22848 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_200
timestamp 1698431365
transform 1 0 23744 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_245
timestamp 1698431365
transform 1 0 28784 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_247
timestamp 1698431365
transform 1 0 29008 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_49_261
timestamp 1698431365
transform 1 0 30576 0 -1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_277
timestamp 1698431365
transform 1 0 32368 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_279
timestamp 1698431365
transform 1 0 32592 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_288
timestamp 1698431365
transform 1 0 33600 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_333
timestamp 1698431365
transform 1 0 38640 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_337
timestamp 1698431365
transform 1 0 39088 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_341
timestamp 1698431365
transform 1 0 39536 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_343
timestamp 1698431365
transform 1 0 39760 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_348
timestamp 1698431365
transform 1 0 40320 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_352
timestamp 1698431365
transform 1 0 40768 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_49_356
timestamp 1698431365
transform 1 0 41216 0 -1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_388
timestamp 1698431365
transform 1 0 44800 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_392
timestamp 1698431365
transform 1 0 45248 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_415
timestamp 1698431365
transform 1 0 47824 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_419
timestamp 1698431365
transform 1 0 48272 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_2
timestamp 1698431365
transform 1 0 1568 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_33
timestamp 1698431365
transform 1 0 5040 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_73
timestamp 1698431365
transform 1 0 9520 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_89
timestamp 1698431365
transform 1 0 11312 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_91
timestamp 1698431365
transform 1 0 11536 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_102
timestamp 1698431365
transform 1 0 12768 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_104
timestamp 1698431365
transform 1 0 12992 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_107
timestamp 1698431365
transform 1 0 13328 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_115
timestamp 1698431365
transform 1 0 14224 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_117
timestamp 1698431365
transform 1 0 14448 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_138
timestamp 1698431365
transform 1 0 16800 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_169
timestamp 1698431365
transform 1 0 20272 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_177
timestamp 1698431365
transform 1 0 21168 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_205
timestamp 1698431365
transform 1 0 24304 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_209
timestamp 1698431365
transform 1 0 24752 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_211
timestamp 1698431365
transform 1 0 24976 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_224
timestamp 1698431365
transform 1 0 26432 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_228
timestamp 1698431365
transform 1 0 26880 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_237
timestamp 1698431365
transform 1 0 27888 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_247
timestamp 1698431365
transform 1 0 29008 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_251
timestamp 1698431365
transform 1 0 29456 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_276
timestamp 1698431365
transform 1 0 32256 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_301
timestamp 1698431365
transform 1 0 35056 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_309
timestamp 1698431365
transform 1 0 35952 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_313
timestamp 1698431365
transform 1 0 36400 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_325
timestamp 1698431365
transform 1 0 37744 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_349
timestamp 1698431365
transform 1 0 40432 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_353
timestamp 1698431365
transform 1 0 40880 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_384
timestamp 1698431365
transform 1 0 44352 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_387
timestamp 1698431365
transform 1 0 44688 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_391
timestamp 1698431365
transform 1 0 45136 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_399
timestamp 1698431365
transform 1 0 46032 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_403
timestamp 1698431365
transform 1 0 46480 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_407
timestamp 1698431365
transform 1 0 46928 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_411
timestamp 1698431365
transform 1 0 47376 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_415
timestamp 1698431365
transform 1 0 47824 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_417
timestamp 1698431365
transform 1 0 48048 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_51_2
timestamp 1698431365
transform 1 0 1568 0 -1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_18
timestamp 1698431365
transform 1 0 3360 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_51_39
timestamp 1698431365
transform 1 0 5712 0 -1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_55
timestamp 1698431365
transform 1 0 7504 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_57
timestamp 1698431365
transform 1 0 7728 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_63
timestamp 1698431365
transform 1 0 8400 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_67
timestamp 1698431365
transform 1 0 8848 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_69
timestamp 1698431365
transform 1 0 9072 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_72
timestamp 1698431365
transform 1 0 9408 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_76
timestamp 1698431365
transform 1 0 9856 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_51_107
timestamp 1698431365
transform 1 0 13328 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_115
timestamp 1698431365
transform 1 0 14224 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_119
timestamp 1698431365
transform 1 0 14672 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_123
timestamp 1698431365
transform 1 0 15120 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_51_191
timestamp 1698431365
transform 1 0 22736 0 -1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_207
timestamp 1698431365
transform 1 0 24528 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_209
timestamp 1698431365
transform 1 0 24752 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_216
timestamp 1698431365
transform 1 0 25536 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_242
timestamp 1698431365
transform 1 0 28448 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_244
timestamp 1698431365
transform 1 0 28672 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_51_267
timestamp 1698431365
transform 1 0 31248 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_275
timestamp 1698431365
transform 1 0 32144 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_279
timestamp 1698431365
transform 1 0 32592 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_319
timestamp 1698431365
transform 1 0 37072 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_323
timestamp 1698431365
transform 1 0 37520 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_327
timestamp 1698431365
transform 1 0 37968 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_340
timestamp 1698431365
transform 1 0 39424 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_344
timestamp 1698431365
transform 1 0 39872 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_348
timestamp 1698431365
transform 1 0 40320 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_356
timestamp 1698431365
transform 1 0 41216 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_51_360
timestamp 1698431365
transform 1 0 41664 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_368
timestamp 1698431365
transform 1 0 42560 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_372
timestamp 1698431365
transform 1 0 43008 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_413
timestamp 1698431365
transform 1 0 47600 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_417
timestamp 1698431365
transform 1 0 48048 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_31
timestamp 1698431365
transform 1 0 4816 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_37
timestamp 1698431365
transform 1 0 5488 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_41
timestamp 1698431365
transform 1 0 5936 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_60
timestamp 1698431365
transform 1 0 8064 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_64
timestamp 1698431365
transform 1 0 8512 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_71
timestamp 1698431365
transform 1 0 9296 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_78
timestamp 1698431365
transform 1 0 10080 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_80
timestamp 1698431365
transform 1 0 10304 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_91
timestamp 1698431365
transform 1 0 11536 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_100
timestamp 1698431365
transform 1 0 12544 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_104
timestamp 1698431365
transform 1 0 12992 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_52_107
timestamp 1698431365
transform 1 0 13328 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_115
timestamp 1698431365
transform 1 0 14224 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_156
timestamp 1698431365
transform 1 0 18816 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_160
timestamp 1698431365
transform 1 0 19264 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_163
timestamp 1698431365
transform 1 0 19600 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_167
timestamp 1698431365
transform 1 0 20048 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_171
timestamp 1698431365
transform 1 0 20496 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_52_177
timestamp 1698431365
transform 1 0 21168 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_185
timestamp 1698431365
transform 1 0 22064 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_189
timestamp 1698431365
transform 1 0 22512 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_193
timestamp 1698431365
transform 1 0 22960 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_195
timestamp 1698431365
transform 1 0 23184 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_239
timestamp 1698431365
transform 1 0 28112 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_243
timestamp 1698431365
transform 1 0 28560 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_52_279
timestamp 1698431365
transform 1 0 32592 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_287
timestamp 1698431365
transform 1 0 33488 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_289
timestamp 1698431365
transform 1 0 33712 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_299
timestamp 1698431365
transform 1 0 34832 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_303
timestamp 1698431365
transform 1 0 35280 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_305
timestamp 1698431365
transform 1 0 35504 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_312
timestamp 1698431365
transform 1 0 36288 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_314
timestamp 1698431365
transform 1 0 36512 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_317
timestamp 1698431365
transform 1 0 36848 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_321
timestamp 1698431365
transform 1 0 37296 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_325
timestamp 1698431365
transform 1 0 37744 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_331
timestamp 1698431365
transform 1 0 38416 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_52_335
timestamp 1698431365
transform 1 0 38864 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_343
timestamp 1698431365
transform 1 0 39760 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_345
timestamp 1698431365
transform 1 0 39984 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_363
timestamp 1698431365
transform 1 0 42000 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_374
timestamp 1698431365
transform 1 0 43232 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_387
timestamp 1698431365
transform 1 0 44688 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_2
timestamp 1698431365
transform 1 0 1568 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_6
timestamp 1698431365
transform 1 0 2016 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_28
timestamp 1698431365
transform 1 0 4480 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_66
timestamp 1698431365
transform 1 0 8736 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_53_92
timestamp 1698431365
transform 1 0 11648 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_100
timestamp 1698431365
transform 1 0 12544 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_131
timestamp 1698431365
transform 1 0 16016 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_171
timestamp 1698431365
transform 1 0 20496 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_175
timestamp 1698431365
transform 1 0 20944 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_179
timestamp 1698431365
transform 1 0 21392 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_53_236
timestamp 1698431365
transform 1 0 27776 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_244
timestamp 1698431365
transform 1 0 28672 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_282
timestamp 1698431365
transform 1 0 32928 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_284
timestamp 1698431365
transform 1 0 33152 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_290
timestamp 1698431365
transform 1 0 33824 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_300
timestamp 1698431365
transform 1 0 34944 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_366
timestamp 1698431365
transform 1 0 42336 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_398
timestamp 1698431365
transform 1 0 45920 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_418
timestamp 1698431365
transform 1 0 48160 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_2
timestamp 1698431365
transform 1 0 1568 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_6
timestamp 1698431365
transform 1 0 2016 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_33
timestamp 1698431365
transform 1 0 5040 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_37
timestamp 1698431365
transform 1 0 5488 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_39
timestamp 1698431365
transform 1 0 5712 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_54_61
timestamp 1698431365
transform 1 0 8176 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_77
timestamp 1698431365
transform 1 0 9968 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_93
timestamp 1698431365
transform 1 0 11760 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_125
timestamp 1698431365
transform 1 0 15344 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_135
timestamp 1698431365
transform 1 0 16464 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_177
timestamp 1698431365
transform 1 0 21168 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_197
timestamp 1698431365
transform 1 0 23408 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_201
timestamp 1698431365
transform 1 0 23856 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_222
timestamp 1698431365
transform 1 0 26208 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_230
timestamp 1698431365
transform 1 0 27104 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_239
timestamp 1698431365
transform 1 0 28112 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_243
timestamp 1698431365
transform 1 0 28560 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_247
timestamp 1698431365
transform 1 0 29008 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_257
timestamp 1698431365
transform 1 0 30128 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_261
timestamp 1698431365
transform 1 0 30576 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_291
timestamp 1698431365
transform 1 0 33936 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_380
timestamp 1698431365
transform 1 0 43904 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_384
timestamp 1698431365
transform 1 0 44352 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_410
timestamp 1698431365
transform 1 0 47264 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_55_2
timestamp 1698431365
transform 1 0 1568 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_10
timestamp 1698431365
transform 1 0 2464 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_24
timestamp 1698431365
transform 1 0 4032 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_26
timestamp 1698431365
transform 1 0 4256 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_55_35
timestamp 1698431365
transform 1 0 5264 0 -1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_51
timestamp 1698431365
transform 1 0 7056 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_55_60
timestamp 1698431365
transform 1 0 8064 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_68
timestamp 1698431365
transform 1 0 8960 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_72
timestamp 1698431365
transform 1 0 9408 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_74
timestamp 1698431365
transform 1 0 9632 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_87
timestamp 1698431365
transform 1 0 11088 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_93
timestamp 1698431365
transform 1 0 11760 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_95
timestamp 1698431365
transform 1 0 11984 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_55_100
timestamp 1698431365
transform 1 0 12544 0 -1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_116
timestamp 1698431365
transform 1 0 14336 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_118
timestamp 1698431365
transform 1 0 14560 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_133
timestamp 1698431365
transform 1 0 16240 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_142
timestamp 1698431365
transform 1 0 17248 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_162
timestamp 1698431365
transform 1 0 19488 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_164
timestamp 1698431365
transform 1 0 19712 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_212
timestamp 1698431365
transform 1 0 25088 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_216
timestamp 1698431365
transform 1 0 25536 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_220
timestamp 1698431365
transform 1 0 25984 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_55_264
timestamp 1698431365
transform 1 0 30912 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_282
timestamp 1698431365
transform 1 0 32928 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_296
timestamp 1698431365
transform 1 0 34496 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_346
timestamp 1698431365
transform 1 0 40096 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_352
timestamp 1698431365
transform 1 0 40768 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_385
timestamp 1698431365
transform 1 0 44464 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_389
timestamp 1698431365
transform 1 0 44912 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_31
timestamp 1698431365
transform 1 0 4816 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_56_37
timestamp 1698431365
transform 1 0 5488 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_45
timestamp 1698431365
transform 1 0 6384 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_75
timestamp 1698431365
transform 1 0 9744 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_77
timestamp 1698431365
transform 1 0 9968 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_84
timestamp 1698431365
transform 1 0 10752 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_86
timestamp 1698431365
transform 1 0 10976 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_107
timestamp 1698431365
transform 1 0 13328 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_137
timestamp 1698431365
transform 1 0 16688 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_141
timestamp 1698431365
transform 1 0 17136 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_145
timestamp 1698431365
transform 1 0 17584 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_149
timestamp 1698431365
transform 1 0 18032 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_156
timestamp 1698431365
transform 1 0 18816 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_182
timestamp 1698431365
transform 1 0 21728 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_204
timestamp 1698431365
transform 1 0 24192 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_243
timestamp 1698431365
transform 1 0 28560 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_277
timestamp 1698431365
transform 1 0 32368 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_287
timestamp 1698431365
transform 1 0 33488 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_291
timestamp 1698431365
transform 1 0 33936 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_308
timestamp 1698431365
transform 1 0 35840 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_312
timestamp 1698431365
transform 1 0 36288 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_314
timestamp 1698431365
transform 1 0 36512 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_317
timestamp 1698431365
transform 1 0 36848 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_325
timestamp 1698431365
transform 1 0 37744 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_362
timestamp 1698431365
transform 1 0 41888 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_374
timestamp 1698431365
transform 1 0 43232 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_378
timestamp 1698431365
transform 1 0 43680 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_382
timestamp 1698431365
transform 1 0 44128 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_395
timestamp 1698431365
transform 1 0 45584 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_418
timestamp 1698431365
transform 1 0 48160 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_2
timestamp 1698431365
transform 1 0 1568 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_4
timestamp 1698431365
transform 1 0 1792 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_34
timestamp 1698431365
transform 1 0 5152 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_67
timestamp 1698431365
transform 1 0 8848 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_69
timestamp 1698431365
transform 1 0 9072 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_85
timestamp 1698431365
transform 1 0 10864 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_87
timestamp 1698431365
transform 1 0 11088 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_57_106
timestamp 1698431365
transform 1 0 13216 0 -1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_122
timestamp 1698431365
transform 1 0 15008 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_124
timestamp 1698431365
transform 1 0 15232 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_206
timestamp 1698431365
transform 1 0 24416 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_232
timestamp 1698431365
transform 1 0 27328 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_234
timestamp 1698431365
transform 1 0 27552 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_275
timestamp 1698431365
transform 1 0 32144 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_279
timestamp 1698431365
transform 1 0 32592 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_57_282
timestamp 1698431365
transform 1 0 32928 0 -1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_298
timestamp 1698431365
transform 1 0 34720 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_302
timestamp 1698431365
transform 1 0 35168 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_352
timestamp 1698431365
transform 1 0 40768 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_362
timestamp 1698431365
transform 1 0 41888 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_373
timestamp 1698431365
transform 1 0 43120 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_377
timestamp 1698431365
transform 1 0 43568 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_383
timestamp 1698431365
transform 1 0 44240 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_387
timestamp 1698431365
transform 1 0 44688 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_58_2
timestamp 1698431365
transform 1 0 1568 0 1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_18
timestamp 1698431365
transform 1 0 3360 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_20
timestamp 1698431365
transform 1 0 3584 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_23
timestamp 1698431365
transform 1 0 3920 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_27
timestamp 1698431365
transform 1 0 4368 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_29
timestamp 1698431365
transform 1 0 4592 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_58
timestamp 1698431365
transform 1 0 7840 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_62
timestamp 1698431365
transform 1 0 8288 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_79
timestamp 1698431365
transform 1 0 10192 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_83
timestamp 1698431365
transform 1 0 10640 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_87
timestamp 1698431365
transform 1 0 11088 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_89
timestamp 1698431365
transform 1 0 11312 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_95
timestamp 1698431365
transform 1 0 11984 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_99
timestamp 1698431365
transform 1 0 12432 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_103
timestamp 1698431365
transform 1 0 12880 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_107
timestamp 1698431365
transform 1 0 13328 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_111
timestamp 1698431365
transform 1 0 13776 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_58_117
timestamp 1698431365
transform 1 0 14448 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_156
timestamp 1698431365
transform 1 0 18816 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_160
timestamp 1698431365
transform 1 0 19264 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_173
timestamp 1698431365
transform 1 0 20720 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_58_177
timestamp 1698431365
transform 1 0 21168 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_185
timestamp 1698431365
transform 1 0 22064 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_187
timestamp 1698431365
transform 1 0 22288 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_194
timestamp 1698431365
transform 1 0 23072 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_198
timestamp 1698431365
transform 1 0 23520 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_210
timestamp 1698431365
transform 1 0 24864 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_247
timestamp 1698431365
transform 1 0 29008 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_283
timestamp 1698431365
transform 1 0 33040 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_299
timestamp 1698431365
transform 1 0 34832 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_301
timestamp 1698431365
transform 1 0 35056 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_312
timestamp 1698431365
transform 1 0 36288 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_314
timestamp 1698431365
transform 1 0 36512 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_317
timestamp 1698431365
transform 1 0 36848 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_321
timestamp 1698431365
transform 1 0 37296 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_58_327
timestamp 1698431365
transform 1 0 37968 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_335
timestamp 1698431365
transform 1 0 38864 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_338
timestamp 1698431365
transform 1 0 39200 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_342
timestamp 1698431365
transform 1 0 39648 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_348
timestamp 1698431365
transform 1 0 40320 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_395
timestamp 1698431365
transform 1 0 45584 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_399
timestamp 1698431365
transform 1 0 46032 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_407
timestamp 1698431365
transform 1 0 46928 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_409
timestamp 1698431365
transform 1 0 47152 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_54
timestamp 1698431365
transform 1 0 7392 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_59_60
timestamp 1698431365
transform 1 0 8064 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_68
timestamp 1698431365
transform 1 0 8960 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_59_72
timestamp 1698431365
transform 1 0 9408 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_80
timestamp 1698431365
transform 1 0 10304 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_98
timestamp 1698431365
transform 1 0 12320 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_102
timestamp 1698431365
transform 1 0 12768 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_59_125
timestamp 1698431365
transform 1 0 15344 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_133
timestamp 1698431365
transform 1 0 16240 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_137
timestamp 1698431365
transform 1 0 16688 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_139
timestamp 1698431365
transform 1 0 16912 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_59_142
timestamp 1698431365
transform 1 0 17248 0 -1 50176
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_59_174
timestamp 1698431365
transform 1 0 20832 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_182
timestamp 1698431365
transform 1 0 21728 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_186
timestamp 1698431365
transform 1 0 22176 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_193
timestamp 1698431365
transform 1 0 22960 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_205
timestamp 1698431365
transform 1 0 24304 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_209
timestamp 1698431365
transform 1 0 24752 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_212
timestamp 1698431365
transform 1 0 25088 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_216
timestamp 1698431365
transform 1 0 25536 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_255
timestamp 1698431365
transform 1 0 29904 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_59_259
timestamp 1698431365
transform 1 0 30352 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_267
timestamp 1698431365
transform 1 0 31248 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_271
timestamp 1698431365
transform 1 0 31696 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_273
timestamp 1698431365
transform 1 0 31920 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_320
timestamp 1698431365
transform 1 0 37184 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_324
timestamp 1698431365
transform 1 0 37632 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_326
timestamp 1698431365
transform 1 0 37856 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_331
timestamp 1698431365
transform 1 0 38416 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_349
timestamp 1698431365
transform 1 0 40432 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_352
timestamp 1698431365
transform 1 0 40768 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_354
timestamp 1698431365
transform 1 0 40992 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_369
timestamp 1698431365
transform 1 0 42672 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_399
timestamp 1698431365
transform 1 0 46032 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_404
timestamp 1698431365
transform 1 0 46592 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_60_10
timestamp 1698431365
transform 1 0 2464 0 1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_26
timestamp 1698431365
transform 1 0 4256 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_30
timestamp 1698431365
transform 1 0 4704 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_33
timestamp 1698431365
transform 1 0 5040 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_55
timestamp 1698431365
transform 1 0 7504 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_59
timestamp 1698431365
transform 1 0 7952 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_81
timestamp 1698431365
transform 1 0 10416 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_107
timestamp 1698431365
transform 1 0 13328 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_133
timestamp 1698431365
transform 1 0 16240 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_140
timestamp 1698431365
transform 1 0 17024 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_144
timestamp 1698431365
transform 1 0 17472 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_148
timestamp 1698431365
transform 1 0 17920 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_150
timestamp 1698431365
transform 1 0 18144 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_157
timestamp 1698431365
transform 1 0 18928 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_236
timestamp 1698431365
transform 1 0 27776 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_247
timestamp 1698431365
transform 1 0 29008 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_260
timestamp 1698431365
transform 1 0 30464 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_307
timestamp 1698431365
transform 1 0 35728 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_314
timestamp 1698431365
transform 1 0 36512 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_321
timestamp 1698431365
transform 1 0 37296 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_360
timestamp 1698431365
transform 1 0 41664 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_410
timestamp 1698431365
transform 1 0 47264 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_414
timestamp 1698431365
transform 1 0 47712 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_418
timestamp 1698431365
transform 1 0 48160 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_2
timestamp 1698431365
transform 1 0 1568 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_61_6
timestamp 1698431365
transform 1 0 2016 0 -1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_61_22
timestamp 1698431365
transform 1 0 3808 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_30
timestamp 1698431365
transform 1 0 4704 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_101
timestamp 1698431365
transform 1 0 12656 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_105
timestamp 1698431365
transform 1 0 13104 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_115
timestamp 1698431365
transform 1 0 14224 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_194
timestamp 1698431365
transform 1 0 23072 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_61_202
timestamp 1698431365
transform 1 0 23968 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_212
timestamp 1698431365
transform 1 0 25088 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_254
timestamp 1698431365
transform 1 0 29792 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_258
timestamp 1698431365
transform 1 0 30240 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_260
timestamp 1698431365
transform 1 0 30464 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_282
timestamp 1698431365
transform 1 0 32928 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_286
timestamp 1698431365
transform 1 0 33376 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_299
timestamp 1698431365
transform 1 0 34832 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_303
timestamp 1698431365
transform 1 0 35280 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_313
timestamp 1698431365
transform 1 0 36400 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_315
timestamp 1698431365
transform 1 0 36624 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_322
timestamp 1698431365
transform 1 0 37408 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_326
timestamp 1698431365
transform 1 0 37856 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_330
timestamp 1698431365
transform 1 0 38304 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_352
timestamp 1698431365
transform 1 0 40768 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_387
timestamp 1698431365
transform 1 0 44688 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_62_2
timestamp 1698431365
transform 1 0 1568 0 1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_34
timestamp 1698431365
transform 1 0 5152 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_45
timestamp 1698431365
transform 1 0 6384 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_63
timestamp 1698431365
transform 1 0 8400 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_67
timestamp 1698431365
transform 1 0 8848 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_76
timestamp 1698431365
transform 1 0 9856 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_78
timestamp 1698431365
transform 1 0 10080 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_85
timestamp 1698431365
transform 1 0 10864 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_62_89
timestamp 1698431365
transform 1 0 11312 0 1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_107
timestamp 1698431365
transform 1 0 13328 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_111
timestamp 1698431365
transform 1 0 13776 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_62_117
timestamp 1698431365
transform 1 0 14448 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_154
timestamp 1698431365
transform 1 0 18592 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_158
timestamp 1698431365
transform 1 0 19040 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_160
timestamp 1698431365
transform 1 0 19264 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_172
timestamp 1698431365
transform 1 0 20608 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_174
timestamp 1698431365
transform 1 0 20832 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_183
timestamp 1698431365
transform 1 0 21840 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_185
timestamp 1698431365
transform 1 0 22064 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_206
timestamp 1698431365
transform 1 0 24416 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_210
timestamp 1698431365
transform 1 0 24864 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_218
timestamp 1698431365
transform 1 0 25760 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_62_235
timestamp 1698431365
transform 1 0 27664 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_243
timestamp 1698431365
transform 1 0 28560 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_259
timestamp 1698431365
transform 1 0 30352 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_62_290
timestamp 1698431365
transform 1 0 33824 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_308
timestamp 1698431365
transform 1 0 35840 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_312
timestamp 1698431365
transform 1 0 36288 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_335
timestamp 1698431365
transform 1 0 38864 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_339
timestamp 1698431365
transform 1 0 39312 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_378
timestamp 1698431365
transform 1 0 43680 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_393
timestamp 1698431365
transform 1 0 45360 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_63_2
timestamp 1698431365
transform 1 0 1568 0 -1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_18
timestamp 1698431365
transform 1 0 3360 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_22
timestamp 1698431365
transform 1 0 3808 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_57
timestamp 1698431365
transform 1 0 7728 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_63_61
timestamp 1698431365
transform 1 0 8176 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_69
timestamp 1698431365
transform 1 0 9072 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_63_72
timestamp 1698431365
transform 1 0 9408 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_80
timestamp 1698431365
transform 1 0 10304 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_84
timestamp 1698431365
transform 1 0 10752 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_86
timestamp 1698431365
transform 1 0 10976 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_116
timestamp 1698431365
transform 1 0 14336 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_120
timestamp 1698431365
transform 1 0 14784 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_142
timestamp 1698431365
transform 1 0 17248 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_63_146
timestamp 1698431365
transform 1 0 17696 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_154
timestamp 1698431365
transform 1 0 18592 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_158
timestamp 1698431365
transform 1 0 19040 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_160
timestamp 1698431365
transform 1 0 19264 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_192
timestamp 1698431365
transform 1 0 22848 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_198
timestamp 1698431365
transform 1 0 23520 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_202
timestamp 1698431365
transform 1 0 23968 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_206
timestamp 1698431365
transform 1 0 24416 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_212
timestamp 1698431365
transform 1 0 25088 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_216
timestamp 1698431365
transform 1 0 25536 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_63_220
timestamp 1698431365
transform 1 0 25984 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_228
timestamp 1698431365
transform 1 0 26880 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_63_234
timestamp 1698431365
transform 1 0 27552 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_242
timestamp 1698431365
transform 1 0 28448 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_246
timestamp 1698431365
transform 1 0 28896 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_63_253
timestamp 1698431365
transform 1 0 29680 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_273
timestamp 1698431365
transform 1 0 31920 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_277
timestamp 1698431365
transform 1 0 32368 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_279
timestamp 1698431365
transform 1 0 32592 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_282
timestamp 1698431365
transform 1 0 32928 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_286
timestamp 1698431365
transform 1 0 33376 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_347
timestamp 1698431365
transform 1 0 40208 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_349
timestamp 1698431365
transform 1 0 40432 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_384
timestamp 1698431365
transform 1 0 44352 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_419
timestamp 1698431365
transform 1 0 48272 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_64_2
timestamp 1698431365
transform 1 0 1568 0 1 53312
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_34
timestamp 1698431365
transform 1 0 5152 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_64_37
timestamp 1698431365
transform 1 0 5488 0 1 53312
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_69
timestamp 1698431365
transform 1 0 9072 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_107
timestamp 1698431365
transform 1 0 13328 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_124
timestamp 1698431365
transform 1 0 15232 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_128
timestamp 1698431365
transform 1 0 15680 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_64_136
timestamp 1698431365
transform 1 0 16576 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_144
timestamp 1698431365
transform 1 0 17472 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_146
timestamp 1698431365
transform 1 0 17696 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_173
timestamp 1698431365
transform 1 0 20720 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_177
timestamp 1698431365
transform 1 0 21168 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_179
timestamp 1698431365
transform 1 0 21392 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_226
timestamp 1698431365
transform 1 0 26656 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_243
timestamp 1698431365
transform 1 0 28560 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_255
timestamp 1698431365
transform 1 0 29904 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_259
timestamp 1698431365
transform 1 0 30352 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_261
timestamp 1698431365
transform 1 0 30576 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_64_270
timestamp 1698431365
transform 1 0 31584 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_278
timestamp 1698431365
transform 1 0 32480 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_280
timestamp 1698431365
transform 1 0 32704 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_283
timestamp 1698431365
transform 1 0 33040 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_313
timestamp 1698431365
transform 1 0 36400 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_326
timestamp 1698431365
transform 1 0 37856 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_387
timestamp 1698431365
transform 1 0 44688 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_65_2
timestamp 1698431365
transform 1 0 1568 0 -1 54880
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_34
timestamp 1698431365
transform 1 0 5152 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_38
timestamp 1698431365
transform 1 0 5600 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_40
timestamp 1698431365
transform 1 0 5824 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_95
timestamp 1698431365
transform 1 0 11984 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_97
timestamp 1698431365
transform 1 0 12208 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_133
timestamp 1698431365
transform 1 0 16240 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_137
timestamp 1698431365
transform 1 0 16688 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_139
timestamp 1698431365
transform 1 0 16912 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_142
timestamp 1698431365
transform 1 0 17248 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_148
timestamp 1698431365
transform 1 0 17920 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_150
timestamp 1698431365
transform 1 0 18144 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_224
timestamp 1698431365
transform 1 0 26432 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_266
timestamp 1698431365
transform 1 0 31136 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_270
timestamp 1698431365
transform 1 0 31584 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_274
timestamp 1698431365
transform 1 0 32032 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_345
timestamp 1698431365
transform 1 0 39984 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_412
timestamp 1698431365
transform 1 0 47488 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_66_2
timestamp 1698431365
transform 1 0 1568 0 1 54880
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_34
timestamp 1698431365
transform 1 0 5152 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_66_37
timestamp 1698431365
transform 1 0 5488 0 1 54880
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_69
timestamp 1698431365
transform 1 0 9072 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_94
timestamp 1698431365
transform 1 0 11872 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_98
timestamp 1698431365
transform 1 0 12320 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_102
timestamp 1698431365
transform 1 0 12768 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_104
timestamp 1698431365
transform 1 0 12992 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_115
timestamp 1698431365
transform 1 0 14224 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_177
timestamp 1698431365
transform 1 0 21168 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_181
timestamp 1698431365
transform 1 0 21616 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_196
timestamp 1698431365
transform 1 0 23296 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_236
timestamp 1698431365
transform 1 0 27776 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_251
timestamp 1698431365
transform 1 0 29456 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_253
timestamp 1698431365
transform 1 0 29680 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_309
timestamp 1698431365
transform 1 0 35952 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_334
timestamp 1698431365
transform 1 0 38752 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_67_2
timestamp 1698431365
transform 1 0 1568 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_18
timestamp 1698431365
transform 1 0 3360 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_20
timestamp 1698431365
transform 1 0 3584 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_67_25
timestamp 1698431365
transform 1 0 4144 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_33
timestamp 1698431365
transform 1 0 5040 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_67_40
timestamp 1698431365
transform 1 0 5824 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_48
timestamp 1698431365
transform 1 0 6720 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_67_53
timestamp 1698431365
transform 1 0 7280 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_61
timestamp 1698431365
transform 1 0 8176 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_67
timestamp 1698431365
transform 1 0 8848 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_70
timestamp 1698431365
transform 1 0 9184 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_74
timestamp 1698431365
transform 1 0 9632 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_76
timestamp 1698431365
transform 1 0 9856 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_67_81
timestamp 1698431365
transform 1 0 10416 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_89
timestamp 1698431365
transform 1 0 11312 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_95
timestamp 1698431365
transform 1 0 11984 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_97
timestamp 1698431365
transform 1 0 12208 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_104
timestamp 1698431365
transform 1 0 12992 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_167
timestamp 1698431365
transform 1 0 20048 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_169
timestamp 1698431365
transform 1 0 20272 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_172
timestamp 1698431365
transform 1 0 20608 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_174
timestamp 1698431365
transform 1 0 20832 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_201
timestamp 1698431365
transform 1 0 23856 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_203
timestamp 1698431365
transform 1 0 24080 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_236
timestamp 1698431365
transform 1 0 27776 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_244
timestamp 1698431365
transform 1 0 28672 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_303
timestamp 1698431365
transform 1 0 35280 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_305
timestamp 1698431365
transform 1 0 35504 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_337
timestamp 1698431365
transform 1 0 39088 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_339
timestamp 1698431365
transform 1 0 39312 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input1
timestamp 1698431365
transform -1 0 48384 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input2
timestamp 1698431365
transform 1 0 43792 0 1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input3
timestamp 1698431365
transform -1 0 48384 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input4
timestamp 1698431365
transform -1 0 48384 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input5
timestamp 1698431365
transform -1 0 48384 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input6
timestamp 1698431365
transform -1 0 48384 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input7
timestamp 1698431365
transform -1 0 48384 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input8
timestamp 1698431365
transform -1 0 48384 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input9
timestamp 1698431365
transform -1 0 48384 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input10
timestamp 1698431365
transform -1 0 48384 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input11
timestamp 1698431365
transform 1 0 1568 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input12
timestamp 1698431365
transform 1 0 1568 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output13
timestamp 1698431365
transform 1 0 19376 0 -1 53312
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output14
timestamp 1698431365
transform 1 0 20944 0 -1 56448
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output15
timestamp 1698431365
transform -1 0 27328 0 -1 56448
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output16
timestamp 1698431365
transform -1 0 31808 0 -1 56448
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output17
timestamp 1698431365
transform 1 0 33040 0 1 54880
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output18
timestamp 1698431365
transform 1 0 33488 0 1 53312
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output19
timestamp 1698431365
transform -1 0 39088 0 -1 54880
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output20
timestamp 1698431365
transform 1 0 39648 0 -1 56448
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output21
timestamp 1698431365
transform 1 0 43456 0 -1 56448
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output22
timestamp 1698431365
transform 1 0 40768 0 -1 53312
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output23
timestamp 1698431365
transform 1 0 41552 0 1 53312
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output24
timestamp 1698431365
transform 1 0 44576 0 -1 54880
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output25
timestamp 1698431365
transform 1 0 44464 0 -1 53312
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output26
timestamp 1698431365
transform 1 0 45472 0 1 51744
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output27
timestamp 1698431365
transform -1 0 16576 0 -1 56448
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output28
timestamp 1698431365
transform 1 0 17808 0 1 53312
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_68 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1698431365
transform -1 0 48608 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_69
timestamp 1698431365
transform 1 0 1344 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1698431365
transform -1 0 48608 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_70
timestamp 1698431365
transform 1 0 1344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1698431365
transform -1 0 48608 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_71
timestamp 1698431365
transform 1 0 1344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1698431365
transform -1 0 48608 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_72
timestamp 1698431365
transform 1 0 1344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1698431365
transform -1 0 48608 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_73
timestamp 1698431365
transform 1 0 1344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1698431365
transform -1 0 48608 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_74
timestamp 1698431365
transform 1 0 1344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1698431365
transform -1 0 48608 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_75
timestamp 1698431365
transform 1 0 1344 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1698431365
transform -1 0 48608 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_76
timestamp 1698431365
transform 1 0 1344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1698431365
transform -1 0 48608 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_77
timestamp 1698431365
transform 1 0 1344 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1698431365
transform -1 0 48608 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_78
timestamp 1698431365
transform 1 0 1344 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1698431365
transform -1 0 48608 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_79
timestamp 1698431365
transform 1 0 1344 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1698431365
transform -1 0 48608 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_80
timestamp 1698431365
transform 1 0 1344 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1698431365
transform -1 0 48608 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_81
timestamp 1698431365
transform 1 0 1344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1698431365
transform -1 0 48608 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_82
timestamp 1698431365
transform 1 0 1344 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1698431365
transform -1 0 48608 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_83
timestamp 1698431365
transform 1 0 1344 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1698431365
transform -1 0 48608 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Left_84
timestamp 1698431365
transform 1 0 1344 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1698431365
transform -1 0 48608 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Left_85
timestamp 1698431365
transform 1 0 1344 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Right_17
timestamp 1698431365
transform -1 0 48608 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Left_86
timestamp 1698431365
transform 1 0 1344 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Right_18
timestamp 1698431365
transform -1 0 48608 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Left_87
timestamp 1698431365
transform 1 0 1344 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Right_19
timestamp 1698431365
transform -1 0 48608 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Left_88
timestamp 1698431365
transform 1 0 1344 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Right_20
timestamp 1698431365
transform -1 0 48608 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Left_89
timestamp 1698431365
transform 1 0 1344 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Right_21
timestamp 1698431365
transform -1 0 48608 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Left_90
timestamp 1698431365
transform 1 0 1344 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Right_22
timestamp 1698431365
transform -1 0 48608 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Left_91
timestamp 1698431365
transform 1 0 1344 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Right_23
timestamp 1698431365
transform -1 0 48608 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Left_92
timestamp 1698431365
transform 1 0 1344 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Right_24
timestamp 1698431365
transform -1 0 48608 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Left_93
timestamp 1698431365
transform 1 0 1344 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Right_25
timestamp 1698431365
transform -1 0 48608 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Left_94
timestamp 1698431365
transform 1 0 1344 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Right_26
timestamp 1698431365
transform -1 0 48608 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Left_95
timestamp 1698431365
transform 1 0 1344 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Right_27
timestamp 1698431365
transform -1 0 48608 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Left_96
timestamp 1698431365
transform 1 0 1344 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Right_28
timestamp 1698431365
transform -1 0 48608 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Left_97
timestamp 1698431365
transform 1 0 1344 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Right_29
timestamp 1698431365
transform -1 0 48608 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Left_98
timestamp 1698431365
transform 1 0 1344 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Right_30
timestamp 1698431365
transform -1 0 48608 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Left_99
timestamp 1698431365
transform 1 0 1344 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Right_31
timestamp 1698431365
transform -1 0 48608 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Left_100
timestamp 1698431365
transform 1 0 1344 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Right_32
timestamp 1698431365
transform -1 0 48608 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Left_101
timestamp 1698431365
transform 1 0 1344 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Right_33
timestamp 1698431365
transform -1 0 48608 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Left_102
timestamp 1698431365
transform 1 0 1344 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Right_34
timestamp 1698431365
transform -1 0 48608 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Left_103
timestamp 1698431365
transform 1 0 1344 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Right_35
timestamp 1698431365
transform -1 0 48608 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Left_104
timestamp 1698431365
transform 1 0 1344 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Right_36
timestamp 1698431365
transform -1 0 48608 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Left_105
timestamp 1698431365
transform 1 0 1344 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Right_37
timestamp 1698431365
transform -1 0 48608 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Left_106
timestamp 1698431365
transform 1 0 1344 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Right_38
timestamp 1698431365
transform -1 0 48608 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Left_107
timestamp 1698431365
transform 1 0 1344 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Right_39
timestamp 1698431365
transform -1 0 48608 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Left_108
timestamp 1698431365
transform 1 0 1344 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Right_40
timestamp 1698431365
transform -1 0 48608 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Left_109
timestamp 1698431365
transform 1 0 1344 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Right_41
timestamp 1698431365
transform -1 0 48608 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Left_110
timestamp 1698431365
transform 1 0 1344 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Right_42
timestamp 1698431365
transform -1 0 48608 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Left_111
timestamp 1698431365
transform 1 0 1344 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Right_43
timestamp 1698431365
transform -1 0 48608 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Left_112
timestamp 1698431365
transform 1 0 1344 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Right_44
timestamp 1698431365
transform -1 0 48608 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_45_Left_113
timestamp 1698431365
transform 1 0 1344 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_45_Right_45
timestamp 1698431365
transform -1 0 48608 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_46_Left_114
timestamp 1698431365
transform 1 0 1344 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_46_Right_46
timestamp 1698431365
transform -1 0 48608 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_47_Left_115
timestamp 1698431365
transform 1 0 1344 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_47_Right_47
timestamp 1698431365
transform -1 0 48608 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_48_Left_116
timestamp 1698431365
transform 1 0 1344 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_48_Right_48
timestamp 1698431365
transform -1 0 48608 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_49_Left_117
timestamp 1698431365
transform 1 0 1344 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_49_Right_49
timestamp 1698431365
transform -1 0 48608 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_50_Left_118
timestamp 1698431365
transform 1 0 1344 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_50_Right_50
timestamp 1698431365
transform -1 0 48608 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_51_Left_119
timestamp 1698431365
transform 1 0 1344 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_51_Right_51
timestamp 1698431365
transform -1 0 48608 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_52_Left_120
timestamp 1698431365
transform 1 0 1344 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_52_Right_52
timestamp 1698431365
transform -1 0 48608 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_53_Left_121
timestamp 1698431365
transform 1 0 1344 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_53_Right_53
timestamp 1698431365
transform -1 0 48608 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_54_Left_122
timestamp 1698431365
transform 1 0 1344 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_54_Right_54
timestamp 1698431365
transform -1 0 48608 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_55_Left_123
timestamp 1698431365
transform 1 0 1344 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_55_Right_55
timestamp 1698431365
transform -1 0 48608 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_56_Left_124
timestamp 1698431365
transform 1 0 1344 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_56_Right_56
timestamp 1698431365
transform -1 0 48608 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_57_Left_125
timestamp 1698431365
transform 1 0 1344 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_57_Right_57
timestamp 1698431365
transform -1 0 48608 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_58_Left_126
timestamp 1698431365
transform 1 0 1344 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_58_Right_58
timestamp 1698431365
transform -1 0 48608 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_59_Left_127
timestamp 1698431365
transform 1 0 1344 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_59_Right_59
timestamp 1698431365
transform -1 0 48608 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_60_Left_128
timestamp 1698431365
transform 1 0 1344 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_60_Right_60
timestamp 1698431365
transform -1 0 48608 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_61_Left_129
timestamp 1698431365
transform 1 0 1344 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_61_Right_61
timestamp 1698431365
transform -1 0 48608 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_62_Left_130
timestamp 1698431365
transform 1 0 1344 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_62_Right_62
timestamp 1698431365
transform -1 0 48608 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_63_Left_131
timestamp 1698431365
transform 1 0 1344 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_63_Right_63
timestamp 1698431365
transform -1 0 48608 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_64_Left_132
timestamp 1698431365
transform 1 0 1344 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_64_Right_64
timestamp 1698431365
transform -1 0 48608 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_65_Left_133
timestamp 1698431365
transform 1 0 1344 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_65_Right_65
timestamp 1698431365
transform -1 0 48608 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_66_Left_134
timestamp 1698431365
transform 1 0 1344 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_66_Right_66
timestamp 1698431365
transform -1 0 48608 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_67_Left_135
timestamp 1698431365
transform 1 0 1344 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_67_Right_67
timestamp 1698431365
transform -1 0 48608 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  rebuffer1
timestamp 1698431365
transform 1 0 47712 0 -1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  rebuffer2
timestamp 1698431365
transform -1 0 11312 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  rebuffer3
timestamp 1698431365
transform 1 0 8512 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  rebuffer4
timestamp 1698431365
transform -1 0 16128 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  rebuffer5
timestamp 1698431365
transform -1 0 16352 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  rebuffer6
timestamp 1698431365
transform 1 0 11424 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  rebuffer7
timestamp 1698431365
transform -1 0 15008 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  rebuffer8
timestamp 1698431365
transform -1 0 15680 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  rebuffer9
timestamp 1698431365
transform 1 0 12096 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  rebuffer10
timestamp 1698431365
transform 1 0 30912 0 1 50176
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  rebuffer11
timestamp 1698431365
transform 1 0 30464 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  rebuffer12
timestamp 1698431365
transform -1 0 45360 0 1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  rebuffer13
timestamp 1698431365
transform -1 0 9408 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  rebuffer14
timestamp 1698431365
transform -1 0 8848 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  rebuffer15
timestamp 1698431365
transform -1 0 13888 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  rebuffer16
timestamp 1698431365
transform 1 0 11872 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  rebuffer17
timestamp 1698431365
transform -1 0 7952 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  rebuffer18
timestamp 1698431365
transform -1 0 3920 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  rebuffer19
timestamp 1698431365
transform 1 0 21280 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  rebuffer20
timestamp 1698431365
transform 1 0 9408 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  rebuffer21
timestamp 1698431365
transform -1 0 48272 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  rebuffer22
timestamp 1698431365
transform -1 0 29904 0 -1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  rebuffer23
timestamp 1698431365
transform 1 0 11760 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  rebuffer24
timestamp 1698431365
transform -1 0 28448 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  rebuffer25
timestamp 1698431365
transform -1 0 29680 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  rebuffer26
timestamp 1698431365
transform -1 0 30352 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  rebuffer27
timestamp 1698431365
transform -1 0 13888 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  rebuffer28
timestamp 1698431365
transform 1 0 11536 0 1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  rebuffer29
timestamp 1698431365
transform 1 0 12320 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  rebuffer30
timestamp 1698431365
transform 1 0 29456 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_136 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5152 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_137
timestamp 1698431365
transform 1 0 8960 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_138
timestamp 1698431365
transform 1 0 12768 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_139
timestamp 1698431365
transform 1 0 16576 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_140
timestamp 1698431365
transform 1 0 20384 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_141
timestamp 1698431365
transform 1 0 24192 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_142
timestamp 1698431365
transform 1 0 28000 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_143
timestamp 1698431365
transform 1 0 31808 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_144
timestamp 1698431365
transform 1 0 35616 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_145
timestamp 1698431365
transform 1 0 39424 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_146
timestamp 1698431365
transform 1 0 43232 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_147
timestamp 1698431365
transform 1 0 47040 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_148
timestamp 1698431365
transform 1 0 9184 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_149
timestamp 1698431365
transform 1 0 17024 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_150
timestamp 1698431365
transform 1 0 24864 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_151
timestamp 1698431365
transform 1 0 32704 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_152
timestamp 1698431365
transform 1 0 40544 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_153
timestamp 1698431365
transform 1 0 5264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_154
timestamp 1698431365
transform 1 0 13104 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_155
timestamp 1698431365
transform 1 0 20944 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_156
timestamp 1698431365
transform 1 0 28784 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_157
timestamp 1698431365
transform 1 0 36624 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_158
timestamp 1698431365
transform 1 0 44464 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_159
timestamp 1698431365
transform 1 0 9184 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_160
timestamp 1698431365
transform 1 0 17024 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_161
timestamp 1698431365
transform 1 0 24864 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_162
timestamp 1698431365
transform 1 0 32704 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_163
timestamp 1698431365
transform 1 0 40544 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_164
timestamp 1698431365
transform 1 0 5264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_165
timestamp 1698431365
transform 1 0 13104 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_166
timestamp 1698431365
transform 1 0 20944 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_167
timestamp 1698431365
transform 1 0 28784 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_168
timestamp 1698431365
transform 1 0 36624 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_169
timestamp 1698431365
transform 1 0 44464 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_170
timestamp 1698431365
transform 1 0 9184 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_171
timestamp 1698431365
transform 1 0 17024 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_172
timestamp 1698431365
transform 1 0 24864 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_173
timestamp 1698431365
transform 1 0 32704 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_174
timestamp 1698431365
transform 1 0 40544 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_175
timestamp 1698431365
transform 1 0 5264 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_176
timestamp 1698431365
transform 1 0 13104 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_177
timestamp 1698431365
transform 1 0 20944 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_178
timestamp 1698431365
transform 1 0 28784 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_179
timestamp 1698431365
transform 1 0 36624 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_180
timestamp 1698431365
transform 1 0 44464 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_181
timestamp 1698431365
transform 1 0 9184 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_182
timestamp 1698431365
transform 1 0 17024 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_183
timestamp 1698431365
transform 1 0 24864 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_184
timestamp 1698431365
transform 1 0 32704 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_185
timestamp 1698431365
transform 1 0 40544 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_186
timestamp 1698431365
transform 1 0 5264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_187
timestamp 1698431365
transform 1 0 13104 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_188
timestamp 1698431365
transform 1 0 20944 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_189
timestamp 1698431365
transform 1 0 28784 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_190
timestamp 1698431365
transform 1 0 36624 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_191
timestamp 1698431365
transform 1 0 44464 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_192
timestamp 1698431365
transform 1 0 9184 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_193
timestamp 1698431365
transform 1 0 17024 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_194
timestamp 1698431365
transform 1 0 24864 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_195
timestamp 1698431365
transform 1 0 32704 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_196
timestamp 1698431365
transform 1 0 40544 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_197
timestamp 1698431365
transform 1 0 5264 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_198
timestamp 1698431365
transform 1 0 13104 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_199
timestamp 1698431365
transform 1 0 20944 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_200
timestamp 1698431365
transform 1 0 28784 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_201
timestamp 1698431365
transform 1 0 36624 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_202
timestamp 1698431365
transform 1 0 44464 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_203
timestamp 1698431365
transform 1 0 9184 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_204
timestamp 1698431365
transform 1 0 17024 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_205
timestamp 1698431365
transform 1 0 24864 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_206
timestamp 1698431365
transform 1 0 32704 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_207
timestamp 1698431365
transform 1 0 40544 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_208
timestamp 1698431365
transform 1 0 5264 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_209
timestamp 1698431365
transform 1 0 13104 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_210
timestamp 1698431365
transform 1 0 20944 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_211
timestamp 1698431365
transform 1 0 28784 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_212
timestamp 1698431365
transform 1 0 36624 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_213
timestamp 1698431365
transform 1 0 44464 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_214
timestamp 1698431365
transform 1 0 9184 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_215
timestamp 1698431365
transform 1 0 17024 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_216
timestamp 1698431365
transform 1 0 24864 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_217
timestamp 1698431365
transform 1 0 32704 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_218
timestamp 1698431365
transform 1 0 40544 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_219
timestamp 1698431365
transform 1 0 5264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_220
timestamp 1698431365
transform 1 0 13104 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_221
timestamp 1698431365
transform 1 0 20944 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_222
timestamp 1698431365
transform 1 0 28784 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_223
timestamp 1698431365
transform 1 0 36624 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_224
timestamp 1698431365
transform 1 0 44464 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_225
timestamp 1698431365
transform 1 0 9184 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_226
timestamp 1698431365
transform 1 0 17024 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_227
timestamp 1698431365
transform 1 0 24864 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_228
timestamp 1698431365
transform 1 0 32704 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_229
timestamp 1698431365
transform 1 0 40544 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_230
timestamp 1698431365
transform 1 0 5264 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_231
timestamp 1698431365
transform 1 0 13104 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_232
timestamp 1698431365
transform 1 0 20944 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_233
timestamp 1698431365
transform 1 0 28784 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_234
timestamp 1698431365
transform 1 0 36624 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_235
timestamp 1698431365
transform 1 0 44464 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_236
timestamp 1698431365
transform 1 0 9184 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_237
timestamp 1698431365
transform 1 0 17024 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_238
timestamp 1698431365
transform 1 0 24864 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_239
timestamp 1698431365
transform 1 0 32704 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_240
timestamp 1698431365
transform 1 0 40544 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_241
timestamp 1698431365
transform 1 0 5264 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_242
timestamp 1698431365
transform 1 0 13104 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_243
timestamp 1698431365
transform 1 0 20944 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_244
timestamp 1698431365
transform 1 0 28784 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_245
timestamp 1698431365
transform 1 0 36624 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_246
timestamp 1698431365
transform 1 0 44464 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_247
timestamp 1698431365
transform 1 0 9184 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_248
timestamp 1698431365
transform 1 0 17024 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_249
timestamp 1698431365
transform 1 0 24864 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_250
timestamp 1698431365
transform 1 0 32704 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_251
timestamp 1698431365
transform 1 0 40544 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_252
timestamp 1698431365
transform 1 0 5264 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_253
timestamp 1698431365
transform 1 0 13104 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_254
timestamp 1698431365
transform 1 0 20944 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_255
timestamp 1698431365
transform 1 0 28784 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_256
timestamp 1698431365
transform 1 0 36624 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_257
timestamp 1698431365
transform 1 0 44464 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_258
timestamp 1698431365
transform 1 0 9184 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_259
timestamp 1698431365
transform 1 0 17024 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_260
timestamp 1698431365
transform 1 0 24864 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_261
timestamp 1698431365
transform 1 0 32704 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_262
timestamp 1698431365
transform 1 0 40544 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_263
timestamp 1698431365
transform 1 0 5264 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_264
timestamp 1698431365
transform 1 0 13104 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_265
timestamp 1698431365
transform 1 0 20944 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_266
timestamp 1698431365
transform 1 0 28784 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_267
timestamp 1698431365
transform 1 0 36624 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_268
timestamp 1698431365
transform 1 0 44464 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_269
timestamp 1698431365
transform 1 0 9184 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_270
timestamp 1698431365
transform 1 0 17024 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_271
timestamp 1698431365
transform 1 0 24864 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_272
timestamp 1698431365
transform 1 0 32704 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_273
timestamp 1698431365
transform 1 0 40544 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_274
timestamp 1698431365
transform 1 0 5264 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_275
timestamp 1698431365
transform 1 0 13104 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_276
timestamp 1698431365
transform 1 0 20944 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_277
timestamp 1698431365
transform 1 0 28784 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_278
timestamp 1698431365
transform 1 0 36624 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_279
timestamp 1698431365
transform 1 0 44464 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_280
timestamp 1698431365
transform 1 0 9184 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_281
timestamp 1698431365
transform 1 0 17024 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_282
timestamp 1698431365
transform 1 0 24864 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_283
timestamp 1698431365
transform 1 0 32704 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_284
timestamp 1698431365
transform 1 0 40544 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_285
timestamp 1698431365
transform 1 0 5264 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_286
timestamp 1698431365
transform 1 0 13104 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_287
timestamp 1698431365
transform 1 0 20944 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_288
timestamp 1698431365
transform 1 0 28784 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_289
timestamp 1698431365
transform 1 0 36624 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_290
timestamp 1698431365
transform 1 0 44464 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_291
timestamp 1698431365
transform 1 0 9184 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_292
timestamp 1698431365
transform 1 0 17024 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_293
timestamp 1698431365
transform 1 0 24864 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_294
timestamp 1698431365
transform 1 0 32704 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_295
timestamp 1698431365
transform 1 0 40544 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_296
timestamp 1698431365
transform 1 0 5264 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_297
timestamp 1698431365
transform 1 0 13104 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_298
timestamp 1698431365
transform 1 0 20944 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_299
timestamp 1698431365
transform 1 0 28784 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_300
timestamp 1698431365
transform 1 0 36624 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_301
timestamp 1698431365
transform 1 0 44464 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_302
timestamp 1698431365
transform 1 0 9184 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_303
timestamp 1698431365
transform 1 0 17024 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_304
timestamp 1698431365
transform 1 0 24864 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_305
timestamp 1698431365
transform 1 0 32704 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_306
timestamp 1698431365
transform 1 0 40544 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_307
timestamp 1698431365
transform 1 0 5264 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_308
timestamp 1698431365
transform 1 0 13104 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_309
timestamp 1698431365
transform 1 0 20944 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_310
timestamp 1698431365
transform 1 0 28784 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_311
timestamp 1698431365
transform 1 0 36624 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_312
timestamp 1698431365
transform 1 0 44464 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_313
timestamp 1698431365
transform 1 0 9184 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_314
timestamp 1698431365
transform 1 0 17024 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_315
timestamp 1698431365
transform 1 0 24864 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_316
timestamp 1698431365
transform 1 0 32704 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_317
timestamp 1698431365
transform 1 0 40544 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_318
timestamp 1698431365
transform 1 0 5264 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_319
timestamp 1698431365
transform 1 0 13104 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_320
timestamp 1698431365
transform 1 0 20944 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_321
timestamp 1698431365
transform 1 0 28784 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_322
timestamp 1698431365
transform 1 0 36624 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_323
timestamp 1698431365
transform 1 0 44464 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_324
timestamp 1698431365
transform 1 0 9184 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_325
timestamp 1698431365
transform 1 0 17024 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_326
timestamp 1698431365
transform 1 0 24864 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_327
timestamp 1698431365
transform 1 0 32704 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_328
timestamp 1698431365
transform 1 0 40544 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_329
timestamp 1698431365
transform 1 0 5264 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_330
timestamp 1698431365
transform 1 0 13104 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_331
timestamp 1698431365
transform 1 0 20944 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_332
timestamp 1698431365
transform 1 0 28784 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_333
timestamp 1698431365
transform 1 0 36624 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_334
timestamp 1698431365
transform 1 0 44464 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_335
timestamp 1698431365
transform 1 0 9184 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_336
timestamp 1698431365
transform 1 0 17024 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_337
timestamp 1698431365
transform 1 0 24864 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_338
timestamp 1698431365
transform 1 0 32704 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_339
timestamp 1698431365
transform 1 0 40544 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_340
timestamp 1698431365
transform 1 0 5264 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_341
timestamp 1698431365
transform 1 0 13104 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_342
timestamp 1698431365
transform 1 0 20944 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_343
timestamp 1698431365
transform 1 0 28784 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_344
timestamp 1698431365
transform 1 0 36624 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_345
timestamp 1698431365
transform 1 0 44464 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_346
timestamp 1698431365
transform 1 0 9184 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_347
timestamp 1698431365
transform 1 0 17024 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_348
timestamp 1698431365
transform 1 0 24864 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_349
timestamp 1698431365
transform 1 0 32704 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_350
timestamp 1698431365
transform 1 0 40544 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_351
timestamp 1698431365
transform 1 0 5264 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_352
timestamp 1698431365
transform 1 0 13104 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_353
timestamp 1698431365
transform 1 0 20944 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_354
timestamp 1698431365
transform 1 0 28784 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_355
timestamp 1698431365
transform 1 0 36624 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_356
timestamp 1698431365
transform 1 0 44464 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_357
timestamp 1698431365
transform 1 0 9184 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_358
timestamp 1698431365
transform 1 0 17024 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_359
timestamp 1698431365
transform 1 0 24864 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_360
timestamp 1698431365
transform 1 0 32704 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_361
timestamp 1698431365
transform 1 0 40544 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_362
timestamp 1698431365
transform 1 0 5264 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_363
timestamp 1698431365
transform 1 0 13104 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_364
timestamp 1698431365
transform 1 0 20944 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_365
timestamp 1698431365
transform 1 0 28784 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_366
timestamp 1698431365
transform 1 0 36624 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_367
timestamp 1698431365
transform 1 0 44464 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_368
timestamp 1698431365
transform 1 0 9184 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_369
timestamp 1698431365
transform 1 0 17024 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_370
timestamp 1698431365
transform 1 0 24864 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_371
timestamp 1698431365
transform 1 0 32704 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_372
timestamp 1698431365
transform 1 0 40544 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_373
timestamp 1698431365
transform 1 0 5264 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_374
timestamp 1698431365
transform 1 0 13104 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_375
timestamp 1698431365
transform 1 0 20944 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_376
timestamp 1698431365
transform 1 0 28784 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_377
timestamp 1698431365
transform 1 0 36624 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_378
timestamp 1698431365
transform 1 0 44464 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_379
timestamp 1698431365
transform 1 0 9184 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_380
timestamp 1698431365
transform 1 0 17024 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_381
timestamp 1698431365
transform 1 0 24864 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_382
timestamp 1698431365
transform 1 0 32704 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_383
timestamp 1698431365
transform 1 0 40544 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_384
timestamp 1698431365
transform 1 0 5264 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_385
timestamp 1698431365
transform 1 0 13104 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_386
timestamp 1698431365
transform 1 0 20944 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_387
timestamp 1698431365
transform 1 0 28784 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_388
timestamp 1698431365
transform 1 0 36624 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_389
timestamp 1698431365
transform 1 0 44464 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_390
timestamp 1698431365
transform 1 0 9184 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_391
timestamp 1698431365
transform 1 0 17024 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_392
timestamp 1698431365
transform 1 0 24864 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_393
timestamp 1698431365
transform 1 0 32704 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_394
timestamp 1698431365
transform 1 0 40544 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_395
timestamp 1698431365
transform 1 0 5264 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_396
timestamp 1698431365
transform 1 0 13104 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_397
timestamp 1698431365
transform 1 0 20944 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_398
timestamp 1698431365
transform 1 0 28784 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_399
timestamp 1698431365
transform 1 0 36624 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_400
timestamp 1698431365
transform 1 0 44464 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_401
timestamp 1698431365
transform 1 0 9184 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_402
timestamp 1698431365
transform 1 0 17024 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_403
timestamp 1698431365
transform 1 0 24864 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_404
timestamp 1698431365
transform 1 0 32704 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_405
timestamp 1698431365
transform 1 0 40544 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_406
timestamp 1698431365
transform 1 0 5264 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_407
timestamp 1698431365
transform 1 0 13104 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_408
timestamp 1698431365
transform 1 0 20944 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_409
timestamp 1698431365
transform 1 0 28784 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_410
timestamp 1698431365
transform 1 0 36624 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_411
timestamp 1698431365
transform 1 0 44464 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_412
timestamp 1698431365
transform 1 0 9184 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_413
timestamp 1698431365
transform 1 0 17024 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_414
timestamp 1698431365
transform 1 0 24864 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_415
timestamp 1698431365
transform 1 0 32704 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_416
timestamp 1698431365
transform 1 0 40544 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_417
timestamp 1698431365
transform 1 0 5264 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_418
timestamp 1698431365
transform 1 0 13104 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_419
timestamp 1698431365
transform 1 0 20944 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_420
timestamp 1698431365
transform 1 0 28784 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_421
timestamp 1698431365
transform 1 0 36624 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_422
timestamp 1698431365
transform 1 0 44464 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_423
timestamp 1698431365
transform 1 0 9184 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_424
timestamp 1698431365
transform 1 0 17024 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_425
timestamp 1698431365
transform 1 0 24864 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_426
timestamp 1698431365
transform 1 0 32704 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_427
timestamp 1698431365
transform 1 0 40544 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_428
timestamp 1698431365
transform 1 0 5264 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_429
timestamp 1698431365
transform 1 0 13104 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_430
timestamp 1698431365
transform 1 0 20944 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_431
timestamp 1698431365
transform 1 0 28784 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_432
timestamp 1698431365
transform 1 0 36624 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_433
timestamp 1698431365
transform 1 0 44464 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_434
timestamp 1698431365
transform 1 0 9184 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_435
timestamp 1698431365
transform 1 0 17024 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_436
timestamp 1698431365
transform 1 0 24864 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_437
timestamp 1698431365
transform 1 0 32704 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_438
timestamp 1698431365
transform 1 0 40544 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_439
timestamp 1698431365
transform 1 0 5264 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_440
timestamp 1698431365
transform 1 0 13104 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_441
timestamp 1698431365
transform 1 0 20944 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_442
timestamp 1698431365
transform 1 0 28784 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_443
timestamp 1698431365
transform 1 0 36624 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_444
timestamp 1698431365
transform 1 0 44464 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_445
timestamp 1698431365
transform 1 0 9184 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_446
timestamp 1698431365
transform 1 0 17024 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_447
timestamp 1698431365
transform 1 0 24864 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_448
timestamp 1698431365
transform 1 0 32704 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_449
timestamp 1698431365
transform 1 0 40544 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_450
timestamp 1698431365
transform 1 0 5264 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_451
timestamp 1698431365
transform 1 0 13104 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_452
timestamp 1698431365
transform 1 0 20944 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_453
timestamp 1698431365
transform 1 0 28784 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_454
timestamp 1698431365
transform 1 0 36624 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_455
timestamp 1698431365
transform 1 0 44464 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_456
timestamp 1698431365
transform 1 0 9184 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_457
timestamp 1698431365
transform 1 0 17024 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_458
timestamp 1698431365
transform 1 0 24864 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_459
timestamp 1698431365
transform 1 0 32704 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_460
timestamp 1698431365
transform 1 0 40544 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_461
timestamp 1698431365
transform 1 0 5264 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_462
timestamp 1698431365
transform 1 0 13104 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_463
timestamp 1698431365
transform 1 0 20944 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_464
timestamp 1698431365
transform 1 0 28784 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_465
timestamp 1698431365
transform 1 0 36624 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_466
timestamp 1698431365
transform 1 0 44464 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_467
timestamp 1698431365
transform 1 0 9184 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_468
timestamp 1698431365
transform 1 0 17024 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_469
timestamp 1698431365
transform 1 0 24864 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_470
timestamp 1698431365
transform 1 0 32704 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_471
timestamp 1698431365
transform 1 0 40544 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_472
timestamp 1698431365
transform 1 0 5264 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_473
timestamp 1698431365
transform 1 0 13104 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_474
timestamp 1698431365
transform 1 0 20944 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_475
timestamp 1698431365
transform 1 0 28784 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_476
timestamp 1698431365
transform 1 0 36624 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_477
timestamp 1698431365
transform 1 0 44464 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_478
timestamp 1698431365
transform 1 0 9184 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_479
timestamp 1698431365
transform 1 0 17024 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_480
timestamp 1698431365
transform 1 0 24864 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_481
timestamp 1698431365
transform 1 0 32704 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_482
timestamp 1698431365
transform 1 0 40544 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_483
timestamp 1698431365
transform 1 0 5264 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_484
timestamp 1698431365
transform 1 0 13104 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_485
timestamp 1698431365
transform 1 0 20944 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_486
timestamp 1698431365
transform 1 0 28784 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_487
timestamp 1698431365
transform 1 0 36624 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_488
timestamp 1698431365
transform 1 0 44464 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_489
timestamp 1698431365
transform 1 0 9184 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_490
timestamp 1698431365
transform 1 0 17024 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_491
timestamp 1698431365
transform 1 0 24864 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_492
timestamp 1698431365
transform 1 0 32704 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_493
timestamp 1698431365
transform 1 0 40544 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_494
timestamp 1698431365
transform 1 0 5264 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_495
timestamp 1698431365
transform 1 0 13104 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_496
timestamp 1698431365
transform 1 0 20944 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_497
timestamp 1698431365
transform 1 0 28784 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_498
timestamp 1698431365
transform 1 0 36624 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_499
timestamp 1698431365
transform 1 0 44464 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_500
timestamp 1698431365
transform 1 0 9184 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_501
timestamp 1698431365
transform 1 0 17024 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_502
timestamp 1698431365
transform 1 0 24864 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_503
timestamp 1698431365
transform 1 0 32704 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_504
timestamp 1698431365
transform 1 0 40544 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_505
timestamp 1698431365
transform 1 0 5264 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_506
timestamp 1698431365
transform 1 0 13104 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_507
timestamp 1698431365
transform 1 0 20944 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_508
timestamp 1698431365
transform 1 0 28784 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_509
timestamp 1698431365
transform 1 0 36624 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_510
timestamp 1698431365
transform 1 0 44464 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_511
timestamp 1698431365
transform 1 0 5152 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_512
timestamp 1698431365
transform 1 0 8960 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_513
timestamp 1698431365
transform 1 0 12768 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_514
timestamp 1698431365
transform 1 0 16576 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_515
timestamp 1698431365
transform 1 0 20384 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_516
timestamp 1698431365
transform 1 0 24192 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_517
timestamp 1698431365
transform 1 0 28000 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_518
timestamp 1698431365
transform 1 0 31808 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_519
timestamp 1698431365
transform 1 0 35616 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_520
timestamp 1698431365
transform 1 0 39424 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_521
timestamp 1698431365
transform 1 0 43232 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_522
timestamp 1698431365
transform 1 0 47040 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_sn76489_29 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 4144 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_sn76489_30
timestamp 1698431365
transform -1 0 5824 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_sn76489_31
timestamp 1698431365
transform -1 0 7280 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_sn76489_32
timestamp 1698431365
transform -1 0 8848 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_sn76489_33
timestamp 1698431365
transform -1 0 10416 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_sn76489_34
timestamp 1698431365
transform -1 0 11984 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_sn76489_35
timestamp 1698431365
transform 1 0 12320 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_sn76489_36
timestamp 1698431365
transform 1 0 13216 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_sn76489_37
timestamp 1698431365
transform 1 0 23520 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_sn76489_38
timestamp 1698431365
transform -1 0 27776 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_sn76489_39
timestamp 1698431365
transform -1 0 28672 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wrapped_sn76489_40
timestamp 1698431365
transform -1 0 29456 0 1 54880
box -86 -86 534 870
<< labels >>
flabel metal3 s 49200 50176 50000 50288 0 FreeSans 448 0 0 0 custom_settings[0]
port 0 nsew signal input
flabel metal3 s 49200 56000 50000 56112 0 FreeSans 448 0 0 0 custom_settings[1]
port 1 nsew signal input
flabel metal3 s 49200 3584 50000 3696 0 FreeSans 448 0 0 0 io_in_1[0]
port 2 nsew signal input
flabel metal3 s 49200 9408 50000 9520 0 FreeSans 448 0 0 0 io_in_1[1]
port 3 nsew signal input
flabel metal3 s 49200 15232 50000 15344 0 FreeSans 448 0 0 0 io_in_1[2]
port 4 nsew signal input
flabel metal3 s 49200 21056 50000 21168 0 FreeSans 448 0 0 0 io_in_1[3]
port 5 nsew signal input
flabel metal3 s 49200 26880 50000 26992 0 FreeSans 448 0 0 0 io_in_1[4]
port 6 nsew signal input
flabel metal3 s 49200 32704 50000 32816 0 FreeSans 448 0 0 0 io_in_1[5]
port 7 nsew signal input
flabel metal3 s 49200 38528 50000 38640 0 FreeSans 448 0 0 0 io_in_1[6]
port 8 nsew signal input
flabel metal3 s 49200 44352 50000 44464 0 FreeSans 448 0 0 0 io_in_1[7]
port 9 nsew signal input
flabel metal3 s 0 49728 800 49840 0 FreeSans 448 0 0 0 io_in_2
port 10 nsew signal input
flabel metal2 s 3584 59200 3696 60000 0 FreeSans 448 90 0 0 io_out[0]
port 11 nsew signal tristate
flabel metal2 s 19264 59200 19376 60000 0 FreeSans 448 90 0 0 io_out[10]
port 12 nsew signal tristate
flabel metal2 s 20832 59200 20944 60000 0 FreeSans 448 90 0 0 io_out[11]
port 13 nsew signal tristate
flabel metal2 s 22400 59200 22512 60000 0 FreeSans 448 90 0 0 io_out[12]
port 14 nsew signal tristate
flabel metal2 s 23968 59200 24080 60000 0 FreeSans 448 90 0 0 io_out[13]
port 15 nsew signal tristate
flabel metal2 s 25536 59200 25648 60000 0 FreeSans 448 90 0 0 io_out[14]
port 16 nsew signal tristate
flabel metal2 s 27104 59200 27216 60000 0 FreeSans 448 90 0 0 io_out[15]
port 17 nsew signal tristate
flabel metal2 s 28672 59200 28784 60000 0 FreeSans 448 90 0 0 io_out[16]
port 18 nsew signal tristate
flabel metal2 s 30240 59200 30352 60000 0 FreeSans 448 90 0 0 io_out[17]
port 19 nsew signal tristate
flabel metal2 s 31808 59200 31920 60000 0 FreeSans 448 90 0 0 io_out[18]
port 20 nsew signal tristate
flabel metal2 s 33376 59200 33488 60000 0 FreeSans 448 90 0 0 io_out[19]
port 21 nsew signal tristate
flabel metal2 s 5152 59200 5264 60000 0 FreeSans 448 90 0 0 io_out[1]
port 22 nsew signal tristate
flabel metal2 s 34944 59200 35056 60000 0 FreeSans 448 90 0 0 io_out[20]
port 23 nsew signal tristate
flabel metal2 s 36512 59200 36624 60000 0 FreeSans 448 90 0 0 io_out[21]
port 24 nsew signal tristate
flabel metal2 s 38080 59200 38192 60000 0 FreeSans 448 90 0 0 io_out[22]
port 25 nsew signal tristate
flabel metal2 s 39648 59200 39760 60000 0 FreeSans 448 90 0 0 io_out[23]
port 26 nsew signal tristate
flabel metal2 s 41216 59200 41328 60000 0 FreeSans 448 90 0 0 io_out[24]
port 27 nsew signal tristate
flabel metal2 s 42784 59200 42896 60000 0 FreeSans 448 90 0 0 io_out[25]
port 28 nsew signal tristate
flabel metal2 s 44352 59200 44464 60000 0 FreeSans 448 90 0 0 io_out[26]
port 29 nsew signal tristate
flabel metal2 s 45920 59200 46032 60000 0 FreeSans 448 90 0 0 io_out[27]
port 30 nsew signal tristate
flabel metal2 s 6720 59200 6832 60000 0 FreeSans 448 90 0 0 io_out[2]
port 31 nsew signal tristate
flabel metal2 s 8288 59200 8400 60000 0 FreeSans 448 90 0 0 io_out[3]
port 32 nsew signal tristate
flabel metal2 s 9856 59200 9968 60000 0 FreeSans 448 90 0 0 io_out[4]
port 33 nsew signal tristate
flabel metal2 s 11424 59200 11536 60000 0 FreeSans 448 90 0 0 io_out[5]
port 34 nsew signal tristate
flabel metal2 s 12992 59200 13104 60000 0 FreeSans 448 90 0 0 io_out[6]
port 35 nsew signal tristate
flabel metal2 s 14560 59200 14672 60000 0 FreeSans 448 90 0 0 io_out[7]
port 36 nsew signal tristate
flabel metal2 s 16128 59200 16240 60000 0 FreeSans 448 90 0 0 io_out[8]
port 37 nsew signal tristate
flabel metal2 s 17696 59200 17808 60000 0 FreeSans 448 90 0 0 io_out[9]
port 38 nsew signal tristate
flabel metal3 s 0 29792 800 29904 0 FreeSans 448 0 0 0 rst_n
port 39 nsew signal input
flabel metal4 s 4448 3076 4768 56508 0 FreeSans 1280 90 0 0 vdd
port 40 nsew power bidirectional
flabel metal4 s 35168 3076 35488 56508 0 FreeSans 1280 90 0 0 vdd
port 40 nsew power bidirectional
flabel metal4 s 19808 3076 20128 56508 0 FreeSans 1280 90 0 0 vss
port 41 nsew ground bidirectional
flabel metal3 s 0 9856 800 9968 0 FreeSans 448 0 0 0 wb_clk_i
port 42 nsew signal input
rlabel metal1 24976 55664 24976 55664 0 vdd
rlabel metal1 24976 56448 24976 56448 0 vss
rlabel metal2 40096 48328 40096 48328 0 _0000_
rlabel metal2 30352 12040 30352 12040 0 _0001_
rlabel metal3 30688 9688 30688 9688 0 _0002_
rlabel metal2 27496 9800 27496 9800 0 _0003_
rlabel metal2 28168 10920 28168 10920 0 _0004_
rlabel metal2 43288 11088 43288 11088 0 _0005_
rlabel metal3 40768 9128 40768 9128 0 _0006_
rlabel metal2 41272 11760 41272 11760 0 _0007_
rlabel metal2 38696 10696 38696 10696 0 _0008_
rlabel metal2 42616 21168 42616 21168 0 _0009_
rlabel metal2 40264 19600 40264 19600 0 _0010_
rlabel metal2 41160 22064 41160 22064 0 _0011_
rlabel metal2 38696 21392 38696 21392 0 _0012_
rlabel metal2 31080 34552 31080 34552 0 _0013_
rlabel metal2 32312 32144 32312 32144 0 _0014_
rlabel metal2 16408 35504 16408 35504 0 _0015_
rlabel metal2 18536 42392 18536 42392 0 _0016_
rlabel metal2 15176 41552 15176 41552 0 _0017_
rlabel metal2 13720 45360 13720 45360 0 _0018_
rlabel metal2 18200 45416 18200 45416 0 _0019_
rlabel metal2 18256 47656 18256 47656 0 _0020_
rlabel metal2 18424 51016 18424 51016 0 _0021_
rlabel metal2 14392 47096 14392 47096 0 _0022_
rlabel metal2 18592 49112 18592 49112 0 _0023_
rlabel metal2 2520 30576 2520 30576 0 _0024_
rlabel metal3 4312 32536 4312 32536 0 _0025_
rlabel metal2 2856 35672 2856 35672 0 _0026_
rlabel metal3 4480 38696 4480 38696 0 _0027_
rlabel metal2 2520 42112 2520 42112 0 _0028_
rlabel metal2 2520 45024 2520 45024 0 _0029_
rlabel metal2 2520 47824 2520 47824 0 _0030_
rlabel metal2 2520 49448 2520 49448 0 _0031_
rlabel metal3 5488 52248 5488 52248 0 _0032_
rlabel metal2 16632 51408 16632 51408 0 _0033_
rlabel metal2 16016 53928 16016 53928 0 _0034_
rlabel metal2 4928 31080 4928 31080 0 _0035_
rlabel metal2 4872 34272 4872 34272 0 _0036_
rlabel metal2 5936 37352 5936 37352 0 _0037_
rlabel metal2 6440 39256 6440 39256 0 _0038_
rlabel metal2 6104 42280 6104 42280 0 _0039_
rlabel metal2 5544 45248 5544 45248 0 _0040_
rlabel metal2 7784 46928 7784 46928 0 _0041_
rlabel metal2 6888 51688 6888 51688 0 _0042_
rlabel metal2 6888 54824 6888 54824 0 _0043_
rlabel metal2 12040 53088 12040 53088 0 _0044_
rlabel metal2 13944 54656 13944 54656 0 _0045_
rlabel metal2 46088 35280 46088 35280 0 _0046_
rlabel metal2 43400 40712 43400 40712 0 _0047_
rlabel metal2 46088 41664 46088 41664 0 _0048_
rlabel metal2 44632 37632 44632 37632 0 _0049_
rlabel metal2 39592 38360 39592 38360 0 _0050_
rlabel metal2 41832 39144 41832 39144 0 _0051_
rlabel metal2 39816 35952 39816 35952 0 _0052_
rlabel metal2 40376 25760 40376 25760 0 _0053_
rlabel metal2 43568 24808 43568 24808 0 _0054_
rlabel metal2 45640 23576 45640 23576 0 _0055_
rlabel metal2 47432 21392 47432 21392 0 _0056_
rlabel metal2 47432 22568 47432 22568 0 _0057_
rlabel metal2 46088 25648 46088 25648 0 _0058_
rlabel metal2 47376 27160 47376 27160 0 _0059_
rlabel metal2 45640 29736 45640 29736 0 _0060_
rlabel metal2 46984 31416 46984 31416 0 _0061_
rlabel metal2 46088 33544 46088 33544 0 _0062_
rlabel metal2 43792 35000 43792 35000 0 _0063_
rlabel metal3 43008 33992 43008 33992 0 _0064_
rlabel metal2 43848 31416 43848 31416 0 _0065_
rlabel metal2 42168 29008 42168 29008 0 _0066_
rlabel metal3 40656 27160 40656 27160 0 _0067_
rlabel metal2 33880 24864 33880 24864 0 _0068_
rlabel metal2 37576 25088 37576 25088 0 _0069_
rlabel metal2 33320 27384 33320 27384 0 _0070_
rlabel metal2 38304 27272 38304 27272 0 _0071_
rlabel metal2 39704 30408 39704 30408 0 _0072_
rlabel metal2 37576 32984 37576 32984 0 _0073_
rlabel metal2 33936 30968 33936 30968 0 _0074_
rlabel metal2 32144 28728 32144 28728 0 _0075_
rlabel metal2 34664 32984 34664 32984 0 _0076_
rlabel metal2 27384 39144 27384 39144 0 _0077_
rlabel metal2 20552 42000 20552 42000 0 _0078_
rlabel metal2 23576 44688 23576 44688 0 _0079_
rlabel metal3 26656 47320 26656 47320 0 _0080_
rlabel metal2 24920 51464 24920 51464 0 _0081_
rlabel metal2 30184 54824 30184 54824 0 _0082_
rlabel metal2 25144 54488 25144 54488 0 _0083_
rlabel metal3 21448 53928 21448 53928 0 _0084_
rlabel metal2 18648 54936 18648 54936 0 _0085_
rlabel metal2 45640 13104 45640 13104 0 _0086_
rlabel metal2 46088 18760 46088 18760 0 _0087_
rlabel metal3 45528 17528 45528 17528 0 _0088_
rlabel metal2 44744 15288 44744 15288 0 _0089_
rlabel metal2 42616 13496 42616 13496 0 _0090_
rlabel metal2 39256 14168 39256 14168 0 _0091_
rlabel metal3 37128 15176 37128 15176 0 _0092_
rlabel metal2 36064 21448 36064 21448 0 _0093_
rlabel metal2 37016 18424 37016 18424 0 _0094_
rlabel metal2 32312 21168 32312 21168 0 _0095_
rlabel metal2 33208 29736 33208 29736 0 _0096_
rlabel metal2 46648 9352 46648 9352 0 _0097_
rlabel metal3 45640 6552 45640 6552 0 _0098_
rlabel metal2 46312 4648 46312 4648 0 _0099_
rlabel metal2 41720 4648 41720 4648 0 _0100_
rlabel metal3 38808 5096 38808 5096 0 _0101_
rlabel metal2 38472 4648 38472 4648 0 _0102_
rlabel metal2 33880 4648 33880 4648 0 _0103_
rlabel metal2 35224 10416 35224 10416 0 _0104_
rlabel metal2 35336 12544 35336 12544 0 _0105_
rlabel metal2 33488 15064 33488 15064 0 _0106_
rlabel metal2 10696 18424 10696 18424 0 _0107_
rlabel metal2 33600 8344 33600 8344 0 _0108_
rlabel metal2 31080 4760 31080 4760 0 _0109_
rlabel metal2 28168 4760 28168 4760 0 _0110_
rlabel metal2 26544 4536 26544 4536 0 _0111_
rlabel metal2 22792 3976 22792 3976 0 _0112_
rlabel metal2 22120 6216 22120 6216 0 _0113_
rlabel metal2 22176 9912 22176 9912 0 _0114_
rlabel metal2 23912 11592 23912 11592 0 _0115_
rlabel metal2 27496 15512 27496 15512 0 _0116_
rlabel metal2 24528 15960 24528 15960 0 _0117_
rlabel metal2 17920 28616 17920 28616 0 _0118_
rlabel metal2 32088 36512 32088 36512 0 _0119_
rlabel metal2 37800 36008 37800 36008 0 _0120_
rlabel metal2 33152 39704 33152 39704 0 _0121_
rlabel metal2 36904 39368 36904 39368 0 _0122_
rlabel metal2 35000 42224 35000 42224 0 _0123_
rlabel metal2 31640 46088 31640 46088 0 _0124_
rlabel metal3 38024 47656 38024 47656 0 _0125_
rlabel metal2 33880 50120 33880 50120 0 _0126_
rlabel metal2 37240 51240 37240 51240 0 _0127_
rlabel metal2 39368 55216 39368 55216 0 _0128_
rlabel metal3 45752 51464 45752 51464 0 _0129_
rlabel metal2 47376 53704 47376 53704 0 _0130_
rlabel metal2 47432 55412 47432 55412 0 _0131_
rlabel metal3 41888 47208 41888 47208 0 _0132_
rlabel metal2 44744 45304 44744 45304 0 _0133_
rlabel metal2 47432 44632 47432 44632 0 _0134_
rlabel metal3 47040 48328 47040 48328 0 _0135_
rlabel metal2 46984 46256 46984 46256 0 _0136_
rlabel metal2 40768 48776 40768 48776 0 _0137_
rlabel metal2 43176 46312 43176 46312 0 _0138_
rlabel metal2 38192 40488 38192 40488 0 _0139_
rlabel metal2 36344 42224 36344 42224 0 _0140_
rlabel metal2 41496 41496 41496 41496 0 _0141_
rlabel metal2 36456 43904 36456 43904 0 _0142_
rlabel metal2 38080 44520 38080 44520 0 _0143_
rlabel metal2 38920 47768 38920 47768 0 _0144_
rlabel metal2 38696 50904 38696 50904 0 _0145_
rlabel metal2 39704 53032 39704 53032 0 _0146_
rlabel metal2 40264 54936 40264 54936 0 _0147_
rlabel metal2 43624 54824 43624 54824 0 _0148_
rlabel metal3 45696 49672 45696 49672 0 _0149_
rlabel metal2 42168 49224 42168 49224 0 _0150_
rlabel metal2 40040 32984 40040 32984 0 _0151_
rlabel metal2 29960 19432 29960 19432 0 _0152_
rlabel metal2 30128 16184 30128 16184 0 _0153_
rlabel metal2 29456 16968 29456 16968 0 _0154_
rlabel metal2 28168 19600 28168 19600 0 _0155_
rlabel metal2 26040 18480 26040 18480 0 _0156_
rlabel metal2 22568 17808 22568 17808 0 _0157_
rlabel metal2 18704 5208 18704 5208 0 _0158_
rlabel metal2 19096 5096 19096 5096 0 _0159_
rlabel metal2 19992 7616 19992 7616 0 _0160_
rlabel metal2 19992 10752 19992 10752 0 _0161_
rlabel metal3 20944 12824 20944 12824 0 _0162_
rlabel metal2 21448 15484 21448 15484 0 _0163_
rlabel metal2 17192 6888 17192 6888 0 _0164_
rlabel metal2 16408 7896 16408 7896 0 _0165_
rlabel metal2 15736 9968 15736 9968 0 _0166_
rlabel metal2 15624 11536 15624 11536 0 _0167_
rlabel metal2 14728 14504 14728 14504 0 _0168_
rlabel metal3 16688 15848 16688 15848 0 _0169_
rlabel metal2 24584 23912 24584 23912 0 _0170_
rlabel metal2 23688 22904 23688 22904 0 _0171_
rlabel metal2 22008 26040 22008 26040 0 _0172_
rlabel metal2 23352 25200 23352 25200 0 _0173_
rlabel metal2 16184 25256 16184 25256 0 _0174_
rlabel metal2 17584 25704 17584 25704 0 _0175_
rlabel metal2 19320 26236 19320 26236 0 _0176_
rlabel metal2 18088 23632 18088 23632 0 _0177_
rlabel metal2 5320 24080 5320 24080 0 _0178_
rlabel metal2 10360 21728 10360 21728 0 _0179_
rlabel metal3 10192 20104 10192 20104 0 _0180_
rlabel metal3 10024 19320 10024 19320 0 _0181_
rlabel metal2 14280 22120 14280 22120 0 _0182_
rlabel metal2 14224 24024 14224 24024 0 _0183_
rlabel metal2 14840 24304 14840 24304 0 _0184_
rlabel metal2 12376 18592 12376 18592 0 _0185_
rlabel metal2 14840 18368 14840 18368 0 _0186_
rlabel metal2 14728 17640 14728 17640 0 _0187_
rlabel metal2 15848 20440 15848 20440 0 _0188_
rlabel metal2 35168 22568 35168 22568 0 _0189_
rlabel metal2 29512 22736 29512 22736 0 _0190_
rlabel metal2 30800 24920 30800 24920 0 _0191_
rlabel metal2 29960 25872 29960 25872 0 _0192_
rlabel metal2 7280 46760 7280 46760 0 _0193_
rlabel metal2 42840 41328 42840 41328 0 _0194_
rlabel metal2 9408 48440 9408 48440 0 _0195_
rlabel metal2 9464 47824 9464 47824 0 _0196_
rlabel metal2 8848 49224 8848 49224 0 _0197_
rlabel metal2 11480 51632 11480 51632 0 _0198_
rlabel metal2 9464 51296 9464 51296 0 _0199_
rlabel metal2 8680 50680 8680 50680 0 _0200_
rlabel metal2 10136 54264 10136 54264 0 _0201_
rlabel metal2 11704 54936 11704 54936 0 _0202_
rlabel metal2 10024 54376 10024 54376 0 _0203_
rlabel metal2 9800 55272 9800 55272 0 _0204_
rlabel metal2 10248 54544 10248 54544 0 _0205_
rlabel metal2 10920 54320 10920 54320 0 _0206_
rlabel metal2 11032 53872 11032 53872 0 _0207_
rlabel metal2 14728 53928 14728 53928 0 _0208_
rlabel metal2 31976 29680 31976 29680 0 _0209_
rlabel metal3 23184 46872 23184 46872 0 _0210_
rlabel metal2 14056 54488 14056 54488 0 _0211_
rlabel metal2 46760 41160 46760 41160 0 _0212_
rlabel metal2 38696 17808 38696 17808 0 _0213_
rlabel metal2 43512 41552 43512 41552 0 _0214_
rlabel metal2 47208 40824 47208 40824 0 _0215_
rlabel metal2 47264 39704 47264 39704 0 _0216_
rlabel metal2 47544 41160 47544 41160 0 _0217_
rlabel metal2 44128 40152 44128 40152 0 _0218_
rlabel metal3 44576 38248 44576 38248 0 _0219_
rlabel metal2 39592 33208 39592 33208 0 _0220_
rlabel metal2 39928 38416 39928 38416 0 _0221_
rlabel metal2 42056 39648 42056 39648 0 _0222_
rlabel metal3 44408 44184 44408 44184 0 _0223_
rlabel metal2 41384 41216 41384 41216 0 _0224_
rlabel metal2 42280 36736 42280 36736 0 _0225_
rlabel metal2 41608 37016 41608 37016 0 _0226_
rlabel metal2 40152 36064 40152 36064 0 _0227_
rlabel metal3 39116 30856 39116 30856 0 _0228_
rlabel metal2 41440 31080 41440 31080 0 _0229_
rlabel metal3 42168 31192 42168 31192 0 _0230_
rlabel metal2 42616 25984 42616 25984 0 _0231_
rlabel metal3 42672 26488 42672 26488 0 _0232_
rlabel metal2 41944 25872 41944 25872 0 _0233_
rlabel metal2 42280 30072 42280 30072 0 _0234_
rlabel metal2 43288 26376 43288 26376 0 _0235_
rlabel metal2 43400 26824 43400 26824 0 _0236_
rlabel metal2 44296 32312 44296 32312 0 _0237_
rlabel metal2 45192 25816 45192 25816 0 _0238_
rlabel metal3 44408 24920 44408 24920 0 _0239_
rlabel metal3 43568 25480 43568 25480 0 _0240_
rlabel metal2 46872 24696 46872 24696 0 _0241_
rlabel metal2 45528 23800 45528 23800 0 _0242_
rlabel metal2 45976 23184 45976 23184 0 _0243_
rlabel metal2 44968 23408 44968 23408 0 _0244_
rlabel metal2 46872 22456 46872 22456 0 _0245_
rlabel metal2 47096 21336 47096 21336 0 _0246_
rlabel metal2 47320 23800 47320 23800 0 _0247_
rlabel metal2 47320 25032 47320 25032 0 _0248_
rlabel metal2 44968 27496 44968 27496 0 _0249_
rlabel metal2 46648 26544 46648 26544 0 _0250_
rlabel metal2 46872 26908 46872 26908 0 _0251_
rlabel metal2 47432 32928 47432 32928 0 _0252_
rlabel metal2 47040 27048 47040 27048 0 _0253_
rlabel metal2 47544 27720 47544 27720 0 _0254_
rlabel metal2 47096 29512 47096 29512 0 _0255_
rlabel metal2 47432 30464 47432 30464 0 _0256_
rlabel metal3 47432 31080 47432 31080 0 _0257_
rlabel metal2 46760 31752 46760 31752 0 _0258_
rlabel metal2 46200 33376 46200 33376 0 _0259_
rlabel metal2 43512 32760 43512 32760 0 _0260_
rlabel metal2 45696 32760 45696 32760 0 _0261_
rlabel metal2 44632 34496 44632 34496 0 _0262_
rlabel metal2 44856 33264 44856 33264 0 _0263_
rlabel metal2 44968 34328 44968 34328 0 _0264_
rlabel metal2 43848 33152 43848 33152 0 _0265_
rlabel metal2 44408 34384 44408 34384 0 _0266_
rlabel metal2 44016 33320 44016 33320 0 _0267_
rlabel metal2 44352 31192 44352 31192 0 _0268_
rlabel metal2 43736 31360 43736 31360 0 _0269_
rlabel metal2 43176 29792 43176 29792 0 _0270_
rlabel metal2 42952 27608 42952 27608 0 _0271_
rlabel metal2 39144 26684 39144 26684 0 _0272_
rlabel metal2 40936 28280 40936 28280 0 _0273_
rlabel metal2 41776 28056 41776 28056 0 _0274_
rlabel metal2 47880 39452 47880 39452 0 _0275_
rlabel metal3 45416 37352 45416 37352 0 _0276_
rlabel metal2 46480 39480 46480 39480 0 _0277_
rlabel metal2 46088 38696 46088 38696 0 _0278_
rlabel metal3 46368 37912 46368 37912 0 _0279_
rlabel metal2 43736 19712 43736 19712 0 _0280_
rlabel metal2 35560 22904 35560 22904 0 _0281_
rlabel metal2 35112 24696 35112 24696 0 _0282_
rlabel metal3 42896 45864 42896 45864 0 _0283_
rlabel metal2 47768 36904 47768 36904 0 _0284_
rlabel metal2 40376 28672 40376 28672 0 _0285_
rlabel metal2 25816 15624 25816 15624 0 _0286_
rlabel metal2 26824 16128 26824 16128 0 _0287_
rlabel metal2 35896 9184 35896 9184 0 _0288_
rlabel metal2 35672 23856 35672 23856 0 _0289_
rlabel metal2 35952 24024 35952 24024 0 _0290_
rlabel metal2 35784 25368 35784 25368 0 _0291_
rlabel metal3 36288 25480 36288 25480 0 _0292_
rlabel metal2 37016 27216 37016 27216 0 _0293_
rlabel metal2 35896 27384 35896 27384 0 _0294_
rlabel metal2 37520 28840 37520 28840 0 _0295_
rlabel metal2 38192 28392 38192 28392 0 _0296_
rlabel metal2 43736 17640 43736 17640 0 _0297_
rlabel metal2 37520 27048 37520 27048 0 _0298_
rlabel metal2 39032 31248 39032 31248 0 _0299_
rlabel metal3 38472 30968 38472 30968 0 _0300_
rlabel metal2 38248 32200 38248 32200 0 _0301_
rlabel metal2 37128 32480 37128 32480 0 _0302_
rlabel metal2 37408 32648 37408 32648 0 _0303_
rlabel metal2 34888 30688 34888 30688 0 _0304_
rlabel metal2 36008 29624 36008 29624 0 _0305_
rlabel metal2 33712 30296 33712 30296 0 _0306_
rlabel metal2 33768 33432 33768 33432 0 _0307_
rlabel metal3 33992 33432 33992 33432 0 _0308_
rlabel metal2 34776 32592 34776 32592 0 _0309_
rlabel metal3 34832 34104 34832 34104 0 _0310_
rlabel metal3 33992 32312 33992 32312 0 _0311_
rlabel metal2 25592 39648 25592 39648 0 _0312_
rlabel metal2 26320 38920 26320 38920 0 _0313_
rlabel metal2 26040 38864 26040 38864 0 _0314_
rlabel metal2 24584 42896 24584 42896 0 _0315_
rlabel metal2 24136 39648 24136 39648 0 _0316_
rlabel metal2 24752 39592 24752 39592 0 _0317_
rlabel metal2 23352 40208 23352 40208 0 _0318_
rlabel metal2 23464 41496 23464 41496 0 _0319_
rlabel metal3 22232 42840 22232 42840 0 _0320_
rlabel metal3 21448 42728 21448 42728 0 _0321_
rlabel metal2 23688 44184 23688 44184 0 _0322_
rlabel metal2 25928 45360 25928 45360 0 _0323_
rlabel metal2 24360 45416 24360 45416 0 _0324_
rlabel metal2 24024 44632 24024 44632 0 _0325_
rlabel metal2 25592 45752 25592 45752 0 _0326_
rlabel metal2 25312 46088 25312 46088 0 _0327_
rlabel metal2 26712 48832 26712 48832 0 _0328_
rlabel metal2 27720 47824 27720 47824 0 _0329_
rlabel metal2 26600 48608 26600 48608 0 _0330_
rlabel metal2 28392 47768 28392 47768 0 _0331_
rlabel metal2 26824 48888 26824 48888 0 _0332_
rlabel metal2 27328 46088 27328 46088 0 _0333_
rlabel metal2 26600 50036 26600 50036 0 _0334_
rlabel metal2 25592 51800 25592 51800 0 _0335_
rlabel metal2 26824 51912 26824 51912 0 _0336_
rlabel metal2 27384 50792 27384 50792 0 _0337_
rlabel metal2 29344 53480 29344 53480 0 _0338_
rlabel metal2 27776 54376 27776 54376 0 _0339_
rlabel metal2 29288 54040 29288 54040 0 _0340_
rlabel metal2 28000 53704 28000 53704 0 _0341_
rlabel metal2 27664 53816 27664 53816 0 _0342_
rlabel metal3 25760 53704 25760 53704 0 _0343_
rlabel metal2 25928 53368 25928 53368 0 _0344_
rlabel metal2 25816 53704 25816 53704 0 _0345_
rlabel metal2 22848 55048 22848 55048 0 _0346_
rlabel metal2 23072 53032 23072 53032 0 _0347_
rlabel metal2 23464 53816 23464 53816 0 _0348_
rlabel metal2 23352 54096 23352 54096 0 _0349_
rlabel metal2 22232 55440 22232 55440 0 _0350_
rlabel metal2 22232 53872 22232 53872 0 _0351_
rlabel metal2 21896 54096 21896 54096 0 _0352_
rlabel metal3 45472 19880 45472 19880 0 _0353_
rlabel metal3 45192 13720 45192 13720 0 _0354_
rlabel metal2 25480 7392 25480 7392 0 _0355_
rlabel metal3 46312 16912 46312 16912 0 _0356_
rlabel metal3 40376 17528 40376 17528 0 _0357_
rlabel metal2 40376 18088 40376 18088 0 _0358_
rlabel metal2 44520 17080 44520 17080 0 _0359_
rlabel metal2 44352 12936 44352 12936 0 _0360_
rlabel metal2 41160 13384 41160 13384 0 _0361_
rlabel metal2 43960 17808 43960 17808 0 _0362_
rlabel metal2 43176 17528 43176 17528 0 _0363_
rlabel metal2 45080 17640 45080 17640 0 _0364_
rlabel metal2 34664 16632 34664 16632 0 _0365_
rlabel metal2 43456 16072 43456 16072 0 _0366_
rlabel metal3 43288 18312 43288 18312 0 _0367_
rlabel metal2 44968 18480 44968 18480 0 _0368_
rlabel metal2 45416 17136 45416 17136 0 _0369_
rlabel metal3 45192 17080 45192 17080 0 _0370_
rlabel metal2 45528 16800 45528 16800 0 _0371_
rlabel metal2 44296 17808 44296 17808 0 _0372_
rlabel metal3 41328 18424 41328 18424 0 _0373_
rlabel metal2 42952 17080 42952 17080 0 _0374_
rlabel metal2 43680 16072 43680 16072 0 _0375_
rlabel metal2 43792 16296 43792 16296 0 _0376_
rlabel metal2 42056 15624 42056 15624 0 _0377_
rlabel metal2 43624 15512 43624 15512 0 _0378_
rlabel metal2 43064 15344 43064 15344 0 _0379_
rlabel metal3 40488 16968 40488 16968 0 _0380_
rlabel metal2 42728 10416 42728 10416 0 _0381_
rlabel metal2 42392 15624 42392 15624 0 _0382_
rlabel metal2 42392 14112 42392 14112 0 _0383_
rlabel metal2 39144 15232 39144 15232 0 _0384_
rlabel metal3 40264 16856 40264 16856 0 _0385_
rlabel metal2 39256 16520 39256 16520 0 _0386_
rlabel metal2 39816 15456 39816 15456 0 _0387_
rlabel metal2 39088 13832 39088 13832 0 _0388_
rlabel metal2 36120 17136 36120 17136 0 _0389_
rlabel metal3 36736 17080 36736 17080 0 _0390_
rlabel metal2 36456 16464 36456 16464 0 _0391_
rlabel metal3 35728 18424 35728 18424 0 _0392_
rlabel metal2 35896 16184 35896 16184 0 _0393_
rlabel metal2 38472 15512 38472 15512 0 _0394_
rlabel metal3 36624 20664 36624 20664 0 _0395_
rlabel metal2 26824 12936 26824 12936 0 _0396_
rlabel metal3 34104 18312 34104 18312 0 _0397_
rlabel metal3 36008 18648 36008 18648 0 _0398_
rlabel metal2 36232 19824 36232 19824 0 _0399_
rlabel metal2 35336 19376 35336 19376 0 _0400_
rlabel metal3 34776 17640 34776 17640 0 _0401_
rlabel metal3 34720 19320 34720 19320 0 _0402_
rlabel metal2 44520 19880 44520 19880 0 _0403_
rlabel metal2 35616 17528 35616 17528 0 _0404_
rlabel metal2 36232 18312 36232 18312 0 _0405_
rlabel metal2 32928 18424 32928 18424 0 _0406_
rlabel metal2 33208 18984 33208 18984 0 _0407_
rlabel metal2 32424 20272 32424 20272 0 _0408_
rlabel metal2 33656 29736 33656 29736 0 _0409_
rlabel metal2 45528 8624 45528 8624 0 _0410_
rlabel metal3 41440 8232 41440 8232 0 _0411_
rlabel metal2 37576 7840 37576 7840 0 _0412_
rlabel metal3 43736 7560 43736 7560 0 _0413_
rlabel metal2 42392 9016 42392 9016 0 _0414_
rlabel metal2 44968 9072 44968 9072 0 _0415_
rlabel metal3 42168 8008 42168 8008 0 _0416_
rlabel metal2 41832 6776 41832 6776 0 _0417_
rlabel metal2 42392 7560 42392 7560 0 _0418_
rlabel metal2 38696 5880 38696 5880 0 _0419_
rlabel metal2 43400 6608 43400 6608 0 _0420_
rlabel metal2 42056 6720 42056 6720 0 _0421_
rlabel metal2 42280 6664 42280 6664 0 _0422_
rlabel metal2 41944 7000 41944 7000 0 _0423_
rlabel metal2 42896 5208 42896 5208 0 _0424_
rlabel metal2 39928 5264 39928 5264 0 _0425_
rlabel metal2 39592 7504 39592 7504 0 _0426_
rlabel metal2 40040 6664 40040 6664 0 _0427_
rlabel metal2 40040 5992 40040 5992 0 _0428_
rlabel metal3 39704 6384 39704 6384 0 _0429_
rlabel metal2 40936 6160 40936 6160 0 _0430_
rlabel metal2 41160 5264 41160 5264 0 _0431_
rlabel metal3 39312 6552 39312 6552 0 _0432_
rlabel metal3 39256 5880 39256 5880 0 _0433_
rlabel metal2 39144 6048 39144 6048 0 _0434_
rlabel metal2 37464 5264 37464 5264 0 _0435_
rlabel metal2 35672 6048 35672 6048 0 _0436_
rlabel metal2 34888 6608 34888 6608 0 _0437_
rlabel metal2 35560 5152 35560 5152 0 _0438_
rlabel metal3 30576 5992 30576 5992 0 _0439_
rlabel metal2 36344 5264 36344 5264 0 _0440_
rlabel metal2 33432 14224 33432 14224 0 _0441_
rlabel metal2 34664 7336 34664 7336 0 _0442_
rlabel metal2 34776 6160 34776 6160 0 _0443_
rlabel metal2 35000 11312 35000 11312 0 _0444_
rlabel metal2 34608 5880 34608 5880 0 _0445_
rlabel metal2 33544 5544 33544 5544 0 _0446_
rlabel metal2 35560 10472 35560 10472 0 _0447_
rlabel metal2 34328 11424 34328 11424 0 _0448_
rlabel metal2 34216 11760 34216 11760 0 _0449_
rlabel metal2 34888 10920 34888 10920 0 _0450_
rlabel metal2 34664 10080 34664 10080 0 _0451_
rlabel metal2 34496 13720 34496 13720 0 _0452_
rlabel metal2 35560 13888 35560 13888 0 _0453_
rlabel metal2 34776 12936 34776 12936 0 _0454_
rlabel metal3 34664 13048 34664 13048 0 _0455_
rlabel metal2 24248 11368 24248 11368 0 _0456_
rlabel metal2 13664 17080 13664 17080 0 _0457_
rlabel metal2 31976 14000 31976 14000 0 _0458_
rlabel metal2 32872 15064 32872 15064 0 _0459_
rlabel metal2 15176 25760 15176 25760 0 _0460_
rlabel metal2 11144 18312 11144 18312 0 _0461_
rlabel metal3 33656 9016 33656 9016 0 _0462_
rlabel metal3 30800 7448 30800 7448 0 _0463_
rlabel metal2 25928 7784 25928 7784 0 _0464_
rlabel metal2 27048 7840 27048 7840 0 _0465_
rlabel metal2 31472 6664 31472 6664 0 _0466_
rlabel metal2 33432 7896 33432 7896 0 _0467_
rlabel metal2 24808 5320 24808 5320 0 _0468_
rlabel metal2 31920 6664 31920 6664 0 _0469_
rlabel metal3 29456 6552 29456 6552 0 _0470_
rlabel metal2 32032 5880 32032 5880 0 _0471_
rlabel metal2 31192 5152 31192 5152 0 _0472_
rlabel metal3 28840 6664 28840 6664 0 _0473_
rlabel metal3 26040 5936 26040 5936 0 _0474_
rlabel metal2 23800 5488 23800 5488 0 _0475_
rlabel metal2 30072 5880 30072 5880 0 _0476_
rlabel metal2 29232 5208 29232 5208 0 _0477_
rlabel metal2 23800 8288 23800 8288 0 _0478_
rlabel metal2 26040 5656 26040 5656 0 _0479_
rlabel metal2 23464 5376 23464 5376 0 _0480_
rlabel metal3 27104 5768 27104 5768 0 _0481_
rlabel metal2 25368 9688 25368 9688 0 _0482_
rlabel metal2 26712 4760 26712 4760 0 _0483_
rlabel metal2 22792 7448 22792 7448 0 _0484_
rlabel metal2 22456 6384 22456 6384 0 _0485_
rlabel metal3 23744 5096 23744 5096 0 _0486_
rlabel metal2 22904 4424 22904 4424 0 _0487_
rlabel metal2 23856 6664 23856 6664 0 _0488_
rlabel metal2 24360 6720 24360 6720 0 _0489_
rlabel metal2 23968 6440 23968 6440 0 _0490_
rlabel metal2 22008 6720 22008 6720 0 _0491_
rlabel metal3 25200 15176 25200 15176 0 _0492_
rlabel metal2 23576 9912 23576 9912 0 _0493_
rlabel metal3 24976 10024 24976 10024 0 _0494_
rlabel metal3 24696 10584 24696 10584 0 _0495_
rlabel metal2 25592 10192 25592 10192 0 _0496_
rlabel metal3 23688 9912 23688 9912 0 _0497_
rlabel metal2 26264 12432 26264 12432 0 _0498_
rlabel metal3 24584 12040 24584 12040 0 _0499_
rlabel metal2 26600 12880 26600 12880 0 _0500_
rlabel metal2 25704 11648 25704 11648 0 _0501_
rlabel metal2 25256 11872 25256 11872 0 _0502_
rlabel metal3 25536 14280 25536 14280 0 _0503_
rlabel metal2 26264 15232 26264 15232 0 _0504_
rlabel metal2 27720 13888 27720 13888 0 _0505_
rlabel metal2 26824 14616 26824 14616 0 _0506_
rlabel metal2 15792 26488 15792 26488 0 _0507_
rlabel metal4 23912 14504 23912 14504 0 _0508_
rlabel metal2 24472 12264 24472 12264 0 _0509_
rlabel metal2 15848 26264 15848 26264 0 _0510_
rlabel metal3 36288 38920 36288 38920 0 _0511_
rlabel metal2 33656 37464 33656 37464 0 _0512_
rlabel metal2 34384 38808 34384 38808 0 _0513_
rlabel metal2 25704 35504 25704 35504 0 _0514_
rlabel metal2 26824 36960 26824 36960 0 _0515_
rlabel metal2 34552 36904 34552 36904 0 _0516_
rlabel metal2 36120 37072 36120 37072 0 _0517_
rlabel metal2 34888 37408 34888 37408 0 _0518_
rlabel metal2 35560 37240 35560 37240 0 _0519_
rlabel metal2 32088 40432 32088 40432 0 _0520_
rlabel metal2 39368 42448 39368 42448 0 _0521_
rlabel metal2 32312 39648 32312 39648 0 _0522_
rlabel metal3 32536 39032 32536 39032 0 _0523_
rlabel metal2 33544 39816 33544 39816 0 _0524_
rlabel metal2 34440 41216 34440 41216 0 _0525_
rlabel metal2 36008 39592 36008 39592 0 _0526_
rlabel metal3 34832 41720 34832 41720 0 _0527_
rlabel metal3 34944 39816 34944 39816 0 _0528_
rlabel metal3 34944 41160 34944 41160 0 _0529_
rlabel metal2 33208 42448 33208 42448 0 _0530_
rlabel metal3 32592 42728 32592 42728 0 _0531_
rlabel metal2 32984 42616 32984 42616 0 _0532_
rlabel metal2 33432 42280 33432 42280 0 _0533_
rlabel metal2 34216 44240 34216 44240 0 _0534_
rlabel metal2 34888 42280 34888 42280 0 _0535_
rlabel metal3 33824 45304 33824 45304 0 _0536_
rlabel metal2 32984 45752 32984 45752 0 _0537_
rlabel metal2 32760 47152 32760 47152 0 _0538_
rlabel metal2 32200 21168 32200 21168 0 _0539_
rlabel metal2 32536 46872 32536 46872 0 _0540_
rlabel metal2 44968 51688 44968 51688 0 _0541_
rlabel metal2 34608 45304 34608 45304 0 _0542_
rlabel metal3 35784 46424 35784 46424 0 _0543_
rlabel metal2 35784 45472 35784 45472 0 _0544_
rlabel metal2 35896 45136 35896 45136 0 _0545_
rlabel metal2 36456 46648 36456 46648 0 _0546_
rlabel metal2 36008 49280 36008 49280 0 _0547_
rlabel metal2 35560 48776 35560 48776 0 _0548_
rlabel metal2 35168 49000 35168 49000 0 _0549_
rlabel metal2 36792 49392 36792 49392 0 _0550_
rlabel metal2 35000 50288 35000 50288 0 _0551_
rlabel metal2 34888 50568 34888 50568 0 _0552_
rlabel metal2 36120 51744 36120 51744 0 _0553_
rlabel metal2 35896 50568 35896 50568 0 _0554_
rlabel metal2 36008 51856 36008 51856 0 _0555_
rlabel metal3 36512 52808 36512 52808 0 _0556_
rlabel metal2 37240 51576 37240 51576 0 _0557_
rlabel metal2 39480 54544 39480 54544 0 _0558_
rlabel metal2 36344 55216 36344 55216 0 _0559_
rlabel metal2 38248 52640 38248 52640 0 _0560_
rlabel metal2 39256 54432 39256 54432 0 _0561_
rlabel metal2 37576 52752 37576 52752 0 _0562_
rlabel metal2 37352 53760 37352 53760 0 _0563_
rlabel metal2 38584 52584 38584 52584 0 _0564_
rlabel metal2 47992 52752 47992 52752 0 _0565_
rlabel metal2 43848 51408 43848 51408 0 _0566_
rlabel metal3 46424 49224 46424 49224 0 _0567_
rlabel metal2 44520 50456 44520 50456 0 _0568_
rlabel metal2 47880 52192 47880 52192 0 _0569_
rlabel metal2 47096 53060 47096 53060 0 _0570_
rlabel metal2 41216 54712 41216 54712 0 _0571_
rlabel metal3 45668 55832 45668 55832 0 _0572_
rlabel metal3 46872 44968 46872 44968 0 _0573_
rlabel metal3 42224 45080 42224 45080 0 _0574_
rlabel metal2 46200 44968 46200 44968 0 _0575_
rlabel metal2 44184 44744 44184 44744 0 _0576_
rlabel metal2 47096 44016 47096 44016 0 _0577_
rlabel metal2 47992 47488 47992 47488 0 _0578_
rlabel metal2 46760 48272 46760 48272 0 _0579_
rlabel metal2 47096 46200 47096 46200 0 _0580_
rlabel metal2 41160 44800 41160 44800 0 _0581_
rlabel metal2 43568 46088 43568 46088 0 _0582_
rlabel metal2 46312 46648 46312 46648 0 _0583_
rlabel metal3 44744 45864 44744 45864 0 _0584_
rlabel metal2 38696 45976 38696 45976 0 _0585_
rlabel metal3 38080 41048 38080 41048 0 _0586_
rlabel metal3 32536 38808 32536 38808 0 _0587_
rlabel metal2 37688 42784 37688 42784 0 _0588_
rlabel metal3 42056 48328 42056 48328 0 _0589_
rlabel metal2 42056 44912 42056 44912 0 _0590_
rlabel metal2 40040 42280 40040 42280 0 _0591_
rlabel metal2 38808 43456 38808 43456 0 _0592_
rlabel metal2 39480 50568 39480 50568 0 _0593_
rlabel metal2 38248 44688 38248 44688 0 _0594_
rlabel metal2 39704 47488 39704 47488 0 _0595_
rlabel metal2 42168 53424 42168 53424 0 _0596_
rlabel metal2 40488 53592 40488 53592 0 _0597_
rlabel metal2 39760 50008 39760 50008 0 _0598_
rlabel metal2 40096 51576 40096 51576 0 _0599_
rlabel metal2 40376 53144 40376 53144 0 _0600_
rlabel metal2 43736 55104 43736 55104 0 _0601_
rlabel metal2 42952 50568 42952 50568 0 _0602_
rlabel metal2 42616 49112 42616 49112 0 _0603_
rlabel metal2 25368 21280 25368 21280 0 _0604_
rlabel metal2 25704 19040 25704 19040 0 _0605_
rlabel metal2 21672 17752 21672 17752 0 _0606_
rlabel metal2 22792 16072 22792 16072 0 _0607_
rlabel metal2 19096 16072 19096 16072 0 _0608_
rlabel metal2 19936 21000 19936 21000 0 _0609_
rlabel metal2 21560 18144 21560 18144 0 _0610_
rlabel metal2 25368 18312 25368 18312 0 _0611_
rlabel metal2 22680 18872 22680 18872 0 _0612_
rlabel metal2 30744 20132 30744 20132 0 _0613_
rlabel metal3 21728 16072 21728 16072 0 _0614_
rlabel metal3 24528 17416 24528 17416 0 _0615_
rlabel metal2 30912 17752 30912 17752 0 _0616_
rlabel metal2 24136 19376 24136 19376 0 _0617_
rlabel metal3 28840 17528 28840 17528 0 _0618_
rlabel metal2 28840 18872 28840 18872 0 _0619_
rlabel metal2 25480 19320 25480 19320 0 _0620_
rlabel metal2 26152 18424 26152 18424 0 _0621_
rlabel metal3 24136 20664 24136 20664 0 _0622_
rlabel metal2 23016 19488 23016 19488 0 _0623_
rlabel metal2 23464 18256 23464 18256 0 _0624_
rlabel metal3 23632 18424 23632 18424 0 _0625_
rlabel metal2 22288 15400 22288 15400 0 _0626_
rlabel metal2 19152 18536 19152 18536 0 _0627_
rlabel metal2 20552 15316 20552 15316 0 _0628_
rlabel metal2 19208 11144 19208 11144 0 _0629_
rlabel metal2 20440 5432 20440 5432 0 _0630_
rlabel metal3 20272 5880 20272 5880 0 _0631_
rlabel metal2 23240 24024 23240 24024 0 _0632_
rlabel metal2 21448 5320 21448 5320 0 _0633_
rlabel metal2 18200 21056 18200 21056 0 _0634_
rlabel metal2 21336 11088 21336 11088 0 _0635_
rlabel metal2 20664 9184 20664 9184 0 _0636_
rlabel metal2 15736 17528 15736 17528 0 _0637_
rlabel metal2 18984 12656 18984 12656 0 _0638_
rlabel metal3 21056 11256 21056 11256 0 _0639_
rlabel metal2 19544 14000 19544 14000 0 _0640_
rlabel metal3 21336 15512 21336 15512 0 _0641_
rlabel metal2 18872 18648 18872 18648 0 _0642_
rlabel metal2 16408 10696 16408 10696 0 _0643_
rlabel via2 17976 8232 17976 8232 0 _0644_
rlabel metal2 18872 8680 18872 8680 0 _0645_
rlabel metal3 18648 15848 18648 15848 0 _0646_
rlabel metal2 16856 7616 16856 7616 0 _0647_
rlabel metal2 17920 10808 17920 10808 0 _0648_
rlabel metal2 16856 10640 16856 10640 0 _0649_
rlabel metal2 16856 12208 16856 12208 0 _0650_
rlabel metal2 16856 15204 16856 15204 0 _0651_
rlabel metal3 22176 17752 22176 17752 0 _0652_
rlabel metal2 18088 15736 18088 15736 0 _0653_
rlabel metal2 19544 24416 19544 24416 0 _0654_
rlabel metal3 21896 21672 21896 21672 0 _0655_
rlabel metal3 22176 21336 22176 21336 0 _0656_
rlabel metal2 20664 20944 20664 20944 0 _0657_
rlabel metal3 19880 20776 19880 20776 0 _0658_
rlabel metal2 20552 21224 20552 21224 0 _0659_
rlabel metal2 21336 22456 21336 22456 0 _0660_
rlabel metal3 22512 23688 22512 23688 0 _0661_
rlabel metal2 23240 23128 23240 23128 0 _0662_
rlabel metal2 24136 24136 24136 24136 0 _0663_
rlabel metal2 23128 24528 23128 24528 0 _0664_
rlabel metal2 21672 25256 21672 25256 0 _0665_
rlabel metal3 22736 25368 22736 25368 0 _0666_
rlabel metal2 23016 23688 23016 23688 0 _0667_
rlabel metal2 20776 19992 20776 19992 0 _0668_
rlabel metal3 19600 19992 19600 19992 0 _0669_
rlabel metal2 20552 20160 20552 20160 0 _0670_
rlabel metal2 19320 23716 19320 23716 0 _0671_
rlabel metal3 18760 23352 18760 23352 0 _0672_
rlabel metal2 20664 24248 20664 24248 0 _0673_
rlabel metal2 19656 25424 19656 25424 0 _0674_
rlabel metal2 18200 25032 18200 25032 0 _0675_
rlabel metal2 17640 23184 17640 23184 0 _0676_
rlabel metal2 19432 25704 19432 25704 0 _0677_
rlabel metal2 20328 24304 20328 24304 0 _0678_
rlabel metal2 20440 21224 20440 21224 0 _0679_
rlabel metal3 20328 21784 20328 21784 0 _0680_
rlabel metal3 20216 22400 20216 22400 0 _0681_
rlabel metal2 12208 19992 12208 19992 0 _0682_
rlabel metal2 15288 21000 15288 21000 0 _0683_
rlabel metal2 11928 21168 11928 21168 0 _0684_
rlabel metal2 14280 20104 14280 20104 0 _0685_
rlabel metal2 10696 21392 10696 21392 0 _0686_
rlabel metal2 14952 20944 14952 20944 0 _0687_
rlabel metal2 12040 19488 12040 19488 0 _0688_
rlabel metal2 22792 20272 22792 20272 0 _0689_
rlabel metal2 14728 20048 14728 20048 0 _0690_
rlabel metal2 14392 23800 14392 23800 0 _0691_
rlabel metal2 15400 20720 15400 20720 0 _0692_
rlabel metal2 14616 21392 14616 21392 0 _0693_
rlabel metal2 13944 25368 13944 25368 0 _0694_
rlabel metal2 15176 23968 15176 23968 0 _0695_
rlabel metal2 14952 23968 14952 23968 0 _0696_
rlabel metal2 15232 19768 15232 19768 0 _0697_
rlabel metal3 16968 20104 16968 20104 0 _0698_
rlabel metal3 17192 18984 17192 18984 0 _0699_
rlabel metal2 16856 18480 16856 18480 0 _0700_
rlabel metal3 16632 19880 16632 19880 0 _0701_
rlabel metal2 30520 23912 30520 23912 0 _0702_
rlabel metal2 30072 23576 30072 23576 0 _0703_
rlabel metal3 30240 22120 30240 22120 0 _0704_
rlabel metal2 31080 24864 31080 24864 0 _0705_
rlabel metal2 30072 25704 30072 25704 0 _0706_
rlabel metal2 29960 25144 29960 25144 0 _0707_
rlabel metal3 18704 30856 18704 30856 0 _0708_
rlabel metal2 23240 34832 23240 34832 0 _0709_
rlabel metal2 21560 31416 21560 31416 0 _0710_
rlabel metal2 20440 30688 20440 30688 0 _0711_
rlabel metal2 21896 30520 21896 30520 0 _0712_
rlabel metal2 22344 30128 22344 30128 0 _0713_
rlabel metal2 23632 35000 23632 35000 0 _0714_
rlabel metal2 20328 27776 20328 27776 0 _0715_
rlabel metal2 20328 25592 20328 25592 0 _0716_
rlabel metal2 19264 32648 19264 32648 0 _0717_
rlabel metal2 19992 34272 19992 34272 0 _0718_
rlabel metal2 22792 35056 22792 35056 0 _0719_
rlabel metal2 17752 33208 17752 33208 0 _0720_
rlabel metal2 23464 36176 23464 36176 0 _0721_
rlabel metal3 24584 35000 24584 35000 0 _0722_
rlabel metal3 19936 26376 19936 26376 0 _0723_
rlabel metal2 19096 26600 19096 26600 0 _0724_
rlabel metal2 24192 35672 24192 35672 0 _0725_
rlabel metal2 16296 34552 16296 34552 0 _0726_
rlabel metal3 18816 37352 18816 37352 0 _0727_
rlabel metal2 25480 34888 25480 34888 0 _0728_
rlabel metal2 28224 26264 28224 26264 0 _0729_
rlabel metal2 24136 29120 24136 29120 0 _0730_
rlabel metal3 25116 27944 25116 27944 0 _0731_
rlabel metal3 24864 26936 24864 26936 0 _0732_
rlabel metal2 26600 26824 26600 26824 0 _0733_
rlabel metal2 26264 25088 26264 25088 0 _0734_
rlabel metal3 22736 26712 22736 26712 0 _0735_
rlabel metal3 27160 26376 27160 26376 0 _0736_
rlabel metal2 24696 28896 24696 28896 0 _0737_
rlabel metal2 33544 27888 33544 27888 0 _0738_
rlabel metal2 39256 29008 39256 29008 0 _0739_
rlabel metal2 26824 33040 26824 33040 0 _0740_
rlabel metal3 28840 27048 28840 27048 0 _0741_
rlabel metal2 24472 29176 24472 29176 0 _0742_
rlabel metal2 25816 35000 25816 35000 0 _0743_
rlabel metal2 26712 26768 26712 26768 0 _0744_
rlabel metal2 25536 25256 25536 25256 0 _0745_
rlabel metal2 24696 31024 24696 31024 0 _0746_
rlabel metal2 23520 31752 23520 31752 0 _0747_
rlabel metal2 26040 35000 26040 35000 0 _0748_
rlabel metal2 28392 35840 28392 35840 0 _0749_
rlabel metal2 16688 35784 16688 35784 0 _0750_
rlabel metal2 16632 31976 16632 31976 0 _0751_
rlabel metal2 17528 32872 17528 32872 0 _0752_
rlabel metal2 13608 31752 13608 31752 0 _0753_
rlabel metal2 15848 22624 15848 22624 0 _0754_
rlabel metal2 12488 29792 12488 29792 0 _0755_
rlabel metal2 11088 30296 11088 30296 0 _0756_
rlabel metal2 12040 30296 12040 30296 0 _0757_
rlabel metal2 15848 30352 15848 30352 0 _0758_
rlabel metal2 13496 31192 13496 31192 0 _0759_
rlabel metal3 11704 30968 11704 30968 0 _0760_
rlabel metal2 9912 31808 9912 31808 0 _0761_
rlabel metal3 16856 32424 16856 32424 0 _0762_
rlabel metal3 14616 30184 14616 30184 0 _0763_
rlabel metal2 15176 32816 15176 32816 0 _0764_
rlabel metal2 11144 31360 11144 31360 0 _0765_
rlabel metal2 11032 32480 11032 32480 0 _0766_
rlabel metal2 11480 24136 11480 24136 0 _0767_
rlabel metal2 6776 19600 6776 19600 0 _0768_
rlabel metal2 7448 22568 7448 22568 0 _0769_
rlabel metal2 6440 27552 6440 27552 0 _0770_
rlabel metal2 7224 23240 7224 23240 0 _0771_
rlabel metal3 5936 26824 5936 26824 0 _0772_
rlabel metal2 12152 24248 12152 24248 0 _0773_
rlabel metal2 8456 23968 8456 23968 0 _0774_
rlabel metal3 13216 23912 13216 23912 0 _0775_
rlabel metal3 7952 26600 7952 26600 0 _0776_
rlabel metal2 11144 22512 11144 22512 0 _0777_
rlabel metal2 9688 22848 9688 22848 0 _0778_
rlabel metal2 8456 28728 8456 28728 0 _0779_
rlabel metal2 12152 23240 12152 23240 0 _0780_
rlabel metal2 6888 22624 6888 22624 0 _0781_
rlabel metal2 10304 25256 10304 25256 0 _0782_
rlabel metal3 5712 25256 5712 25256 0 _0783_
rlabel metal3 7672 30744 7672 30744 0 _0784_
rlabel metal3 9072 35672 9072 35672 0 _0785_
rlabel metal2 24808 37912 24808 37912 0 _0786_
rlabel metal2 27832 36904 27832 36904 0 _0787_
rlabel metal3 28672 34888 28672 34888 0 _0788_
rlabel metal2 33544 29400 33544 29400 0 _0789_
rlabel metal2 27608 36904 27608 36904 0 _0790_
rlabel metal2 28056 37744 28056 37744 0 _0791_
rlabel metal3 21168 31864 21168 31864 0 _0792_
rlabel metal2 23240 33264 23240 33264 0 _0793_
rlabel metal2 23464 32760 23464 32760 0 _0794_
rlabel metal2 24584 24752 24584 24752 0 _0795_
rlabel metal2 27944 32480 27944 32480 0 _0796_
rlabel metal3 25732 32536 25732 32536 0 _0797_
rlabel metal2 30184 29568 30184 29568 0 _0798_
rlabel metal2 28280 31024 28280 31024 0 _0799_
rlabel metal2 28056 31192 28056 31192 0 _0800_
rlabel metal2 28504 32984 28504 32984 0 _0801_
rlabel metal3 29232 35784 29232 35784 0 _0802_
rlabel metal3 13608 26376 13608 26376 0 _0803_
rlabel metal2 9520 26264 9520 26264 0 _0804_
rlabel metal2 12992 34888 12992 34888 0 _0805_
rlabel metal2 16744 33992 16744 33992 0 _0806_
rlabel metal2 17304 34552 17304 34552 0 _0807_
rlabel metal2 11312 36232 11312 36232 0 _0808_
rlabel metal2 15736 34216 15736 34216 0 _0809_
rlabel metal2 15624 34440 15624 34440 0 _0810_
rlabel metal2 9128 33432 9128 33432 0 _0811_
rlabel metal2 14392 25312 14392 25312 0 _0812_
rlabel metal2 18368 28392 18368 28392 0 _0813_
rlabel metal2 8120 25984 8120 25984 0 _0814_
rlabel metal2 9352 23072 9352 23072 0 _0815_
rlabel metal2 12712 23128 12712 23128 0 _0816_
rlabel metal2 4984 21448 4984 21448 0 _0817_
rlabel metal3 9632 34888 9632 34888 0 _0818_
rlabel metal3 21672 35000 21672 35000 0 _0819_
rlabel metal2 30184 37352 30184 37352 0 _0820_
rlabel metal3 29344 39480 29344 39480 0 _0821_
rlabel metal2 29512 32760 29512 32760 0 _0822_
rlabel metal2 28840 33544 28840 33544 0 _0823_
rlabel metal2 29736 39648 29736 39648 0 _0824_
rlabel metal2 10584 25032 10584 25032 0 _0825_
rlabel metal2 9016 33880 9016 33880 0 _0826_
rlabel metal2 11032 36736 11032 36736 0 _0827_
rlabel metal2 9016 34328 9016 34328 0 _0828_
rlabel metal3 11368 38024 11368 38024 0 _0829_
rlabel metal2 15176 38304 15176 38304 0 _0830_
rlabel metal2 4760 25424 4760 25424 0 _0831_
rlabel metal2 4872 27888 4872 27888 0 _0832_
rlabel metal2 12600 22344 12600 22344 0 _0833_
rlabel metal2 7056 25032 7056 25032 0 _0834_
rlabel metal3 7784 29176 7784 29176 0 _0835_
rlabel metal2 12040 25284 12040 25284 0 _0836_
rlabel metal3 10080 28392 10080 28392 0 _0837_
rlabel metal2 9800 25032 9800 25032 0 _0838_
rlabel metal2 10584 40376 10584 40376 0 _0839_
rlabel metal2 12376 33936 12376 33936 0 _0840_
rlabel metal2 15288 34776 15288 34776 0 _0841_
rlabel metal2 15624 26600 15624 26600 0 _0842_
rlabel metal2 17640 36064 17640 36064 0 _0843_
rlabel metal2 17304 36288 17304 36288 0 _0844_
rlabel metal2 11368 34048 11368 34048 0 _0845_
rlabel metal2 15288 35896 15288 35896 0 _0846_
rlabel metal2 13608 40488 13608 40488 0 _0847_
rlabel metal2 16072 39984 16072 39984 0 _0848_
rlabel metal3 29904 30072 29904 30072 0 _0849_
rlabel metal2 27944 28112 27944 28112 0 _0850_
rlabel metal2 25200 31864 25200 31864 0 _0851_
rlabel metal2 24808 29848 24808 29848 0 _0852_
rlabel metal2 25984 24920 25984 24920 0 _0853_
rlabel metal2 26712 29904 26712 29904 0 _0854_
rlabel metal2 23128 37968 23128 37968 0 _0855_
rlabel metal2 21560 36400 21560 36400 0 _0856_
rlabel metal2 20664 35504 20664 35504 0 _0857_
rlabel metal2 20776 34664 20776 34664 0 _0858_
rlabel metal2 22904 36064 22904 36064 0 _0859_
rlabel metal2 20328 36960 20328 36960 0 _0860_
rlabel metal2 21896 35896 21896 35896 0 _0861_
rlabel metal2 22120 38668 22120 38668 0 _0862_
rlabel metal3 18872 38696 18872 38696 0 _0863_
rlabel metal2 16632 39424 16632 39424 0 _0864_
rlabel metal2 28056 39984 28056 39984 0 _0865_
rlabel metal2 28952 39312 28952 39312 0 _0866_
rlabel metal2 28952 40488 28952 40488 0 _0867_
rlabel metal2 22344 39536 22344 39536 0 _0868_
rlabel metal3 23912 38808 23912 38808 0 _0869_
rlabel metal3 21112 38808 21112 38808 0 _0870_
rlabel metal2 22680 39256 22680 39256 0 _0871_
rlabel metal2 27160 40040 27160 40040 0 _0872_
rlabel metal2 25592 28280 25592 28280 0 _0873_
rlabel metal2 23688 28112 23688 28112 0 _0874_
rlabel metal2 24584 29456 24584 29456 0 _0875_
rlabel metal2 22456 39760 22456 39760 0 _0876_
rlabel metal2 21504 34664 21504 34664 0 _0877_
rlabel metal2 19432 34944 19432 34944 0 _0878_
rlabel metal2 14056 33656 14056 33656 0 _0879_
rlabel metal3 17360 34776 17360 34776 0 _0880_
rlabel metal2 19544 39816 19544 39816 0 _0881_
rlabel metal2 19656 38808 19656 38808 0 _0882_
rlabel metal2 9352 27160 9352 27160 0 _0883_
rlabel metal2 9408 24920 9408 24920 0 _0884_
rlabel metal2 11816 39312 11816 39312 0 _0885_
rlabel metal2 14112 39032 14112 39032 0 _0886_
rlabel metal2 11256 31360 11256 31360 0 _0887_
rlabel metal2 15848 35616 15848 35616 0 _0888_
rlabel metal3 11816 38864 11816 38864 0 _0889_
rlabel metal2 17976 39480 17976 39480 0 _0890_
rlabel metal2 9912 40488 9912 40488 0 _0891_
rlabel metal3 10864 40488 10864 40488 0 _0892_
rlabel metal2 14392 39200 14392 39200 0 _0893_
rlabel metal2 19544 39368 19544 39368 0 _0894_
rlabel metal2 20104 39760 20104 39760 0 _0895_
rlabel metal2 29064 40376 29064 40376 0 _0896_
rlabel metal2 27832 41216 27832 41216 0 _0897_
rlabel metal2 30184 41720 30184 41720 0 _0898_
rlabel metal2 21336 40432 21336 40432 0 _0899_
rlabel metal3 21000 42616 21000 42616 0 _0900_
rlabel metal2 17640 41440 17640 41440 0 _0901_
rlabel metal2 20888 40768 20888 40768 0 _0902_
rlabel metal2 27384 41104 27384 41104 0 _0903_
rlabel metal3 19992 37912 19992 37912 0 _0904_
rlabel metal2 23856 40488 23856 40488 0 _0905_
rlabel metal2 20664 31080 20664 31080 0 _0906_
rlabel metal2 24584 40656 24584 40656 0 _0907_
rlabel metal2 25536 41272 25536 41272 0 _0908_
rlabel metal2 11256 39984 11256 39984 0 _0909_
rlabel metal3 9352 40936 9352 40936 0 _0910_
rlabel metal2 11592 40824 11592 40824 0 _0911_
rlabel metal2 12600 40208 12600 40208 0 _0912_
rlabel metal2 2856 40096 2856 40096 0 _0913_
rlabel metal2 10920 40768 10920 40768 0 _0914_
rlabel metal2 11816 41104 11816 41104 0 _0915_
rlabel metal2 13944 40488 13944 40488 0 _0916_
rlabel metal2 25928 42112 25928 42112 0 _0917_
rlabel metal2 27440 42728 27440 42728 0 _0918_
rlabel metal2 29848 41888 29848 41888 0 _0919_
rlabel metal2 31080 43848 31080 43848 0 _0920_
rlabel metal3 28504 41944 28504 41944 0 _0921_
rlabel metal2 30856 44016 30856 44016 0 _0922_
rlabel metal2 25592 41888 25592 41888 0 _0923_
rlabel metal3 25032 41944 25032 41944 0 _0924_
rlabel metal2 26040 41664 26040 41664 0 _0925_
rlabel metal2 26488 42504 26488 42504 0 _0926_
rlabel metal2 23352 37016 23352 37016 0 _0927_
rlabel metal2 26376 42560 26376 42560 0 _0928_
rlabel metal2 21000 31360 21000 31360 0 _0929_
rlabel metal2 26712 43568 26712 43568 0 _0930_
rlabel metal2 26824 43652 26824 43652 0 _0931_
rlabel metal2 11816 42672 11816 42672 0 _0932_
rlabel metal2 12040 41608 12040 41608 0 _0933_
rlabel metal3 12320 33320 12320 33320 0 _0934_
rlabel metal2 10472 42504 10472 42504 0 _0935_
rlabel metal2 11144 29344 11144 29344 0 _0936_
rlabel metal2 7672 30240 7672 30240 0 _0937_
rlabel metal2 8008 29680 8008 29680 0 _0938_
rlabel metal2 10920 42448 10920 42448 0 _0939_
rlabel metal3 11984 42952 11984 42952 0 _0940_
rlabel metal2 12152 43960 12152 43960 0 _0941_
rlabel metal2 12768 42504 12768 42504 0 _0942_
rlabel metal2 27720 43904 27720 43904 0 _0943_
rlabel metal2 29400 44800 29400 44800 0 _0944_
rlabel metal2 30408 44296 30408 44296 0 _0945_
rlabel metal2 34776 44744 34776 44744 0 _0946_
rlabel metal3 22792 26488 22792 26488 0 _0947_
rlabel metal2 22232 28336 22232 28336 0 _0948_
rlabel metal3 23296 28728 23296 28728 0 _0949_
rlabel metal2 22960 30184 22960 30184 0 _0950_
rlabel metal2 22848 44072 22848 44072 0 _0951_
rlabel metal2 21448 28952 21448 28952 0 _0952_
rlabel metal3 21448 37240 21448 37240 0 _0953_
rlabel metal2 24696 36960 24696 36960 0 _0954_
rlabel metal2 21784 37016 21784 37016 0 _0955_
rlabel metal3 20552 35784 20552 35784 0 _0956_
rlabel metal2 22120 42728 22120 42728 0 _0957_
rlabel metal3 22288 46648 22288 46648 0 _0958_
rlabel metal3 15232 38024 15232 38024 0 _0959_
rlabel metal2 16520 36288 16520 36288 0 _0960_
rlabel metal2 17528 35504 17528 35504 0 _0961_
rlabel metal2 16520 39816 16520 39816 0 _0962_
rlabel metal2 18984 28504 18984 28504 0 _0963_
rlabel metal2 13160 22120 13160 22120 0 _0964_
rlabel metal2 12096 29400 12096 29400 0 _0965_
rlabel metal2 11144 44632 11144 44632 0 _0966_
rlabel metal3 13160 45864 13160 45864 0 _0967_
rlabel metal2 11480 43848 11480 43848 0 _0968_
rlabel metal2 12880 45752 12880 45752 0 _0969_
rlabel metal2 21336 46648 21336 46648 0 _0970_
rlabel metal2 29624 46480 29624 46480 0 _0971_
rlabel metal2 26600 45136 26600 45136 0 _0972_
rlabel metal2 27608 44856 27608 44856 0 _0973_
rlabel metal2 26600 43792 26600 43792 0 _0974_
rlabel metal2 30408 46032 30408 46032 0 _0975_
rlabel metal2 30744 47880 30744 47880 0 _0976_
rlabel metal2 29736 44296 29736 44296 0 _0977_
rlabel metal3 30800 45080 30800 45080 0 _0978_
rlabel metal2 29736 46088 29736 46088 0 _0979_
rlabel metal3 33600 47432 33600 47432 0 _0980_
rlabel metal2 29960 47488 29960 47488 0 _0981_
rlabel metal2 29512 47152 29512 47152 0 _0982_
rlabel metal2 24696 47040 24696 47040 0 _0983_
rlabel metal2 20216 46144 20216 46144 0 _0984_
rlabel metal2 23464 47264 23464 47264 0 _0985_
rlabel metal3 22624 47432 22624 47432 0 _0986_
rlabel metal2 27944 47936 27944 47936 0 _0987_
rlabel metal2 4984 29512 4984 29512 0 _0988_
rlabel metal2 9856 46536 9856 46536 0 _0989_
rlabel metal2 15456 35448 15456 35448 0 _0990_
rlabel metal2 10192 47320 10192 47320 0 _0991_
rlabel metal2 11368 46872 11368 46872 0 _0992_
rlabel metal2 10080 48776 10080 48776 0 _0993_
rlabel metal2 10584 47768 10584 47768 0 _0994_
rlabel metal3 12376 48328 12376 48328 0 _0995_
rlabel metal2 12152 47488 12152 47488 0 _0996_
rlabel metal2 9576 47488 9576 47488 0 _0997_
rlabel metal2 10696 46592 10696 46592 0 _0998_
rlabel metal3 11872 46760 11872 46760 0 _0999_
rlabel metal2 12376 46144 12376 46144 0 _1000_
rlabel metal2 12824 46704 12824 46704 0 _1001_
rlabel metal3 20244 49112 20244 49112 0 _1002_
rlabel metal2 21000 33152 21000 33152 0 _1003_
rlabel metal2 24528 49000 24528 49000 0 _1004_
rlabel metal2 20328 26096 20328 26096 0 _1005_
rlabel metal2 24696 47768 24696 47768 0 _1006_
rlabel metal2 26264 48440 26264 48440 0 _1007_
rlabel metal2 27944 49336 27944 49336 0 _1008_
rlabel metal3 30408 49000 30408 49000 0 _1009_
rlabel metal3 33320 49112 33320 49112 0 _1010_
rlabel metal2 30296 50960 30296 50960 0 _1011_
rlabel metal3 30520 50456 30520 50456 0 _1012_
rlabel metal2 33992 51016 33992 51016 0 _1013_
rlabel metal3 25424 48776 25424 48776 0 _1014_
rlabel metal2 26320 49000 26320 49000 0 _1015_
rlabel metal2 26488 49504 26488 49504 0 _1016_
rlabel metal3 29008 50456 29008 50456 0 _1017_
rlabel metal3 21896 45528 21896 45528 0 _1018_
rlabel metal2 21896 50904 21896 50904 0 _1019_
rlabel metal2 21336 40040 21336 40040 0 _1020_
rlabel metal2 22344 52640 22344 52640 0 _1021_
rlabel metal2 21336 51744 21336 51744 0 _1022_
rlabel metal2 21728 50456 21728 50456 0 _1023_
rlabel metal2 22680 52416 22680 52416 0 _1024_
rlabel metal3 12376 48776 12376 48776 0 _1025_
rlabel metal2 10360 54656 10360 54656 0 _1026_
rlabel metal3 12768 48888 12768 48888 0 _1027_
rlabel metal2 7672 44100 7672 44100 0 _1028_
rlabel metal2 3192 44912 3192 44912 0 _1029_
rlabel metal2 10528 44296 10528 44296 0 _1030_
rlabel metal2 9352 43120 9352 43120 0 _1031_
rlabel metal2 3304 42672 3304 42672 0 _1032_
rlabel metal2 10360 43904 10360 43904 0 _1033_
rlabel metal2 11928 47488 11928 47488 0 _1034_
rlabel metal2 12152 47992 12152 47992 0 _1035_
rlabel metal2 12656 48440 12656 48440 0 _1036_
rlabel metal2 22904 51464 22904 51464 0 _1037_
rlabel metal2 29288 52528 29288 52528 0 _1038_
rlabel metal2 34328 51968 34328 51968 0 _1039_
rlabel metal2 34664 51744 34664 51744 0 _1040_
rlabel metal3 30408 50792 30408 50792 0 _1041_
rlabel metal2 29624 52472 29624 52472 0 _1042_
rlabel metal2 31080 52192 31080 52192 0 _1043_
rlabel metal2 22792 51576 22792 51576 0 _1044_
rlabel metal2 23800 45920 23800 45920 0 _1045_
rlabel metal2 22456 45920 22456 45920 0 _1046_
rlabel metal3 24136 49896 24136 49896 0 _1047_
rlabel metal2 2128 50008 2128 50008 0 _1048_
rlabel metal2 13552 49560 13552 49560 0 _1049_
rlabel metal3 14504 50008 14504 50008 0 _1050_
rlabel metal2 16184 52920 16184 52920 0 _1051_
rlabel metal2 14560 50008 14560 50008 0 _1052_
rlabel metal2 15176 50148 15176 50148 0 _1053_
rlabel metal2 14840 50288 14840 50288 0 _1054_
rlabel metal3 7392 50344 7392 50344 0 _1055_
rlabel metal2 11704 48440 11704 48440 0 _1056_
rlabel metal2 12040 49168 12040 49168 0 _1057_
rlabel metal3 12824 50120 12824 50120 0 _1058_
rlabel metal3 19488 50568 19488 50568 0 _1059_
rlabel metal2 28952 50960 28952 50960 0 _1060_
rlabel metal3 30296 52808 30296 52808 0 _1061_
rlabel metal2 39480 53200 39480 53200 0 _1062_
rlabel metal2 22680 49392 22680 49392 0 _1063_
rlabel metal2 22120 48552 22120 48552 0 _1064_
rlabel metal2 23184 49896 23184 49896 0 _1065_
rlabel metal2 23576 49672 23576 49672 0 _1066_
rlabel metal2 23464 49616 23464 49616 0 _1067_
rlabel metal2 14392 49784 14392 49784 0 _1068_
rlabel metal3 21476 50680 21476 50680 0 _1069_
rlabel metal2 32312 50232 32312 50232 0 _1070_
rlabel metal2 28616 52192 28616 52192 0 _1071_
rlabel metal2 32144 49896 32144 49896 0 _1072_
rlabel metal2 44240 51352 44240 51352 0 _1073_
rlabel metal3 33040 50568 33040 50568 0 _1074_
rlabel metal2 43736 51520 43736 51520 0 _1075_
rlabel metal2 43960 44800 43960 44800 0 _1076_
rlabel metal2 44072 45136 44072 45136 0 _1077_
rlabel metal2 42392 44632 42392 44632 0 _1078_
rlabel metal2 41496 47768 41496 47768 0 _1079_
rlabel metal3 31136 12264 31136 12264 0 _1080_
rlabel metal2 24920 20776 24920 20776 0 _1081_
rlabel metal2 26600 21784 26600 21784 0 _1082_
rlabel metal2 22120 20776 22120 20776 0 _1083_
rlabel metal2 17752 22176 17752 22176 0 _1084_
rlabel metal2 22512 20664 22512 20664 0 _1085_
rlabel metal2 21896 20440 21896 20440 0 _1086_
rlabel metal2 27496 19264 27496 19264 0 _1087_
rlabel metal2 30800 12152 30800 12152 0 _1088_
rlabel metal2 29176 11704 29176 11704 0 _1089_
rlabel metal2 30968 12040 30968 12040 0 _1090_
rlabel metal3 32368 23912 32368 23912 0 _1091_
rlabel metal2 21672 23968 21672 23968 0 _1092_
rlabel metal2 24248 23688 24248 23688 0 _1093_
rlabel metal2 47544 11256 47544 11256 0 _1094_
rlabel metal2 25928 21056 25928 21056 0 _1095_
rlabel metal2 41160 19880 41160 19880 0 _1096_
rlabel metal3 21616 15960 21616 15960 0 _1097_
rlabel metal2 36736 17192 36736 17192 0 _1098_
rlabel metal2 40824 10640 40824 10640 0 _1099_
rlabel metal2 31416 10696 31416 10696 0 _1100_
rlabel metal2 17640 22456 17640 22456 0 _1101_
rlabel metal2 41160 21056 41160 21056 0 _1102_
rlabel metal2 29792 10584 29792 10584 0 _1103_
rlabel metal2 16240 21560 16240 21560 0 _1104_
rlabel metal2 39480 10976 39480 10976 0 _1105_
rlabel metal2 29288 11032 29288 11032 0 _1106_
rlabel metal3 43680 11144 43680 11144 0 _1107_
rlabel metal2 26152 21336 26152 21336 0 _1108_
rlabel metal2 31416 21616 31416 21616 0 _1109_
rlabel metal2 39368 13160 39368 13160 0 _1110_
rlabel metal2 41160 11424 41160 11424 0 _1111_
rlabel metal2 40040 11816 40040 11816 0 _1112_
rlabel metal2 42280 10864 42280 10864 0 _1113_
rlabel metal3 40824 10584 40824 10584 0 _1114_
rlabel metal2 42280 19824 42280 19824 0 _1115_
rlabel metal3 42616 11256 42616 11256 0 _1116_
rlabel metal2 39536 11368 39536 11368 0 _1117_
rlabel metal2 42952 20496 42952 20496 0 _1118_
rlabel metal3 25004 21672 25004 21672 0 _1119_
rlabel metal2 38808 20132 38808 20132 0 _1120_
rlabel metal2 40824 21112 40824 21112 0 _1121_
rlabel metal3 41608 22176 41608 22176 0 _1122_
rlabel metal2 43064 21392 43064 21392 0 _1123_
rlabel metal3 41664 19992 41664 19992 0 _1124_
rlabel metal2 41608 21672 41608 21672 0 _1125_
rlabel metal2 8456 32368 8456 32368 0 _1126_
rlabel metal2 16800 40376 16800 40376 0 _1127_
rlabel metal2 39368 21224 39368 21224 0 _1128_
rlabel metal2 31584 34216 31584 34216 0 _1129_
rlabel metal2 40824 43988 40824 43988 0 _1130_
rlabel metal2 38864 34776 38864 34776 0 _1131_
rlabel metal2 44184 20328 44184 20328 0 _1132_
rlabel metal2 31080 33600 31080 33600 0 _1133_
rlabel metal2 31920 32424 31920 32424 0 _1134_
rlabel metal2 30184 33712 30184 33712 0 _1135_
rlabel metal2 29624 33712 29624 33712 0 _1136_
rlabel metal2 20216 37800 20216 37800 0 _1137_
rlabel metal2 18592 37240 18592 37240 0 _1138_
rlabel metal2 18424 36792 18424 36792 0 _1139_
rlabel metal2 38416 38920 38416 38920 0 _1140_
rlabel metal2 18536 39088 18536 39088 0 _1141_
rlabel metal2 18312 40488 18312 40488 0 _1142_
rlabel metal2 18816 38808 18816 38808 0 _1143_
rlabel metal3 19040 37464 19040 37464 0 _1144_
rlabel metal2 17920 40376 17920 40376 0 _1145_
rlabel metal2 18760 41328 18760 41328 0 _1146_
rlabel metal2 17752 41104 17752 41104 0 _1147_
rlabel metal2 19096 41048 19096 41048 0 _1148_
rlabel metal2 16184 40712 16184 40712 0 _1149_
rlabel metal2 16408 41272 16408 41272 0 _1150_
rlabel metal2 15288 41440 15288 41440 0 _1151_
rlabel metal2 15848 41160 15848 41160 0 _1152_
rlabel metal2 15064 43120 15064 43120 0 _1153_
rlabel metal2 15624 43008 15624 43008 0 _1154_
rlabel metal2 15624 46256 15624 46256 0 _1155_
rlabel metal3 16296 43456 16296 43456 0 _1156_
rlabel metal2 2632 42448 2632 42448 0 _1157_
rlabel metal2 16408 43652 16408 43652 0 _1158_
rlabel metal2 16352 45080 16352 45080 0 _1159_
rlabel metal2 16352 44856 16352 44856 0 _1160_
rlabel metal2 19208 45472 19208 45472 0 _1161_
rlabel metal2 20328 43680 20328 43680 0 _1162_
rlabel metal2 18760 46648 18760 46648 0 _1163_
rlabel metal2 19656 46144 19656 46144 0 _1164_
rlabel metal3 20496 47432 20496 47432 0 _1165_
rlabel metal2 18648 47880 18648 47880 0 _1166_
rlabel metal2 19656 48328 19656 48328 0 _1167_
rlabel metal2 20552 48104 20552 48104 0 _1168_
rlabel metal2 19432 48860 19432 48860 0 _1169_
rlabel metal2 18760 51016 18760 51016 0 _1170_
rlabel metal2 2968 34720 2968 34720 0 _1171_
rlabel metal2 19656 52080 19656 52080 0 _1172_
rlabel metal2 19432 51240 19432 51240 0 _1173_
rlabel metal2 20552 51016 20552 51016 0 _1174_
rlabel metal2 18760 49672 18760 49672 0 _1175_
rlabel metal2 16072 47152 16072 47152 0 _1176_
rlabel metal2 15736 47992 15736 47992 0 _1177_
rlabel metal2 16744 48664 16744 48664 0 _1178_
rlabel metal2 3304 30912 3304 30912 0 _1179_
rlabel metal2 2968 31136 2968 31136 0 _1180_
rlabel metal2 3752 32480 3752 32480 0 _1181_
rlabel metal2 3640 32368 3640 32368 0 _1182_
rlabel metal3 3136 33432 3136 33432 0 _1183_
rlabel metal2 3304 33992 3304 33992 0 _1184_
rlabel metal2 2968 35504 2968 35504 0 _1185_
rlabel metal2 2856 37296 2856 37296 0 _1186_
rlabel metal2 4200 37408 4200 37408 0 _1187_
rlabel metal2 3080 36288 3080 36288 0 _1188_
rlabel metal2 2632 35336 2632 35336 0 _1189_
rlabel metal2 4928 36680 4928 36680 0 _1190_
rlabel metal2 3808 39592 3808 39592 0 _1191_
rlabel metal2 4088 38136 4088 38136 0 _1192_
rlabel metal2 3640 39648 3640 39648 0 _1193_
rlabel metal2 4536 39704 4536 39704 0 _1194_
rlabel metal2 3976 41160 3976 41160 0 _1195_
rlabel metal2 4312 43568 4312 43568 0 _1196_
rlabel metal2 2856 42560 2856 42560 0 _1197_
rlabel metal2 3640 42728 3640 42728 0 _1198_
rlabel metal3 5040 42728 5040 42728 0 _1199_
rlabel metal2 4872 42952 4872 42952 0 _1200_
rlabel metal2 3304 45360 3304 45360 0 _1201_
rlabel metal2 2352 45192 2352 45192 0 _1202_
rlabel metal2 5824 44072 5824 44072 0 _1203_
rlabel metal2 2856 45528 2856 45528 0 _1204_
rlabel metal2 4760 45808 4760 45808 0 _1205_
rlabel metal3 4256 45752 4256 45752 0 _1206_
rlabel metal3 2800 48216 2800 48216 0 _1207_
rlabel metal2 2800 48216 2800 48216 0 _1208_
rlabel metal2 2184 48328 2184 48328 0 _1209_
rlabel metal2 17192 39200 17192 39200 0 _1210_
rlabel metal2 17416 39816 17416 39816 0 _1211_
rlabel metal2 4536 46928 4536 46928 0 _1212_
rlabel metal2 4536 46424 4536 46424 0 _1213_
rlabel metal2 6328 47936 6328 47936 0 _1214_
rlabel metal2 7336 49448 7336 49448 0 _1215_
rlabel metal2 5880 49728 5880 49728 0 _1216_
rlabel metal3 5152 49000 5152 49000 0 _1217_
rlabel via2 5992 51352 5992 51352 0 _1218_
rlabel metal2 7560 51856 7560 51856 0 _1219_
rlabel metal3 5992 51576 5992 51576 0 _1220_
rlabel metal2 5656 51800 5656 51800 0 _1221_
rlabel metal2 6944 52136 6944 52136 0 _1222_
rlabel metal2 7224 52248 7224 52248 0 _1223_
rlabel metal2 15400 52696 15400 52696 0 _1224_
rlabel metal2 16520 50960 16520 50960 0 _1225_
rlabel metal2 15848 53424 15848 53424 0 _1226_
rlabel metal2 33880 21448 33880 21448 0 _1227_
rlabel metal2 1624 35896 1624 35896 0 _1228_
rlabel metal2 16408 53368 16408 53368 0 _1229_
rlabel metal2 7560 32312 7560 32312 0 _1230_
rlabel metal2 6216 31528 6216 31528 0 _1231_
rlabel metal2 6440 34216 6440 34216 0 _1232_
rlabel metal2 4368 35112 4368 35112 0 _1233_
rlabel metal3 5432 34888 5432 34888 0 _1234_
rlabel metal2 7224 34608 7224 34608 0 _1235_
rlabel metal2 6552 36568 6552 36568 0 _1236_
rlabel metal2 6216 37296 6216 37296 0 _1237_
rlabel metal2 7336 44184 7336 44184 0 _1238_
rlabel metal2 7112 38024 7112 38024 0 _1239_
rlabel metal2 8848 40152 8848 40152 0 _1240_
rlabel metal2 8680 37464 8680 37464 0 _1241_
rlabel metal2 9576 39200 9576 39200 0 _1242_
rlabel metal2 6552 39144 6552 39144 0 _1243_
rlabel metal3 8848 38696 8848 38696 0 _1244_
rlabel metal3 8904 40152 8904 40152 0 _1245_
rlabel metal2 8120 43288 8120 43288 0 _1246_
rlabel metal2 8120 41944 8120 41944 0 _1247_
rlabel metal2 6552 41888 6552 41888 0 _1248_
rlabel metal2 5768 42672 5768 42672 0 _1249_
rlabel metal2 9016 43120 9016 43120 0 _1250_
rlabel metal2 7784 43120 7784 43120 0 _1251_
rlabel metal2 8400 45192 8400 45192 0 _1252_
rlabel via2 6440 45640 6440 45640 0 _1253_
rlabel metal2 6776 45864 6776 45864 0 _1254_
rlabel metal2 7840 44520 7840 44520 0 _1255_
rlabel metal2 8120 45528 8120 45528 0 _1256_
rlabel metal3 8008 47432 8008 47432 0 _1257_
rlabel metal2 7784 47320 7784 47320 0 _1258_
rlabel metal2 40376 46200 40376 46200 0 clknet_0_wb_clk_i
rlabel metal2 15064 10304 15064 10304 0 clknet_4_0_0_wb_clk_i
rlabel metal2 1848 48608 1848 48608 0 clknet_4_10_0_wb_clk_i
rlabel metal2 17584 48216 17584 48216 0 clknet_4_11_0_wb_clk_i
rlabel metal2 38920 41104 38920 41104 0 clknet_4_12_0_wb_clk_i
rlabel metal2 45416 40768 45416 40768 0 clknet_4_13_0_wb_clk_i
rlabel metal2 38696 44688 38696 44688 0 clknet_4_14_0_wb_clk_i
rlabel metal2 48104 54488 48104 54488 0 clknet_4_15_0_wb_clk_i
rlabel metal2 24584 12208 24584 12208 0 clknet_4_1_0_wb_clk_i
rlabel metal2 15400 25872 15400 25872 0 clknet_4_2_0_wb_clk_i
rlabel metal2 17080 18928 17080 18928 0 clknet_4_3_0_wb_clk_i
rlabel metal2 39256 15848 39256 15848 0 clknet_4_4_0_wb_clk_i
rlabel metal2 46760 16240 46760 16240 0 clknet_4_5_0_wb_clk_i
rlabel metal2 40992 22456 40992 22456 0 clknet_4_6_0_wb_clk_i
rlabel metal2 47768 23968 47768 23968 0 clknet_4_7_0_wb_clk_i
rlabel metal2 1848 36568 1848 36568 0 clknet_4_8_0_wb_clk_i
rlabel metal2 1848 30576 1848 30576 0 clknet_4_9_0_wb_clk_i
rlabel metal2 48272 48776 48272 48776 0 custom_settings[0]
rlabel metal3 46088 53480 46088 53480 0 custom_settings[1]
rlabel metal3 48818 3640 48818 3640 0 io_in_1[0]
rlabel metal2 48216 9576 48216 9576 0 io_in_1[1]
rlabel metal2 48216 15624 48216 15624 0 io_in_1[2]
rlabel metal2 48216 21336 48216 21336 0 io_in_1[3]
rlabel metal3 48818 26936 48818 26936 0 io_in_1[4]
rlabel metal2 48216 32928 48216 32928 0 io_in_1[5]
rlabel metal2 48216 39032 48216 39032 0 io_in_1[6]
rlabel metal3 48762 44408 48762 44408 0 io_in_1[7]
rlabel metal2 1736 50120 1736 50120 0 io_in_2
rlabel metal2 19320 56210 19320 56210 0 io_out[10]
rlabel metal2 20888 57778 20888 57778 0 io_out[11]
rlabel metal2 22456 57722 22456 57722 0 io_out[12]
rlabel metal2 30240 55944 30240 55944 0 io_out[17]
rlabel metal2 31864 57330 31864 57330 0 io_out[18]
rlabel metal2 33432 56378 33432 56378 0 io_out[19]
rlabel metal2 35000 56938 35000 56938 0 io_out[20]
rlabel metal2 36568 57778 36568 57778 0 io_out[21]
rlabel metal2 44632 56672 44632 56672 0 io_out[22]
rlabel metal3 40880 53144 40880 53144 0 io_out[23]
rlabel metal2 41440 54152 41440 54152 0 io_out[24]
rlabel metal3 44632 54712 44632 54712 0 io_out[25]
rlabel metal2 45416 53144 45416 53144 0 io_out[26]
rlabel metal2 46312 52360 46312 52360 0 io_out[27]
rlabel metal3 15792 56280 15792 56280 0 io_out[8]
rlabel metal2 17752 57778 17752 57778 0 io_out[9]
rlabel metal3 47040 49000 47040 49000 0 net1
rlabel metal3 46368 45528 46368 45528 0 net10
rlabel metal3 1904 48776 1904 48776 0 net11
rlabel metal2 2296 28448 2296 28448 0 net12
rlabel metal2 19880 55496 19880 55496 0 net13
rlabel metal2 20776 55720 20776 55720 0 net14
rlabel metal3 44492 55384 44492 55384 0 net15
rlabel metal2 41328 46536 41328 46536 0 net16
rlabel metal2 32872 55328 32872 55328 0 net17
rlabel metal2 32200 55720 32200 55720 0 net18
rlabel metal4 38696 52920 38696 52920 0 net19
rlabel metal2 45640 53368 45640 53368 0 net2
rlabel metal2 38808 47936 38808 47936 0 net20
rlabel metal2 44408 51296 44408 51296 0 net21
rlabel metal3 40320 51576 40320 51576 0 net22
rlabel metal2 40264 52808 40264 52808 0 net23
rlabel metal2 42504 54768 42504 54768 0 net24
rlabel metal2 45080 50344 45080 50344 0 net25
rlabel metal2 45192 51688 45192 51688 0 net26
rlabel metal2 16072 55216 16072 55216 0 net27
rlabel metal2 17528 54544 17528 54544 0 net28
rlabel metal2 3752 56280 3752 56280 0 net29
rlabel metal2 42616 21896 42616 21896 0 net3
rlabel metal2 5544 57008 5544 57008 0 net30
rlabel metal2 6888 56280 6888 56280 0 net31
rlabel metal2 8456 56280 8456 56280 0 net32
rlabel metal2 10024 56280 10024 56280 0 net33
rlabel metal2 11592 56280 11592 56280 0 net34
rlabel metal2 12600 57008 12600 57008 0 net35
rlabel metal2 13496 56672 13496 56672 0 net36
rlabel metal2 23800 54264 23800 54264 0 net37
rlabel metal2 25592 57778 25592 57778 0 net38
rlabel metal2 28392 56672 28392 56672 0 net39
rlabel metal2 47880 10080 47880 10080 0 net4
rlabel metal2 29176 56224 29176 56224 0 net40
rlabel metal2 48216 55384 48216 55384 0 net41
rlabel metal2 10024 35672 10024 35672 0 net42
rlabel metal2 24080 37912 24080 37912 0 net43
rlabel metal2 15344 40264 15344 40264 0 net44
rlabel metal2 15848 39536 15848 39536 0 net45
rlabel metal2 11928 36904 11928 36904 0 net46
rlabel metal2 14504 36176 14504 36176 0 net47
rlabel metal2 12376 37296 12376 37296 0 net48
rlabel metal2 17416 36120 17416 36120 0 net49
rlabel metal2 47880 16072 47880 16072 0 net5
rlabel metal2 31584 50792 31584 50792 0 net50
rlabel metal2 30968 37968 30968 37968 0 net51
rlabel metal2 44856 52640 44856 52640 0 net52
rlabel metal2 7560 34384 7560 34384 0 net53
rlabel metal2 8344 35896 8344 35896 0 net54
rlabel metal2 12824 39144 12824 39144 0 net55
rlabel metal2 12376 40824 12376 40824 0 net56
rlabel metal2 2744 33824 2744 33824 0 net57
rlabel metal2 2632 32424 2632 32424 0 net58
rlabel metal2 21784 39536 21784 39536 0 net59
rlabel metal2 47880 20888 47880 20888 0 net6
rlabel metal2 9968 31192 9968 31192 0 net60
rlabel metal2 43624 51688 43624 51688 0 net61
rlabel metal3 29064 49784 29064 49784 0 net62
rlabel metal2 12208 41160 12208 41160 0 net63
rlabel metal2 29512 29008 29512 29008 0 net64
rlabel metal2 20888 30744 20888 30744 0 net65
rlabel metal3 29232 30184 29232 30184 0 net66
rlabel metal3 12040 32648 12040 32648 0 net67
rlabel metal3 13104 38808 13104 38808 0 net68
rlabel metal2 17416 28280 17416 28280 0 net69
rlabel metal3 26712 21504 26712 21504 0 net7
rlabel metal2 30128 45752 30128 45752 0 net70
rlabel metal2 25200 20776 25200 20776 0 net8
rlabel metal3 45472 39592 45472 39592 0 net9
rlabel metal2 1736 29736 1736 29736 0 rst_n
rlabel metal2 16408 22400 16408 22400 0 tt_um_rejunity_sn76489.chan\[0\].attenuation.control\[0\]
rlabel metal3 17416 29344 17416 29344 0 tt_um_rejunity_sn76489.chan\[0\].attenuation.control\[1\]
rlabel metal2 16632 26152 16632 26152 0 tt_um_rejunity_sn76489.chan\[0\].attenuation.control\[2\]
rlabel metal2 16296 20104 16296 20104 0 tt_um_rejunity_sn76489.chan\[0\].attenuation.control\[3\]
rlabel metal2 14168 29064 14168 29064 0 tt_um_rejunity_sn76489.chan\[0\].attenuation.in
rlabel metal3 3276 24584 3276 24584 0 tt_um_rejunity_sn76489.chan\[1\].attenuation.control\[0\]
rlabel metal2 4984 22680 4984 22680 0 tt_um_rejunity_sn76489.chan\[1\].attenuation.control\[1\]
rlabel metal2 8232 23184 8232 23184 0 tt_um_rejunity_sn76489.chan\[1\].attenuation.control\[2\]
rlabel metal2 5768 19488 5768 19488 0 tt_um_rejunity_sn76489.chan\[1\].attenuation.control\[3\]
rlabel metal2 10248 18816 10248 18816 0 tt_um_rejunity_sn76489.chan\[1\].attenuation.in
rlabel metal2 18368 25592 18368 25592 0 tt_um_rejunity_sn76489.chan\[2\].attenuation.control\[0\]
rlabel metal2 19208 27636 19208 27636 0 tt_um_rejunity_sn76489.chan\[2\].attenuation.control\[1\]
rlabel metal2 21000 29456 21000 29456 0 tt_um_rejunity_sn76489.chan\[2\].attenuation.control\[2\]
rlabel metal2 15960 24416 15960 24416 0 tt_um_rejunity_sn76489.chan\[2\].attenuation.control\[3\]
rlabel metal2 19320 27720 19320 27720 0 tt_um_rejunity_sn76489.chan\[2\].attenuation.in
rlabel metal2 27720 25872 27720 25872 0 tt_um_rejunity_sn76489.chan\[3\].attenuation.control\[0\]
rlabel metal2 26824 25312 26824 25312 0 tt_um_rejunity_sn76489.chan\[3\].attenuation.control\[1\]
rlabel metal2 24360 28000 24360 28000 0 tt_um_rejunity_sn76489.chan\[3\].attenuation.control\[2\]
rlabel metal2 23240 23408 23240 23408 0 tt_um_rejunity_sn76489.chan\[3\].attenuation.control\[3\]
rlabel metal3 35224 26600 35224 26600 0 tt_um_rejunity_sn76489.chan\[3\].attenuation.in
rlabel metal3 47600 36232 47600 36232 0 tt_um_rejunity_sn76489.clk_counter\[0\]
rlabel metal2 47432 39200 47432 39200 0 tt_um_rejunity_sn76489.clk_counter\[1\]
rlabel metal3 46144 39480 46144 39480 0 tt_um_rejunity_sn76489.clk_counter\[2\]
rlabel metal3 46368 38808 46368 38808 0 tt_um_rejunity_sn76489.clk_counter\[3\]
rlabel metal2 42616 39480 42616 39480 0 tt_um_rejunity_sn76489.clk_counter\[4\]
rlabel metal2 42952 39088 42952 39088 0 tt_um_rejunity_sn76489.clk_counter\[5\]
rlabel metal2 42952 36456 42952 36456 0 tt_um_rejunity_sn76489.clk_counter\[6\]
rlabel metal3 30688 23016 30688 23016 0 tt_um_rejunity_sn76489.control_noise\[0\]\[0\]
rlabel metal2 33656 25648 33656 25648 0 tt_um_rejunity_sn76489.control_noise\[0\]\[1\]
rlabel metal2 32088 26264 32088 26264 0 tt_um_rejunity_sn76489.control_noise\[0\]\[2\]
rlabel metal2 30520 9940 30520 9940 0 tt_um_rejunity_sn76489.control_tone_freq\[0\]\[0\]
rlabel metal2 32424 9968 32424 9968 0 tt_um_rejunity_sn76489.control_tone_freq\[0\]\[1\]
rlabel metal2 29624 8960 29624 8960 0 tt_um_rejunity_sn76489.control_tone_freq\[0\]\[2\]
rlabel metal2 28728 10472 28728 10472 0 tt_um_rejunity_sn76489.control_tone_freq\[0\]\[3\]
rlabel metal3 21504 8232 21504 8232 0 tt_um_rejunity_sn76489.control_tone_freq\[0\]\[4\]
rlabel metal3 21056 7448 21056 7448 0 tt_um_rejunity_sn76489.control_tone_freq\[0\]\[5\]
rlabel metal2 17864 9464 17864 9464 0 tt_um_rejunity_sn76489.control_tone_freq\[0\]\[6\]
rlabel metal3 20496 11480 20496 11480 0 tt_um_rejunity_sn76489.control_tone_freq\[0\]\[7\]
rlabel metal2 18032 13720 18032 13720 0 tt_um_rejunity_sn76489.control_tone_freq\[0\]\[8\]
rlabel metal2 18200 14280 18200 14280 0 tt_um_rejunity_sn76489.control_tone_freq\[0\]\[9\]
rlabel metal2 45416 10416 45416 10416 0 tt_um_rejunity_sn76489.control_tone_freq\[1\]\[0\]
rlabel metal2 42504 9128 42504 9128 0 tt_um_rejunity_sn76489.control_tone_freq\[1\]\[1\]
rlabel metal2 43624 10360 43624 10360 0 tt_um_rejunity_sn76489.control_tone_freq\[1\]\[2\]
rlabel metal2 40096 9912 40096 9912 0 tt_um_rejunity_sn76489.control_tone_freq\[1\]\[3\]
rlabel metal2 21560 6328 21560 6328 0 tt_um_rejunity_sn76489.control_tone_freq\[1\]\[4\]
rlabel metal3 21896 4984 21896 4984 0 tt_um_rejunity_sn76489.control_tone_freq\[1\]\[5\]
rlabel metal2 22120 7560 22120 7560 0 tt_um_rejunity_sn76489.control_tone_freq\[1\]\[6\]
rlabel metal2 22120 10360 22120 10360 0 tt_um_rejunity_sn76489.control_tone_freq\[1\]\[7\]
rlabel metal2 24248 13272 24248 13272 0 tt_um_rejunity_sn76489.control_tone_freq\[1\]\[8\]
rlabel metal2 23016 15260 23016 15260 0 tt_um_rejunity_sn76489.control_tone_freq\[1\]\[9\]
rlabel metal2 44744 21056 44744 21056 0 tt_um_rejunity_sn76489.control_tone_freq\[2\]\[0\]
rlabel metal2 42392 19600 42392 19600 0 tt_um_rejunity_sn76489.control_tone_freq\[2\]\[1\]
rlabel metal2 43792 23016 43792 23016 0 tt_um_rejunity_sn76489.control_tone_freq\[2\]\[2\]
rlabel via2 40264 20552 40264 20552 0 tt_um_rejunity_sn76489.control_tone_freq\[2\]\[3\]
rlabel metal2 42056 17304 42056 17304 0 tt_um_rejunity_sn76489.control_tone_freq\[2\]\[4\]
rlabel metal2 32312 16464 32312 16464 0 tt_um_rejunity_sn76489.control_tone_freq\[2\]\[5\]
rlabel metal2 28392 17192 28392 17192 0 tt_um_rejunity_sn76489.control_tone_freq\[2\]\[6\]
rlabel metal2 28952 18144 28952 18144 0 tt_um_rejunity_sn76489.control_tone_freq\[2\]\[7\]
rlabel metal2 28168 17976 28168 17976 0 tt_um_rejunity_sn76489.control_tone_freq\[2\]\[8\]
rlabel metal2 24696 18088 24696 18088 0 tt_um_rejunity_sn76489.control_tone_freq\[2\]\[9\]
rlabel metal2 6216 32144 6216 32144 0 tt_um_rejunity_sn76489.genblk4\[0\].pwm.accumulator\[0\]
rlabel via2 7000 34328 7000 34328 0 tt_um_rejunity_sn76489.genblk4\[0\].pwm.accumulator\[1\]
rlabel metal2 8512 39928 8512 39928 0 tt_um_rejunity_sn76489.genblk4\[0\].pwm.accumulator\[2\]
rlabel metal2 8568 39592 8568 39592 0 tt_um_rejunity_sn76489.genblk4\[0\].pwm.accumulator\[3\]
rlabel metal3 8960 41832 8960 41832 0 tt_um_rejunity_sn76489.genblk4\[0\].pwm.accumulator\[4\]
rlabel metal2 7784 44016 7784 44016 0 tt_um_rejunity_sn76489.genblk4\[0\].pwm.accumulator\[5\]
rlabel metal2 8680 48216 8680 48216 0 tt_um_rejunity_sn76489.genblk4\[0\].pwm.accumulator\[6\]
rlabel metal2 9016 51184 9016 51184 0 tt_um_rejunity_sn76489.genblk4\[0\].pwm.accumulator\[7\]
rlabel metal2 9800 53816 9800 53816 0 tt_um_rejunity_sn76489.genblk4\[0\].pwm.accumulator\[8\]
rlabel metal3 13328 53592 13328 53592 0 tt_um_rejunity_sn76489.genblk4\[0\].pwm.accumulator\[9\]
rlabel metal2 4424 31136 4424 31136 0 tt_um_rejunity_sn76489.genblk4\[1\].pwm.accumulator\[0\]
rlabel metal2 2072 31780 2072 31780 0 tt_um_rejunity_sn76489.genblk4\[1\].pwm.accumulator\[1\]
rlabel metal2 4480 36568 4480 36568 0 tt_um_rejunity_sn76489.genblk4\[1\].pwm.accumulator\[2\]
rlabel metal2 3080 39984 3080 39984 0 tt_um_rejunity_sn76489.genblk4\[1\].pwm.accumulator\[3\]
rlabel metal2 4424 41160 4424 41160 0 tt_um_rejunity_sn76489.genblk4\[1\].pwm.accumulator\[4\]
rlabel metal2 3080 45024 3080 45024 0 tt_um_rejunity_sn76489.genblk4\[1\].pwm.accumulator\[5\]
rlabel metal2 3304 47040 3304 47040 0 tt_um_rejunity_sn76489.genblk4\[1\].pwm.accumulator\[6\]
rlabel metal3 5152 49672 5152 49672 0 tt_um_rejunity_sn76489.genblk4\[1\].pwm.accumulator\[7\]
rlabel metal2 8232 52472 8232 52472 0 tt_um_rejunity_sn76489.genblk4\[1\].pwm.accumulator\[8\]
rlabel metal3 16128 52920 16128 52920 0 tt_um_rejunity_sn76489.genblk4\[1\].pwm.accumulator\[9\]
rlabel metal2 31304 34944 31304 34944 0 tt_um_rejunity_sn76489.genblk4\[2\].pwm.accumulator\[0\]
rlabel metal2 30184 32256 30184 32256 0 tt_um_rejunity_sn76489.genblk4\[2\].pwm.accumulator\[1\]
rlabel metal2 18088 37240 18088 37240 0 tt_um_rejunity_sn76489.genblk4\[2\].pwm.accumulator\[2\]
rlabel metal2 17752 42056 17752 42056 0 tt_um_rejunity_sn76489.genblk4\[2\].pwm.accumulator\[3\]
rlabel metal2 16296 40936 16296 40936 0 tt_um_rejunity_sn76489.genblk4\[2\].pwm.accumulator\[4\]
rlabel metal2 16128 45864 16128 45864 0 tt_um_rejunity_sn76489.genblk4\[2\].pwm.accumulator\[5\]
rlabel metal2 20272 44968 20272 44968 0 tt_um_rejunity_sn76489.genblk4\[2\].pwm.accumulator\[6\]
rlabel metal2 20328 48216 20328 48216 0 tt_um_rejunity_sn76489.genblk4\[2\].pwm.accumulator\[7\]
rlabel metal2 20328 51128 20328 51128 0 tt_um_rejunity_sn76489.genblk4\[2\].pwm.accumulator\[8\]
rlabel metal2 16576 48216 16576 48216 0 tt_um_rejunity_sn76489.genblk4\[2\].pwm.accumulator\[9\]
rlabel metal2 34216 28896 34216 28896 0 tt_um_rejunity_sn76489.genblk4\[3\].pwm.accumulator\[0\]
rlabel metal2 35896 33040 35896 33040 0 tt_um_rejunity_sn76489.genblk4\[3\].pwm.accumulator\[1\]
rlabel metal2 24024 39144 24024 39144 0 tt_um_rejunity_sn76489.genblk4\[3\].pwm.accumulator\[2\]
rlabel metal2 21672 42224 21672 42224 0 tt_um_rejunity_sn76489.genblk4\[3\].pwm.accumulator\[3\]
rlabel metal2 25256 43652 25256 43652 0 tt_um_rejunity_sn76489.genblk4\[3\].pwm.accumulator\[4\]
rlabel metal2 27440 46648 27440 46648 0 tt_um_rejunity_sn76489.genblk4\[3\].pwm.accumulator\[5\]
rlabel metal3 27608 51464 27608 51464 0 tt_um_rejunity_sn76489.genblk4\[3\].pwm.accumulator\[6\]
rlabel metal2 28056 54432 28056 54432 0 tt_um_rejunity_sn76489.genblk4\[3\].pwm.accumulator\[7\]
rlabel metal2 25816 54936 25816 54936 0 tt_um_rejunity_sn76489.genblk4\[3\].pwm.accumulator\[8\]
rlabel metal2 22568 54040 22568 54040 0 tt_um_rejunity_sn76489.genblk4\[3\].pwm.accumulator\[9\]
rlabel metal2 19208 19824 19208 19824 0 tt_um_rejunity_sn76489.latch_control_reg\[0\]
rlabel metal3 17752 16968 17752 16968 0 tt_um_rejunity_sn76489.latch_control_reg\[1\]
rlabel metal2 17752 21056 17752 21056 0 tt_um_rejunity_sn76489.latch_control_reg\[2\]
rlabel metal2 36064 24584 36064 24584 0 tt_um_rejunity_sn76489.noise\[0\].gen.counter\[0\]
rlabel metal3 36176 24584 36176 24584 0 tt_um_rejunity_sn76489.noise\[0\].gen.counter\[1\]
rlabel metal2 36008 26712 36008 26712 0 tt_um_rejunity_sn76489.noise\[0\].gen.counter\[2\]
rlabel metal2 36176 27720 36176 27720 0 tt_um_rejunity_sn76489.noise\[0\].gen.counter\[3\]
rlabel metal2 38808 31024 38808 31024 0 tt_um_rejunity_sn76489.noise\[0\].gen.counter\[4\]
rlabel metal2 37016 32312 37016 32312 0 tt_um_rejunity_sn76489.noise\[0\].gen.counter\[5\]
rlabel metal2 35560 30520 35560 30520 0 tt_um_rejunity_sn76489.noise\[0\].gen.counter\[6\]
rlabel metal3 45304 33208 45304 33208 0 tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[10\]
rlabel metal2 43848 34048 43848 34048 0 tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[11\]
rlabel metal2 44184 31920 44184 31920 0 tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[12\]
rlabel metal2 43848 29960 43848 29960 0 tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[13\]
rlabel via2 42504 27944 42504 27944 0 tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[14\]
rlabel metal3 40712 25480 40712 25480 0 tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[1\]
rlabel metal2 45080 24416 45080 24416 0 tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[2\]
rlabel metal2 44744 22904 44744 22904 0 tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[3\]
rlabel metal3 45976 21784 45976 21784 0 tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[4\]
rlabel metal2 47656 25256 47656 25256 0 tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[5\]
rlabel metal2 46480 26936 46480 26936 0 tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[6\]
rlabel metal2 47656 28896 47656 28896 0 tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[7\]
rlabel metal2 48216 32200 48216 32200 0 tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[8\]
rlabel metal2 46872 33600 46872 33600 0 tt_um_rejunity_sn76489.noise\[0\].gen.lfsr\[9\]
rlabel metal2 40768 24024 40768 24024 0 tt_um_rejunity_sn76489.noise\[0\].gen.restart_noise
rlabel metal2 41272 33040 41272 33040 0 tt_um_rejunity_sn76489.noise\[0\].gen.signal_edge.previous_signal_state_0
rlabel metal3 33880 38024 33880 38024 0 tt_um_rejunity_sn76489.pwm.accumulator\[0\]
rlabel metal2 45304 50120 45304 50120 0 tt_um_rejunity_sn76489.pwm.accumulator\[10\]
rlabel metal3 45192 53816 45192 53816 0 tt_um_rejunity_sn76489.pwm.accumulator\[11\]
rlabel metal2 34720 36344 34720 36344 0 tt_um_rejunity_sn76489.pwm.accumulator\[1\]
rlabel metal2 33320 39872 33320 39872 0 tt_um_rejunity_sn76489.pwm.accumulator\[2\]
rlabel metal2 35784 40768 35784 40768 0 tt_um_rejunity_sn76489.pwm.accumulator\[3\]
rlabel metal2 33096 43344 33096 43344 0 tt_um_rejunity_sn76489.pwm.accumulator\[4\]
rlabel metal2 33768 45864 33768 45864 0 tt_um_rejunity_sn76489.pwm.accumulator\[5\]
rlabel metal2 35224 47152 35224 47152 0 tt_um_rejunity_sn76489.pwm.accumulator\[6\]
rlabel metal3 37128 49672 37128 49672 0 tt_um_rejunity_sn76489.pwm.accumulator\[7\]
rlabel metal2 37240 54264 37240 54264 0 tt_um_rejunity_sn76489.pwm.accumulator\[8\]
rlabel metal2 38024 55384 38024 55384 0 tt_um_rejunity_sn76489.pwm.accumulator\[9\]
rlabel metal2 45640 45136 45640 45136 0 tt_um_rejunity_sn76489.spi_dac_i_2.counter\[0\]
rlabel metal3 45864 45080 45864 45080 0 tt_um_rejunity_sn76489.spi_dac_i_2.counter\[1\]
rlabel metal2 46648 44744 46648 44744 0 tt_um_rejunity_sn76489.spi_dac_i_2.counter\[2\]
rlabel metal2 46648 47376 46648 47376 0 tt_um_rejunity_sn76489.spi_dac_i_2.counter\[3\]
rlabel metal3 46256 47432 46256 47432 0 tt_um_rejunity_sn76489.spi_dac_i_2.counter\[4\]
rlabel metal2 40376 40600 40376 40600 0 tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff\[0\]
rlabel metal2 43064 49672 43064 49672 0 tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff\[10\]
rlabel metal2 44296 48888 44296 48888 0 tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff\[11\]
rlabel metal2 38416 41832 38416 41832 0 tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff\[1\]
rlabel metal2 39256 43232 39256 43232 0 tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff\[2\]
rlabel metal2 38864 43736 38864 43736 0 tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff\[3\]
rlabel metal2 39648 45976 39648 45976 0 tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff\[4\]
rlabel metal2 39872 46648 39872 46648 0 tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff\[5\]
rlabel metal2 40824 51016 40824 51016 0 tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff\[6\]
rlabel metal2 41272 52976 41272 52976 0 tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff\[7\]
rlabel metal2 43064 53648 43064 53648 0 tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff\[8\]
rlabel metal2 41496 54880 41496 54880 0 tt_um_rejunity_sn76489.spi_dac_i_2.spi_dat_buff\[9\]
rlabel metal2 31528 8736 31528 8736 0 tt_um_rejunity_sn76489.tone\[0\].gen.counter\[0\]
rlabel metal2 31080 5544 31080 5544 0 tt_um_rejunity_sn76489.tone\[0\].gen.counter\[1\]
rlabel metal3 29680 5880 29680 5880 0 tt_um_rejunity_sn76489.tone\[0\].gen.counter\[2\]
rlabel metal2 27720 6720 27720 6720 0 tt_um_rejunity_sn76489.tone\[0\].gen.counter\[3\]
rlabel metal3 24920 8232 24920 8232 0 tt_um_rejunity_sn76489.tone\[0\].gen.counter\[4\]
rlabel via2 25256 7448 25256 7448 0 tt_um_rejunity_sn76489.tone\[0\].gen.counter\[5\]
rlabel metal2 24192 9016 24192 9016 0 tt_um_rejunity_sn76489.tone\[0\].gen.counter\[6\]
rlabel metal2 25816 11984 25816 11984 0 tt_um_rejunity_sn76489.tone\[0\].gen.counter\[7\]
rlabel metal2 25704 14056 25704 14056 0 tt_um_rejunity_sn76489.tone\[0\].gen.counter\[8\]
rlabel metal2 26488 14952 26488 14952 0 tt_um_rejunity_sn76489.tone\[0\].gen.counter\[9\]
rlabel metal2 43568 8456 43568 8456 0 tt_um_rejunity_sn76489.tone\[1\].gen.counter\[0\]
rlabel metal2 43848 8176 43848 8176 0 tt_um_rejunity_sn76489.tone\[1\].gen.counter\[1\]
rlabel metal3 44240 7448 44240 7448 0 tt_um_rejunity_sn76489.tone\[1\].gen.counter\[2\]
rlabel metal2 43792 4200 43792 4200 0 tt_um_rejunity_sn76489.tone\[1\].gen.counter\[3\]
rlabel metal2 37352 6944 37352 6944 0 tt_um_rejunity_sn76489.tone\[1\].gen.counter\[4\]
rlabel metal2 36960 5880 36960 5880 0 tt_um_rejunity_sn76489.tone\[1\].gen.counter\[5\]
rlabel metal2 36680 7616 36680 7616 0 tt_um_rejunity_sn76489.tone\[1\].gen.counter\[6\]
rlabel metal2 37352 10416 37352 10416 0 tt_um_rejunity_sn76489.tone\[1\].gen.counter\[7\]
rlabel metal2 37464 10136 37464 10136 0 tt_um_rejunity_sn76489.tone\[1\].gen.counter\[8\]
rlabel metal2 31304 15204 31304 15204 0 tt_um_rejunity_sn76489.tone\[1\].gen.counter\[9\]
rlabel metal2 46760 17920 46760 17920 0 tt_um_rejunity_sn76489.tone\[2\].gen.counter\[0\]
rlabel metal3 44240 18424 44240 18424 0 tt_um_rejunity_sn76489.tone\[2\].gen.counter\[1\]
rlabel metal3 43904 17640 43904 17640 0 tt_um_rejunity_sn76489.tone\[2\].gen.counter\[2\]
rlabel metal2 42952 16352 42952 16352 0 tt_um_rejunity_sn76489.tone\[2\].gen.counter\[3\]
rlabel metal2 42392 17080 42392 17080 0 tt_um_rejunity_sn76489.tone\[2\].gen.counter\[4\]
rlabel metal2 38696 15904 38696 15904 0 tt_um_rejunity_sn76489.tone\[2\].gen.counter\[5\]
rlabel metal2 37912 16016 37912 16016 0 tt_um_rejunity_sn76489.tone\[2\].gen.counter\[6\]
rlabel metal2 37128 20384 37128 20384 0 tt_um_rejunity_sn76489.tone\[2\].gen.counter\[7\]
rlabel metal2 39088 18312 39088 18312 0 tt_um_rejunity_sn76489.tone\[2\].gen.counter\[8\]
rlabel metal2 39144 16688 39144 16688 0 tt_um_rejunity_sn76489.tone\[2\].gen.counter\[9\]
rlabel metal3 3374 9912 3374 9912 0 wb_clk_i
<< properties >>
string FIXED_BBOX 0 0 50000 60000
<< end >>
