VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO wrapped_tholin_riscv
  CLASS BLOCK ;
  FOREIGN wrapped_tholin_riscv ;
  ORIGIN 0.000 0.000 ;
  SIZE 1100.000 BY 1150.000 ;
  PIN custom_settings[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 90.720 4.000 91.280 ;
    END
  END custom_settings[0]
  PIN custom_settings[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 120.960 4.000 121.520 ;
    END
  END custom_settings[1]
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 151.200 4.000 151.760 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 453.600 4.000 454.160 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 483.840 4.000 484.400 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 514.080 4.000 514.640 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 544.320 4.000 544.880 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 574.560 4.000 575.120 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 604.800 4.000 605.360 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 635.040 4.000 635.600 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 665.280 4.000 665.840 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 695.520 4.000 696.080 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 725.760 4.000 726.320 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 181.440 4.000 182.000 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 756.000 4.000 756.560 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 786.240 4.000 786.800 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 816.480 4.000 817.040 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 846.720 4.000 847.280 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 876.960 4.000 877.520 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 907.200 4.000 907.760 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 937.440 4.000 938.000 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 967.680 4.000 968.240 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 997.920 4.000 998.480 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1028.160 4.000 1028.720 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 211.680 4.000 212.240 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1058.400 4.000 1058.960 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1088.640 4.000 1089.200 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1118.880 4.000 1119.440 ;
    END
  END io_in[32]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 241.920 4.000 242.480 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 272.160 4.000 272.720 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 302.400 4.000 302.960 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 332.640 4.000 333.200 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 362.880 4.000 363.440 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 393.120 4.000 393.680 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 423.360 4.000 423.920 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 29.120 1146.000 29.680 1150.000 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 353.920 1146.000 354.480 1150.000 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 386.400 1146.000 386.960 1150.000 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 418.880 1146.000 419.440 1150.000 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 451.360 1146.000 451.920 1150.000 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 483.840 1146.000 484.400 1150.000 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 516.320 1146.000 516.880 1150.000 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 548.800 1146.000 549.360 1150.000 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 581.280 1146.000 581.840 1150.000 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 613.760 1146.000 614.320 1150.000 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 646.240 1146.000 646.800 1150.000 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 61.600 1146.000 62.160 1150.000 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 678.720 1146.000 679.280 1150.000 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 711.200 1146.000 711.760 1150.000 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 743.680 1146.000 744.240 1150.000 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 776.160 1146.000 776.720 1150.000 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 808.640 1146.000 809.200 1150.000 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 841.120 1146.000 841.680 1150.000 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 873.600 1146.000 874.160 1150.000 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 906.080 1146.000 906.640 1150.000 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 938.560 1146.000 939.120 1150.000 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 971.040 1146.000 971.600 1150.000 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 94.080 1146.000 94.640 1150.000 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1003.520 1146.000 1004.080 1150.000 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1036.000 1146.000 1036.560 1150.000 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1068.480 1146.000 1069.040 1150.000 ;
    END
  END io_oeb[32]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 126.560 1146.000 127.120 1150.000 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 159.040 1146.000 159.600 1150.000 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 191.520 1146.000 192.080 1150.000 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 224.000 1146.000 224.560 1150.000 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 256.480 1146.000 257.040 1150.000 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 288.960 1146.000 289.520 1150.000 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 321.440 1146.000 322.000 1150.000 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 29.120 0.000 29.680 4.000 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 353.920 0.000 354.480 4.000 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 386.400 0.000 386.960 4.000 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 418.880 0.000 419.440 4.000 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 451.360 0.000 451.920 4.000 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 483.840 0.000 484.400 4.000 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 516.320 0.000 516.880 4.000 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 548.800 0.000 549.360 4.000 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 581.280 0.000 581.840 4.000 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 613.760 0.000 614.320 4.000 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 646.240 0.000 646.800 4.000 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 61.600 0.000 62.160 4.000 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 678.720 0.000 679.280 4.000 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 711.200 0.000 711.760 4.000 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 743.680 0.000 744.240 4.000 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 776.160 0.000 776.720 4.000 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 808.640 0.000 809.200 4.000 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 841.120 0.000 841.680 4.000 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 873.600 0.000 874.160 4.000 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 906.080 0.000 906.640 4.000 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 938.560 0.000 939.120 4.000 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 971.040 0.000 971.600 4.000 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 94.080 0.000 94.640 4.000 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1003.520 0.000 1004.080 4.000 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1036.000 0.000 1036.560 4.000 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1068.480 0.000 1069.040 4.000 ;
    END
  END io_out[32]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 126.560 0.000 127.120 4.000 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 159.040 0.000 159.600 4.000 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 191.520 0.000 192.080 4.000 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 224.000 0.000 224.560 4.000 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 256.480 0.000 257.040 4.000 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 288.960 0.000 289.520 4.000 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 321.440 0.000 322.000 4.000 ;
    END
  END io_out[9]
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 60.480 4.000 61.040 ;
    END
  END rst_n
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 22.240 15.380 23.840 1133.180 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 175.840 15.380 177.440 1133.180 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 329.440 15.380 331.040 1133.180 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 483.040 15.380 484.640 1133.180 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 636.640 15.380 638.240 1133.180 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 790.240 15.380 791.840 1133.180 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 943.840 15.380 945.440 1133.180 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 99.040 15.380 100.640 1133.180 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 252.640 15.380 254.240 1133.180 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 406.240 15.380 407.840 1133.180 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 559.840 15.380 561.440 1133.180 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 713.440 15.380 715.040 1133.180 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 867.040 15.380 868.640 1133.180 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1020.640 15.380 1022.240 1133.180 ;
    END
  END vss
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.738000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 30.240 4.000 30.800 ;
    END
  END wb_clk_i
  OBS
      LAYER Metal1 ;
        RECT 6.720 15.380 1093.120 1133.850 ;
      LAYER Metal2 ;
        RECT 4.620 1145.700 28.820 1146.740 ;
        RECT 29.980 1145.700 61.300 1146.740 ;
        RECT 62.460 1145.700 93.780 1146.740 ;
        RECT 94.940 1145.700 126.260 1146.740 ;
        RECT 127.420 1145.700 158.740 1146.740 ;
        RECT 159.900 1145.700 191.220 1146.740 ;
        RECT 192.380 1145.700 223.700 1146.740 ;
        RECT 224.860 1145.700 256.180 1146.740 ;
        RECT 257.340 1145.700 288.660 1146.740 ;
        RECT 289.820 1145.700 321.140 1146.740 ;
        RECT 322.300 1145.700 353.620 1146.740 ;
        RECT 354.780 1145.700 386.100 1146.740 ;
        RECT 387.260 1145.700 418.580 1146.740 ;
        RECT 419.740 1145.700 451.060 1146.740 ;
        RECT 452.220 1145.700 483.540 1146.740 ;
        RECT 484.700 1145.700 516.020 1146.740 ;
        RECT 517.180 1145.700 548.500 1146.740 ;
        RECT 549.660 1145.700 580.980 1146.740 ;
        RECT 582.140 1145.700 613.460 1146.740 ;
        RECT 614.620 1145.700 645.940 1146.740 ;
        RECT 647.100 1145.700 678.420 1146.740 ;
        RECT 679.580 1145.700 710.900 1146.740 ;
        RECT 712.060 1145.700 743.380 1146.740 ;
        RECT 744.540 1145.700 775.860 1146.740 ;
        RECT 777.020 1145.700 808.340 1146.740 ;
        RECT 809.500 1145.700 840.820 1146.740 ;
        RECT 841.980 1145.700 873.300 1146.740 ;
        RECT 874.460 1145.700 905.780 1146.740 ;
        RECT 906.940 1145.700 938.260 1146.740 ;
        RECT 939.420 1145.700 970.740 1146.740 ;
        RECT 971.900 1145.700 1003.220 1146.740 ;
        RECT 1004.380 1145.700 1035.700 1146.740 ;
        RECT 1036.860 1145.700 1068.180 1146.740 ;
        RECT 1069.340 1145.700 1092.420 1146.740 ;
        RECT 4.620 4.300 1092.420 1145.700 ;
        RECT 4.620 2.890 28.820 4.300 ;
        RECT 29.980 2.890 61.300 4.300 ;
        RECT 62.460 2.890 93.780 4.300 ;
        RECT 94.940 2.890 126.260 4.300 ;
        RECT 127.420 2.890 158.740 4.300 ;
        RECT 159.900 2.890 191.220 4.300 ;
        RECT 192.380 2.890 223.700 4.300 ;
        RECT 224.860 2.890 256.180 4.300 ;
        RECT 257.340 2.890 288.660 4.300 ;
        RECT 289.820 2.890 321.140 4.300 ;
        RECT 322.300 2.890 353.620 4.300 ;
        RECT 354.780 2.890 386.100 4.300 ;
        RECT 387.260 2.890 418.580 4.300 ;
        RECT 419.740 2.890 451.060 4.300 ;
        RECT 452.220 2.890 483.540 4.300 ;
        RECT 484.700 2.890 516.020 4.300 ;
        RECT 517.180 2.890 548.500 4.300 ;
        RECT 549.660 2.890 580.980 4.300 ;
        RECT 582.140 2.890 613.460 4.300 ;
        RECT 614.620 2.890 645.940 4.300 ;
        RECT 647.100 2.890 678.420 4.300 ;
        RECT 679.580 2.890 710.900 4.300 ;
        RECT 712.060 2.890 743.380 4.300 ;
        RECT 744.540 2.890 775.860 4.300 ;
        RECT 777.020 2.890 808.340 4.300 ;
        RECT 809.500 2.890 840.820 4.300 ;
        RECT 841.980 2.890 873.300 4.300 ;
        RECT 874.460 2.890 905.780 4.300 ;
        RECT 906.940 2.890 938.260 4.300 ;
        RECT 939.420 2.890 970.740 4.300 ;
        RECT 971.900 2.890 1003.220 4.300 ;
        RECT 1004.380 2.890 1035.700 4.300 ;
        RECT 1036.860 2.890 1068.180 4.300 ;
        RECT 1069.340 2.890 1092.420 4.300 ;
      LAYER Metal3 ;
        RECT 4.000 1119.740 1091.910 1135.540 ;
        RECT 4.300 1118.580 1091.910 1119.740 ;
        RECT 4.000 1089.500 1091.910 1118.580 ;
        RECT 4.300 1088.340 1091.910 1089.500 ;
        RECT 4.000 1059.260 1091.910 1088.340 ;
        RECT 4.300 1058.100 1091.910 1059.260 ;
        RECT 4.000 1029.020 1091.910 1058.100 ;
        RECT 4.300 1027.860 1091.910 1029.020 ;
        RECT 4.000 998.780 1091.910 1027.860 ;
        RECT 4.300 997.620 1091.910 998.780 ;
        RECT 4.000 968.540 1091.910 997.620 ;
        RECT 4.300 967.380 1091.910 968.540 ;
        RECT 4.000 938.300 1091.910 967.380 ;
        RECT 4.300 937.140 1091.910 938.300 ;
        RECT 4.000 908.060 1091.910 937.140 ;
        RECT 4.300 906.900 1091.910 908.060 ;
        RECT 4.000 877.820 1091.910 906.900 ;
        RECT 4.300 876.660 1091.910 877.820 ;
        RECT 4.000 847.580 1091.910 876.660 ;
        RECT 4.300 846.420 1091.910 847.580 ;
        RECT 4.000 817.340 1091.910 846.420 ;
        RECT 4.300 816.180 1091.910 817.340 ;
        RECT 4.000 787.100 1091.910 816.180 ;
        RECT 4.300 785.940 1091.910 787.100 ;
        RECT 4.000 756.860 1091.910 785.940 ;
        RECT 4.300 755.700 1091.910 756.860 ;
        RECT 4.000 726.620 1091.910 755.700 ;
        RECT 4.300 725.460 1091.910 726.620 ;
        RECT 4.000 696.380 1091.910 725.460 ;
        RECT 4.300 695.220 1091.910 696.380 ;
        RECT 4.000 666.140 1091.910 695.220 ;
        RECT 4.300 664.980 1091.910 666.140 ;
        RECT 4.000 635.900 1091.910 664.980 ;
        RECT 4.300 634.740 1091.910 635.900 ;
        RECT 4.000 605.660 1091.910 634.740 ;
        RECT 4.300 604.500 1091.910 605.660 ;
        RECT 4.000 575.420 1091.910 604.500 ;
        RECT 4.300 574.260 1091.910 575.420 ;
        RECT 4.000 545.180 1091.910 574.260 ;
        RECT 4.300 544.020 1091.910 545.180 ;
        RECT 4.000 514.940 1091.910 544.020 ;
        RECT 4.300 513.780 1091.910 514.940 ;
        RECT 4.000 484.700 1091.910 513.780 ;
        RECT 4.300 483.540 1091.910 484.700 ;
        RECT 4.000 454.460 1091.910 483.540 ;
        RECT 4.300 453.300 1091.910 454.460 ;
        RECT 4.000 424.220 1091.910 453.300 ;
        RECT 4.300 423.060 1091.910 424.220 ;
        RECT 4.000 393.980 1091.910 423.060 ;
        RECT 4.300 392.820 1091.910 393.980 ;
        RECT 4.000 363.740 1091.910 392.820 ;
        RECT 4.300 362.580 1091.910 363.740 ;
        RECT 4.000 333.500 1091.910 362.580 ;
        RECT 4.300 332.340 1091.910 333.500 ;
        RECT 4.000 303.260 1091.910 332.340 ;
        RECT 4.300 302.100 1091.910 303.260 ;
        RECT 4.000 273.020 1091.910 302.100 ;
        RECT 4.300 271.860 1091.910 273.020 ;
        RECT 4.000 242.780 1091.910 271.860 ;
        RECT 4.300 241.620 1091.910 242.780 ;
        RECT 4.000 212.540 1091.910 241.620 ;
        RECT 4.300 211.380 1091.910 212.540 ;
        RECT 4.000 182.300 1091.910 211.380 ;
        RECT 4.300 181.140 1091.910 182.300 ;
        RECT 4.000 152.060 1091.910 181.140 ;
        RECT 4.300 150.900 1091.910 152.060 ;
        RECT 4.000 121.820 1091.910 150.900 ;
        RECT 4.300 120.660 1091.910 121.820 ;
        RECT 4.000 91.580 1091.910 120.660 ;
        RECT 4.300 90.420 1091.910 91.580 ;
        RECT 4.000 61.340 1091.910 90.420 ;
        RECT 4.300 60.180 1091.910 61.340 ;
        RECT 4.000 31.100 1091.910 60.180 ;
        RECT 4.300 29.940 1091.910 31.100 ;
        RECT 4.000 2.940 1091.910 29.940 ;
      LAYER Metal4 ;
        RECT 11.340 1133.480 1077.860 1135.590 ;
        RECT 11.340 15.080 21.940 1133.480 ;
        RECT 24.140 15.080 98.740 1133.480 ;
        RECT 100.940 15.080 175.540 1133.480 ;
        RECT 177.740 15.080 252.340 1133.480 ;
        RECT 254.540 15.080 329.140 1133.480 ;
        RECT 331.340 15.080 405.940 1133.480 ;
        RECT 408.140 15.080 482.740 1133.480 ;
        RECT 484.940 15.080 559.540 1133.480 ;
        RECT 561.740 15.080 636.340 1133.480 ;
        RECT 638.540 15.080 713.140 1133.480 ;
        RECT 715.340 15.080 789.940 1133.480 ;
        RECT 792.140 15.080 866.740 1133.480 ;
        RECT 868.940 15.080 943.540 1133.480 ;
        RECT 945.740 15.080 1020.340 1133.480 ;
        RECT 1022.540 15.080 1077.860 1133.480 ;
        RECT 11.340 2.890 1077.860 15.080 ;
  END
END wrapped_tholin_riscv
END LIBRARY

