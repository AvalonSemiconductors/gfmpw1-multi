magic
tech gf180mcuD
magscale 1 10
timestamp 1702247295
<< nwell >>
rect 1258 45849 48694 46342
rect 1258 45824 21581 45849
rect 1258 45095 12440 45120
rect 1258 44281 48694 45095
rect 1258 44256 9528 44281
rect 1258 43527 6685 43552
rect 1258 42713 48694 43527
rect 1258 42688 14301 42713
rect 1258 41959 6909 41984
rect 1258 41145 48694 41959
rect 1258 41120 23640 41145
rect 1258 40391 3592 40416
rect 1258 39577 48694 40391
rect 1258 39552 7581 39577
rect 1258 38823 3592 38848
rect 1258 38009 48694 38823
rect 1258 37984 15197 38009
rect 1258 37255 5789 37280
rect 1258 36441 48694 37255
rect 1258 36416 3592 36441
rect 1258 35687 12776 35712
rect 1258 34873 48694 35687
rect 1258 34848 9493 34873
rect 1258 34119 2541 34144
rect 1258 33305 48694 34119
rect 1258 33280 15464 33305
rect 1258 32551 11165 32576
rect 1258 31737 48694 32551
rect 1258 31712 2541 31737
rect 1258 30983 4445 31008
rect 1258 30169 48694 30983
rect 1258 30144 2541 30169
rect 1258 29415 2541 29440
rect 1258 28601 48694 29415
rect 1258 28576 24045 28601
rect 1258 27847 11725 27872
rect 1258 27033 48694 27847
rect 1258 27008 2541 27033
rect 1258 26279 3592 26304
rect 1258 25465 48694 26279
rect 1258 25440 14301 25465
rect 1258 24711 2541 24736
rect 1258 23897 48694 24711
rect 1258 23872 11880 23897
rect 1258 23143 29352 23168
rect 1258 22329 48694 23143
rect 1258 22304 2541 22329
rect 1258 21575 11501 21600
rect 1258 20761 48694 21575
rect 1258 20736 2541 20761
rect 1258 20007 37261 20032
rect 1258 19193 48694 20007
rect 1258 19168 2541 19193
rect 1258 18439 6125 18464
rect 1258 17625 48694 18439
rect 1258 17600 2541 17625
rect 1258 16871 6909 16896
rect 1258 16057 48694 16871
rect 1258 16032 26061 16057
rect 1258 15303 2541 15328
rect 1258 14489 48694 15303
rect 1258 14464 16653 14489
rect 1258 13735 2541 13760
rect 1258 12921 48694 13735
rect 1258 12896 9149 12921
rect 1258 12167 2541 12192
rect 1258 11353 48694 12167
rect 1258 11328 8141 11353
rect 1258 10599 3592 10624
rect 1258 9785 48694 10599
rect 1258 9760 6461 9785
rect 1258 9031 12397 9056
rect 1258 8217 48694 9031
rect 1258 8192 2541 8217
rect 1258 7463 6237 7488
rect 1258 6649 48694 7463
rect 1258 6624 2541 6649
rect 1258 5895 22477 5920
rect 1258 5081 48694 5895
rect 1258 5056 7581 5081
rect 1258 4327 5005 4352
rect 1258 3513 48694 4327
rect 1258 3488 33005 3513
<< pwell >>
rect 1258 45120 48694 45824
rect 1258 43552 48694 44256
rect 1258 41984 48694 42688
rect 1258 40416 48694 41120
rect 1258 38848 48694 39552
rect 1258 37280 48694 37984
rect 1258 35712 48694 36416
rect 1258 34144 48694 34848
rect 1258 32576 48694 33280
rect 1258 31008 48694 31712
rect 1258 29440 48694 30144
rect 1258 27872 48694 28576
rect 1258 26304 48694 27008
rect 1258 24736 48694 25440
rect 1258 23168 48694 23872
rect 1258 21600 48694 22304
rect 1258 20032 48694 20736
rect 1258 18464 48694 19168
rect 1258 16896 48694 17600
rect 1258 15328 48694 16032
rect 1258 13760 48694 14464
rect 1258 12192 48694 12896
rect 1258 10624 48694 11328
rect 1258 9056 48694 9760
rect 1258 7488 48694 8192
rect 1258 5920 48694 6624
rect 1258 4352 48694 5056
rect 1258 3050 48694 3488
<< obsm1 >>
rect 1344 1710 48608 46450
<< metal2 >>
rect 6272 49200 6384 50000
rect 18592 49200 18704 50000
rect 30912 49200 31024 50000
rect 43232 49200 43344 50000
rect 3584 0 3696 800
rect 5152 0 5264 800
rect 6720 0 6832 800
rect 8288 0 8400 800
rect 9856 0 9968 800
rect 11424 0 11536 800
rect 12992 0 13104 800
rect 14560 0 14672 800
rect 16128 0 16240 800
rect 17696 0 17808 800
rect 19264 0 19376 800
rect 20832 0 20944 800
rect 22400 0 22512 800
rect 23968 0 24080 800
rect 25536 0 25648 800
rect 27104 0 27216 800
rect 28672 0 28784 800
rect 30240 0 30352 800
rect 31808 0 31920 800
rect 33376 0 33488 800
rect 34944 0 35056 800
rect 36512 0 36624 800
rect 38080 0 38192 800
rect 39648 0 39760 800
rect 41216 0 41328 800
rect 42784 0 42896 800
rect 44352 0 44464 800
rect 45920 0 46032 800
<< obsm2 >>
rect 1708 49140 6212 49200
rect 6444 49140 18532 49200
rect 18764 49140 30852 49200
rect 31084 49140 43172 49200
rect 43404 49140 48580 49200
rect 1708 860 48580 49140
rect 1708 700 3524 860
rect 3756 700 5092 860
rect 5324 700 6660 860
rect 6892 700 8228 860
rect 8460 700 9796 860
rect 10028 700 11364 860
rect 11596 700 12932 860
rect 13164 700 14500 860
rect 14732 700 16068 860
rect 16300 700 17636 860
rect 17868 700 19204 860
rect 19436 700 20772 860
rect 21004 700 22340 860
rect 22572 700 23908 860
rect 24140 700 25476 860
rect 25708 700 27044 860
rect 27276 700 28612 860
rect 28844 700 30180 860
rect 30412 700 31748 860
rect 31980 700 33316 860
rect 33548 700 34884 860
rect 35116 700 36452 860
rect 36684 700 38020 860
rect 38252 700 39588 860
rect 39820 700 41156 860
rect 41388 700 42724 860
rect 42956 700 44292 860
rect 44524 700 45860 860
rect 46092 700 48580 860
<< metal3 >>
rect 49200 47040 50000 47152
rect 49200 42112 50000 42224
rect 49200 37184 50000 37296
rect 49200 32256 50000 32368
rect 49200 27328 50000 27440
rect 49200 22400 50000 22512
rect 49200 17472 50000 17584
rect 49200 12544 50000 12656
rect 49200 7616 50000 7728
rect 49200 2688 50000 2800
<< obsm3 >>
rect 1698 46980 49140 47124
rect 1698 42284 49200 46980
rect 1698 42052 49140 42284
rect 1698 37356 49200 42052
rect 1698 37124 49140 37356
rect 1698 32428 49200 37124
rect 1698 32196 49140 32428
rect 1698 27500 49200 32196
rect 1698 27268 49140 27500
rect 1698 22572 49200 27268
rect 1698 22340 49140 22572
rect 1698 17644 49200 22340
rect 1698 17412 49140 17644
rect 1698 12716 49200 17412
rect 1698 12484 49140 12716
rect 1698 7788 49200 12484
rect 1698 7556 49140 7788
rect 1698 2860 49200 7556
rect 1698 2628 49140 2860
rect 1698 1708 49200 2628
<< metal4 >>
rect 4448 3076 4768 46316
rect 19808 3076 20128 46316
rect 35168 3076 35488 46316
<< obsm4 >>
rect 16044 4498 19748 44110
rect 20188 4498 35108 44110
rect 35548 4498 47124 44110
<< labels >>
rlabel metal3 s 49200 42112 50000 42224 6 custom_settings[0]
port 1 nsew signal input
rlabel metal3 s 49200 47040 50000 47152 6 custom_settings[1]
port 2 nsew signal input
rlabel metal3 s 49200 2688 50000 2800 6 io_in_1[0]
port 3 nsew signal input
rlabel metal3 s 49200 7616 50000 7728 6 io_in_1[1]
port 4 nsew signal input
rlabel metal3 s 49200 12544 50000 12656 6 io_in_1[2]
port 5 nsew signal input
rlabel metal3 s 49200 17472 50000 17584 6 io_in_1[3]
port 6 nsew signal input
rlabel metal3 s 49200 22400 50000 22512 6 io_in_1[4]
port 7 nsew signal input
rlabel metal3 s 49200 27328 50000 27440 6 io_in_1[5]
port 8 nsew signal input
rlabel metal3 s 49200 32256 50000 32368 6 io_in_1[6]
port 9 nsew signal input
rlabel metal3 s 49200 37184 50000 37296 6 io_in_1[7]
port 10 nsew signal input
rlabel metal2 s 30912 49200 31024 50000 6 io_in_2[0]
port 11 nsew signal input
rlabel metal2 s 43232 49200 43344 50000 6 io_in_2[1]
port 12 nsew signal input
rlabel metal2 s 3584 0 3696 800 6 io_out[0]
port 13 nsew signal output
rlabel metal2 s 19264 0 19376 800 6 io_out[10]
port 14 nsew signal output
rlabel metal2 s 20832 0 20944 800 6 io_out[11]
port 15 nsew signal output
rlabel metal2 s 22400 0 22512 800 6 io_out[12]
port 16 nsew signal output
rlabel metal2 s 23968 0 24080 800 6 io_out[13]
port 17 nsew signal output
rlabel metal2 s 25536 0 25648 800 6 io_out[14]
port 18 nsew signal output
rlabel metal2 s 27104 0 27216 800 6 io_out[15]
port 19 nsew signal output
rlabel metal2 s 28672 0 28784 800 6 io_out[16]
port 20 nsew signal output
rlabel metal2 s 30240 0 30352 800 6 io_out[17]
port 21 nsew signal output
rlabel metal2 s 31808 0 31920 800 6 io_out[18]
port 22 nsew signal output
rlabel metal2 s 33376 0 33488 800 6 io_out[19]
port 23 nsew signal output
rlabel metal2 s 5152 0 5264 800 6 io_out[1]
port 24 nsew signal output
rlabel metal2 s 34944 0 35056 800 6 io_out[20]
port 25 nsew signal output
rlabel metal2 s 36512 0 36624 800 6 io_out[21]
port 26 nsew signal output
rlabel metal2 s 38080 0 38192 800 6 io_out[22]
port 27 nsew signal output
rlabel metal2 s 39648 0 39760 800 6 io_out[23]
port 28 nsew signal output
rlabel metal2 s 41216 0 41328 800 6 io_out[24]
port 29 nsew signal output
rlabel metal2 s 42784 0 42896 800 6 io_out[25]
port 30 nsew signal output
rlabel metal2 s 44352 0 44464 800 6 io_out[26]
port 31 nsew signal output
rlabel metal2 s 45920 0 46032 800 6 io_out[27]
port 32 nsew signal output
rlabel metal2 s 6720 0 6832 800 6 io_out[2]
port 33 nsew signal output
rlabel metal2 s 8288 0 8400 800 6 io_out[3]
port 34 nsew signal output
rlabel metal2 s 9856 0 9968 800 6 io_out[4]
port 35 nsew signal output
rlabel metal2 s 11424 0 11536 800 6 io_out[5]
port 36 nsew signal output
rlabel metal2 s 12992 0 13104 800 6 io_out[6]
port 37 nsew signal output
rlabel metal2 s 14560 0 14672 800 6 io_out[7]
port 38 nsew signal output
rlabel metal2 s 16128 0 16240 800 6 io_out[8]
port 39 nsew signal output
rlabel metal2 s 17696 0 17808 800 6 io_out[9]
port 40 nsew signal output
rlabel metal2 s 18592 49200 18704 50000 6 rst_n
port 41 nsew signal input
rlabel metal4 s 4448 3076 4768 46316 6 vdd
port 42 nsew power bidirectional
rlabel metal4 s 35168 3076 35488 46316 6 vdd
port 42 nsew power bidirectional
rlabel metal4 s 19808 3076 20128 46316 6 vss
port 43 nsew ground bidirectional
rlabel metal2 s 6272 49200 6384 50000 6 wb_clk_i
port 44 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 50000 50000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 2177630
string GDS_FILE /run/media/tholin/fbc90f8f-67e9-406d-9872-54f02ad6a2d8/gfmpw1-multi/openlane/wrapped_ay8913/runs/23_12_10_23_25/results/signoff/wrapped_ay8913.magic.gds
string GDS_START 286528
<< end >>

