* NGSPICE file created from wrapped_mc14500.ext - technology: gf180mcuD

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__antenna abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__antenna I VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__filltie abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__filltie VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_1 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_1 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_2 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_1 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and3_1 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_2 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_1 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_1 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_1 D CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_1 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_8 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__endcap abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__endcap VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_2 D CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_1 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_1 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_1 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_1 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_1 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__tiel abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__tiel ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_1 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_1 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_2 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_1 A1 A2 A3 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_1 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_2 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_1 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_1 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_1 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_2 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_2 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_4 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or4_1 A1 A2 A3 A4 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffnq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffnq_1 D CLKN Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_2 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and4_1 A1 A2 A3 A4 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux2_2 I0 I1 S Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_2 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or3_1 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_1 A1 A2 A3 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_32 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_4 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_2 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_2 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_1 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor2_1 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_2 A1 A2 A3 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_1 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

.subckt wrapped_mc14500 SDI clk_i custom_setting io_in[0] io_in[1] io_in[2] io_in[3]
+ io_in[4] io_in[5] io_in[6] io_in[7] io_out[10] io_out[11] io_out[12] io_out[13]
+ io_out[14] io_out[15] io_out[16] io_out[17] io_out[18] io_out[19] io_out[20] io_out[21]
+ io_out[22] io_out[23] io_out[24] io_out[25] io_out[26] io_out[27] io_out[28] io_out[29]
+ io_out[2] io_out[30] io_out[7] io_out[8] io_out[9] rst_n sram_addr[0] sram_addr[1]
+ sram_addr[2] sram_addr[3] sram_addr[4] sram_addr[5] sram_gwe sram_in[0] sram_in[1]
+ sram_in[2] sram_in[3] sram_in[4] sram_in[5] sram_in[6] sram_in[7] sram_out[0] sram_out[1]
+ sram_out[2] sram_out[3] sram_out[4] sram_out[5] sram_out[6] sram_out[7] vdd vss
+ io_out[1] io_out[0] io_out[6] io_out[5] io_out[4] io_out[3]
XANTENNA__0738__I _0280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_9_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_15_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output37_I net37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0985_ _0480_ _0481_ _0324_ _0482_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_20_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0770_ _0286_ _0308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_11_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_34_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0968_ _0154_ _0465_ _0467_ _0468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA_clkbuf_3_3__f_clk_i_I clknet_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0899_ _0116_ _0408_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__0661__I _0217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0822_ _0120_ _0164_ _0216_ _0351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_0753_ _0248_ _0293_ _0294_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_0684_ _0234_ _0235_ _0231_ _0019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_10_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1098_ _0070_ clknet_3_3__leaf_clk_i net26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_19_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1021_ net46 _0500_ _0509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_0805_ _0116_ _0337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_0736_ dia\[6\] _0263_ _0278_ _0279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_0667_ net52 _0218_ _0223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_0598_ _0158_ _0111_ scratch\[2\] _0159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_1_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0521_ _0088_ _0091_ _0093_ _0094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_1004_ _0203_ _0495_ _0496_ _0078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_12_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0719_ _0264_ _0249_ _0265_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xoutput31 net31 io_out[21] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput53 net53 sram_in[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput20 net20 io_out[10] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput42 net42 io_out[9] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XTAP_TAPCELL_ROW_18_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_26_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0664__I _0131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0839__I _0351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0984_ _0327_ _0462_ _0481_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_1_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1079__CLK clknet_3_2__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_11_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_34_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0967_ _0429_ _0460_ _0466_ _0467_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_12_Right_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_0898_ _0404_ _0407_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_21_Right_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_30_Right_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_29_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0752_ _0284_ _0293_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_9_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0821_ dest\[15\] _0349_ _0350_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_0683_ net55 _0228_ _0235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_34_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1097_ _0069_ clknet_3_3__leaf_clk_i net25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_18_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1020_ _0499_ _0507_ _0508_ _0082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__1008__I _0202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_28_Left_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_0735_ _0277_ _0243_ _0278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_12_Left_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_16_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_0804_ net34 _0326_ _0335_ _0336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_0666_ _0219_ _0220_ _0222_ _0014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_0597_ net8 _0158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__0834__I0 _0185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0520_ mc14500.skip _0092_ _0093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1003_ mar\[0\] _0206_ _0318_ _0496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_8_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0816__I0 _0185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_6_Right_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_0718_ net16 _0264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_0649_ net44 _0204_ _0208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input11_I rst_n vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput43 net43 sram_addr[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput54 net54 sram_in[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_9_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xoutput21 net21 io_out[11] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput32 net32 io_out[22] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XTAP_TAPCELL_ROW_18_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_26_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input3_I io_in[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_15_Left_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_31_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0983_ net30 _0480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__0590__I _0131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_3_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_0_Left_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_13_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_11_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_34_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0617__A1 net10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0966_ net27 _0466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_6_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0897_ net41 _0406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0751_ _0287_ _0290_ _0292_ _0029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_9_29 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0820_ _0348_ _0349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0682_ net56 _0217_ _0234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_10_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1096_ _0068_ clknet_3_3__leaf_clk_i net24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__0838__A1 _0210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0949_ _0338_ _0449_ _0451_ net24 _0452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__0829__A1 _0210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0734_ net19 _0277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_0665_ _0221_ _0222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_24_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0803_ _0331_ _0335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_0596_ _0151_ _0155_ _0157_ _0001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1079_ _0051_ clknet_3_2__leaf_clk_i dest\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_21_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1002_ mc14500.DATA_OUT _0204_ _0495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_16_20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0717_ _0242_ _0263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0648_ _0203_ _0205_ _0207_ _0011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_12_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0579_ _0142_ _0143_ _0144_ _0003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_35_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput55 net55 sram_in[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput44 net44 sram_addr[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput33 net33 io_out[23] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput22 net22 io_out[12] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_26_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_26_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0588__I net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0653__A2 _0171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_3_3__f_clk_i clknet_0_clk_i clknet_3_3__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_13_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0982_ _0475_ _0479_ _0073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_3_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0580__A1 _0125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_20_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output35_I net35 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0626__A2 _0185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_11_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_34_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0896_ _0404_ _0405_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0965_ _0462_ _0405_ _0463_ _0464_ _0465_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__0553__A1 _0109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0750_ dib\[0\] _0291_ _0281_ _0292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_0681_ _0232_ _0233_ _0231_ _0018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1095_ _0067_ clknet_3_2__leaf_clk_i net23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0948_ _0425_ _0450_ _0451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_0879_ _0390_ _0391_ _0392_ _0057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__0829__A2 _0355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_3_2__f_clk_i_I clknet_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0802_ _0332_ _0333_ _0334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_0733_ _0262_ _0275_ _0276_ _0027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_0664_ _0131_ _0221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_0595_ mc14500.OEN_l _0156_ _0157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1078_ _0050_ clknet_3_2__leaf_clk_i dest\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_15_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xwrapped_mc14500_70 io_out[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_16_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1001_ _0420_ _0493_ _0494_ _0230_ _0077_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_TAPCELL_ROW_29_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0647_ net44 _0206_ _0138_ _0207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_12_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0716_ _0240_ _0262_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0578_ mc14500.DATA_OUT _0143_ _0144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_25_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__0968__A1 _0154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput34 net34 io_out[24] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput23 net23 io_out[13] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput45 net45 sram_addr[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput56 net56 sram_in[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__0869__I _0351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_14_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0981_ net29 _0476_ _0478_ _0338_ _0479_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__0599__I _0110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_20_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0964_ _0337_ _0464_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0895_ _0403_ _0404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1092__CLK clknet_3_2__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0680_ net54 _0228_ _0233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_10_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1094_ _0066_ clknet_3_2__leaf_clk_i net22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0947_ _0333_ _0447_ _0450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_0878_ _0343_ _0392_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_18_140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0801_ _0323_ _0333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0663_ net50 _0213_ _0220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_0732_ dia\[6\] _0267_ _0260_ _0276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_0594_ _0151_ _0155_ _0156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_1077_ _0049_ clknet_3_2__leaf_clk_i dest\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xwrapped_mc14500_71 io_out[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_21_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1000_ _0464_ _0489_ net33 _0494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_8_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_29_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0715_ _0241_ _0259_ _0261_ _0024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__1000__B net33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0646_ _0202_ _0206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_12_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0577_ _0126_ _0108_ _0121_ _0143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
Xoutput24 net24 io_out[14] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput35 net35 io_out[25] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput46 net46 sram_addr[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput57 net57 sram_in[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XPHY_EDGE_ROW_19_Right_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_28_Right_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_27_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0629_ _0188_ _0189_ _0190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_13_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_14_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0980_ net29 _0407_ _0469_ _0477_ _0478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA_input1_I SDI vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_19_Left_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_9_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_20_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0562__A3 _0131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0894_ _0088_ _0101_ _0403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_0963_ dest\[9\] _0440_ _0463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_5_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_0_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1093_ _0065_ clknet_3_2__leaf_clk_i net21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1003__B _0318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0877_ dest\[10\] _0383_ _0391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_0946_ _0446_ _0448_ _0449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_0731_ dia\[5\] _0263_ _0274_ _0275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_21_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1082__CLK clknet_3_2__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0800_ _0326_ _0331_ net34 _0332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_0662_ net51 _0218_ _0219_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_0593_ _0088_ _0155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__0837__B _0318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1076_ _0048_ clknet_3_0__leaf_clk_i dest\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_15_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0929_ _0434_ _0065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XPHY_EDGE_ROW_7_Left_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xwrapped_mc14500_72 io_out[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_16_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_29_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0645_ net45 _0204_ _0205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_0714_ dia\[3\] _0246_ _0260_ _0261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_12_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0576_ _0138_ scratch\[0\] _0142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1059_ net6 net64 mc14500.instr_l\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_7_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_33_Left_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xoutput47 net47 sram_addr[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_11_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput36 net36 io_out[26] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput25 net25 io_out[15] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_27_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0628_ _0114_ _0189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_0559_ _0126_ _0128_ _0129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_30_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_8_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0574__A1 mc14500.DATA_OUT vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_14_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1006__B _0318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_20_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1039__CLK clknet_3_4__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_20_Left_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_0962_ _0330_ _0462_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_6_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0893_ _0400_ _0401_ _0402_ _0061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_4_77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output33_I net33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout60 net23 net60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_0_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_11 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1092_ _0064_ clknet_3_2__leaf_clk_i net20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0876_ dest\[11\] _0385_ _0390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_0945_ _0333_ _0441_ _0447_ _0448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_33_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0730_ _0273_ _0243_ _0274_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_0661_ _0217_ _0218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_24_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0592_ _0150_ _0152_ _0154_ _0115_ _0002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_1075_ _0047_ clknet_3_0__leaf_clk_i dest\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0859_ dest\[5\] _0372_ _0378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_0928_ net21 _0430_ _0433_ _0154_ _0434_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
Xwrapped_mc14500_73 io_out[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_21_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_3_6__f_clk_i clknet_0_clk_i clknet_3_6__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_29_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0644_ _0198_ _0204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0713_ _0153_ _0260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_12_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_20_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0575_ _0139_ _0140_ _0141_ _0004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1058_ net5 net63 mc14500.instr_l\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xoutput26 net26 io_out[16] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA_clkbuf_3_1__f_clk_i_I clknet_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput48 net48 sram_addr[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XPHY_EDGE_ROW_1_Right_1 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xoutput37 net37 io_out[27] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_4_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0627_ _0091_ _0188_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_0558_ _0127_ _0128_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__1095__CLK clknet_3_2__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_23_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_8_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_14_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0961_ _0457_ _0341_ _0458_ _0461_ _0230_ _0070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_0892_ _0230_ _0402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_10_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout61 net20 net61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_0_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1091_ _0063_ clknet_3_2__leaf_clk_i net42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0944_ net24 _0441_ _0447_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_2_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0875_ _0388_ _0389_ _0381_ _0056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_0660_ _0119_ _0216_ _0211_ _0217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_21_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0591_ _0153_ _0154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_1_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1074_ _0046_ clknet_3_1__leaf_clk_i dest\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_15_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0927_ _0431_ _0421_ _0432_ _0425_ _0433_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_0858_ dest\[6\] _0374_ _0377_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_0789_ rst_latency\[1\] rst_latency\[0\] _0322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xwrapped_mc14500_74 io_out[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_21_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0643_ _0202_ _0203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0712_ dia\[2\] _0244_ _0258_ _0259_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_20_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0574_ mc14500.DATA_OUT _0140_ _0141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1057_ net4 net63 mc14500.instr_l\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_22_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput27 net27 io_out[17] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_11_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput38 net38 io_out[28] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput49 net49 sram_gwe vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XTAP_TAPCELL_ROW_17_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_15_Right_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_0626_ mc14500.IEN_l _0185_ _0186_ _0187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_0557_ net9 _0127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1109_ _0081_ clknet_3_0__leaf_clk_i net47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_16_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_24_Right_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_23_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_33_Right_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_16_285 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1062__CLK clknet_3_4__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0609_ net38 _0170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_5_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1085__CLK clknet_3_3__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0960_ net59 _0459_ _0460_ _0429_ _0461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_0891_ dest\[14\] _0394_ _0401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_30_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout62 net66 net62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_0_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1090_ _0062_ clknet_3_2__leaf_clk_i net41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_0874_ dest\[9\] _0383_ _0389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_0943_ dest\[6\] _0440_ _0446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_2_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1100__CLK clknet_3_3__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0590_ _0131_ _0153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1073_ _0045_ net62 mc14500.OEN_l vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_11_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0857_ _0375_ _0376_ _0370_ _0051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_0926_ dest\[3\] _0416_ _0432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_0788_ _0320_ rst_latency\[0\] _0321_ _0037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_input18_I sram_out[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0711_ _0257_ _0249_ _0258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_32_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0642_ _0198_ _0200_ _0201_ _0202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_0573_ _0126_ _0108_ _0132_ _0140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_7_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1056_ net3 net65 mc14500.instr_l\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0909_ dest\[1\] _0416_ _0417_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_22_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput39 net39 io_out[29] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput28 net28 io_out[18] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_27_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_17_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0625_ _0151_ _0149_ _0099_ _0186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_0556_ _0125_ _0126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1108_ _0080_ clknet_3_0__leaf_clk_i net48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1039_ _0026_ clknet_3_4__leaf_clk_i dia\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_17_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0608_ _0160_ _0167_ _0168_ _0158_ _0169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_0539_ net7 _0110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0890_ dest\[15\] _0352_ _0400_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_33_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout63 net64 net63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_0_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0873_ dest\[10\] _0385_ _0388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_0942_ _0444_ _0445_ _0067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_33_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1072_ _0044_ clknet_3_7__leaf_clk_i net40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0787_ _0123_ _0321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0925_ _0328_ _0431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0856_ dest\[4\] _0372_ _0376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1098__CLK clknet_3_3__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0710_ net15 _0257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_0641_ _0095_ _0115_ _0201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_0572_ _0138_ scratch\[1\] _0139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_27_Left_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_11_Left_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1055_ _0040_ net62 mc14500.IEN_l vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_7_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0839_ _0351_ _0363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_0908_ _0403_ _0416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput29 net29 io_out[19] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_34_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0537__I net9 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_17_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0624_ _0166_ _0174_ _0182_ _0184_ _0185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_0555_ net8 _0125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1107_ _0079_ clknet_3_0__leaf_clk_i mar\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_5_Right_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1038_ _0025_ clknet_3_4__leaf_clk_i dia\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_16_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_3_0__f_clk_i_I clknet_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0538_ _0107_ _0108_ _0109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_0607_ _0110_ scratch\[4\] _0168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_21_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_14_Left_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_5_4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_33_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout64 net65 net64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__0622__A1 net10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_0_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0941_ net60 _0411_ _0412_ _0445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_0872_ _0386_ _0387_ _0381_ _0055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_24_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1071_ _0043_ clknet_3_7__leaf_clk_i net39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0924_ _0428_ _0325_ _0429_ _0430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_11_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_0855_ dest\[5\] _0374_ _0375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_0786_ rst_latency\[1\] _0320_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__1002__A1 mc14500.DATA_OUT vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0823__I _0351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0640_ _0158_ _0111_ _0199_ _0178_ _0200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or4_1
X_0571_ _0113_ _0138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_20_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1054_ _0000_ net62 net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_22_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0907_ _0406_ _0333_ _0415_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_0769_ dib\[3\] _0305_ _0306_ _0307_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_0838_ _0210_ _0361_ _0362_ _0046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__0908__I _0403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0643__I _0202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_17_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1088__CLK clknet_3_3__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0623_ _0163_ _0183_ _0184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_0554_ _0105_ _0109_ _0122_ _0124_ _0007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_1106_ _0078_ clknet_3_0__leaf_clk_i mar\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1037_ _0024_ clknet_3_4__leaf_clk_i dia\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_17_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_11_Right_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_3_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_20_Right_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_0537_ net9 _0108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_0606_ scratch\[5\] _0167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_5_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0631__A2 _0185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0622__A2 net9 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout65 net66 net65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_0_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0689__A2 net35 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0940_ dest\[5\] _0405_ _0443_ _0429_ _0444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_27_114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0871_ dest\[8\] _0383_ _0387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_33_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0646__I _0202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__0556__I _0125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1070_ _0008_ clknet_3_7__leaf_clk_i scratch\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0854_ _0351_ _0374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0923_ _0238_ _0429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0785_ _0304_ _0317_ _0319_ _0036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_11_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xwrapped_mc14500_67 io_out[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_14_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0570_ _0105_ _0122_ _0129_ _0137_ _0005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_1053_ _0002_ net66 mc14500.skip vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_0906_ net42 _0414_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0837_ dest\[0\] _0349_ _0318_ _0362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_0768_ _0264_ _0293_ _0306_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_0699_ net13 _0248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__0743__A1 net35 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_input16_I sram_out[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0553_ _0109_ _0122_ _0123_ scratch\[4\] _0124_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA_input8_I io_in[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0622_ net10 net9 _0183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_17_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1105_ _0077_ clknet_3_6__leaf_clk_i net33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_33_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1036_ _0023_ clknet_3_1__leaf_clk_i dia\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_16_223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_3_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0605_ _0159_ _0161_ _0162_ _0165_ _0166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_28_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0536_ _0106_ _0107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1019_ net46 _0502_ _0503_ _0508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__1078__CLK clknet_3_2__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0519_ net6 mc14500.instr_l\[3\] _0085_ _0092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xfanout66 mc14500.X1 net66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_0_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_17 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0870_ dest\[9\] _0385_ _0386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_0_clk_i clk_i clknet_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_0999_ dest\[15\] _0325_ _0492_ _0493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_11_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0853_ _0371_ _0373_ _0370_ _0050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_0922_ net61 _0414_ _0406_ _0428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_0784_ dib\[7\] _0308_ _0318_ _0319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xinput1 SDI net1 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xwrapped_mc14500_68 io_out[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_1052_ _0039_ clknet_3_6__leaf_clk_i net34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XTAP_TAPCELL_ROW_28_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0767_ _0284_ _0305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0836_ _0348_ _0361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0905_ _0410_ _0413_ _0062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_0698_ _0241_ _0245_ _0247_ _0021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_6_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1011__I _0202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0621_ _0176_ _0181_ _0175_ _0182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_0552_ _0113_ _0123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1035_ _0022_ clknet_3_1__leaf_clk_i dia\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1104_ _0076_ clknet_3_6__leaf_clk_i net32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_33_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0819_ _0201_ _0199_ _0184_ _0348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XTAP_TAPCELL_ROW_13_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_9_Right_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_0604_ scratch\[0\] _0164_ _0108_ _0165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_0535_ net8 _0106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1018_ net47 _0500_ _0507_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_5_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0518_ _0089_ _0090_ _0091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_18_Left_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__0607__A1 _0110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0998_ _0326_ _0335_ _0404_ _0492_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XPHY_EDGE_ROW_3_Left_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__0828__A1 net39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0921_ _0427_ _0064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_0783_ _0280_ _0318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_0852_ dest\[3\] _0372_ _0373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_23_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput2 custom_setting net2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__0763__I _0280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xwrapped_mc14500_69 io_out[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__1009__I _0198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1051_ _0038_ clknet_3_7__leaf_clk_i rst_latency\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_3_2__f_clk_i clknet_0_clk_i clknet_3_2__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_7_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0904_ _0406_ _0411_ _0412_ _0413_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_28_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0697_ dia\[0\] _0246_ _0214_ _0247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_0766_ _0286_ _0304_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0835_ _0360_ _0045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__0743__A3 _0211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_6_Left_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_0620_ _0177_ _0178_ _0179_ _0180_ _0145_ _0181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_0551_ _0121_ _0122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1034_ _0021_ clknet_3_1__leaf_clk_i dia\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1103_ _0075_ clknet_3_6__leaf_clk_i net31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_0749_ _0286_ _0291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0818_ _0095_ _0222_ _0041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__0951__I _0403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_32_Left_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_22_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_13_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0603_ _0163_ _0164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_0534_ _0104_ _0105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1017_ _0499_ _0505_ _0506_ _0081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_8_211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_283 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0517_ net5 mc14500.instr_l\[2\] _0085_ _0090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_12_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_35_19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_35_Left_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_25_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0997_ _0488_ _0341_ _0491_ _0475_ _0076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__0828__A2 _0355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0920_ net61 _0420_ _0426_ _0154_ _0427_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_0782_ dib\[6\] _0305_ _0316_ _0317_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_0851_ _0349_ _0372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_23_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_1_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_18_Right_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xinput3 io_in[0] net3 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_27_Right_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_14_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1050_ _0037_ clknet_3_6__leaf_clk_i rst_latency\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0834_ _0185_ mc14500.OEN_l _0359_ _0360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_22_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0903_ _0153_ _0412_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0765_ _0287_ _0301_ _0303_ _0032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_0696_ _0240_ _0246_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_11_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_19_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0550_ _0111_ _0112_ _0113_ _0120_ _0121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_1102_ _0074_ clknet_3_6__leaf_clk_i net30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_33_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1033_ _0020_ clknet_3_1__leaf_clk_i net57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_16_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0817_ _0347_ _0040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_8_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0748_ net12 _0289_ _0290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_0679_ net55 _0217_ _0232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input14_I sram_out[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_0_Right_0 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_22_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0602_ net8 net7 _0163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_21_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0533_ mc14500.DATA_OUT _0104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA_input6_I io_in[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1016_ net47 _0502_ _0503_ _0506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_12_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0516_ _0087_ _0089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout58 net28 net58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__1091__CLK clknet_3_2__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0996_ dest\[14\] _0421_ _0490_ _0238_ _0491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_0850_ dest\[4\] _0363_ _0371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_0781_ _0277_ _0288_ _0316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_11_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput4 io_in[1] net4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_1_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0979_ dest\[11\] _0453_ _0477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_7_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0833_ _0100_ _0345_ _0359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_0902_ _0337_ _0411_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0695_ net12 _0244_ _0245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_0764_ dib\[3\] _0291_ _0302_ _0303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_6_184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1101_ _0073_ clknet_3_6__leaf_clk_i net29 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_1032_ _0019_ clknet_3_1__leaf_clk_i net56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_17_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_16_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_8_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0747_ _0288_ _0289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_3_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0816_ _0185_ mc14500.IEN_l _0346_ _0347_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_35_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0678_ _0227_ _0229_ _0231_ _0017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_22_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_15_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0601_ _0107_ _0160_ scratch\[1\] _0162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_0532_ _0103_ net49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_28_20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1015_ net48 _0500_ _0505_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__0619__A1 _0171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_285 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_4_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0515_ _0084_ _0086_ _0087_ _0088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xfanout59 net26 net59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_26_141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0995_ _0488_ _0335_ _0489_ _0490_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_17_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0636__C _0136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0780_ _0304_ _0314_ _0315_ _0035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_11_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_23_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_1_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput5 io_in[2] net5 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_14_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1081__CLK clknet_3_2__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0978_ _0464_ _0470_ _0476_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__0682__A2 _0217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0647__B _0138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0832_ _0210_ _0357_ _0358_ _0321_ _0044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_0763_ _0280_ _0302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_22_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0901_ dest\[0\] _0405_ _0409_ _0410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_0694_ _0243_ _0244_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_11_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1100_ _0072_ clknet_3_3__leaf_clk_i net28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1031_ _0018_ clknet_3_1__leaf_clk_i net55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_17_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_16_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0746_ _0284_ _0288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_0815_ _0149_ _0099_ _0345_ _0346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_0677_ _0230_ _0231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__0582__A1 _0132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_15_250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_22_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0531_ _0096_ _0100_ _0102_ _0103_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_0600_ _0125_ _0160_ scratch\[3\] _0161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_1014_ _0499_ _0501_ _0504_ _0080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_8_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0729_ net18 _0273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__0794__A1 net33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_4_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0514_ mc14500.skip _0087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__1038__CLK clknet_3_4__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_3_5__f_clk_i clknet_0_clk_i clknet_3_5__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_0994_ _0488_ _0331_ _0324_ _0489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_10_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_17_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_23_Left_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_1_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput6 io_in[3] net6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_0977_ _0221_ _0475_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_9_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_14_Right_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_20_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_23_Right_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_32_Right_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_0900_ _0406_ _0407_ _0408_ _0409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_0693_ _0242_ _0243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0762_ dib\[2\] _0289_ _0300_ _0301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_11_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0831_ net40 _0357_ _0358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_10_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_25_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1030_ _0017_ clknet_3_1__leaf_clk_i net54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_17_56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0814_ _0188_ _0189_ _0345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_16_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1001__C _0230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_26_Left_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_0745_ _0286_ _0287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_10_Left_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_0676_ _0221_ _0230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__1094__CLK clknet_3_2__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0530_ _0101_ _0102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_28_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1013_ net48 _0502_ _0503_ _0504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_8_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_4_Right_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_0728_ _0262_ _0271_ _0272_ _0026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_0659_ _0183_ _0216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA_input12_I sram_out[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_10_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_33_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_4_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0513_ net3 mc14500.instr_l\[0\] _0085_ _0086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_input4_I io_in[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0993_ net32 _0488_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_26_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput7 io_in[4] net7 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_0976_ _0474_ _0072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_14_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0600__A1 _0125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0658__A1 _0210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0928__C _0154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0830__A1 _0211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0830_ _0211_ _0354_ _0357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_0761_ _0257_ _0293_ _0300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_11_105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0692_ _0158_ _0130_ _0183_ _0242_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_TAPCELL_ROW_19_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0959_ net59 _0459_ _0453_ _0460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_27_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_25_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput10 io_in[7] net10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_0813_ _0339_ _0342_ _0344_ _0039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_0675_ net53 _0228_ _0229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_0744_ _0284_ _0285_ _0201_ _0286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__0584__B _0136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1089_ _0061_ clknet_3_3__leaf_clk_i dest\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_15_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0573__A3 _0132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1012_ _0280_ _0503_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0727_ dia\[5\] _0267_ _0260_ _0272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_12_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_0658_ _0210_ _0213_ _0215_ _0013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_0589_ _0151_ _0102_ _0152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_7_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_10_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_33_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_4_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0512_ net63 _0085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__1084__CLK clknet_3_2__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0992_ _0420_ _0486_ _0487_ _0475_ _0075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_5_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0592__B _0154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0685__A2 _0217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output36_I net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput8 io_in[5] net8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_0975_ net58 _0411_ _0473_ _0412_ _0474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_0760_ _0287_ _0298_ _0299_ _0031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_0691_ _0240_ _0241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_11_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_19_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0889_ _0398_ _0399_ _0392_ _0060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_0958_ _0431_ _0329_ _0459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_10_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_25_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0576__A1 _0138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput11 rst_n net11 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_0743_ net35 _0216_ _0211_ _0285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_0812_ _0343_ _0344_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0674_ _0212_ _0228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__0584__C net37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1088_ _0060_ clknet_3_3__leaf_clk_i dest\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_21_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1011_ _0202_ _0502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_28_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0726_ dia\[4\] _0263_ _0270_ _0271_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_0657_ net50 _0212_ _0214_ _0215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_0588_ net36 _0151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XTAP_TAPCELL_ROW_10_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0614__I net10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__0524__I _0095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0511_ net4 mc14500.instr_l\[1\] net63 _0084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_30_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0709_ _0241_ _0255_ _0256_ _0023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_35_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0991_ _0464_ _0482_ net31 _0487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_1_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput9 io_in[6] net9 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_14_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0974_ _0470_ _0471_ _0408_ _0472_ _0473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_22_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1097__CLK clknet_3_3__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0690_ _0238_ _0239_ _0240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_EDGE_ROW_10_Right_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_19_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0888_ dest\[13\] _0394_ _0399_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_0957_ dest\[8\] _0405_ _0458_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_25_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0567__A2 _0109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0673_ net54 _0218_ _0227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xinput12 sram_out[0] net12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_0811_ _0221_ _0343_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_0742_ _0164_ _0283_ _0284_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_1087_ _0059_ clknet_3_3__leaf_clk_i dest\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_15_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_21_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1010_ mar\[1\] _0500_ _0501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_0725_ _0269_ _0243_ _0270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_0656_ _0153_ _0214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0587_ _0149_ _0099_ _0150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_19_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_10_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0540__I _0110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_8_Right_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__0630__A1 net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0708_ dia\[2\] _0246_ _0214_ _0256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_0639_ _0091_ _0114_ _0118_ _0199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA_input10_I io_in[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_25_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0990_ dest\[13\] _0325_ _0485_ _0486_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_5_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input2_I custom_setting vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_17_Left_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_0973_ dest\[10\] _0440_ _0472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_2_Left_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_28_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_19_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0956_ net59 _0457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_0887_ dest\[14\] _0352_ _0398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_10_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput13 sram_out[1] net13 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_0810_ net34 _0340_ _0341_ _0342_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_0672_ _0225_ _0226_ _0222_ _0016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_0741_ _0112_ _0128_ _0283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_24_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1086_ _0058_ clknet_3_3__leaf_clk_i dest\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_15_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1087__CLK clknet_3_3__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0939_ _0440_ _0441_ _0442_ _0443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XTAP_TAPCELL_ROW_7_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_13_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_5_Left_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_21_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0655_ _0212_ _0213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0724_ net17 _0269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_0586_ _0098_ _0149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_12_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_35_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1069_ _0006_ clknet_3_7__leaf_clk_i scratch\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_31_Left_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_0707_ dia\[1\] _0244_ _0254_ _0255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_20_71 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0638_ _0097_ _0098_ _0086_ _0102_ _0198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_0569_ _0121_ _0129_ _0136_ scratch\[2\] _0137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_29_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0679__A2 _0217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_34_Left_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_0972_ net58 _0462_ _0471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_22_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_28_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0886_ _0396_ _0397_ _0392_ _0059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_0955_ _0402_ _0456_ _0069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_33_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput14 sram_out[2] net14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_0740_ _0262_ _0279_ _0282_ _0028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_0671_ net52 _0213_ _0226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1085_ _0057_ clknet_3_3__leaf_clk_i dest\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_23_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0869_ _0351_ _0385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_23_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0938_ _0435_ _0431_ net60 _0442_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_7_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0644__I _0198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_13_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_21_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0723_ _0262_ _0266_ _0268_ _0025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_0654_ _0119_ _0183_ _0211_ _0212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_0585_ _0104_ _0122_ _0146_ _0148_ _0009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA_clkbuf_3_7__f_clk_i_I clknet_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_35_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1068_ _0007_ clknet_3_7__leaf_clk_i scratch\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_30_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1077__CLK clknet_3_2__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0706_ _0253_ _0249_ _0254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_0637_ _0187_ _0196_ _0197_ _0000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_0568_ _0113_ _0136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_35_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0971_ _0324_ _0469_ _0470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_22_140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0737__I _0131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0557__I net9 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0885_ dest\[12\] _0394_ _0397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_0954_ net25 _0451_ _0455_ _0338_ _0456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_33_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0670_ net53 _0218_ _0225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xinput15 sram_out[3] net15 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1084_ _0056_ clknet_3_2__leaf_clk_i dest\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_15_246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0868_ _0382_ _0384_ _0381_ _0054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_30_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0799_ net31 net30 _0327_ _0330_ _0331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_0937_ net60 _0435_ _0328_ _0441_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XTAP_TAPCELL_ROW_7_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_21_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0642__A1 _0198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0722_ dia\[4\] _0267_ _0260_ _0268_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_0653_ _0106_ _0171_ _0211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_0584_ _0121_ _0146_ _0136_ net37 _0148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_1067_ _0009_ clknet_3_7__leaf_clk_i net37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_35_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0655__I _0212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0705_ net14 _0253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_0636_ net36 _0194_ _0115_ _0136_ _0197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_0567_ _0105_ _0109_ _0133_ _0135_ _0008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_17_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_17_Right_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_26_Right_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_25_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_35_Right_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1044__CLK clknet_3_4__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_3_1__f_clk_i clknet_0_clk_i clknet_3_1__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_0_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0619_ _0171_ net1 _0180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__0818__A1 _0095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0970_ net58 _0462_ _0469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_22_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0884_ dest\[13\] _0352_ _0396_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_0953_ net25 _0407_ _0447_ _0454_ _0455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_10_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_10_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput16 sram_out[4] net16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_24_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1083_ _0055_ clknet_3_2__leaf_clk_i dest\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_23_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0936_ _0403_ _0440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_0798_ net27 net59 _0328_ _0329_ _0330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XTAP_TAPCELL_ROW_7_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0867_ dest\[7\] _0383_ _0384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_30_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input19_I sram_out[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1012__I _0280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0721_ _0240_ _0267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0652_ _0104_ _0210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_0583_ _0104_ _0133_ _0146_ _0147_ _0010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_20_283 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_35_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1066_ _0010_ clknet_3_7__leaf_clk_i net38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_7_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0919_ _0421_ _0423_ _0424_ _0425_ _0426_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_11_250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_9_Left_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__0936__I _0403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_32_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0704_ _0241_ _0251_ _0252_ _0022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_0635_ _0192_ _0195_ _0196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_20_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0566_ _0109_ _0132_ _0123_ scratch\[5\] _0135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_29_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1049_ _0036_ clknet_3_5__leaf_clk_i dib\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_26_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_31_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0549_ _0119_ _0120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_0618_ _0125_ _0171_ _0179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_23_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_22_Left_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__0854__I _0351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0952_ dest\[7\] _0453_ _0454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_10_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0883_ _0393_ _0395_ _0392_ _0058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__0674__I _0212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_24_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput17 sram_out[5] net17 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1082_ _0054_ clknet_3_2__leaf_clk_i dest\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__0660__A3 _0211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0866_ _0349_ _0383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0935_ _0439_ _0066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_30_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0797_ net25 net24 net60 net22 _0329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_21_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0720_ dia\[3\] _0263_ _0265_ _0266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_0651_ _0203_ _0208_ _0209_ _0012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_0582_ _0132_ _0146_ _0136_ net38 _0147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XPHY_EDGE_ROW_25_Left_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1065_ _0042_ clknet_3_6__leaf_clk_i dest\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0849_ _0368_ _0369_ _0370_ _0049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_0918_ _0337_ _0425_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_32_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0703_ dia\[1\] _0246_ _0214_ _0252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_20_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_20_75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0565_ _0105_ _0129_ _0133_ _0134_ _0006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_0634_ _0100_ _0156_ _0193_ _0194_ _0195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_1048_ _0035_ clknet_3_5__leaf_clk_i dib\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_3_Right_3 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_9_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_3_6__f_clk_i_I clknet_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1090__CLK clknet_3_2__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0548_ _0091_ _0114_ _0116_ _0118_ _0119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_0617_ net10 _0127_ _0178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_22_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_16_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0677__I _0230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0882_ dest\[11\] _0394_ _0395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_0951_ _0403_ _0453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_10_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput18 sram_out[6] net18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_24_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1081_ _0053_ clknet_3_2__leaf_clk_i dest\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0865_ dest\[8\] _0374_ _0382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_0934_ _0435_ _0420_ _0438_ _0412_ _0439_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_TAPCELL_ROW_30_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0796_ net21 net61 net42 net41 _0328_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_23_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0636__A1 net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0650_ net43 _0206_ _0138_ _0209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_20_285 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0581_ _0145_ _0146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_18_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1064_ _0005_ clknet_3_6__leaf_clk_i scratch\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__0618__A1 _0125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0779_ dib\[6\] _0308_ _0302_ _0315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_0917_ dest\[2\] _0416_ _0424_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_0848_ _0343_ _0370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_32_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0702_ dia\[0\] _0244_ _0250_ _0251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_0633_ _0155_ _0188_ _0189_ _0194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_20_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0564_ _0129_ _0133_ _0123_ scratch\[3\] _0134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_1047_ _0034_ clknet_3_5__leaf_clk_i dib\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_13_Right_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_15_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_22_Right_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_31_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0616_ dia\[7\] _0177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_0547_ _0097_ _0084_ _0117_ _0118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XPHY_EDGE_ROW_31_Right_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__0783__I _0280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_6_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1080__CLK clknet_3_2__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0950_ _0402_ _0452_ _0068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_12_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0881_ _0348_ _0394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_18_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput19 sram_out[7] net19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_24_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1080_ _0052_ clknet_3_2__leaf_clk_i dest\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0864_ _0379_ _0380_ _0381_ _0053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_0933_ _0407_ _0436_ _0437_ _0425_ _0438_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_30_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0795_ net29 net58 _0327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_2_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0572__A1 _0138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0650__B _0138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0580_ _0125_ _0127_ _0145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__0618__A2 _0171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1063_ _0004_ clknet_3_6__leaf_clk_i scratch\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0916_ net61 _0422_ _0423_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_0778_ dib\[5\] _0305_ _0313_ _0314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xclkbuf_3_4__f_clk_i clknet_0_clk_i clknet_3_4__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_0847_ dest\[2\] _0361_ _0369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input17_I sram_out[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0545__A1 _0095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_32_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0563_ _0132_ _0133_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0701_ _0248_ _0249_ _0250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_0632_ _0188_ _0189_ _0193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA_input9_I io_in[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1046_ _0033_ clknet_3_5__leaf_clk_i dib\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_9_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1037__CLK clknet_3_4__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0546_ mc14500.OEN_l _0117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_0615_ dib\[7\] _0175_ _0127_ _0164_ _0176_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_1029_ _0016_ clknet_3_1__leaf_clk_i net53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_16_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0529_ _0089_ _0090_ _0092_ _0101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_8_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_27_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0880_ dest\[12\] _0385_ _0393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_18_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0654__A3 _0211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0920__C _0154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0932_ dest\[4\] _0416_ _0437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_23_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0863_ _0343_ _0381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_0794_ net33 net32 _0326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_6_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_12_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1093__CLK clknet_3_2__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_35_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0892__I _0230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1062_ _0003_ clknet_3_4__leaf_clk_i scratch\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0915_ _0414_ net41 _0422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_0777_ _0273_ _0288_ _0313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_0846_ dest\[3\] _0363_ _0368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__0554__A2 _0109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0700_ _0242_ _0249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_29_Left_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_0631_ mc14500.IEN_l _0185_ _0191_ _0150_ _0192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_0562_ _0130_ _0112_ _0131_ _0120_ _0132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XPHY_EDGE_ROW_13_Left_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1045_ _0032_ clknet_3_5__leaf_clk_i dib\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_28_151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0829_ _0210_ _0355_ _0356_ _0321_ _0043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_19_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_7_Right_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_0545_ _0095_ _0115_ _0116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_0614_ net10 _0175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1028_ _0015_ clknet_3_0__leaf_clk_i net52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_26_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_3_5__f_clk_i_I clknet_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0528_ _0098_ _0099_ _0100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XPHY_EDGE_ROW_16_Left_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_8_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_27_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0895__I _0403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_1_Left_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_17_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0862_ dest\[6\] _0372_ _0380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_0931_ _0435_ _0431_ _0436_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_0793_ _0324_ _0325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_6_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_12_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_35_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1061_ _0041_ clknet_3_0__leaf_clk_i mc14500.X1 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0845_ _0366_ _0367_ _0344_ _0048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_0914_ _0404_ _0421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0776_ _0304_ _0311_ _0312_ _0034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__0569__B _0136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_4_Left_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_0561_ net11 _0131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_0630_ net36 _0100_ _0156_ _0190_ _0191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_20_79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1044_ _0031_ clknet_3_4__leaf_clk_i dib\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_28_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0828_ net39 _0355_ _0356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_0759_ dib\[2\] _0291_ _0281_ _0299_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_9_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1083__CLK clknet_3_2__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_30_Left_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_15_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0613_ _0128_ _0169_ _0173_ _0112_ _0174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_0_25_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0544_ rst_latency\[1\] rst_latency\[0\] _0115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_0_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1027_ _0014_ clknet_3_1__leaf_clk_i net51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__0582__B _0136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0527_ _0097_ _0086_ _0099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_13_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_8_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0657__A2 _0212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_27_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_2_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0930_ net22 _0435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0861_ dest\[7\] _0374_ _0379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_23_79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0792_ _0323_ _0324_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__0566__A1 _0109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_6_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_29_Right_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_12_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1060_ _0001_ net62 mc14500.DATA_OUT vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_35_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_0_clk_i_I clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0775_ dib\[5\] _0308_ _0302_ _0312_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_11_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0844_ dest\[1\] _0361_ _0367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_0913_ _0408_ _0420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_4_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0560_ _0110_ _0130_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1043_ _0030_ clknet_3_4__leaf_clk_i dib\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_9_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0758_ dib\[1\] _0289_ _0297_ _0298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_0827_ _0107_ _0130_ _0354_ _0355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_0689_ _0126_ net35 _0216_ _0130_ _0239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA_input15_I sram_out[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_31_35 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0612_ _0160_ _0170_ _0172_ _0107_ _0173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XANTENNA_input7_I io_in[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0543_ _0089_ _0092_ _0114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1026_ _0013_ clknet_3_0__leaf_clk_i net50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_16_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_26_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0526_ _0097_ _0084_ _0098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_1009_ _0198_ _0500_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_12_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_27_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_2_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1096__CLK clknet_3_3__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_3_7__f_clk_i clknet_0_clk_i clknet_3_7__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_2_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0860_ _0377_ _0378_ _0370_ _0052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_0791_ _0155_ _0102_ _0323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__0566__A2 _0132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0989_ _0335_ _0453_ _0485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_TAPCELL_ROW_6_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_12_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_35_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0912_ _0402_ _0419_ _0063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_0774_ dib\[4\] _0305_ _0310_ _0311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_0843_ dest\[2\] _0363_ _0366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1042_ _0029_ clknet_3_1__leaf_clk_i dib\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1111_ _0083_ clknet_3_0__leaf_clk_i net45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_0_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_31_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0757_ _0253_ _0293_ _0297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_10_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0688_ _0201_ _0238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0826_ _0120_ _0283_ _0354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_19_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_5_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0542_ net11 _0113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_0611_ _0171_ net37 _0172_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__0611__A1 _0171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1025_ _0012_ clknet_3_0__leaf_clk_i net43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_16_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0809_ _0238_ _0341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__0832__A1 _0210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0525_ _0089_ _0097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_21_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1008_ _0202_ _0499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_29_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0784__B _0318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output39_I net39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_285 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_2_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_9_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_3_4__f_clk_i_I clknet_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_15_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0961__C _0230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0533__I mc14500.DATA_OUT vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0790_ _0321_ _0322_ _0038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_3_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0988_ _0480_ _0341_ _0484_ _0475_ _0074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_1_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1086__CLK clknet_3_3__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0842_ _0364_ _0365_ _0344_ _0047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_0911_ _0414_ _0409_ _0418_ _0411_ _0419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_0773_ _0269_ _0288_ _0310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1110_ _0082_ clknet_3_0__leaf_clk_i net46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_29_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1041_ _0028_ clknet_3_5__leaf_clk_i dia\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0825_ _0350_ _0353_ _0344_ _0042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_31_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0687_ _0236_ _0237_ _0231_ _0020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_0756_ _0287_ _0295_ _0296_ _0030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_19_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_34_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_8_Left_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_15_38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0541__I net10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_5_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0611__A2 net37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0610_ net7 _0171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_0541_ net10 _0112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_1024_ _0011_ clknet_3_0__leaf_clk_i net44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0808_ net2 _0340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_31_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0739_ dia\[7\] _0267_ _0281_ _0282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_26_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0524_ _0095_ _0096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1007_ _0203_ _0497_ _0498_ _0079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_8_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__0578__A1 mc14500.DATA_OUT vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_2_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput50 net50 sram_in[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_5_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_27_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_9_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_15_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_21_Left_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_23_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0987_ dest\[12\] _0421_ _0483_ _0484_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_0_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_16_Right_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_7_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0772_ _0304_ _0307_ _0309_ _0033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_0841_ dest\[0\] _0361_ _0365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_25_Right_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_0910_ _0414_ _0415_ _0417_ _0418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_34_Right_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_6_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1040_ _0027_ clknet_3_5__leaf_clk_i dia\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_31_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0755_ dib\[1\] _0291_ _0281_ _0296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_9_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0824_ _0340_ dest\[16\] _0352_ _0353_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XPHY_EDGE_ROW_24_Left_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_0686_ net56 _0228_ _0237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_10_83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_5_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0540_ _0110_ _0111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__1099__CLK clknet_3_3__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1023_ _0499_ _0509_ _0510_ _0083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_16_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0738_ _0280_ _0281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0807_ dest\[16\] _0325_ _0334_ _0336_ _0338_ _0339_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_0669_ _0223_ _0224_ _0222_ _0015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XPHY_EDGE_ROW_2_Right_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_input13_I sram_out[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input5_I io_in[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0523_ _0085_ _0095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1006_ mar\[1\] _0206_ _0318_ _0498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xoutput51 net51 sram_in[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput40 net40 io_out[30] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XTAP_TAPCELL_ROW_9_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_15_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_23_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0986_ _0480_ _0481_ _0482_ _0408_ _0483_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_0771_ dib\[4\] _0308_ _0302_ _0309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_0840_ dest\[1\] _0363_ _0364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__0641__A1 _0095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0560__I _0110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0969_ _0468_ _0071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_10_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_3_0__f_clk_i clknet_0_clk_i clknet_3_0__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_28_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_31_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0754_ dib\[0\] _0289_ _0294_ _0295_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_3_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0685_ net57 _0217_ _0236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_0823_ _0351_ _0352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_19_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1099_ _0071_ clknet_3_3__leaf_clk_i net27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_19_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_5_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1022_ net45 _0502_ _0503_ _0510_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_21_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0668_ net51 _0213_ _0224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1043__CLK clknet_3_4__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0737_ _0131_ _0280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0806_ _0337_ _0338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_34_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0599_ _0110_ _0160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_13_108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0522_ _0094_ net35 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1005_ mar\[0\] _0204_ _0497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_8_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_32_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1089__CLK clknet_3_3__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput30 net30 io_out[20] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput41 net41 io_out[8] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput52 net52 sram_in[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XTAP_TAPCELL_ROW_26_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0563__I _0132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
.ends

