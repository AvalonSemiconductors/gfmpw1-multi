magic
tech gf180mcuD
magscale 1 10
timestamp 1753965783
<< metal1 >>
rect 1344 32170 34608 32204
rect 1344 32118 5372 32170
rect 5424 32118 5476 32170
rect 5528 32118 5580 32170
rect 5632 32118 13688 32170
rect 13740 32118 13792 32170
rect 13844 32118 13896 32170
rect 13948 32118 22004 32170
rect 22056 32118 22108 32170
rect 22160 32118 22212 32170
rect 22264 32118 30320 32170
rect 30372 32118 30424 32170
rect 30476 32118 30528 32170
rect 30580 32118 34608 32170
rect 1344 32084 34608 32118
rect 13122 31838 13134 31890
rect 13186 31838 13198 31890
rect 19618 31838 19630 31890
rect 19682 31838 19694 31890
rect 16158 31778 16210 31790
rect 13458 31726 13470 31778
rect 13522 31726 13534 31778
rect 19170 31726 19182 31778
rect 19234 31726 19246 31778
rect 13290 31670 13302 31722
rect 13354 31670 13366 31722
rect 16158 31714 16210 31726
rect 19450 31670 19462 31722
rect 19514 31670 19526 31722
rect 15822 31554 15874 31566
rect 15822 31490 15874 31502
rect 1344 31386 34768 31420
rect 1344 31334 9530 31386
rect 9582 31334 9634 31386
rect 9686 31334 9738 31386
rect 9790 31334 17846 31386
rect 17898 31334 17950 31386
rect 18002 31334 18054 31386
rect 18106 31334 26162 31386
rect 26214 31334 26266 31386
rect 26318 31334 26370 31386
rect 26422 31334 34478 31386
rect 34530 31334 34582 31386
rect 34634 31334 34686 31386
rect 34738 31334 34768 31386
rect 1344 31300 34768 31334
rect 13918 30994 13970 31006
rect 13122 30942 13134 30994
rect 13186 30942 13198 30994
rect 13918 30930 13970 30942
rect 14030 30994 14082 31006
rect 21310 30994 21362 31006
rect 14802 30942 14814 30994
rect 14866 30942 14878 30994
rect 20514 30942 20526 30994
rect 20578 30942 20590 30994
rect 14030 30930 14082 30942
rect 21310 30930 21362 30942
rect 21870 30994 21922 31006
rect 21870 30930 21922 30942
rect 25678 30994 25730 31006
rect 25678 30930 25730 30942
rect 27246 30994 27298 31006
rect 27246 30930 27298 30942
rect 25342 30882 25394 30894
rect 11218 30830 11230 30882
rect 11282 30830 11294 30882
rect 16706 30830 16718 30882
rect 16770 30830 16782 30882
rect 18610 30830 18622 30882
rect 18674 30830 18686 30882
rect 22642 30830 22654 30882
rect 22706 30830 22718 30882
rect 24546 30830 24558 30882
rect 24610 30830 24622 30882
rect 25342 30818 25394 30830
rect 27582 30770 27634 30782
rect 27582 30706 27634 30718
rect 1344 30602 34608 30636
rect 1344 30550 5372 30602
rect 5424 30550 5476 30602
rect 5528 30550 5580 30602
rect 5632 30550 13688 30602
rect 13740 30550 13792 30602
rect 13844 30550 13896 30602
rect 13948 30550 22004 30602
rect 22056 30550 22108 30602
rect 22160 30550 22212 30602
rect 22264 30550 30320 30602
rect 30372 30550 30424 30602
rect 30476 30550 30528 30602
rect 30580 30550 34608 30602
rect 1344 30516 34608 30550
rect 19966 30434 20018 30446
rect 17826 30326 17838 30378
rect 17890 30326 17902 30378
rect 19966 30370 20018 30382
rect 27906 30270 27918 30322
rect 27970 30270 27982 30322
rect 9662 30210 9714 30222
rect 13582 30210 13634 30222
rect 10434 30158 10446 30210
rect 10498 30158 10510 30210
rect 9662 30146 9714 30158
rect 13582 30146 13634 30158
rect 14702 30210 14754 30222
rect 16382 30210 16434 30222
rect 15698 30158 15710 30210
rect 15762 30158 15774 30210
rect 12350 30098 12402 30110
rect 13813 30102 13825 30154
rect 13877 30102 13889 30154
rect 14702 30146 14754 30158
rect 16034 30102 16046 30154
rect 16098 30102 16110 30154
rect 16382 30146 16434 30158
rect 16830 30210 16882 30222
rect 16830 30146 16882 30158
rect 17054 30210 17106 30222
rect 18846 30210 18898 30222
rect 17714 30158 17726 30210
rect 17778 30158 17790 30210
rect 18050 30158 18062 30210
rect 18114 30158 18126 30210
rect 17054 30146 17106 30158
rect 18846 30146 18898 30158
rect 20302 30210 20354 30222
rect 19710 30102 19722 30154
rect 19774 30102 19786 30154
rect 20302 30146 20354 30158
rect 21646 30210 21698 30222
rect 24670 30210 24722 30222
rect 22418 30158 22430 30210
rect 22482 30158 22494 30210
rect 21646 30146 21698 30158
rect 24670 30146 24722 30158
rect 24894 30210 24946 30222
rect 24894 30146 24946 30158
rect 28702 30210 28754 30222
rect 28702 30146 28754 30158
rect 29318 30210 29370 30222
rect 29318 30146 29370 30158
rect 20638 30098 20690 30110
rect 17322 30046 17334 30098
rect 17386 30046 17398 30098
rect 12350 30034 12402 30046
rect 12966 29986 13018 29998
rect 16258 29990 16270 30042
rect 16322 29990 16334 30042
rect 20638 30034 20690 30046
rect 24334 30098 24386 30110
rect 26014 30098 26066 30110
rect 25162 30046 25174 30098
rect 25226 30046 25238 30098
rect 24334 30034 24386 30046
rect 26014 30034 26066 30046
rect 12966 29922 13018 29934
rect 1344 29818 34768 29852
rect 1344 29766 9530 29818
rect 9582 29766 9634 29818
rect 9686 29766 9738 29818
rect 9790 29766 17846 29818
rect 17898 29766 17950 29818
rect 18002 29766 18054 29818
rect 18106 29766 26162 29818
rect 26214 29766 26266 29818
rect 26318 29766 26370 29818
rect 26422 29766 34478 29818
rect 34530 29766 34582 29818
rect 34634 29766 34686 29818
rect 34738 29766 34768 29818
rect 1344 29732 34768 29766
rect 12786 29542 12798 29594
rect 12850 29542 12862 29594
rect 16034 29542 16046 29594
rect 16098 29542 16110 29594
rect 19618 29542 19630 29594
rect 19682 29542 19694 29594
rect 23426 29542 23438 29594
rect 23490 29542 23502 29594
rect 25778 29542 25790 29594
rect 25842 29542 25854 29594
rect 27682 29542 27694 29594
rect 27746 29542 27758 29594
rect 14634 29486 14646 29538
rect 14698 29486 14710 29538
rect 20458 29486 20470 29538
rect 20522 29486 20534 29538
rect 11778 29418 11790 29470
rect 11842 29418 11854 29470
rect 12114 29374 12126 29426
rect 12178 29374 12190 29426
rect 12674 29389 12686 29441
rect 12738 29389 12750 29441
rect 13358 29426 13410 29438
rect 12898 29374 12910 29426
rect 12962 29374 12974 29426
rect 13358 29362 13410 29374
rect 13470 29426 13522 29438
rect 13470 29362 13522 29374
rect 14254 29426 14306 29438
rect 14254 29362 14306 29374
rect 14366 29426 14418 29438
rect 15922 29418 15934 29470
rect 15986 29418 15998 29470
rect 16258 29374 16270 29426
rect 16322 29374 16334 29426
rect 18162 29374 18174 29426
rect 18226 29374 18238 29426
rect 18386 29418 18398 29470
rect 18450 29418 18462 29470
rect 18946 29374 18958 29426
rect 19010 29374 19022 29426
rect 19170 29401 19182 29453
rect 19234 29401 19246 29453
rect 19518 29426 19570 29438
rect 14366 29362 14418 29374
rect 19518 29362 19570 29374
rect 19966 29426 20018 29438
rect 19966 29362 20018 29374
rect 20190 29426 20242 29438
rect 20190 29362 20242 29374
rect 20750 29426 20802 29438
rect 22642 29374 22654 29426
rect 22706 29374 22718 29426
rect 22866 29418 22878 29470
rect 22930 29418 22942 29470
rect 23314 29374 23326 29426
rect 23378 29374 23390 29426
rect 23650 29401 23662 29453
rect 23714 29401 23726 29453
rect 23998 29426 24050 29438
rect 25218 29374 25230 29426
rect 25282 29374 25294 29426
rect 25554 29401 25566 29453
rect 25618 29401 25630 29453
rect 25902 29426 25954 29438
rect 26898 29374 26910 29426
rect 26962 29374 26974 29426
rect 27234 29401 27246 29453
rect 27298 29401 27310 29453
rect 27582 29426 27634 29438
rect 20750 29362 20802 29374
rect 23998 29362 24050 29374
rect 25902 29362 25954 29374
rect 27582 29362 27634 29374
rect 11666 29262 11678 29314
rect 11730 29262 11742 29314
rect 18498 29262 18510 29314
rect 18562 29262 18574 29314
rect 22978 29262 22990 29314
rect 23042 29262 23054 29314
rect 21086 29202 21138 29214
rect 13738 29150 13750 29202
rect 13802 29150 13814 29202
rect 21086 29138 21138 29150
rect 1344 29034 34608 29068
rect 1344 28982 5372 29034
rect 5424 28982 5476 29034
rect 5528 28982 5580 29034
rect 5632 28982 13688 29034
rect 13740 28982 13792 29034
rect 13844 28982 13896 29034
rect 13948 28982 22004 29034
rect 22056 28982 22108 29034
rect 22160 28982 22212 29034
rect 22264 28982 30320 29034
rect 30372 28982 30424 29034
rect 30476 28982 30528 29034
rect 30580 28982 34608 29034
rect 1344 28948 34608 28982
rect 14198 28866 14250 28878
rect 22990 28866 23042 28878
rect 14198 28802 14250 28814
rect 15038 28810 15090 28822
rect 15418 28814 15430 28866
rect 15482 28814 15494 28866
rect 25722 28814 25734 28866
rect 25786 28814 25798 28866
rect 12966 28754 13018 28766
rect 12338 28702 12350 28754
rect 12402 28702 12414 28754
rect 22990 28802 23042 28814
rect 15038 28746 15090 28758
rect 18162 28702 18174 28754
rect 18226 28702 18238 28754
rect 20066 28702 20078 28754
rect 20130 28702 20142 28754
rect 23986 28702 23998 28754
rect 24050 28702 24062 28754
rect 27122 28702 27134 28754
rect 27186 28702 27198 28754
rect 12966 28690 13018 28702
rect 9662 28642 9714 28654
rect 13470 28642 13522 28654
rect 10434 28590 10446 28642
rect 10498 28590 10510 28642
rect 9662 28578 9714 28590
rect 13470 28578 13522 28590
rect 13638 28642 13690 28654
rect 13918 28642 13970 28654
rect 15710 28642 15762 28654
rect 13794 28590 13806 28642
rect 13858 28590 13870 28642
rect 14690 28590 14702 28642
rect 14754 28590 14766 28642
rect 14914 28590 14926 28642
rect 14978 28590 14990 28642
rect 13638 28578 13690 28590
rect 13918 28578 13970 28590
rect 15710 28578 15762 28590
rect 15822 28642 15874 28654
rect 15822 28578 15874 28590
rect 17614 28642 17666 28654
rect 17614 28578 17666 28590
rect 17838 28642 17890 28654
rect 17838 28578 17890 28590
rect 20862 28642 20914 28654
rect 20862 28578 20914 28590
rect 23326 28642 23378 28654
rect 24446 28642 24498 28654
rect 23762 28590 23774 28642
rect 23826 28590 23838 28642
rect 23326 28578 23378 28590
rect 24098 28563 24110 28615
rect 24162 28563 24174 28615
rect 24446 28578 24498 28590
rect 24782 28642 24834 28654
rect 24782 28578 24834 28590
rect 25230 28642 25282 28654
rect 25230 28578 25282 28590
rect 25454 28642 25506 28654
rect 27358 28642 27410 28654
rect 26674 28590 26686 28642
rect 26738 28590 26750 28642
rect 25454 28578 25506 28590
rect 27010 28546 27022 28598
rect 27074 28546 27086 28598
rect 27358 28578 27410 28590
rect 27582 28642 27634 28654
rect 27582 28578 27634 28590
rect 17322 28478 17334 28530
rect 17386 28478 17398 28530
rect 27850 28478 27862 28530
rect 27914 28478 27926 28530
rect 1344 28250 34768 28284
rect 1344 28198 9530 28250
rect 9582 28198 9634 28250
rect 9686 28198 9738 28250
rect 9790 28198 17846 28250
rect 17898 28198 17950 28250
rect 18002 28198 18054 28250
rect 18106 28198 26162 28250
rect 26214 28198 26266 28250
rect 26318 28198 26370 28250
rect 26422 28198 34478 28250
rect 34530 28198 34582 28250
rect 34634 28198 34686 28250
rect 34738 28198 34768 28250
rect 1344 28164 34768 28198
rect 11118 28082 11170 28094
rect 11118 28018 11170 28030
rect 12338 27974 12350 28026
rect 12402 27974 12414 28026
rect 16718 27970 16770 27982
rect 27010 27974 27022 28026
rect 27074 27974 27086 28026
rect 28074 27918 28086 27970
rect 28138 27918 28150 27970
rect 29194 27918 29206 27970
rect 29258 27918 29270 27970
rect 12686 27897 12738 27909
rect 16718 27906 16770 27918
rect 8094 27858 8146 27870
rect 8094 27794 8146 27806
rect 11454 27858 11506 27870
rect 12226 27806 12238 27858
rect 12290 27806 12302 27858
rect 12686 27833 12738 27845
rect 12910 27858 12962 27870
rect 11454 27794 11506 27806
rect 12910 27794 12962 27806
rect 14030 27858 14082 27870
rect 14030 27794 14082 27806
rect 21198 27858 21250 27870
rect 21198 27794 21250 27806
rect 23774 27858 23826 27870
rect 23774 27794 23826 27806
rect 23886 27858 23938 27870
rect 25498 27862 25510 27914
rect 25562 27862 25574 27914
rect 27246 27897 27298 27909
rect 25218 27806 25230 27858
rect 25282 27806 25294 27858
rect 26786 27806 26798 27858
rect 26850 27806 26862 27858
rect 27246 27833 27298 27845
rect 27470 27858 27522 27870
rect 23886 27794 23938 27806
rect 27470 27794 27522 27806
rect 28366 27858 28418 27870
rect 28366 27794 28418 27806
rect 28478 27858 28530 27870
rect 28478 27794 28530 27806
rect 28702 27858 28754 27870
rect 28702 27794 28754 27806
rect 28926 27858 28978 27870
rect 28926 27794 28978 27806
rect 14802 27694 14814 27746
rect 14866 27694 14878 27746
rect 25666 27694 25678 27746
rect 25730 27694 25742 27746
rect 8430 27634 8482 27646
rect 8430 27570 8482 27582
rect 21534 27634 21586 27646
rect 23482 27582 23494 27634
rect 23546 27582 23558 27634
rect 21534 27570 21586 27582
rect 1344 27466 34608 27500
rect 1344 27414 5372 27466
rect 5424 27414 5476 27466
rect 5528 27414 5580 27466
rect 5632 27414 13688 27466
rect 13740 27414 13792 27466
rect 13844 27414 13896 27466
rect 13948 27414 22004 27466
rect 22056 27414 22108 27466
rect 22160 27414 22212 27466
rect 22264 27414 30320 27466
rect 30372 27414 30424 27466
rect 30476 27414 30528 27466
rect 30580 27414 34608 27466
rect 1344 27380 34608 27414
rect 14478 27242 14530 27254
rect 8306 27134 8318 27186
rect 8370 27134 8382 27186
rect 14478 27178 14530 27190
rect 14802 27134 14814 27186
rect 14866 27134 14878 27186
rect 17602 27134 17614 27186
rect 17666 27134 17678 27186
rect 21970 27134 21982 27186
rect 22034 27134 22046 27186
rect 23874 27134 23886 27186
rect 23938 27134 23950 27186
rect 27794 27134 27806 27186
rect 27858 27134 27870 27186
rect 7310 27074 7362 27086
rect 7310 27010 7362 27022
rect 7534 27074 7586 27086
rect 16718 27074 16770 27086
rect 14018 27022 14030 27074
rect 14082 27022 14094 27074
rect 14354 27022 14366 27074
rect 14418 27022 14430 27074
rect 7534 27010 7586 27022
rect 14914 27007 14926 27059
rect 14978 27007 14990 27059
rect 15250 27022 15262 27074
rect 15314 27022 15326 27074
rect 16718 27010 16770 27022
rect 16942 27074 16994 27086
rect 20190 27074 20242 27086
rect 17154 27022 17166 27074
rect 17218 27022 17230 27074
rect 16942 27010 16994 27022
rect 17490 27007 17502 27059
rect 17554 27007 17566 27059
rect 20190 27010 20242 27022
rect 20414 27074 20466 27086
rect 20414 27010 20466 27022
rect 21198 27074 21250 27086
rect 21198 27010 21250 27022
rect 25118 27074 25170 27086
rect 25890 27022 25902 27074
rect 25954 27022 25966 27074
rect 25118 27010 25170 27022
rect 6974 26962 7026 26974
rect 6974 26898 7026 26910
rect 10222 26962 10274 26974
rect 16426 26910 16438 26962
rect 16490 26910 16502 26962
rect 20682 26910 20694 26962
rect 20746 26910 20758 26962
rect 10222 26898 10274 26910
rect 5798 26850 5850 26862
rect 5798 26786 5850 26798
rect 10838 26850 10890 26862
rect 10838 26786 10890 26798
rect 1344 26682 34768 26716
rect 1344 26630 9530 26682
rect 9582 26630 9634 26682
rect 9686 26630 9738 26682
rect 9790 26630 17846 26682
rect 17898 26630 17950 26682
rect 18002 26630 18054 26682
rect 18106 26630 26162 26682
rect 26214 26630 26266 26682
rect 26318 26630 26370 26682
rect 26422 26630 34478 26682
rect 34530 26630 34582 26682
rect 34634 26630 34686 26682
rect 34738 26630 34768 26682
rect 1344 26596 34768 26630
rect 23214 26514 23266 26526
rect 23214 26450 23266 26462
rect 26574 26514 26626 26526
rect 26574 26450 26626 26462
rect 21242 26350 21254 26402
rect 21306 26350 21318 26402
rect 2270 26290 2322 26302
rect 2270 26226 2322 26238
rect 5294 26290 5346 26302
rect 8766 26290 8818 26302
rect 6066 26238 6078 26290
rect 6130 26238 6142 26290
rect 5294 26226 5346 26238
rect 8766 26226 8818 26238
rect 8878 26290 8930 26302
rect 9650 26253 9662 26305
rect 9714 26253 9726 26305
rect 11566 26290 11618 26302
rect 9986 26238 9998 26290
rect 10050 26238 10062 26290
rect 8878 26226 8930 26238
rect 11566 26226 11618 26238
rect 12574 26290 12626 26302
rect 12574 26226 12626 26238
rect 12686 26290 12738 26302
rect 12686 26226 12738 26238
rect 17278 26290 17330 26302
rect 17278 26226 17330 26238
rect 20862 26290 20914 26302
rect 20862 26226 20914 26238
rect 20974 26290 21026 26302
rect 20974 26226 21026 26238
rect 22878 26290 22930 26302
rect 23874 26253 23886 26305
rect 23938 26253 23950 26305
rect 26910 26290 26962 26302
rect 24098 26238 24110 26290
rect 24162 26238 24174 26290
rect 27570 26253 27582 26305
rect 27634 26253 27646 26305
rect 27794 26238 27806 26290
rect 27858 26238 27870 26290
rect 28578 26282 28590 26334
rect 28642 26282 28654 26334
rect 29262 26290 29314 26302
rect 28914 26238 28926 26290
rect 28978 26238 28990 26290
rect 22878 26226 22930 26238
rect 26910 26226 26962 26238
rect 29262 26226 29314 26238
rect 29374 26290 29426 26302
rect 29374 26226 29426 26238
rect 10502 26178 10554 26190
rect 3042 26126 3054 26178
rect 3106 26126 3118 26178
rect 4946 26126 4958 26178
rect 5010 26126 5022 26178
rect 7970 26126 7982 26178
rect 8034 26126 8046 26178
rect 9538 26126 9550 26178
rect 9602 26126 9614 26178
rect 10502 26114 10554 26126
rect 11958 26178 12010 26190
rect 11958 26114 12010 26126
rect 13190 26178 13242 26190
rect 13190 26114 13242 26126
rect 15990 26178 16042 26190
rect 15990 26114 16042 26126
rect 16438 26178 16490 26190
rect 18050 26126 18062 26178
rect 18114 26126 18126 26178
rect 19954 26126 19966 26178
rect 20018 26126 20030 26178
rect 23762 26126 23774 26178
rect 23826 26126 23838 26178
rect 27458 26126 27470 26178
rect 27522 26126 27534 26178
rect 28466 26126 28478 26178
rect 28530 26126 28542 26178
rect 16438 26114 16490 26126
rect 11230 26066 11282 26078
rect 8474 26014 8486 26066
rect 8538 26014 8550 26066
rect 12282 26014 12294 26066
rect 12346 26014 12358 26066
rect 29642 26014 29654 26066
rect 29706 26014 29718 26066
rect 11230 26002 11282 26014
rect 1344 25898 34608 25932
rect 1344 25846 5372 25898
rect 5424 25846 5476 25898
rect 5528 25846 5580 25898
rect 5632 25846 13688 25898
rect 13740 25846 13792 25898
rect 13844 25846 13896 25898
rect 13948 25846 22004 25898
rect 22056 25846 22108 25898
rect 22160 25846 22212 25898
rect 22264 25846 30320 25898
rect 30372 25846 30424 25898
rect 30476 25846 30528 25898
rect 30580 25846 34608 25898
rect 1344 25812 34608 25846
rect 4846 25730 4898 25742
rect 4846 25666 4898 25678
rect 7814 25730 7866 25742
rect 7814 25666 7866 25678
rect 17502 25730 17554 25742
rect 17502 25666 17554 25678
rect 5798 25618 5850 25630
rect 15598 25618 15650 25630
rect 19170 25622 19182 25674
rect 19234 25622 19246 25674
rect 10882 25566 10894 25618
rect 10946 25566 10958 25618
rect 12786 25566 12798 25618
rect 12850 25566 12862 25618
rect 5798 25554 5850 25566
rect 15598 25554 15650 25566
rect 20414 25618 20466 25630
rect 28130 25566 28142 25618
rect 28194 25566 28206 25618
rect 20414 25554 20466 25566
rect 1598 25506 1650 25518
rect 5182 25506 5234 25518
rect 2370 25454 2382 25506
rect 2434 25454 2446 25506
rect 1598 25442 1650 25454
rect 5182 25442 5234 25454
rect 6526 25506 6578 25518
rect 6526 25442 6578 25454
rect 6750 25506 6802 25518
rect 6750 25442 6802 25454
rect 7310 25506 7362 25518
rect 7310 25442 7362 25454
rect 7422 25506 7474 25518
rect 7422 25442 7474 25454
rect 8094 25506 8146 25518
rect 8094 25442 8146 25454
rect 8542 25506 8594 25518
rect 10110 25506 10162 25518
rect 14478 25506 14530 25518
rect 8754 25454 8766 25506
rect 8818 25454 8830 25506
rect 13346 25454 13358 25506
rect 13410 25454 13422 25506
rect 4286 25394 4338 25406
rect 8206 25394 8258 25406
rect 8362 25398 8374 25450
rect 8426 25398 8438 25450
rect 8542 25442 8594 25454
rect 10110 25442 10162 25454
rect 14478 25442 14530 25454
rect 14590 25506 14642 25518
rect 14590 25442 14642 25454
rect 15262 25506 15314 25518
rect 16886 25506 16938 25518
rect 16158 25478 16210 25490
rect 15262 25442 15314 25454
rect 16046 25450 16098 25462
rect 16158 25414 16210 25426
rect 16370 25398 16382 25450
rect 16434 25398 16446 25450
rect 16594 25398 16606 25450
rect 16658 25398 16670 25450
rect 16886 25442 16938 25454
rect 17166 25506 17218 25518
rect 23998 25506 24050 25518
rect 18946 25454 18958 25506
rect 19010 25454 19022 25506
rect 19282 25454 19294 25506
rect 19346 25454 19358 25506
rect 19854 25468 19906 25480
rect 17166 25442 17218 25454
rect 19742 25450 19794 25462
rect 19854 25404 19906 25416
rect 20582 25450 20634 25462
rect 6234 25342 6246 25394
rect 6298 25342 6310 25394
rect 7018 25342 7030 25394
rect 7082 25342 7094 25394
rect 16046 25386 16098 25398
rect 19742 25386 19794 25398
rect 23998 25442 24050 25454
rect 24110 25506 24162 25518
rect 24110 25442 24162 25454
rect 24446 25506 24498 25518
rect 24446 25442 24498 25454
rect 24558 25506 24610 25518
rect 24558 25442 24610 25454
rect 27358 25506 27410 25518
rect 27358 25442 27410 25454
rect 27694 25506 27746 25518
rect 31950 25506 32002 25518
rect 28354 25454 28366 25506
rect 28418 25454 28430 25506
rect 31154 25454 31166 25506
rect 31218 25454 31230 25506
rect 27694 25442 27746 25454
rect 28018 25398 28030 25450
rect 28082 25398 28094 25450
rect 31950 25442 32002 25454
rect 32342 25506 32394 25518
rect 32342 25442 32394 25454
rect 20582 25386 20634 25398
rect 29262 25394 29314 25406
rect 4286 25330 4338 25342
rect 8206 25330 8258 25342
rect 13526 25338 13578 25350
rect 23706 25342 23718 25394
rect 23770 25342 23782 25394
rect 24826 25342 24838 25394
rect 24890 25342 24902 25394
rect 9830 25282 9882 25294
rect 29262 25330 29314 25342
rect 13526 25274 13578 25286
rect 14142 25282 14194 25294
rect 9830 25218 9882 25230
rect 14142 25218 14194 25230
rect 14926 25282 14978 25294
rect 14926 25218 14978 25230
rect 23382 25282 23434 25294
rect 23382 25218 23434 25230
rect 1344 25114 34768 25148
rect 1344 25062 9530 25114
rect 9582 25062 9634 25114
rect 9686 25062 9738 25114
rect 9790 25062 17846 25114
rect 17898 25062 17950 25114
rect 18002 25062 18054 25114
rect 18106 25062 26162 25114
rect 26214 25062 26266 25114
rect 26318 25062 26370 25114
rect 26422 25062 34478 25114
rect 34530 25062 34582 25114
rect 34634 25062 34686 25114
rect 34738 25062 34768 25114
rect 1344 25028 34768 25062
rect 2718 24946 2770 24958
rect 2718 24882 2770 24894
rect 17614 24946 17666 24958
rect 17614 24882 17666 24894
rect 29710 24946 29762 24958
rect 19070 24834 19122 24846
rect 24434 24838 24446 24890
rect 24498 24838 24510 24890
rect 29026 24838 29038 24890
rect 29090 24838 29102 24890
rect 29710 24882 29762 24894
rect 12730 24782 12742 24834
rect 12794 24782 12806 24834
rect 16090 24782 16102 24834
rect 16154 24782 16166 24834
rect 27850 24782 27862 24834
rect 27914 24782 27926 24834
rect 3054 24722 3106 24734
rect 3054 24658 3106 24670
rect 4398 24722 4450 24734
rect 4398 24658 4450 24670
rect 4510 24722 4562 24734
rect 4510 24658 4562 24670
rect 5182 24722 5234 24734
rect 5182 24658 5234 24670
rect 5294 24722 5346 24734
rect 5294 24658 5346 24670
rect 6638 24722 6690 24734
rect 6638 24658 6690 24670
rect 6862 24722 6914 24734
rect 6862 24658 6914 24670
rect 7534 24722 7586 24734
rect 7690 24726 7702 24778
rect 7754 24726 7766 24778
rect 19070 24770 19122 24782
rect 7982 24722 8034 24734
rect 7858 24670 7870 24722
rect 7922 24670 7934 24722
rect 7534 24658 7586 24670
rect 7982 24658 8034 24670
rect 8262 24722 8314 24734
rect 11890 24697 11902 24749
rect 11954 24697 11966 24749
rect 12238 24722 12290 24734
rect 8262 24658 8314 24670
rect 12238 24658 12290 24670
rect 12462 24722 12514 24734
rect 13234 24697 13246 24749
rect 13298 24697 13310 24749
rect 16382 24722 16434 24734
rect 12462 24658 12514 24670
rect 16382 24658 16434 24670
rect 16494 24722 16546 24734
rect 16494 24658 16546 24670
rect 17278 24722 17330 24734
rect 21758 24722 21810 24734
rect 18386 24670 18398 24722
rect 18450 24670 18462 24722
rect 20962 24670 20974 24722
rect 21026 24670 21038 24722
rect 22082 24670 22094 24722
rect 22146 24670 22158 24722
rect 22418 24670 22430 24722
rect 22482 24670 22494 24722
rect 22978 24714 22990 24766
rect 23042 24714 23054 24766
rect 23314 24670 23326 24722
rect 23378 24670 23390 24722
rect 23650 24670 23662 24722
rect 23714 24670 23726 24722
rect 23986 24697 23998 24749
rect 24050 24697 24062 24749
rect 24334 24722 24386 24734
rect 17278 24658 17330 24670
rect 21758 24658 21810 24670
rect 24334 24658 24386 24670
rect 25118 24722 25170 24734
rect 25118 24658 25170 24670
rect 27358 24722 27410 24734
rect 27358 24658 27410 24670
rect 27582 24722 27634 24734
rect 28578 24726 28590 24778
rect 28642 24726 28654 24778
rect 28926 24722 28978 24734
rect 28242 24670 28254 24722
rect 28306 24670 28318 24722
rect 27582 24658 27634 24670
rect 28926 24658 28978 24670
rect 29374 24722 29426 24734
rect 29374 24658 29426 24670
rect 26742 24610 26794 24622
rect 21982 24554 22034 24566
rect 22866 24558 22878 24610
rect 22930 24558 22942 24610
rect 10334 24498 10386 24510
rect 4106 24446 4118 24498
rect 4170 24446 4182 24498
rect 4890 24446 4902 24498
rect 4954 24446 4966 24498
rect 7130 24446 7142 24498
rect 7194 24446 7206 24498
rect 10334 24434 10386 24446
rect 14254 24498 14306 24510
rect 14254 24434 14306 24446
rect 18566 24498 18618 24510
rect 26742 24546 26794 24558
rect 27190 24610 27242 24622
rect 27190 24546 27242 24558
rect 21982 24490 22034 24502
rect 25454 24498 25506 24510
rect 18566 24434 18618 24446
rect 25454 24434 25506 24446
rect 1344 24330 34608 24364
rect 1344 24278 5372 24330
rect 5424 24278 5476 24330
rect 5528 24278 5580 24330
rect 5632 24278 13688 24330
rect 13740 24278 13792 24330
rect 13844 24278 13896 24330
rect 13948 24278 22004 24330
rect 22056 24278 22108 24330
rect 22160 24278 22212 24330
rect 22264 24278 30320 24330
rect 30372 24278 30424 24330
rect 30476 24278 30528 24330
rect 30580 24278 34608 24330
rect 1344 24244 34608 24278
rect 4342 24162 4394 24174
rect 4342 24098 4394 24110
rect 6582 24162 6634 24174
rect 6582 24098 6634 24110
rect 12798 24162 12850 24174
rect 20694 24162 20746 24174
rect 16314 24110 16326 24162
rect 16378 24110 16390 24162
rect 12798 24098 12850 24110
rect 20694 24098 20746 24110
rect 11678 24050 11730 24062
rect 4902 23994 4954 24006
rect 3838 23938 3890 23950
rect 3838 23874 3890 23886
rect 3950 23938 4002 23950
rect 3950 23874 4002 23886
rect 4622 23938 4674 23950
rect 7142 23994 7194 24006
rect 4902 23930 4954 23942
rect 5070 23938 5122 23950
rect 6078 23938 6130 23950
rect 4622 23874 4674 23886
rect 5786 23886 5798 23938
rect 5850 23886 5862 23938
rect 5070 23874 5122 23886
rect 6078 23874 6130 23886
rect 6302 23938 6354 23950
rect 6302 23874 6354 23886
rect 6862 23938 6914 23950
rect 7142 23930 7194 23942
rect 7310 23938 7362 23950
rect 6862 23874 6914 23886
rect 7310 23874 7362 23886
rect 7870 23938 7922 23950
rect 9326 23938 9378 23950
rect 7870 23874 7922 23886
rect 8194 23859 8206 23911
rect 8258 23859 8270 23911
rect 8530 23886 8542 23938
rect 8594 23886 8606 23938
rect 9326 23874 9378 23886
rect 9550 23938 9602 23950
rect 10110 23938 10162 23950
rect 9818 23886 9830 23938
rect 9882 23886 9894 23938
rect 9550 23874 9602 23886
rect 10110 23874 10162 23886
rect 10222 23938 10274 23950
rect 10994 23942 11006 23994
rect 11058 23942 11070 23994
rect 11678 23986 11730 23998
rect 11846 23994 11898 24006
rect 18790 23994 18842 24006
rect 20134 23994 20186 24006
rect 24322 23998 24334 24050
rect 24386 23998 24398 24050
rect 26226 23998 26238 24050
rect 26290 23998 26302 24050
rect 11846 23930 11898 23942
rect 12126 23938 12178 23950
rect 12404 23938 12456 23950
rect 10222 23874 10274 23886
rect 11218 23858 11230 23910
rect 11282 23858 11294 23910
rect 12226 23886 12238 23938
rect 12290 23886 12302 23938
rect 16606 23938 16658 23950
rect 12126 23874 12178 23886
rect 12404 23874 12456 23886
rect 13794 23858 13806 23910
rect 13858 23858 13870 23910
rect 16606 23874 16658 23886
rect 16718 23938 16770 23950
rect 16718 23874 16770 23886
rect 16942 23938 16994 23950
rect 16942 23874 16994 23886
rect 18174 23938 18226 23950
rect 19618 23942 19630 23994
rect 19682 23942 19694 23994
rect 18790 23930 18842 23942
rect 19966 23938 20018 23950
rect 18174 23874 18226 23886
rect 19518 23900 19570 23912
rect 20134 23930 20186 23942
rect 20414 23938 20466 23950
rect 19966 23874 20018 23886
rect 20414 23874 20466 23886
rect 22654 23938 22706 23950
rect 22654 23874 22706 23886
rect 23550 23938 23602 23950
rect 28366 23938 28418 23950
rect 23550 23874 23602 23886
rect 27010 23871 27022 23923
rect 27074 23871 27086 23923
rect 27234 23886 27246 23938
rect 27298 23886 27310 23938
rect 27682 23886 27694 23938
rect 27746 23886 27758 23938
rect 4734 23826 4786 23838
rect 3546 23774 3558 23826
rect 3610 23774 3622 23826
rect 4734 23762 4786 23774
rect 6974 23826 7026 23838
rect 17838 23826 17890 23838
rect 6974 23762 7026 23774
rect 8206 23770 8258 23782
rect 9034 23774 9046 23826
rect 9098 23774 9110 23826
rect 17838 23762 17890 23774
rect 18958 23826 19010 23838
rect 19518 23836 19570 23848
rect 18958 23762 19010 23774
rect 20302 23826 20354 23838
rect 27962 23830 27974 23882
rect 28026 23830 28038 23882
rect 28366 23874 28418 23886
rect 29038 23938 29090 23950
rect 29038 23874 29090 23886
rect 20302 23762 20354 23774
rect 8206 23706 8258 23718
rect 17278 23714 17330 23726
rect 17278 23650 17330 23662
rect 22990 23714 23042 23726
rect 27234 23718 27246 23770
rect 27298 23718 27310 23770
rect 28466 23718 28478 23770
rect 28530 23718 28542 23770
rect 22990 23650 23042 23662
rect 29374 23714 29426 23726
rect 29374 23650 29426 23662
rect 1344 23546 34768 23580
rect 1344 23494 9530 23546
rect 9582 23494 9634 23546
rect 9686 23494 9738 23546
rect 9790 23494 17846 23546
rect 17898 23494 17950 23546
rect 18002 23494 18054 23546
rect 18106 23494 26162 23546
rect 26214 23494 26266 23546
rect 26318 23494 26370 23546
rect 26422 23494 34478 23546
rect 34530 23494 34582 23546
rect 34634 23494 34686 23546
rect 34738 23494 34768 23546
rect 1344 23460 34768 23494
rect 20134 23378 20186 23390
rect 20134 23314 20186 23326
rect 20638 23378 20690 23390
rect 20638 23314 20690 23326
rect 26182 23378 26234 23390
rect 26182 23314 26234 23326
rect 29878 23378 29930 23390
rect 29878 23314 29930 23326
rect 4286 23266 4338 23278
rect 4286 23202 4338 23214
rect 8318 23266 8370 23278
rect 1598 23154 1650 23166
rect 1598 23090 1650 23102
rect 4734 23154 4786 23166
rect 5598 23158 5610 23210
rect 5662 23158 5674 23210
rect 8318 23202 8370 23214
rect 10110 23266 10162 23278
rect 10110 23202 10162 23214
rect 13358 23266 13410 23278
rect 13358 23202 13410 23214
rect 26798 23266 26850 23278
rect 6290 23102 6302 23154
rect 6354 23102 6366 23154
rect 6626 23146 6638 23198
rect 6690 23146 6702 23198
rect 18510 23192 18562 23204
rect 26798 23202 26850 23214
rect 8206 23154 8258 23166
rect 8654 23154 8706 23166
rect 4734 23090 4786 23102
rect 8206 23090 8258 23102
rect 8486 23098 8538 23110
rect 8654 23090 8706 23102
rect 12798 23154 12850 23166
rect 12798 23090 12850 23102
rect 13022 23154 13074 23166
rect 13470 23154 13522 23166
rect 13022 23090 13074 23102
rect 13190 23098 13242 23110
rect 2370 22990 2382 23042
rect 2434 22990 2446 23042
rect 6738 22990 6750 23042
rect 6802 22990 6814 23042
rect 8486 23034 8538 23046
rect 13470 23090 13522 23102
rect 14030 23154 14082 23166
rect 14802 23102 14814 23154
rect 14866 23102 14878 23154
rect 14030 23090 14082 23102
rect 17782 23098 17834 23110
rect 18162 23102 18174 23154
rect 18226 23102 18238 23154
rect 20302 23154 20354 23166
rect 18510 23128 18562 23140
rect 19282 23102 19294 23154
rect 19346 23102 19358 23154
rect 19618 23102 19630 23154
rect 19682 23102 19694 23154
rect 22194 23129 22206 23181
rect 22258 23129 22270 23181
rect 25566 23154 25618 23166
rect 12002 22990 12014 23042
rect 12066 22990 12078 23042
rect 13190 23034 13242 23046
rect 20302 23090 20354 23102
rect 25566 23090 25618 23102
rect 25790 23154 25842 23166
rect 29486 23154 29538 23166
rect 28690 23102 28702 23154
rect 28754 23102 28766 23154
rect 25790 23090 25842 23102
rect 29486 23090 29538 23102
rect 30942 23154 30994 23166
rect 30942 23090 30994 23102
rect 16706 22990 16718 23042
rect 16770 22990 16782 23042
rect 17782 23034 17834 23046
rect 17950 23042 18002 23054
rect 21926 23042 21978 23054
rect 17950 22978 18002 22990
rect 19182 22986 19234 22998
rect 5854 22930 5906 22942
rect 5854 22866 5906 22878
rect 7926 22930 7978 22942
rect 7926 22866 7978 22878
rect 13750 22930 13802 22942
rect 21926 22978 21978 22990
rect 19182 22922 19234 22934
rect 23214 22930 23266 22942
rect 30606 22930 30658 22942
rect 13750 22866 13802 22878
rect 25274 22878 25286 22930
rect 25338 22878 25350 22930
rect 23214 22866 23266 22878
rect 30606 22866 30658 22878
rect 1344 22762 34608 22796
rect 1344 22710 5372 22762
rect 5424 22710 5476 22762
rect 5528 22710 5580 22762
rect 5632 22710 13688 22762
rect 13740 22710 13792 22762
rect 13844 22710 13896 22762
rect 13948 22710 22004 22762
rect 22056 22710 22108 22762
rect 22160 22710 22212 22762
rect 22264 22710 30320 22762
rect 30372 22710 30424 22762
rect 30476 22710 30528 22762
rect 30580 22710 34608 22762
rect 1344 22676 34608 22710
rect 2718 22594 2770 22606
rect 2718 22530 2770 22542
rect 9886 22594 9938 22606
rect 9886 22530 9938 22542
rect 12070 22594 12122 22606
rect 12070 22530 12122 22542
rect 14366 22594 14418 22606
rect 14366 22530 14418 22542
rect 22878 22538 22930 22550
rect 5014 22482 5066 22494
rect 5014 22418 5066 22430
rect 9270 22482 9322 22494
rect 9270 22418 9322 22430
rect 12798 22482 12850 22494
rect 12798 22418 12850 22430
rect 18510 22482 18562 22494
rect 22878 22474 22930 22486
rect 32118 22482 32170 22494
rect 18510 22418 18562 22430
rect 32118 22418 32170 22430
rect 3054 22370 3106 22382
rect 3054 22306 3106 22318
rect 3726 22370 3778 22382
rect 4174 22370 4226 22382
rect 4050 22318 4062 22370
rect 4114 22318 4126 22370
rect 3726 22306 3778 22318
rect 3882 22262 3894 22314
rect 3946 22262 3958 22314
rect 4174 22306 4226 22318
rect 4454 22370 4506 22382
rect 8094 22370 8146 22382
rect 4454 22306 4506 22318
rect 7534 22332 7586 22344
rect 7858 22318 7870 22370
rect 7922 22318 7934 22370
rect 8542 22370 8594 22382
rect 8094 22306 8146 22318
rect 8262 22314 8314 22326
rect 7534 22268 7586 22280
rect 8542 22306 8594 22318
rect 8710 22370 8762 22382
rect 8710 22306 8762 22318
rect 8990 22370 9042 22382
rect 8990 22306 9042 22318
rect 9550 22370 9602 22382
rect 12462 22370 12514 22382
rect 9550 22306 9602 22318
rect 11162 22302 11174 22354
rect 11226 22302 11238 22354
rect 11398 22335 11450 22347
rect 11398 22271 11450 22283
rect 8262 22250 8314 22262
rect 8878 22258 8930 22270
rect 11554 22262 11566 22314
rect 11618 22262 11630 22314
rect 11778 22262 11790 22314
rect 11842 22262 11854 22314
rect 12462 22306 12514 22318
rect 13806 22370 13858 22382
rect 13806 22306 13858 22318
rect 14030 22370 14082 22382
rect 14030 22306 14082 22318
rect 14702 22370 14754 22382
rect 17838 22370 17890 22382
rect 19182 22370 19234 22382
rect 23102 22370 23154 22382
rect 17154 22318 17166 22370
rect 17218 22318 17230 22370
rect 17614 22331 17666 22343
rect 14702 22306 14754 22318
rect 19058 22318 19070 22370
rect 19122 22318 19134 22370
rect 22418 22318 22430 22370
rect 22482 22318 22494 22370
rect 22754 22318 22766 22370
rect 22818 22318 22830 22370
rect 23874 22318 23886 22370
rect 23938 22318 23950 22370
rect 17838 22306 17890 22318
rect 17614 22267 17666 22279
rect 18892 22262 18904 22314
rect 18956 22262 18968 22314
rect 19182 22306 19234 22318
rect 23102 22306 23154 22318
rect 29474 22290 29486 22342
rect 29538 22290 29550 22342
rect 25790 22258 25842 22270
rect 13514 22206 13526 22258
rect 13578 22206 13590 22258
rect 8878 22194 8930 22206
rect 10950 22146 11002 22158
rect 10950 22082 11002 22094
rect 15990 22146 16042 22158
rect 17266 22150 17278 22202
rect 17330 22150 17342 22202
rect 25790 22194 25842 22206
rect 15990 22082 16042 22094
rect 1344 21978 34768 22012
rect 1344 21926 9530 21978
rect 9582 21926 9634 21978
rect 9686 21926 9738 21978
rect 9790 21926 17846 21978
rect 17898 21926 17950 21978
rect 18002 21926 18054 21978
rect 18106 21926 26162 21978
rect 26214 21926 26266 21978
rect 26318 21926 26370 21978
rect 26422 21926 34478 21978
rect 34530 21926 34582 21978
rect 34634 21926 34686 21978
rect 34738 21926 34768 21978
rect 1344 21892 34768 21926
rect 11790 21810 11842 21822
rect 11790 21746 11842 21758
rect 18062 21810 18114 21822
rect 18062 21746 18114 21758
rect 18566 21810 18618 21822
rect 18566 21746 18618 21758
rect 21870 21810 21922 21822
rect 21870 21746 21922 21758
rect 23326 21698 23378 21710
rect 4218 21646 4230 21698
rect 4282 21646 4294 21698
rect 23158 21642 23210 21654
rect 4510 21586 4562 21598
rect 4510 21522 4562 21534
rect 4734 21586 4786 21598
rect 8318 21586 8370 21598
rect 4834 21534 4846 21586
rect 4898 21534 4910 21586
rect 4734 21522 4786 21534
rect 8318 21522 8370 21534
rect 8654 21586 8706 21598
rect 8654 21522 8706 21534
rect 12126 21586 12178 21598
rect 17726 21586 17778 21598
rect 21422 21586 21474 21598
rect 13122 21534 13134 21586
rect 13186 21534 13198 21586
rect 18722 21534 18734 21586
rect 18786 21534 18798 21586
rect 12126 21522 12178 21534
rect 17726 21522 17778 21534
rect 21422 21522 21474 21534
rect 21534 21586 21586 21598
rect 23326 21634 23378 21646
rect 33238 21698 33290 21710
rect 33238 21634 33290 21646
rect 23158 21578 23210 21590
rect 23538 21534 23550 21586
rect 23602 21534 23614 21586
rect 23762 21562 23774 21614
rect 23826 21562 23838 21614
rect 29374 21586 29426 21598
rect 21534 21522 21586 21534
rect 29374 21522 29426 21534
rect 29486 21586 29538 21598
rect 29486 21522 29538 21534
rect 32622 21586 32674 21598
rect 32622 21522 32674 21534
rect 9046 21474 9098 21486
rect 9046 21410 9098 21422
rect 22934 21474 22986 21486
rect 29922 21422 29934 21474
rect 29986 21422 29998 21474
rect 31826 21422 31838 21474
rect 31890 21422 31902 21474
rect 22934 21410 22986 21422
rect 5014 21362 5066 21374
rect 5014 21298 5066 21310
rect 13302 21362 13354 21374
rect 13302 21298 13354 21310
rect 21086 21362 21138 21374
rect 29082 21310 29094 21362
rect 29146 21310 29158 21362
rect 21086 21298 21138 21310
rect 1344 21194 34608 21228
rect 1344 21142 5372 21194
rect 5424 21142 5476 21194
rect 5528 21142 5580 21194
rect 5632 21142 13688 21194
rect 13740 21142 13792 21194
rect 13844 21142 13896 21194
rect 13948 21142 22004 21194
rect 22056 21142 22108 21194
rect 22160 21142 22212 21194
rect 22264 21142 30320 21194
rect 30372 21142 30424 21194
rect 30476 21142 30528 21194
rect 30580 21142 34608 21194
rect 1344 21108 34608 21142
rect 6358 21026 6410 21038
rect 6358 20962 6410 20974
rect 7646 20970 7698 20982
rect 32330 20974 32342 21026
rect 32394 20974 32406 21026
rect 3658 20862 3670 20914
rect 3722 20862 3734 20914
rect 7646 20906 7698 20918
rect 12674 20862 12686 20914
rect 12738 20862 12750 20914
rect 15026 20862 15038 20914
rect 15090 20862 15102 20914
rect 3950 20802 4002 20814
rect 3950 20738 4002 20750
rect 4062 20802 4114 20814
rect 4062 20738 4114 20750
rect 5630 20802 5682 20814
rect 6078 20802 6130 20814
rect 11790 20802 11842 20814
rect 5954 20750 5966 20802
rect 6018 20750 6030 20802
rect 7186 20750 7198 20802
rect 7250 20750 7262 20802
rect 7522 20750 7534 20802
rect 7586 20750 7598 20802
rect 5630 20738 5682 20750
rect 5786 20694 5798 20746
rect 5850 20694 5862 20746
rect 6078 20738 6130 20750
rect 11790 20738 11842 20750
rect 12014 20802 12066 20814
rect 20078 20802 20130 20814
rect 12226 20750 12238 20802
rect 12290 20750 12302 20802
rect 14018 20750 14030 20802
rect 14082 20750 14094 20802
rect 14422 20772 14474 20784
rect 12014 20738 12066 20750
rect 12506 20694 12518 20746
rect 12570 20694 12582 20746
rect 14422 20708 14474 20720
rect 15138 20706 15150 20758
rect 15202 20706 15214 20758
rect 15474 20750 15486 20802
rect 15538 20750 15550 20802
rect 16146 20750 16158 20802
rect 16210 20750 16222 20802
rect 20078 20738 20130 20750
rect 20302 20802 20354 20814
rect 20302 20738 20354 20750
rect 20414 20802 20466 20814
rect 20414 20738 20466 20750
rect 21366 20802 21418 20814
rect 21366 20738 21418 20750
rect 21646 20802 21698 20814
rect 22094 20802 22146 20814
rect 21746 20750 21758 20802
rect 21810 20750 21822 20802
rect 21646 20738 21698 20750
rect 21914 20694 21926 20746
rect 21978 20694 21990 20746
rect 22094 20738 22146 20750
rect 22430 20802 22482 20814
rect 22430 20738 22482 20750
rect 22598 20802 22650 20814
rect 22598 20738 22650 20750
rect 22878 20802 22930 20814
rect 22878 20738 22930 20750
rect 23438 20802 23490 20814
rect 26126 20802 26178 20814
rect 24210 20750 24222 20802
rect 24274 20750 24286 20802
rect 23438 20738 23490 20750
rect 26126 20738 26178 20750
rect 26462 20802 26514 20814
rect 26462 20738 26514 20750
rect 26686 20802 26738 20814
rect 26686 20738 26738 20750
rect 27750 20802 27802 20814
rect 27750 20738 27802 20750
rect 28478 20802 28530 20814
rect 31838 20802 31890 20814
rect 28478 20738 28530 20750
rect 29138 20722 29150 20774
rect 29202 20722 29214 20774
rect 31378 20750 31390 20802
rect 31442 20750 31454 20802
rect 31838 20738 31890 20750
rect 32062 20802 32114 20814
rect 32062 20738 32114 20750
rect 22766 20690 22818 20702
rect 11498 20638 11510 20690
rect 11562 20638 11574 20690
rect 14366 20634 14418 20646
rect 20682 20638 20694 20690
rect 20746 20638 20758 20690
rect 22766 20626 22818 20638
rect 23158 20690 23210 20702
rect 26954 20638 26966 20690
rect 27018 20638 27030 20690
rect 23158 20626 23210 20638
rect 14366 20570 14418 20582
rect 15990 20578 16042 20590
rect 15990 20514 16042 20526
rect 19742 20578 19794 20590
rect 19742 20514 19794 20526
rect 28142 20578 28194 20590
rect 28142 20514 28194 20526
rect 1344 20410 34768 20444
rect 1344 20358 9530 20410
rect 9582 20358 9634 20410
rect 9686 20358 9738 20410
rect 9790 20358 17846 20410
rect 17898 20358 17950 20410
rect 18002 20358 18054 20410
rect 18106 20358 26162 20410
rect 26214 20358 26266 20410
rect 26318 20358 26370 20410
rect 26422 20358 34478 20410
rect 34530 20358 34582 20410
rect 34634 20358 34686 20410
rect 34738 20358 34768 20410
rect 1344 20324 34768 20358
rect 23886 20242 23938 20254
rect 23886 20178 23938 20190
rect 30830 20130 30882 20142
rect 4442 20078 4454 20130
rect 4506 20078 4518 20130
rect 12518 20074 12570 20086
rect 22362 20078 22374 20130
rect 22426 20078 22438 20130
rect 3054 20018 3106 20030
rect 3726 20018 3778 20030
rect 3054 19954 3106 19966
rect 3222 19962 3274 19974
rect 3726 19954 3778 19966
rect 3968 20018 4020 20030
rect 3968 19954 4020 19966
rect 4734 20018 4786 20030
rect 4734 19954 4786 19966
rect 4846 20018 4898 20030
rect 5506 20022 5518 20074
rect 5570 20022 5582 20074
rect 7310 20057 7362 20069
rect 5854 20018 5906 20030
rect 5170 19966 5182 20018
rect 5234 19966 5246 20018
rect 6850 19966 6862 20018
rect 6914 19966 6926 20018
rect 7310 19993 7362 20005
rect 7534 20018 7586 20030
rect 4846 19954 4898 19966
rect 5854 19954 5906 19966
rect 7534 19954 7586 19966
rect 7870 20018 7922 20030
rect 7870 19954 7922 19966
rect 8318 20018 8370 20030
rect 8318 19954 8370 19966
rect 8542 20018 8594 20030
rect 9438 20018 9490 20030
rect 8810 19966 8822 20018
rect 8874 19966 8886 20018
rect 30270 20056 30322 20068
rect 30830 20066 30882 20078
rect 12518 20010 12570 20022
rect 12898 19966 12910 20018
rect 12962 19966 12974 20018
rect 13122 19994 13134 20046
rect 13186 19994 13198 20046
rect 13862 20018 13914 20030
rect 8542 19954 8594 19966
rect 9438 19954 9490 19966
rect 13862 19954 13914 19966
rect 14030 20018 14082 20030
rect 18174 20018 18226 20030
rect 14802 19966 14814 20018
rect 14866 19966 14878 20018
rect 14030 19954 14082 19966
rect 18174 19954 18226 19966
rect 18398 20018 18450 20030
rect 18398 19954 18450 19966
rect 18846 20018 18898 20030
rect 21870 20018 21922 20030
rect 19618 19966 19630 20018
rect 19682 19966 19694 20018
rect 18846 19954 18898 19966
rect 21870 19954 21922 19966
rect 22094 20018 22146 20030
rect 22094 19954 22146 19966
rect 23550 20018 23602 20030
rect 23550 19954 23602 19966
rect 26910 20018 26962 20030
rect 26910 19954 26962 19966
rect 27022 20018 27074 20030
rect 27794 19966 27806 20018
rect 27858 19966 27870 20018
rect 30270 19992 30322 20004
rect 30594 19966 30606 20018
rect 30658 19966 30670 20018
rect 31938 19981 31950 20033
rect 32002 19981 32014 20033
rect 32958 20018 33010 20030
rect 27022 19954 27074 19966
rect 30998 19962 31050 19974
rect 32274 19966 32286 20018
rect 32338 19966 32350 20018
rect 3222 19898 3274 19910
rect 5518 19906 5570 19918
rect 12686 19906 12738 19918
rect 32958 19954 33010 19966
rect 6962 19854 6974 19906
rect 7026 19854 7038 19906
rect 10210 19854 10222 19906
rect 10274 19854 10286 19906
rect 12114 19854 12126 19906
rect 12178 19854 12190 19906
rect 16706 19854 16718 19906
rect 16770 19854 16782 19906
rect 21522 19854 21534 19906
rect 21586 19854 21598 19906
rect 29698 19854 29710 19906
rect 29762 19854 29774 19906
rect 30998 19898 31050 19910
rect 31826 19854 31838 19906
rect 31890 19854 31902 19906
rect 5518 19842 5570 19854
rect 12686 19842 12738 19854
rect 26574 19794 26626 19806
rect 17882 19742 17894 19794
rect 17946 19742 17958 19794
rect 26574 19730 26626 19742
rect 33294 19794 33346 19806
rect 33294 19730 33346 19742
rect 1344 19626 34608 19660
rect 1344 19574 5372 19626
rect 5424 19574 5476 19626
rect 5528 19574 5580 19626
rect 5632 19574 13688 19626
rect 13740 19574 13792 19626
rect 13844 19574 13896 19626
rect 13948 19574 22004 19626
rect 22056 19574 22108 19626
rect 22160 19574 22212 19626
rect 22264 19574 30320 19626
rect 30372 19574 30424 19626
rect 30476 19574 30528 19626
rect 30580 19574 34608 19626
rect 1344 19540 34608 19574
rect 7590 19458 7642 19470
rect 2942 19402 2994 19414
rect 4958 19402 5010 19414
rect 10670 19458 10722 19470
rect 2942 19338 2994 19350
rect 3838 19346 3890 19358
rect 5842 19350 5854 19402
rect 5906 19350 5918 19402
rect 7590 19394 7642 19406
rect 7982 19402 8034 19414
rect 4958 19338 5010 19350
rect 7982 19338 8034 19350
rect 9214 19402 9266 19414
rect 10670 19394 10722 19406
rect 15280 19458 15332 19470
rect 15280 19394 15332 19406
rect 9214 19338 9266 19350
rect 17614 19346 17666 19358
rect 31222 19346 31274 19358
rect 3838 19282 3890 19294
rect 14534 19290 14586 19302
rect 3502 19234 3554 19246
rect 6862 19234 6914 19246
rect 2594 19182 2606 19234
rect 2658 19182 2670 19234
rect 2818 19182 2830 19234
rect 2882 19182 2894 19234
rect 4162 19182 4174 19234
rect 4226 19182 4238 19234
rect 4498 19182 4510 19234
rect 4562 19182 4574 19234
rect 4834 19182 4846 19234
rect 4898 19182 4910 19234
rect 5730 19182 5742 19234
rect 5794 19182 5806 19234
rect 3502 19170 3554 19182
rect 3826 19126 3838 19178
rect 3890 19126 3902 19178
rect 6406 19144 6418 19196
rect 6470 19144 6482 19196
rect 6862 19170 6914 19182
rect 7030 19234 7082 19246
rect 7310 19234 7362 19246
rect 11006 19234 11058 19246
rect 11566 19234 11618 19246
rect 7186 19182 7198 19234
rect 7250 19182 7262 19234
rect 8082 19182 8094 19234
rect 8146 19182 8158 19234
rect 8418 19182 8430 19234
rect 8482 19182 8494 19234
rect 8754 19182 8766 19234
rect 8818 19182 8830 19234
rect 9090 19182 9102 19234
rect 9154 19182 9166 19234
rect 11274 19182 11286 19234
rect 11338 19182 11350 19234
rect 7030 19170 7082 19182
rect 7310 19170 7362 19182
rect 11006 19170 11058 19182
rect 11566 19170 11618 19182
rect 11790 19234 11842 19246
rect 12114 19238 12126 19290
rect 12178 19238 12190 19290
rect 12966 19234 13018 19246
rect 13806 19234 13858 19246
rect 11790 19170 11842 19182
rect 12238 19196 12290 19208
rect 13514 19182 13526 19234
rect 13578 19182 13590 19234
rect 12966 19170 13018 19182
rect 13806 19170 13858 19182
rect 13918 19234 13970 19246
rect 13918 19170 13970 19182
rect 14366 19234 14418 19246
rect 16326 19290 16378 19302
rect 14534 19226 14586 19238
rect 15038 19234 15090 19246
rect 14366 19170 14418 19182
rect 15038 19170 15090 19182
rect 16158 19234 16210 19246
rect 21970 19294 21982 19346
rect 22034 19294 22046 19346
rect 25890 19294 25902 19346
rect 25954 19294 25966 19346
rect 29138 19294 29150 19346
rect 29202 19294 29214 19346
rect 33506 19294 33518 19346
rect 33570 19294 33582 19346
rect 17614 19282 17666 19294
rect 31222 19282 31274 19294
rect 16326 19226 16378 19238
rect 16606 19234 16658 19246
rect 16482 19182 16494 19234
rect 16546 19182 16558 19234
rect 16158 19170 16210 19182
rect 16606 19170 16658 19182
rect 16886 19234 16938 19246
rect 17950 19234 18002 19246
rect 17266 19182 17278 19234
rect 17330 19182 17342 19234
rect 16886 19170 16938 19182
rect 12238 19132 12290 19144
rect 12798 19122 12850 19134
rect 17714 19126 17726 19178
rect 17778 19126 17790 19178
rect 17950 19170 18002 19182
rect 18286 19234 18338 19246
rect 19966 19234 20018 19246
rect 24670 19234 24722 19246
rect 18286 19170 18338 19182
rect 19394 19167 19406 19219
rect 19458 19167 19470 19219
rect 19730 19182 19742 19234
rect 19794 19182 19806 19234
rect 21522 19182 21534 19234
rect 21586 19182 21598 19234
rect 23874 19182 23886 19234
rect 23938 19182 23950 19234
rect 19966 19170 20018 19182
rect 24670 19170 24722 19182
rect 25118 19234 25170 19246
rect 34302 19234 34354 19246
rect 29586 19182 29598 19234
rect 29650 19182 29662 19234
rect 25118 19170 25170 19182
rect 27806 19122 27858 19134
rect 29306 19126 29318 19178
rect 29370 19126 29382 19178
rect 34302 19170 34354 19182
rect 12798 19058 12850 19070
rect 21366 19066 21418 19078
rect 19618 19014 19630 19066
rect 19682 19014 19694 19066
rect 20302 19010 20354 19022
rect 27806 19058 27858 19070
rect 31614 19122 31666 19134
rect 31614 19058 31666 19070
rect 21366 19002 21418 19014
rect 30102 19010 30154 19022
rect 20302 18946 20354 18958
rect 30102 18946 30154 18958
rect 1344 18842 34768 18876
rect 1344 18790 9530 18842
rect 9582 18790 9634 18842
rect 9686 18790 9738 18842
rect 9790 18790 17846 18842
rect 17898 18790 17950 18842
rect 18002 18790 18054 18842
rect 18106 18790 26162 18842
rect 26214 18790 26266 18842
rect 26318 18790 26370 18842
rect 26422 18790 34478 18842
rect 34530 18790 34582 18842
rect 34634 18790 34686 18842
rect 34738 18790 34768 18842
rect 1344 18756 34768 18790
rect 7086 18562 7138 18574
rect 8530 18566 8542 18618
rect 8594 18566 8606 18618
rect 4890 18510 4902 18562
rect 4954 18510 4966 18562
rect 6682 18510 6694 18562
rect 6746 18510 6758 18562
rect 7086 18498 7138 18510
rect 14048 18562 14100 18574
rect 5182 18450 5234 18462
rect 3266 18398 3278 18450
rect 3330 18398 3342 18450
rect 3602 18398 3614 18450
rect 3666 18398 3678 18450
rect 4050 18398 4062 18450
rect 4114 18398 4126 18450
rect 4386 18398 4398 18450
rect 4450 18398 4462 18450
rect 5182 18386 5234 18398
rect 5294 18450 5346 18462
rect 5294 18386 5346 18398
rect 6302 18450 6354 18462
rect 6302 18386 6354 18398
rect 6414 18450 6466 18462
rect 7242 18454 7254 18506
rect 7306 18454 7318 18506
rect 14048 18498 14100 18510
rect 14814 18562 14866 18574
rect 14814 18498 14866 18510
rect 15934 18562 15986 18574
rect 27122 18566 27134 18618
rect 27186 18566 27198 18618
rect 28914 18566 28926 18618
rect 28978 18566 28990 18618
rect 32162 18566 32174 18618
rect 32226 18566 32238 18618
rect 15934 18498 15986 18510
rect 21232 18487 21284 18499
rect 6414 18386 6466 18398
rect 7758 18450 7810 18462
rect 8418 18398 8430 18450
rect 8482 18398 8494 18450
rect 8754 18413 8766 18465
rect 8818 18413 8830 18465
rect 12238 18450 12290 18462
rect 7758 18386 7810 18398
rect 12238 18386 12290 18398
rect 12462 18450 12514 18462
rect 12462 18386 12514 18398
rect 13134 18450 13186 18462
rect 13806 18450 13858 18462
rect 13134 18386 13186 18398
rect 13302 18394 13354 18406
rect 8000 18338 8052 18350
rect 3490 18286 3502 18338
rect 3554 18286 3566 18338
rect 13806 18386 13858 18398
rect 14478 18450 14530 18462
rect 14926 18450 14978 18462
rect 14478 18386 14530 18398
rect 14646 18394 14698 18406
rect 13302 18330 13354 18342
rect 14926 18386 14978 18398
rect 15206 18450 15258 18462
rect 15206 18386 15258 18398
rect 15598 18450 15650 18462
rect 16046 18450 16098 18462
rect 15598 18386 15650 18398
rect 15766 18394 15818 18406
rect 14646 18330 14698 18342
rect 17490 18398 17502 18450
rect 17554 18398 17566 18450
rect 17714 18398 17726 18450
rect 17778 18398 17790 18450
rect 18162 18425 18174 18477
rect 18226 18425 18238 18477
rect 20974 18450 21026 18462
rect 21074 18398 21086 18450
rect 21138 18398 21150 18450
rect 22766 18488 22818 18500
rect 21232 18423 21284 18435
rect 22038 18450 22090 18462
rect 16046 18386 16098 18398
rect 20974 18386 21026 18398
rect 22038 18386 22090 18398
rect 22206 18450 22258 18462
rect 22418 18398 22430 18450
rect 22482 18398 22494 18450
rect 27470 18489 27522 18501
rect 22766 18424 22818 18436
rect 27122 18398 27134 18450
rect 27186 18398 27198 18450
rect 27470 18425 27522 18437
rect 27694 18450 27746 18462
rect 22206 18386 22258 18398
rect 27694 18386 27746 18398
rect 28478 18450 28530 18462
rect 28802 18425 28814 18477
rect 28866 18425 28878 18477
rect 30046 18450 30098 18462
rect 29026 18398 29038 18450
rect 29090 18398 29102 18450
rect 28478 18386 28530 18398
rect 30046 18386 30098 18398
rect 30158 18450 30210 18462
rect 30706 18398 30718 18450
rect 30770 18398 30782 18450
rect 30930 18413 30942 18465
rect 30994 18413 31006 18465
rect 31826 18454 31838 18506
rect 31890 18454 31902 18506
rect 32062 18450 32114 18462
rect 31378 18398 31390 18450
rect 31442 18398 31454 18450
rect 33282 18398 33294 18450
rect 33346 18398 33358 18450
rect 30158 18386 30210 18398
rect 32062 18386 32114 18398
rect 15766 18330 15818 18342
rect 21646 18338 21698 18350
rect 8000 18274 8052 18286
rect 17838 18282 17890 18294
rect 16326 18226 16378 18238
rect 12730 18174 12742 18226
rect 12794 18174 12806 18226
rect 31042 18286 31054 18338
rect 31106 18286 31118 18338
rect 21646 18274 21698 18286
rect 17838 18218 17890 18230
rect 19518 18226 19570 18238
rect 33126 18226 33178 18238
rect 16326 18162 16378 18174
rect 29754 18174 29766 18226
rect 29818 18174 29830 18226
rect 19518 18162 19570 18174
rect 33126 18162 33178 18174
rect 1344 18058 34608 18092
rect 1344 18006 5372 18058
rect 5424 18006 5476 18058
rect 5528 18006 5580 18058
rect 5632 18006 13688 18058
rect 13740 18006 13792 18058
rect 13844 18006 13896 18058
rect 13948 18006 22004 18058
rect 22056 18006 22108 18058
rect 22160 18006 22212 18058
rect 22264 18006 30320 18058
rect 30372 18006 30424 18058
rect 30476 18006 30528 18058
rect 30580 18006 34608 18058
rect 1344 17972 34608 18006
rect 3166 17890 3218 17902
rect 4734 17890 4786 17902
rect 3770 17838 3782 17890
rect 3834 17838 3846 17890
rect 12144 17890 12196 17902
rect 3166 17826 3218 17838
rect 4734 17826 4786 17838
rect 6078 17834 6130 17846
rect 6078 17770 6130 17782
rect 7422 17834 7474 17846
rect 19350 17890 19402 17902
rect 12144 17826 12196 17838
rect 12630 17834 12682 17846
rect 7422 17770 7474 17782
rect 12630 17770 12682 17782
rect 15822 17778 15874 17790
rect 18610 17782 18622 17834
rect 18674 17782 18686 17834
rect 19350 17826 19402 17838
rect 20638 17890 20690 17902
rect 20638 17826 20690 17838
rect 13750 17722 13802 17734
rect 3502 17666 3554 17678
rect 3502 17602 3554 17614
rect 4062 17666 4114 17678
rect 4062 17602 4114 17614
rect 4286 17666 4338 17678
rect 4286 17602 4338 17614
rect 4398 17666 4450 17678
rect 10894 17666 10946 17678
rect 5730 17614 5742 17666
rect 5794 17614 5806 17666
rect 5954 17614 5966 17666
rect 6018 17614 6030 17666
rect 6962 17614 6974 17666
rect 7026 17614 7038 17666
rect 7298 17614 7310 17666
rect 7362 17614 7374 17666
rect 7634 17614 7646 17666
rect 7698 17614 7710 17666
rect 4398 17602 4450 17614
rect 10894 17602 10946 17614
rect 11230 17666 11282 17678
rect 11230 17602 11282 17614
rect 11902 17666 11954 17678
rect 13582 17666 13634 17678
rect 12786 17614 12798 17666
rect 12850 17614 12862 17666
rect 15822 17714 15874 17726
rect 22094 17778 22146 17790
rect 30830 17778 30882 17790
rect 27794 17726 27806 17778
rect 27858 17726 27870 17778
rect 31602 17726 31614 17778
rect 31666 17726 31678 17778
rect 22094 17714 22146 17726
rect 30830 17714 30882 17726
rect 13750 17658 13802 17670
rect 14254 17666 14306 17678
rect 11386 17558 11398 17610
rect 11450 17558 11462 17610
rect 11902 17602 11954 17614
rect 13582 17602 13634 17614
rect 14254 17602 14306 17614
rect 15262 17666 15314 17678
rect 15262 17602 15314 17614
rect 15486 17666 15538 17678
rect 15486 17602 15538 17614
rect 16158 17666 16210 17678
rect 16158 17602 16210 17614
rect 17054 17666 17106 17678
rect 17054 17602 17106 17614
rect 17390 17666 17442 17678
rect 19630 17666 19682 17678
rect 18498 17614 18510 17666
rect 18562 17614 18574 17666
rect 18834 17614 18846 17666
rect 18898 17614 18910 17666
rect 17390 17602 17442 17614
rect 19630 17602 19682 17614
rect 20078 17666 20130 17678
rect 14496 17554 14548 17566
rect 19742 17554 19794 17566
rect 19898 17558 19910 17610
rect 19962 17558 19974 17610
rect 20078 17602 20130 17614
rect 20302 17666 20354 17678
rect 22766 17666 22818 17678
rect 29486 17666 29538 17678
rect 22642 17614 22654 17666
rect 22706 17614 22718 17666
rect 23314 17614 23326 17666
rect 23378 17614 23390 17666
rect 20302 17602 20354 17614
rect 22474 17558 22486 17610
rect 22538 17558 22550 17610
rect 22766 17602 22818 17614
rect 26674 17558 26686 17610
rect 26738 17558 26750 17610
rect 27122 17558 27134 17610
rect 27186 17558 27198 17610
rect 27570 17577 27582 17629
rect 27634 17577 27646 17629
rect 27768 17574 27780 17626
rect 27832 17574 27844 17626
rect 28466 17614 28478 17666
rect 28530 17614 28542 17666
rect 29486 17602 29538 17614
rect 29598 17666 29650 17678
rect 29598 17602 29650 17614
rect 30158 17666 30210 17678
rect 30158 17602 30210 17614
rect 30494 17666 30546 17678
rect 34302 17666 34354 17678
rect 30494 17602 30546 17614
rect 30718 17627 30770 17639
rect 31154 17614 31166 17666
rect 31218 17614 31230 17666
rect 33506 17614 33518 17666
rect 33570 17614 33582 17666
rect 34302 17602 34354 17614
rect 30718 17563 30770 17575
rect 14970 17502 14982 17554
rect 15034 17502 15046 17554
rect 14496 17490 14548 17502
rect 19742 17490 19794 17502
rect 23158 17498 23210 17510
rect 29194 17502 29206 17554
rect 29258 17502 29270 17554
rect 7814 17442 7866 17454
rect 7814 17378 7866 17390
rect 10558 17442 10610 17454
rect 10558 17378 10610 17390
rect 17894 17442 17946 17454
rect 23158 17434 23210 17446
rect 28310 17442 28362 17454
rect 17894 17378 17946 17390
rect 28310 17378 28362 17390
rect 1344 17274 34768 17308
rect 1344 17222 9530 17274
rect 9582 17222 9634 17274
rect 9686 17222 9738 17274
rect 9790 17222 17846 17274
rect 17898 17222 17950 17274
rect 18002 17222 18054 17274
rect 18106 17222 26162 17274
rect 26214 17222 26266 17274
rect 26318 17222 26370 17274
rect 26422 17222 34478 17274
rect 34530 17222 34582 17274
rect 34634 17222 34686 17274
rect 34738 17222 34768 17274
rect 1344 17188 34768 17222
rect 4958 17106 5010 17118
rect 4958 17042 5010 17054
rect 8710 17106 8762 17118
rect 8710 17042 8762 17054
rect 17838 17106 17890 17118
rect 17838 17042 17890 17054
rect 23606 17050 23658 17062
rect 8094 16994 8146 17006
rect 8094 16930 8146 16942
rect 12126 16994 12178 17006
rect 12126 16930 12178 16942
rect 12686 16994 12738 17006
rect 23102 16994 23154 17006
rect 12686 16930 12738 16942
rect 20190 16938 20242 16950
rect 18696 16920 18748 16932
rect 4174 16882 4226 16894
rect 4174 16818 4226 16830
rect 4510 16882 4562 16894
rect 4510 16818 4562 16830
rect 4622 16882 4674 16894
rect 4622 16818 4674 16830
rect 5406 16882 5458 16894
rect 5406 16818 5458 16830
rect 9438 16882 9490 16894
rect 13806 16882 13858 16894
rect 10210 16830 10222 16882
rect 10274 16830 10286 16882
rect 12917 16830 12929 16882
rect 12981 16830 12993 16882
rect 9438 16818 9490 16830
rect 13806 16818 13858 16830
rect 14590 16882 14642 16894
rect 14590 16818 14642 16830
rect 14814 16882 14866 16894
rect 15374 16882 15426 16894
rect 15082 16830 15094 16882
rect 15146 16830 15158 16882
rect 14814 16818 14866 16830
rect 15374 16818 15426 16830
rect 18174 16882 18226 16894
rect 18174 16818 18226 16830
rect 18398 16882 18450 16894
rect 18498 16830 18510 16882
rect 18562 16830 18574 16882
rect 18696 16856 18748 16868
rect 19462 16882 19514 16894
rect 21702 16938 21754 16950
rect 19842 16830 19854 16882
rect 19906 16830 19918 16882
rect 20190 16874 20242 16886
rect 20974 16920 21026 16932
rect 28802 16998 28814 17050
rect 28866 16998 28878 17050
rect 29586 16998 29598 17050
rect 29650 16998 29662 17050
rect 32050 16998 32062 17050
rect 32114 16998 32126 17050
rect 23606 16986 23658 16998
rect 23102 16930 23154 16942
rect 20974 16856 21026 16868
rect 21298 16830 21310 16882
rect 21362 16830 21374 16882
rect 21702 16874 21754 16886
rect 21982 16882 22034 16894
rect 28030 16882 28082 16894
rect 28578 16886 28590 16938
rect 28642 16886 28654 16938
rect 28926 16882 28978 16894
rect 29754 16886 29766 16938
rect 29818 16886 29830 16938
rect 30158 16882 30210 16894
rect 31714 16886 31726 16938
rect 31778 16886 31790 16938
rect 31950 16882 32002 16894
rect 22846 16830 22858 16882
rect 22910 16830 22922 16882
rect 23426 16830 23438 16882
rect 23490 16830 23502 16882
rect 28354 16830 28366 16882
rect 28418 16830 28430 16882
rect 29474 16830 29486 16882
rect 29538 16830 29550 16882
rect 31042 16830 31054 16882
rect 31106 16830 31118 16882
rect 31266 16830 31278 16882
rect 31330 16830 31342 16882
rect 18398 16818 18450 16830
rect 19462 16818 19514 16830
rect 21982 16818 22034 16830
rect 28030 16818 28082 16830
rect 28926 16818 28978 16830
rect 30158 16818 30210 16830
rect 31950 16818 32002 16830
rect 32958 16882 33010 16894
rect 32958 16818 33010 16830
rect 33182 16882 33234 16894
rect 33182 16818 33234 16830
rect 19070 16770 19122 16782
rect 6178 16718 6190 16770
rect 6242 16718 6254 16770
rect 19070 16706 19122 16718
rect 19630 16770 19682 16782
rect 19630 16706 19682 16718
rect 21534 16770 21586 16782
rect 25330 16718 25342 16770
rect 25394 16718 25406 16770
rect 27234 16718 27246 16770
rect 27298 16718 27310 16770
rect 21534 16706 21586 16718
rect 15710 16658 15762 16670
rect 15710 16594 15762 16606
rect 30886 16658 30938 16670
rect 33450 16606 33462 16658
rect 33514 16606 33526 16658
rect 30886 16594 30938 16606
rect 1344 16490 34608 16524
rect 1344 16438 5372 16490
rect 5424 16438 5476 16490
rect 5528 16438 5580 16490
rect 5632 16438 13688 16490
rect 13740 16438 13792 16490
rect 13844 16438 13896 16490
rect 13948 16438 22004 16490
rect 22056 16438 22108 16490
rect 22160 16438 22212 16490
rect 22264 16438 30320 16490
rect 30372 16438 30424 16490
rect 30476 16438 30528 16490
rect 30580 16438 34608 16490
rect 1344 16404 34608 16438
rect 19854 16322 19906 16334
rect 19854 16258 19906 16270
rect 26294 16322 26346 16334
rect 32834 16270 32846 16322
rect 32898 16319 32910 16322
rect 33450 16319 33462 16322
rect 32898 16273 33462 16319
rect 32898 16270 32910 16273
rect 33450 16270 33462 16273
rect 33514 16270 33526 16322
rect 26294 16258 26346 16270
rect 27358 16210 27410 16222
rect 4498 16158 4510 16210
rect 4562 16158 4574 16210
rect 10546 16158 10558 16210
rect 10610 16158 10622 16210
rect 14242 16158 14254 16210
rect 14306 16158 14318 16210
rect 16146 16158 16158 16210
rect 16210 16158 16222 16210
rect 19282 16158 19294 16210
rect 19346 16158 19358 16210
rect 22306 16158 22318 16210
rect 22370 16158 22382 16210
rect 24210 16158 24222 16210
rect 24274 16158 24286 16210
rect 27358 16146 27410 16158
rect 29318 16210 29370 16222
rect 29318 16146 29370 16158
rect 31222 16210 31274 16222
rect 31222 16146 31274 16158
rect 32286 16210 32338 16222
rect 1822 16098 1874 16110
rect 5126 16098 5178 16110
rect 2594 16046 2606 16098
rect 2658 16046 2670 16098
rect 1822 16034 1874 16046
rect 5126 16034 5178 16046
rect 7870 16098 7922 16110
rect 16942 16098 16994 16110
rect 19518 16098 19570 16110
rect 8642 16046 8654 16098
rect 8706 16046 8718 16098
rect 18834 16046 18846 16098
rect 18898 16046 18910 16098
rect 19126 16068 19178 16080
rect 7870 16034 7922 16046
rect 16942 16034 16994 16046
rect 19518 16034 19570 16046
rect 21534 16098 21586 16110
rect 27806 16098 27858 16110
rect 26114 16046 26126 16098
rect 26178 16046 26190 16098
rect 21534 16034 21586 16046
rect 26898 16018 26910 16070
rect 26962 16018 26974 16070
rect 27122 16046 27134 16098
rect 27186 16046 27198 16098
rect 27526 16042 27578 16054
rect 19126 16004 19178 16016
rect 27806 16034 27858 16046
rect 27974 16098 28026 16110
rect 27974 16034 28026 16046
rect 28254 16098 28306 16110
rect 31602 16102 31614 16154
rect 31666 16102 31678 16154
rect 32286 16146 32338 16158
rect 32454 16154 32506 16166
rect 32454 16090 32506 16102
rect 28254 16034 28306 16046
rect 31826 16018 31838 16070
rect 31890 16018 31902 16070
rect 27526 15978 27578 15990
rect 28142 15986 28194 15998
rect 28142 15922 28194 15934
rect 28534 15986 28586 15998
rect 28534 15922 28586 15934
rect 11174 15874 11226 15886
rect 11174 15810 11226 15822
rect 12518 15874 12570 15886
rect 12518 15810 12570 15822
rect 24838 15874 24890 15886
rect 24838 15810 24890 15822
rect 1344 15706 34768 15740
rect 1344 15654 9530 15706
rect 9582 15654 9634 15706
rect 9686 15654 9738 15706
rect 9790 15654 17846 15706
rect 17898 15654 17950 15706
rect 18002 15654 18054 15706
rect 18106 15654 26162 15706
rect 26214 15654 26266 15706
rect 26318 15654 26370 15706
rect 26422 15654 34478 15706
rect 34530 15654 34582 15706
rect 34634 15654 34686 15706
rect 34738 15654 34768 15706
rect 1344 15620 34768 15654
rect 4902 15538 4954 15550
rect 4902 15474 4954 15486
rect 12518 15538 12570 15550
rect 12518 15474 12570 15486
rect 17838 15538 17890 15550
rect 28926 15538 28978 15550
rect 17838 15474 17890 15486
rect 18342 15482 18394 15494
rect 4286 15426 4338 15438
rect 4286 15362 4338 15374
rect 6302 15426 6354 15438
rect 6302 15362 6354 15374
rect 14814 15426 14866 15438
rect 1598 15314 1650 15326
rect 1598 15250 1650 15262
rect 8990 15314 9042 15326
rect 9762 15262 9774 15314
rect 9826 15262 9838 15314
rect 12002 15289 12014 15341
rect 12066 15289 12078 15341
rect 14478 15314 14530 15326
rect 14634 15318 14646 15370
rect 14698 15318 14710 15370
rect 14814 15362 14866 15374
rect 15206 15426 15258 15438
rect 28926 15474 28978 15486
rect 30494 15538 30546 15550
rect 30494 15474 30546 15486
rect 18342 15418 18394 15430
rect 21758 15426 21810 15438
rect 15206 15362 15258 15374
rect 21758 15362 21810 15374
rect 8990 15250 9042 15262
rect 14478 15250 14530 15262
rect 14926 15314 14978 15326
rect 14926 15250 14978 15262
rect 16382 15314 16434 15326
rect 16382 15250 16434 15262
rect 17502 15314 17554 15326
rect 19070 15314 19122 15326
rect 28186 15318 28198 15370
rect 28250 15318 28262 15370
rect 29262 15314 29314 15326
rect 18498 15262 18510 15314
rect 18562 15262 18574 15314
rect 19842 15262 19854 15314
rect 19906 15262 19918 15314
rect 27234 15262 27246 15314
rect 27298 15262 27310 15314
rect 27570 15262 27582 15314
rect 27634 15262 27646 15314
rect 28466 15262 28478 15314
rect 28530 15262 28542 15314
rect 17502 15250 17554 15262
rect 19070 15250 19122 15262
rect 29262 15250 29314 15262
rect 30158 15314 30210 15326
rect 30158 15250 30210 15262
rect 31614 15314 31666 15326
rect 31614 15250 31666 15262
rect 31726 15314 31778 15326
rect 31726 15250 31778 15262
rect 16718 15202 16770 15214
rect 2370 15150 2382 15202
rect 2434 15150 2446 15202
rect 8194 15150 8206 15202
rect 8258 15150 8270 15202
rect 16718 15138 16770 15150
rect 22374 15202 22426 15214
rect 28018 15150 28030 15202
rect 28082 15150 28094 15202
rect 22374 15138 22426 15150
rect 27346 15094 27358 15146
rect 27410 15094 27422 15146
rect 31994 15038 32006 15090
rect 32058 15038 32070 15090
rect 1344 14922 34608 14956
rect 1344 14870 5372 14922
rect 5424 14870 5476 14922
rect 5528 14870 5580 14922
rect 5632 14870 13688 14922
rect 13740 14870 13792 14922
rect 13844 14870 13896 14922
rect 13948 14870 22004 14922
rect 22056 14870 22108 14922
rect 22160 14870 22212 14922
rect 22264 14870 30320 14922
rect 30372 14870 30424 14922
rect 30476 14870 30528 14922
rect 30580 14870 34608 14922
rect 1344 14836 34608 14870
rect 3054 14754 3106 14766
rect 3054 14690 3106 14702
rect 6750 14754 6802 14766
rect 6750 14690 6802 14702
rect 7310 14754 7362 14766
rect 7310 14690 7362 14702
rect 31154 14590 31166 14642
rect 31218 14590 31230 14642
rect 3390 14530 3442 14542
rect 3390 14466 3442 14478
rect 6414 14530 6466 14542
rect 6414 14466 6466 14478
rect 7646 14530 7698 14542
rect 12238 14530 12290 14542
rect 7858 14478 7870 14530
rect 7922 14478 7934 14530
rect 11442 14478 11454 14530
rect 11506 14478 11518 14530
rect 7646 14466 7698 14478
rect 12238 14466 12290 14478
rect 17838 14530 17890 14542
rect 26910 14530 26962 14542
rect 26021 14478 26033 14530
rect 26085 14478 26097 14530
rect 17838 14466 17890 14478
rect 26910 14466 26962 14478
rect 27694 14530 27746 14542
rect 29150 14530 29202 14542
rect 27694 14466 27746 14478
rect 28018 14451 28030 14503
rect 28082 14451 28094 14503
rect 28354 14478 28366 14530
rect 28418 14478 28430 14530
rect 29150 14466 29202 14478
rect 29262 14530 29314 14542
rect 30438 14530 30490 14542
rect 34302 14530 34354 14542
rect 29530 14478 29542 14530
rect 29594 14478 29606 14530
rect 30706 14478 30718 14530
rect 30770 14478 30782 14530
rect 29262 14466 29314 14478
rect 30438 14466 30490 14478
rect 31042 14434 31054 14486
rect 31106 14434 31118 14486
rect 33506 14478 33518 14530
rect 33570 14478 33582 14530
rect 34302 14466 34354 14478
rect 9550 14418 9602 14430
rect 9550 14354 9602 14366
rect 25790 14418 25842 14430
rect 25790 14354 25842 14366
rect 31614 14418 31666 14430
rect 14646 14306 14698 14318
rect 14646 14242 14698 14254
rect 18174 14306 18226 14318
rect 28242 14310 28254 14362
rect 28306 14310 28318 14362
rect 31614 14354 31666 14366
rect 18174 14242 18226 14254
rect 1344 14138 34768 14172
rect 1344 14086 9530 14138
rect 9582 14086 9634 14138
rect 9686 14086 9738 14138
rect 9790 14086 17846 14138
rect 17898 14086 17950 14138
rect 18002 14086 18054 14138
rect 18106 14086 26162 14138
rect 26214 14086 26266 14138
rect 26318 14086 26370 14138
rect 26422 14086 34478 14138
rect 34530 14086 34582 14138
rect 34634 14086 34686 14138
rect 34738 14086 34768 14138
rect 1344 14052 34768 14086
rect 9046 13970 9098 13982
rect 9046 13906 9098 13918
rect 9718 13970 9770 13982
rect 9718 13906 9770 13918
rect 15150 13970 15202 13982
rect 15150 13906 15202 13918
rect 22934 13970 22986 13982
rect 22934 13906 22986 13918
rect 29878 13970 29930 13982
rect 29878 13906 29930 13918
rect 30326 13970 30378 13982
rect 30326 13906 30378 13918
rect 33294 13970 33346 13982
rect 17838 13858 17890 13870
rect 31042 13862 31054 13914
rect 31106 13862 31118 13914
rect 33294 13906 33346 13918
rect 2942 13746 2994 13758
rect 2942 13682 2994 13694
rect 3054 13746 3106 13758
rect 3602 13750 3614 13802
rect 3666 13750 3678 13802
rect 5182 13784 5234 13796
rect 17838 13794 17890 13806
rect 3826 13694 3838 13746
rect 3890 13694 3902 13746
rect 3054 13682 3106 13694
rect 4230 13690 4282 13702
rect 4062 13634 4114 13646
rect 4230 13626 4282 13638
rect 4454 13690 4506 13702
rect 4834 13694 4846 13746
rect 4898 13694 4910 13746
rect 5182 13720 5234 13732
rect 11790 13746 11842 13758
rect 11790 13682 11842 13694
rect 14814 13746 14866 13758
rect 14814 13682 14866 13694
rect 16382 13746 16434 13758
rect 16662 13746 16714 13758
rect 16482 13694 16494 13746
rect 16546 13694 16558 13746
rect 16382 13682 16434 13694
rect 16662 13682 16714 13694
rect 16830 13746 16882 13758
rect 16830 13682 16882 13694
rect 17726 13746 17778 13758
rect 17726 13682 17778 13694
rect 18006 13746 18058 13758
rect 18006 13682 18058 13694
rect 18174 13746 18226 13758
rect 18174 13682 18226 13694
rect 18846 13746 18898 13758
rect 18846 13682 18898 13694
rect 18958 13746 19010 13758
rect 18958 13682 19010 13694
rect 21086 13746 21138 13758
rect 21086 13682 21138 13694
rect 21310 13746 21362 13758
rect 21870 13746 21922 13758
rect 21578 13694 21590 13746
rect 21642 13694 21654 13746
rect 23202 13694 23214 13746
rect 23266 13694 23278 13746
rect 23538 13694 23550 13746
rect 23602 13694 23614 13746
rect 25330 13738 25342 13790
rect 25394 13738 25406 13790
rect 31222 13775 31274 13787
rect 26126 13746 26178 13758
rect 25666 13694 25678 13746
rect 25730 13694 25742 13746
rect 21310 13682 21362 13694
rect 21870 13682 21922 13694
rect 26126 13682 26178 13694
rect 26462 13746 26514 13758
rect 26462 13682 26514 13694
rect 26574 13746 26626 13758
rect 30930 13694 30942 13746
rect 30994 13694 31006 13746
rect 31938 13750 31950 13802
rect 32002 13750 32014 13802
rect 32286 13746 32338 13758
rect 31222 13711 31274 13723
rect 31714 13694 31726 13746
rect 31778 13694 31790 13746
rect 26574 13682 26626 13694
rect 32286 13682 32338 13694
rect 32958 13746 33010 13758
rect 32958 13682 33010 13694
rect 4454 13626 4506 13638
rect 4622 13634 4674 13646
rect 24166 13634 24218 13646
rect 31950 13634 32002 13646
rect 4062 13570 4114 13582
rect 12562 13582 12574 13634
rect 12626 13582 12638 13634
rect 14466 13582 14478 13634
rect 14530 13582 14542 13634
rect 25218 13582 25230 13634
rect 25282 13582 25294 13634
rect 27346 13582 27358 13634
rect 27410 13582 27422 13634
rect 29250 13582 29262 13634
rect 29314 13582 29326 13634
rect 4622 13570 4674 13582
rect 16102 13522 16154 13534
rect 2650 13470 2662 13522
rect 2714 13470 2726 13522
rect 16102 13458 16154 13470
rect 17446 13522 17498 13534
rect 22206 13522 22258 13534
rect 23314 13526 23326 13578
rect 23378 13526 23390 13578
rect 24166 13570 24218 13582
rect 31950 13570 32002 13582
rect 18554 13470 18566 13522
rect 18618 13470 18630 13522
rect 17446 13458 17498 13470
rect 22206 13458 22258 13470
rect 1344 13354 34608 13388
rect 1344 13302 5372 13354
rect 5424 13302 5476 13354
rect 5528 13302 5580 13354
rect 5632 13302 13688 13354
rect 13740 13302 13792 13354
rect 13844 13302 13896 13354
rect 13948 13302 22004 13354
rect 22056 13302 22108 13354
rect 22160 13302 22212 13354
rect 22264 13302 30320 13354
rect 30372 13302 30424 13354
rect 30476 13302 30528 13354
rect 30580 13302 34608 13354
rect 1344 13268 34608 13302
rect 6470 13186 6522 13198
rect 2718 13130 2770 13142
rect 4622 13130 4674 13142
rect 2718 13066 2770 13078
rect 3614 13074 3666 13086
rect 22654 13186 22706 13198
rect 27694 13186 27746 13198
rect 6470 13122 6522 13134
rect 7646 13130 7698 13142
rect 4622 13066 4674 13078
rect 11006 13130 11058 13142
rect 5618 13022 5630 13074
rect 5682 13022 5694 13074
rect 7646 13066 7698 13078
rect 9774 13074 9826 13086
rect 26954 13134 26966 13186
rect 27018 13134 27030 13186
rect 22654 13122 22706 13134
rect 27694 13122 27746 13134
rect 29374 13186 29426 13198
rect 29374 13122 29426 13134
rect 11006 13066 11058 13078
rect 17502 13074 17554 13086
rect 15810 13022 15822 13074
rect 15874 13022 15886 13074
rect 23874 13022 23886 13074
rect 23938 13022 23950 13074
rect 25778 13022 25790 13074
rect 25842 13022 25854 13074
rect 33058 13022 33070 13074
rect 33122 13022 33134 13074
rect 3614 13010 3666 13022
rect 9774 13010 9826 13022
rect 17502 13010 17554 13022
rect 10166 12962 10218 12974
rect 10446 12962 10498 12974
rect 13358 12962 13410 12974
rect 16270 12962 16322 12974
rect 2370 12910 2382 12962
rect 2434 12910 2446 12962
rect 2594 12910 2606 12962
rect 2658 12910 2670 12962
rect 3042 12910 3054 12962
rect 3106 12910 3118 12962
rect 3378 12910 3390 12962
rect 3442 12910 3454 12962
rect 3826 12910 3838 12962
rect 3890 12910 3902 12962
rect 4274 12910 4286 12962
rect 4338 12910 4350 12962
rect 4722 12910 4734 12962
rect 4786 12910 4798 12962
rect 5058 12910 5070 12962
rect 5122 12910 5134 12962
rect 5730 12895 5742 12947
rect 5794 12895 5806 12947
rect 5954 12910 5966 12962
rect 6018 12910 6030 12962
rect 6974 12934 7026 12946
rect 6738 12854 6750 12906
rect 6802 12854 6814 12906
rect 6974 12870 7026 12882
rect 7186 12854 7198 12906
rect 7250 12854 7262 12906
rect 7354 12875 7366 12927
rect 7418 12875 7430 12927
rect 7746 12910 7758 12962
rect 7810 12910 7822 12962
rect 8422 12872 8434 12924
rect 8486 12872 8498 12924
rect 10322 12910 10334 12962
rect 10386 12910 10398 12962
rect 11106 12910 11118 12962
rect 11170 12910 11182 12962
rect 11330 12910 11342 12962
rect 11394 12910 11406 12962
rect 12002 12910 12014 12962
rect 12066 12910 12078 12962
rect 14354 12910 14366 12962
rect 14418 12910 14430 12962
rect 15026 12910 15038 12962
rect 15090 12910 15102 12962
rect 15586 12910 15598 12962
rect 15650 12910 15662 12962
rect 10166 12898 10218 12910
rect 10446 12898 10498 12910
rect 13358 12898 13410 12910
rect 15922 12883 15934 12935
rect 15986 12883 15998 12935
rect 16270 12898 16322 12910
rect 16606 12962 16658 12974
rect 18174 12962 18226 12974
rect 18050 12910 18062 12962
rect 18114 12910 18126 12962
rect 16606 12898 16658 12910
rect 17882 12854 17894 12906
rect 17946 12854 17958 12906
rect 18174 12898 18226 12910
rect 18510 12962 18562 12974
rect 18958 12962 19010 12974
rect 21534 12962 21586 12974
rect 23102 12962 23154 12974
rect 18834 12910 18846 12962
rect 18898 12910 18910 12962
rect 19506 12910 19518 12962
rect 19570 12910 19582 12962
rect 22398 12910 22410 12962
rect 22462 12910 22474 12962
rect 18510 12898 18562 12910
rect 18666 12854 18678 12906
rect 18730 12854 18742 12906
rect 18958 12898 19010 12910
rect 21534 12898 21586 12910
rect 23102 12898 23154 12910
rect 26462 12962 26514 12974
rect 26462 12898 26514 12910
rect 26686 12962 26738 12974
rect 26686 12898 26738 12910
rect 28030 12962 28082 12974
rect 28030 12898 28082 12910
rect 28702 12962 28754 12974
rect 28702 12898 28754 12910
rect 29038 12962 29090 12974
rect 29038 12898 29090 12910
rect 29934 12962 29986 12974
rect 29934 12898 29986 12910
rect 30270 12962 30322 12974
rect 30270 12898 30322 12910
rect 30382 12962 30434 12974
rect 31154 12910 31166 12962
rect 31218 12910 31230 12962
rect 30382 12898 30434 12910
rect 33618 12895 33630 12947
rect 33682 12895 33694 12947
rect 33842 12910 33854 12962
rect 33906 12910 33918 12962
rect 19238 12850 19290 12862
rect 15206 12794 15258 12806
rect 13694 12738 13746 12750
rect 13694 12674 13746 12686
rect 14198 12738 14250 12750
rect 14198 12674 14250 12686
rect 14870 12738 14922 12750
rect 19238 12786 19290 12798
rect 19686 12794 19738 12806
rect 15206 12730 15258 12742
rect 33630 12794 33682 12806
rect 19686 12730 19738 12742
rect 28366 12738 28418 12750
rect 14870 12674 14922 12686
rect 33630 12730 33682 12742
rect 28366 12674 28418 12686
rect 1344 12570 34768 12604
rect 1344 12518 9530 12570
rect 9582 12518 9634 12570
rect 9686 12518 9738 12570
rect 9790 12518 17846 12570
rect 17898 12518 17950 12570
rect 18002 12518 18054 12570
rect 18106 12518 26162 12570
rect 26214 12518 26266 12570
rect 26318 12518 26370 12570
rect 26422 12518 34478 12570
rect 34530 12518 34582 12570
rect 34634 12518 34686 12570
rect 34738 12518 34768 12570
rect 1344 12484 34768 12518
rect 15318 12402 15370 12414
rect 15318 12338 15370 12350
rect 2830 12290 2882 12302
rect 6974 12290 7026 12302
rect 2830 12226 2882 12238
rect 6302 12234 6354 12246
rect 2662 12178 2714 12190
rect 3042 12126 3054 12178
rect 3106 12126 3118 12178
rect 3266 12154 3278 12206
rect 3330 12154 3342 12206
rect 3838 12178 3890 12190
rect 3994 12182 4006 12234
rect 4058 12182 4070 12234
rect 2662 12114 2714 12126
rect 3838 12114 3890 12126
rect 4510 12178 4562 12190
rect 6514 12182 6526 12234
rect 6578 12182 6590 12234
rect 6974 12226 7026 12238
rect 8766 12290 8818 12302
rect 8766 12226 8818 12238
rect 10782 12290 10834 12302
rect 10782 12226 10834 12238
rect 16494 12290 16546 12302
rect 17490 12294 17502 12346
rect 17554 12294 17566 12346
rect 31266 12294 31278 12346
rect 31330 12294 31342 12346
rect 11756 12215 11808 12227
rect 16494 12226 16546 12238
rect 5282 12126 5294 12178
rect 5346 12126 5358 12178
rect 5506 12126 5518 12178
rect 5570 12126 5582 12178
rect 6302 12170 6354 12182
rect 7522 12159 7534 12211
rect 7586 12159 7598 12211
rect 7970 12162 7982 12214
rect 8034 12162 8046 12214
rect 8306 12159 8318 12211
rect 8370 12159 8382 12211
rect 8616 12159 8628 12211
rect 8680 12159 8692 12211
rect 10322 12154 10334 12206
rect 10386 12154 10398 12206
rect 10950 12178 11002 12190
rect 4510 12114 4562 12126
rect 7142 12122 7194 12134
rect 10546 12126 10558 12178
rect 10610 12126 10622 12178
rect 12014 12178 12066 12190
rect 11756 12151 11808 12163
rect 11890 12126 11902 12178
rect 11954 12126 11966 12178
rect 12450 12153 12462 12205
rect 12514 12153 12526 12205
rect 16382 12178 16434 12190
rect 16650 12182 16662 12234
rect 16714 12182 16726 12234
rect 14578 12126 14590 12178
rect 14642 12126 14654 12178
rect 4752 12066 4804 12078
rect 10950 12114 11002 12126
rect 12014 12114 12066 12126
rect 16382 12114 16434 12126
rect 16830 12178 16882 12190
rect 17714 12182 17726 12234
rect 17778 12182 17790 12234
rect 18062 12178 18114 12190
rect 22654 12178 22706 12190
rect 24210 12182 24222 12234
rect 24274 12182 24286 12234
rect 24446 12178 24498 12190
rect 17378 12126 17390 12178
rect 17442 12126 17454 12178
rect 18610 12126 18622 12178
rect 18674 12126 18686 12178
rect 18946 12126 18958 12178
rect 19010 12126 19022 12178
rect 21858 12126 21870 12178
rect 21922 12126 21934 12178
rect 22866 12126 22878 12178
rect 22930 12126 22942 12178
rect 23762 12126 23774 12178
rect 23826 12126 23838 12178
rect 25442 12153 25454 12205
rect 25506 12153 25518 12205
rect 28018 12153 28030 12205
rect 28082 12153 28094 12205
rect 31602 12182 31614 12234
rect 31666 12182 31678 12234
rect 31838 12178 31890 12190
rect 30258 12126 30270 12178
rect 30322 12126 30334 12178
rect 31154 12126 31166 12178
rect 31218 12126 31230 12178
rect 16830 12114 16882 12126
rect 18062 12114 18114 12126
rect 22654 12114 22706 12126
rect 24446 12114 24498 12126
rect 31838 12114 31890 12126
rect 7142 12058 7194 12070
rect 11342 12066 11394 12078
rect 4752 12002 4804 12014
rect 5182 12010 5234 12022
rect 19954 12014 19966 12066
rect 20018 12014 20030 12066
rect 23874 12014 23886 12066
rect 23938 12014 23950 12066
rect 11342 12002 11394 12014
rect 5182 11946 5234 11958
rect 16102 11954 16154 11966
rect 18722 11958 18734 12010
rect 18786 11958 18798 12010
rect 16102 11890 16154 11902
rect 26238 11954 26290 11966
rect 26238 11890 26290 11902
rect 1344 11786 34608 11820
rect 1344 11734 5372 11786
rect 5424 11734 5476 11786
rect 5528 11734 5580 11786
rect 5632 11734 13688 11786
rect 13740 11734 13792 11786
rect 13844 11734 13896 11786
rect 13948 11734 22004 11786
rect 22056 11734 22108 11786
rect 22160 11734 22212 11786
rect 22264 11734 30320 11786
rect 30372 11734 30424 11786
rect 30476 11734 30528 11786
rect 30580 11734 34608 11786
rect 1344 11700 34608 11734
rect 3558 11618 3610 11630
rect 3558 11554 3610 11566
rect 11902 11618 11954 11630
rect 11902 11554 11954 11566
rect 12574 11618 12626 11630
rect 12574 11554 12626 11566
rect 14982 11618 15034 11630
rect 18734 11618 18786 11630
rect 14982 11554 15034 11566
rect 16046 11562 16098 11574
rect 31994 11566 32006 11618
rect 32058 11566 32070 11618
rect 18734 11554 18786 11566
rect 16046 11498 16098 11510
rect 29318 11506 29370 11518
rect 4118 11450 4170 11462
rect 24322 11454 24334 11506
rect 24386 11454 24398 11506
rect 25330 11454 25342 11506
rect 25394 11454 25406 11506
rect 3838 11394 3890 11406
rect 29318 11442 29370 11454
rect 29766 11506 29818 11518
rect 29766 11442 29818 11454
rect 30214 11506 30266 11518
rect 32722 11454 32734 11506
rect 32786 11454 32798 11506
rect 30214 11442 30266 11454
rect 4118 11386 4170 11398
rect 4286 11394 4338 11406
rect 3838 11330 3890 11342
rect 9102 11394 9154 11406
rect 10558 11394 10610 11406
rect 4286 11330 4338 11342
rect 6974 11359 7026 11371
rect 7310 11366 7362 11378
rect 6974 11295 7026 11307
rect 3950 11282 4002 11294
rect 7074 11286 7086 11338
rect 7138 11286 7150 11338
rect 7310 11302 7362 11314
rect 7522 11286 7534 11338
rect 7586 11286 7598 11338
rect 9102 11330 9154 11342
rect 9326 11355 9378 11367
rect 9650 11342 9662 11394
rect 9714 11342 9726 11394
rect 10558 11330 10610 11342
rect 11230 11394 11282 11406
rect 11230 11330 11282 11342
rect 11454 11394 11506 11406
rect 11454 11330 11506 11342
rect 12238 11394 12290 11406
rect 12238 11330 12290 11342
rect 12910 11394 12962 11406
rect 14478 11394 14530 11406
rect 13682 11342 13694 11394
rect 13746 11342 13758 11394
rect 12910 11330 12962 11342
rect 14478 11330 14530 11342
rect 15262 11394 15314 11406
rect 15262 11330 15314 11342
rect 15542 11394 15594 11406
rect 15542 11330 15594 11342
rect 15710 11394 15762 11406
rect 15710 11330 15762 11342
rect 16102 11394 16154 11406
rect 17950 11394 18002 11406
rect 16102 11330 16154 11342
rect 16886 11304 16898 11356
rect 16950 11304 16962 11356
rect 17658 11342 17670 11394
rect 17722 11342 17734 11394
rect 17950 11330 18002 11342
rect 18062 11394 18114 11406
rect 18062 11330 18114 11342
rect 19070 11394 19122 11406
rect 19070 11330 19122 11342
rect 22430 11394 22482 11406
rect 22430 11330 22482 11342
rect 25118 11394 25170 11406
rect 26742 11394 26794 11406
rect 25118 11330 25170 11342
rect 3950 11218 4002 11230
rect 7814 11282 7866 11294
rect 9326 11291 9378 11303
rect 25442 11298 25454 11350
rect 25506 11298 25518 11350
rect 25778 11342 25790 11394
rect 25842 11342 25854 11394
rect 26742 11330 26794 11342
rect 27470 11394 27522 11406
rect 27470 11330 27522 11342
rect 27582 11394 27634 11406
rect 27582 11330 27634 11342
rect 32286 11394 32338 11406
rect 32286 11330 32338 11342
rect 32398 11394 32450 11406
rect 33170 11342 33182 11394
rect 33234 11342 33246 11394
rect 32398 11330 32450 11342
rect 15374 11282 15426 11294
rect 32890 11286 32902 11338
rect 32954 11286 32966 11338
rect 10938 11230 10950 11282
rect 11002 11230 11014 11282
rect 7814 11218 7866 11230
rect 3222 11170 3274 11182
rect 9202 11174 9214 11226
rect 9266 11174 9278 11226
rect 15374 11218 15426 11230
rect 3222 11106 3274 11118
rect 10222 11170 10274 11182
rect 10222 11106 10274 11118
rect 13526 11170 13578 11182
rect 13526 11106 13578 11118
rect 14142 11170 14194 11182
rect 14142 11106 14194 11118
rect 22038 11170 22090 11182
rect 22038 11106 22090 11118
rect 26294 11170 26346 11182
rect 26294 11106 26346 11118
rect 27134 11170 27186 11182
rect 27134 11106 27186 11118
rect 1344 11002 34768 11036
rect 1344 10950 9530 11002
rect 9582 10950 9634 11002
rect 9686 10950 9738 11002
rect 9790 10950 17846 11002
rect 17898 10950 17950 11002
rect 18002 10950 18054 11002
rect 18106 10950 26162 11002
rect 26214 10950 26266 11002
rect 26318 10950 26370 11002
rect 26422 10950 34478 11002
rect 34530 10950 34582 11002
rect 34634 10950 34686 11002
rect 34738 10950 34768 11002
rect 1344 10916 34768 10950
rect 24726 10834 24778 10846
rect 15362 10782 15374 10834
rect 15426 10831 15438 10834
rect 15810 10831 15822 10834
rect 15426 10785 15822 10831
rect 15426 10782 15438 10785
rect 15810 10782 15822 10785
rect 15874 10782 15886 10834
rect 24726 10770 24778 10782
rect 31950 10778 32002 10790
rect 4734 10722 4786 10734
rect 4734 10658 4786 10670
rect 7590 10722 7642 10734
rect 31950 10714 32002 10726
rect 33450 10670 33462 10722
rect 33514 10670 33526 10722
rect 3054 10610 3106 10622
rect 3054 10546 3106 10558
rect 3614 10610 3666 10622
rect 3614 10546 3666 10558
rect 3838 10610 3890 10622
rect 3838 10546 3890 10558
rect 4510 10610 4562 10622
rect 4860 10591 4872 10643
rect 4924 10591 4936 10643
rect 5170 10614 5182 10666
rect 5234 10614 5246 10666
rect 5618 10591 5630 10643
rect 5682 10591 5694 10643
rect 5842 10614 5854 10666
rect 5906 10614 5918 10666
rect 7590 10658 7642 10670
rect 7870 10610 7922 10622
rect 8138 10614 8150 10666
rect 8202 10614 8214 10666
rect 8318 10610 8370 10622
rect 4510 10546 4562 10558
rect 7970 10558 7982 10610
rect 8034 10558 8046 10610
rect 7870 10546 7922 10558
rect 8318 10546 8370 10558
rect 10110 10610 10162 10622
rect 12002 10558 12014 10610
rect 12066 10558 12078 10610
rect 12786 10602 12798 10654
rect 12850 10602 12862 10654
rect 29822 10649 29874 10661
rect 13918 10610 13970 10622
rect 13122 10558 13134 10610
rect 13186 10558 13198 10610
rect 10110 10546 10162 10558
rect 13918 10546 13970 10558
rect 14702 10610 14754 10622
rect 14702 10546 14754 10558
rect 14814 10610 14866 10622
rect 14814 10546 14866 10558
rect 21310 10610 21362 10622
rect 23998 10610 24050 10622
rect 23109 10558 23121 10610
rect 23173 10558 23185 10610
rect 25330 10573 25342 10625
rect 25394 10573 25406 10625
rect 25902 10610 25954 10622
rect 29262 10610 29314 10622
rect 25666 10558 25678 10610
rect 25730 10558 25742 10610
rect 26674 10558 26686 10610
rect 26738 10558 26750 10610
rect 21310 10546 21362 10558
rect 23998 10546 24050 10558
rect 25902 10546 25954 10558
rect 29262 10546 29314 10558
rect 29598 10610 29650 10622
rect 29822 10585 29874 10597
rect 30258 10558 30270 10610
rect 30322 10558 30334 10610
rect 30930 10573 30942 10625
rect 30994 10573 31006 10625
rect 32050 10614 32062 10666
rect 32114 10614 32126 10666
rect 32286 10610 32338 10622
rect 31266 10558 31278 10610
rect 31330 10558 31342 10610
rect 31714 10558 31726 10610
rect 31778 10558 31790 10610
rect 29598 10546 29650 10558
rect 32286 10546 32338 10558
rect 32958 10610 33010 10622
rect 32958 10546 33010 10558
rect 33182 10610 33234 10622
rect 33182 10546 33234 10558
rect 29934 10498 29986 10510
rect 12182 10442 12234 10454
rect 12674 10446 12686 10498
rect 12738 10446 12750 10498
rect 25218 10446 25230 10498
rect 25282 10446 25294 10498
rect 28578 10446 28590 10498
rect 28642 10446 28654 10498
rect 30818 10446 30830 10498
rect 30882 10446 30894 10498
rect 2718 10386 2770 10398
rect 4174 10386 4226 10398
rect 3322 10334 3334 10386
rect 3386 10334 3398 10386
rect 2718 10322 2770 10334
rect 4174 10322 4226 10334
rect 9774 10386 9826 10398
rect 29934 10434 29986 10446
rect 12182 10378 12234 10390
rect 13582 10386 13634 10398
rect 20974 10386 21026 10398
rect 9774 10322 9826 10334
rect 14410 10334 14422 10386
rect 14474 10334 14486 10386
rect 13582 10322 13634 10334
rect 20974 10322 21026 10334
rect 22878 10386 22930 10398
rect 22878 10322 22930 10334
rect 1344 10218 34608 10252
rect 1344 10166 5372 10218
rect 5424 10166 5476 10218
rect 5528 10166 5580 10218
rect 5632 10166 13688 10218
rect 13740 10166 13792 10218
rect 13844 10166 13896 10218
rect 13948 10166 22004 10218
rect 22056 10166 22108 10218
rect 22160 10166 22212 10218
rect 22264 10166 30320 10218
rect 30372 10166 30424 10218
rect 30476 10166 30528 10218
rect 30580 10166 34608 10218
rect 1344 10132 34608 10166
rect 3110 10050 3162 10062
rect 27302 10050 27354 10062
rect 3110 9986 3162 9998
rect 4734 9994 4786 10006
rect 8026 9998 8038 10050
rect 8090 9998 8102 10050
rect 10558 9994 10610 10006
rect 5730 9942 5742 9994
rect 5794 9942 5806 9994
rect 27302 9986 27354 9998
rect 4734 9930 4786 9942
rect 10558 9930 10610 9942
rect 16046 9938 16098 9950
rect 23942 9938 23994 9950
rect 13570 9886 13582 9938
rect 13634 9935 13646 9938
rect 14410 9935 14422 9938
rect 13634 9889 14422 9935
rect 13634 9886 13646 9889
rect 14410 9886 14422 9889
rect 14474 9886 14486 9938
rect 17826 9886 17838 9938
rect 17890 9886 17902 9938
rect 19730 9886 19742 9938
rect 19794 9886 19806 9938
rect 25666 9886 25678 9938
rect 25730 9886 25742 9938
rect 30370 9886 30382 9938
rect 30434 9886 30446 9938
rect 34066 9886 34078 9938
rect 34130 9886 34142 9938
rect 16046 9874 16098 9886
rect 23942 9874 23994 9886
rect 7086 9826 7138 9838
rect 3558 9791 3610 9803
rect 3378 9718 3390 9770
rect 3442 9718 3454 9770
rect 3558 9727 3610 9739
rect 3838 9798 3890 9810
rect 3994 9758 4006 9810
rect 4058 9758 4070 9810
rect 4274 9774 4286 9826
rect 4338 9774 4350 9826
rect 4610 9774 4622 9826
rect 4674 9774 4686 9826
rect 5730 9774 5742 9826
rect 5794 9774 5806 9826
rect 5954 9774 5966 9826
rect 6018 9774 6030 9826
rect 7086 9762 7138 9774
rect 7310 9826 7362 9838
rect 7310 9762 7362 9774
rect 8318 9826 8370 9838
rect 8318 9762 8370 9774
rect 8430 9826 8482 9838
rect 11678 9826 11730 9838
rect 10658 9774 10670 9826
rect 10722 9774 10734 9826
rect 10882 9774 10894 9826
rect 10946 9774 10958 9826
rect 11386 9774 11398 9826
rect 11450 9774 11462 9826
rect 8430 9762 8482 9774
rect 11678 9762 11730 9774
rect 11790 9826 11842 9838
rect 11790 9762 11842 9774
rect 12462 9826 12514 9838
rect 12462 9762 12514 9774
rect 12686 9826 12738 9838
rect 12686 9762 12738 9774
rect 15710 9826 15762 9838
rect 17054 9826 17106 9838
rect 22766 9826 22818 9838
rect 24782 9826 24834 9838
rect 26238 9826 26290 9838
rect 15710 9762 15762 9774
rect 15934 9787 15986 9799
rect 3838 9734 3890 9746
rect 16370 9774 16382 9826
rect 16434 9774 16446 9826
rect 17054 9762 17106 9774
rect 15934 9723 15986 9735
rect 21858 9730 21870 9782
rect 21922 9730 21934 9782
rect 22194 9774 22206 9826
rect 22258 9774 22270 9826
rect 22766 9762 22818 9774
rect 23090 9747 23102 9799
rect 23154 9747 23166 9799
rect 23314 9774 23326 9826
rect 23378 9774 23390 9826
rect 25554 9774 25566 9826
rect 25618 9774 25630 9826
rect 26014 9787 26066 9799
rect 24782 9762 24834 9774
rect 26238 9762 26290 9774
rect 26574 9826 26626 9838
rect 28366 9826 28418 9838
rect 27458 9774 27470 9826
rect 27522 9774 27534 9826
rect 27794 9774 27806 9826
rect 27858 9774 27870 9826
rect 26574 9762 26626 9774
rect 26014 9723 26066 9735
rect 27962 9718 27974 9770
rect 28026 9718 28038 9770
rect 28366 9762 28418 9774
rect 29374 9826 29426 9838
rect 31390 9826 31442 9838
rect 29374 9762 29426 9774
rect 29598 9787 29650 9799
rect 29922 9774 29934 9826
rect 29986 9774 29998 9826
rect 29598 9723 29650 9735
rect 30482 9730 30494 9782
rect 30546 9730 30558 9782
rect 30706 9774 30718 9826
rect 30770 9774 30782 9826
rect 32162 9774 32174 9826
rect 32226 9774 32238 9826
rect 31390 9762 31442 9774
rect 7578 9662 7590 9714
rect 7642 9662 7654 9714
rect 12170 9662 12182 9714
rect 12234 9662 12246 9714
rect 2774 9602 2826 9614
rect 21970 9606 21982 9658
rect 22034 9606 22046 9658
rect 22642 9606 22654 9658
rect 22706 9606 22718 9658
rect 2774 9538 2826 9550
rect 25118 9602 25170 9614
rect 28466 9606 28478 9658
rect 28530 9606 28542 9658
rect 29250 9606 29262 9658
rect 29314 9606 29326 9658
rect 25118 9538 25170 9550
rect 1344 9434 34768 9468
rect 1344 9382 9530 9434
rect 9582 9382 9634 9434
rect 9686 9382 9738 9434
rect 9790 9382 17846 9434
rect 17898 9382 17950 9434
rect 18002 9382 18054 9434
rect 18106 9382 26162 9434
rect 26214 9382 26266 9434
rect 26318 9382 26370 9434
rect 26422 9382 34478 9434
rect 34530 9382 34582 9434
rect 34634 9382 34686 9434
rect 34738 9382 34768 9434
rect 1344 9348 34768 9382
rect 33294 9266 33346 9278
rect 33294 9202 33346 9214
rect 3670 9098 3722 9110
rect 6694 9098 6746 9110
rect 3042 9018 3054 9070
rect 3106 9018 3118 9070
rect 3266 8990 3278 9042
rect 3330 8990 3342 9042
rect 3670 9034 3722 9046
rect 4162 9005 4174 9057
rect 4226 9005 4238 9057
rect 6066 9046 6078 9098
rect 6130 9046 6142 9098
rect 6526 9042 6578 9054
rect 4498 8990 4510 9042
rect 4562 8990 4574 9042
rect 6290 8990 6302 9042
rect 6354 8990 6366 9042
rect 8038 9098 8090 9110
rect 23034 9102 23046 9154
rect 23098 9102 23110 9154
rect 6694 9034 6746 9046
rect 7310 9080 7362 9092
rect 13436 9079 13488 9091
rect 7310 9016 7362 9028
rect 7634 8990 7646 9042
rect 7698 8990 7710 9042
rect 8038 9034 8090 9046
rect 12462 9042 12514 9054
rect 8418 8990 8430 9042
rect 8482 8990 8494 9042
rect 8642 8990 8654 9042
rect 8706 8990 8718 9042
rect 11106 8990 11118 9042
rect 11170 8990 11182 9042
rect 6526 8978 6578 8990
rect 12462 8978 12514 8990
rect 12686 9042 12738 9054
rect 13694 9042 13746 9054
rect 13436 9015 13488 9027
rect 13570 8990 13582 9042
rect 13634 8990 13646 9042
rect 12686 8978 12738 8990
rect 13694 8978 13746 8990
rect 14198 9042 14250 9054
rect 14198 8978 14250 8990
rect 14366 9042 14418 9054
rect 15586 9046 15598 9098
rect 15650 9046 15662 9098
rect 15822 9042 15874 9054
rect 15138 8990 15150 9042
rect 15202 8990 15214 9042
rect 14366 8978 14418 8990
rect 15822 8978 15874 8990
rect 19518 9042 19570 9054
rect 22654 9042 22706 9054
rect 20290 8990 20302 9042
rect 20354 8990 20366 9042
rect 19518 8978 19570 8990
rect 22654 8978 22706 8990
rect 22766 9042 22818 9054
rect 25330 8990 25342 9042
rect 25394 8990 25406 9042
rect 25554 9005 25566 9057
rect 25618 9005 25630 9057
rect 28018 8990 28030 9042
rect 28082 8990 28094 9042
rect 28242 9005 28254 9057
rect 28306 9005 28318 9057
rect 28914 9018 28926 9070
rect 28978 9018 28990 9070
rect 29710 9042 29762 9054
rect 29138 8990 29150 9042
rect 29202 8990 29214 9042
rect 22766 8978 22818 8990
rect 29542 8986 29594 8998
rect 3502 8930 3554 8942
rect 7870 8930 7922 8942
rect 4050 8878 4062 8930
rect 4114 8878 4126 8930
rect 13022 8930 13074 8942
rect 23606 8930 23658 8942
rect 29374 8930 29426 8942
rect 3502 8866 3554 8878
rect 7870 8866 7922 8878
rect 8318 8874 8370 8886
rect 15250 8878 15262 8930
rect 15314 8878 15326 8930
rect 22194 8878 22206 8930
rect 22258 8878 22270 8930
rect 25666 8878 25678 8930
rect 25730 8878 25742 8930
rect 28354 8878 28366 8930
rect 28418 8878 28430 8930
rect 29710 8978 29762 8990
rect 32958 9042 33010 9054
rect 32958 8978 33010 8990
rect 29542 8922 29594 8934
rect 30482 8878 30494 8930
rect 30546 8878 30558 8930
rect 32386 8878 32398 8930
rect 32450 8878 32462 8930
rect 13022 8866 13074 8878
rect 23606 8866 23658 8878
rect 29374 8866 29426 8878
rect 8318 8810 8370 8822
rect 11286 8818 11338 8830
rect 14702 8818 14754 8830
rect 12170 8766 12182 8818
rect 12234 8766 12246 8818
rect 11286 8754 11338 8766
rect 14702 8754 14754 8766
rect 1344 8650 34608 8684
rect 1344 8598 5372 8650
rect 5424 8598 5476 8650
rect 5528 8598 5580 8650
rect 5632 8598 13688 8650
rect 13740 8598 13792 8650
rect 13844 8598 13896 8650
rect 13948 8598 22004 8650
rect 22056 8598 22108 8650
rect 22160 8598 22212 8650
rect 22264 8598 30320 8650
rect 30372 8598 30424 8650
rect 30476 8598 30528 8650
rect 30580 8598 34608 8650
rect 1344 8564 34608 8598
rect 31894 8482 31946 8494
rect 4174 8426 4226 8438
rect 29530 8430 29542 8482
rect 29594 8430 29606 8482
rect 31894 8418 31946 8430
rect 4174 8362 4226 8374
rect 7086 8370 7138 8382
rect 15150 8370 15202 8382
rect 22766 8370 22818 8382
rect 3894 8314 3946 8326
rect 9538 8318 9550 8370
rect 9602 8318 9614 8370
rect 13906 8318 13918 8370
rect 13970 8318 13982 8370
rect 18946 8318 18958 8370
rect 19010 8318 19022 8370
rect 21298 8318 21310 8370
rect 21362 8318 21374 8370
rect 7086 8306 7138 8318
rect 15150 8306 15202 8318
rect 22766 8306 22818 8318
rect 28478 8370 28530 8382
rect 28478 8306 28530 8318
rect 30102 8370 30154 8382
rect 30102 8306 30154 8318
rect 3894 8250 3946 8262
rect 7422 8258 7474 8270
rect 8430 8258 8482 8270
rect 10110 8258 10162 8270
rect 3054 8202 3106 8214
rect 3266 8178 3278 8230
rect 3330 8178 3342 8230
rect 4274 8206 4286 8258
rect 4338 8206 4350 8258
rect 4498 8206 4510 8258
rect 4562 8206 4574 8258
rect 7858 8206 7870 8258
rect 7922 8206 7934 8258
rect 8194 8206 8206 8258
rect 8258 8206 8270 8258
rect 8642 8206 8654 8258
rect 8706 8206 8718 8258
rect 9090 8206 9102 8258
rect 9154 8206 9166 8258
rect 9426 8206 9438 8258
rect 9490 8206 9502 8258
rect 7422 8194 7474 8206
rect 8430 8194 8482 8206
rect 3054 8138 3106 8150
rect 3726 8146 3778 8158
rect 9762 8150 9774 8202
rect 9826 8150 9838 8202
rect 10110 8194 10162 8206
rect 11566 8258 11618 8270
rect 15598 8258 15650 8270
rect 13570 8206 13582 8258
rect 13634 8206 13646 8258
rect 11106 8150 11118 8202
rect 11170 8150 11182 8202
rect 11566 8194 11618 8206
rect 12114 8150 12126 8202
rect 12178 8150 12190 8202
rect 12562 8150 12574 8202
rect 12626 8150 12638 8202
rect 13794 8162 13806 8214
rect 13858 8162 13870 8214
rect 15486 8202 15538 8214
rect 15598 8194 15650 8206
rect 15934 8258 15986 8270
rect 15934 8194 15986 8206
rect 16270 8258 16322 8270
rect 23102 8258 23154 8270
rect 17042 8206 17054 8258
rect 17106 8206 17118 8258
rect 16270 8194 16322 8206
rect 21410 8162 21422 8214
rect 21474 8162 21486 8214
rect 21746 8206 21758 8258
rect 21810 8206 21822 8258
rect 22418 8206 22430 8258
rect 22482 8206 22494 8258
rect 22754 8150 22766 8202
rect 22818 8150 22830 8202
rect 23102 8194 23154 8206
rect 23438 8258 23490 8270
rect 27918 8258 27970 8270
rect 23438 8194 23490 8206
rect 24098 8162 24110 8214
rect 24162 8162 24174 8214
rect 24322 8206 24334 8258
rect 24386 8206 24398 8258
rect 27918 8194 27970 8206
rect 28142 8258 28194 8270
rect 28142 8194 28194 8206
rect 29038 8258 29090 8270
rect 29038 8194 29090 8206
rect 29262 8258 29314 8270
rect 32050 8206 32062 8258
rect 32114 8206 32126 8258
rect 29262 8194 29314 8206
rect 15486 8138 15538 8150
rect 3726 8082 3778 8094
rect 24210 8038 24222 8090
rect 24274 8038 24286 8090
rect 27582 8034 27634 8046
rect 27582 7970 27634 7982
rect 31222 8034 31274 8046
rect 31222 7970 31274 7982
rect 1344 7866 34768 7900
rect 1344 7814 9530 7866
rect 9582 7814 9634 7866
rect 9686 7814 9738 7866
rect 9790 7814 17846 7866
rect 17898 7814 17950 7866
rect 18002 7814 18054 7866
rect 18106 7814 26162 7866
rect 26214 7814 26266 7866
rect 26318 7814 26370 7866
rect 26422 7814 34478 7866
rect 34530 7814 34582 7866
rect 34634 7814 34686 7866
rect 34738 7814 34768 7866
rect 1344 7780 34768 7814
rect 4498 7646 4510 7698
rect 4562 7695 4574 7698
rect 4722 7695 4734 7698
rect 4562 7649 4734 7695
rect 4562 7646 4574 7649
rect 4722 7646 4734 7649
rect 4786 7646 4798 7698
rect 11554 7590 11566 7642
rect 11618 7590 11630 7642
rect 14870 7586 14922 7598
rect 7354 7534 7366 7586
rect 7418 7534 7430 7586
rect 11678 7513 11730 7525
rect 3726 7474 3778 7486
rect 7646 7474 7698 7486
rect 3154 7422 3166 7474
rect 3218 7422 3230 7474
rect 4274 7422 4286 7474
rect 4338 7471 4350 7474
rect 4610 7471 4622 7474
rect 4338 7425 4622 7471
rect 4338 7422 4350 7425
rect 4610 7422 4622 7425
rect 4674 7422 4686 7474
rect 3726 7410 3778 7422
rect 7646 7410 7698 7422
rect 7870 7474 7922 7486
rect 7870 7410 7922 7422
rect 10392 7474 10444 7486
rect 10670 7474 10722 7486
rect 10546 7422 10558 7474
rect 10610 7422 10622 7474
rect 10392 7410 10444 7422
rect 10670 7410 10722 7422
rect 11454 7474 11506 7486
rect 14030 7509 14082 7521
rect 12462 7474 12514 7486
rect 11678 7449 11730 7461
rect 12002 7422 12014 7474
rect 12066 7422 12078 7474
rect 11454 7410 11506 7422
rect 12462 7410 12514 7422
rect 12630 7474 12682 7486
rect 12910 7474 12962 7486
rect 12786 7422 12798 7474
rect 12850 7422 12862 7474
rect 14030 7445 14082 7457
rect 14198 7509 14250 7521
rect 14198 7445 14250 7457
rect 14366 7502 14418 7514
rect 14578 7478 14590 7530
rect 14642 7478 14654 7530
rect 14870 7522 14922 7534
rect 22094 7586 22146 7598
rect 22094 7522 22146 7534
rect 23214 7586 23266 7598
rect 29754 7534 29766 7586
rect 29818 7534 29830 7586
rect 14366 7438 14418 7450
rect 15766 7474 15818 7486
rect 16046 7474 16098 7486
rect 12630 7410 12682 7422
rect 12910 7410 12962 7422
rect 15922 7422 15934 7474
rect 15986 7422 15998 7474
rect 15766 7410 15818 7422
rect 16046 7410 16098 7422
rect 19406 7474 19458 7486
rect 22878 7474 22930 7486
rect 23034 7478 23046 7530
rect 23098 7478 23110 7530
rect 23214 7522 23266 7534
rect 27302 7503 27354 7515
rect 20178 7422 20190 7474
rect 20242 7422 20254 7474
rect 19406 7410 19458 7422
rect 22878 7410 22930 7422
rect 23326 7474 23378 7486
rect 23326 7410 23378 7422
rect 23606 7474 23658 7486
rect 24098 7422 24110 7474
rect 24162 7422 24174 7474
rect 24434 7422 24446 7474
rect 24498 7422 24510 7474
rect 26898 7422 26910 7474
rect 26962 7422 26974 7474
rect 27302 7439 27354 7451
rect 29262 7474 29314 7486
rect 23606 7410 23658 7422
rect 29262 7410 29314 7422
rect 29486 7474 29538 7486
rect 31602 7422 31614 7474
rect 31666 7422 31678 7474
rect 31938 7437 31950 7489
rect 32002 7437 32014 7489
rect 32958 7474 33010 7486
rect 29486 7410 29538 7422
rect 32958 7410 33010 7422
rect 9998 7362 10050 7374
rect 2930 7254 2942 7306
rect 2994 7254 3006 7306
rect 9998 7298 10050 7310
rect 23998 7306 24050 7318
rect 27346 7310 27358 7362
rect 27410 7310 27422 7362
rect 32050 7310 32062 7362
rect 32114 7310 32126 7362
rect 13190 7250 13242 7262
rect 13190 7186 13242 7198
rect 15374 7250 15426 7262
rect 23998 7242 24050 7254
rect 33294 7250 33346 7262
rect 15374 7186 15426 7198
rect 33294 7186 33346 7198
rect 1344 7082 34608 7116
rect 1344 7030 5372 7082
rect 5424 7030 5476 7082
rect 5528 7030 5580 7082
rect 5632 7030 13688 7082
rect 13740 7030 13792 7082
rect 13844 7030 13896 7082
rect 13948 7030 22004 7082
rect 22056 7030 22108 7082
rect 22160 7030 22212 7082
rect 22264 7030 30320 7082
rect 30372 7030 30424 7082
rect 30476 7030 30528 7082
rect 30580 7030 34608 7082
rect 1344 6996 34608 7030
rect 5854 6914 5906 6926
rect 5854 6850 5906 6862
rect 8654 6914 8706 6926
rect 8654 6850 8706 6862
rect 11174 6914 11226 6926
rect 15710 6914 15762 6926
rect 13850 6862 13862 6914
rect 13914 6862 13926 6914
rect 11174 6850 11226 6862
rect 15710 6850 15762 6862
rect 22206 6914 22258 6926
rect 17378 6806 17390 6858
rect 17442 6806 17454 6858
rect 22206 6850 22258 6862
rect 23874 6750 23886 6802
rect 23938 6750 23950 6802
rect 25778 6750 25790 6802
rect 25842 6750 25854 6802
rect 28018 6750 28030 6802
rect 28082 6750 28094 6802
rect 32162 6750 32174 6802
rect 32226 6750 32238 6802
rect 2774 6690 2826 6702
rect 2774 6626 2826 6638
rect 3110 6690 3162 6702
rect 4230 6690 4282 6702
rect 5058 6694 5070 6746
rect 5122 6694 5134 6746
rect 3110 6626 3162 6638
rect 3390 6662 3442 6674
rect 3950 6634 4002 6646
rect 3390 6598 3442 6610
rect 3602 6582 3614 6634
rect 3666 6582 3678 6634
rect 3826 6582 3838 6634
rect 3890 6582 3902 6634
rect 5518 6690 5570 6702
rect 8094 6690 8146 6702
rect 4230 6626 4282 6638
rect 4958 6652 5010 6664
rect 5518 6626 5570 6638
rect 7534 6634 7586 6646
rect 7858 6638 7870 6690
rect 7922 6638 7934 6690
rect 8990 6690 9042 6702
rect 3950 6570 4002 6582
rect 4398 6578 4450 6590
rect 4958 6588 5010 6600
rect 8094 6626 8146 6638
rect 8262 6634 8314 6646
rect 7534 6570 7586 6582
rect 8990 6626 9042 6638
rect 11454 6690 11506 6702
rect 11454 6626 11506 6638
rect 11902 6690 11954 6702
rect 8262 6570 8314 6582
rect 11566 6578 11618 6590
rect 11722 6582 11734 6634
rect 11786 6582 11798 6634
rect 11902 6626 11954 6638
rect 13358 6690 13410 6702
rect 13358 6626 13410 6638
rect 13582 6690 13634 6702
rect 13582 6626 13634 6638
rect 14366 6690 14418 6702
rect 14366 6626 14418 6638
rect 14590 6690 14642 6702
rect 14590 6626 14642 6638
rect 15374 6690 15426 6702
rect 15374 6626 15426 6638
rect 16606 6690 16658 6702
rect 18006 6690 18058 6702
rect 22542 6690 22594 6702
rect 17042 6638 17054 6690
rect 17106 6638 17118 6690
rect 17266 6638 17278 6690
rect 17330 6638 17342 6690
rect 17602 6638 17614 6690
rect 17666 6638 17678 6690
rect 18386 6638 18398 6690
rect 18450 6638 18462 6690
rect 16606 6626 16658 6638
rect 18006 6626 18058 6638
rect 18734 6634 18786 6646
rect 16270 6578 16322 6590
rect 4398 6514 4450 6526
rect 14858 6526 14870 6578
rect 14922 6526 14934 6578
rect 11566 6514 11618 6526
rect 16270 6514 16322 6526
rect 18174 6578 18226 6590
rect 22542 6626 22594 6638
rect 22934 6690 22986 6702
rect 22934 6626 22986 6638
rect 23102 6690 23154 6702
rect 23102 6626 23154 6638
rect 26406 6690 26458 6702
rect 29486 6690 29538 6702
rect 31390 6690 31442 6702
rect 26406 6626 26458 6638
rect 28130 6594 28142 6646
rect 28194 6594 28206 6646
rect 28466 6638 28478 6690
rect 28530 6638 28542 6690
rect 30350 6638 30362 6690
rect 30414 6638 30426 6690
rect 29486 6626 29538 6638
rect 31390 6626 31442 6638
rect 34078 6690 34130 6702
rect 34078 6626 34130 6638
rect 18734 6570 18786 6582
rect 30606 6578 30658 6590
rect 29026 6526 29038 6578
rect 29090 6575 29102 6578
rect 29250 6575 29262 6578
rect 29090 6529 29262 6575
rect 29090 6526 29102 6529
rect 29250 6526 29262 6529
rect 29314 6526 29326 6578
rect 18174 6514 18226 6526
rect 30606 6514 30658 6526
rect 16886 6466 16938 6478
rect 12338 6414 12350 6466
rect 12402 6463 12414 6466
rect 12730 6463 12742 6466
rect 12402 6417 12742 6463
rect 12402 6414 12414 6417
rect 12730 6414 12742 6417
rect 12794 6414 12806 6466
rect 16886 6402 16938 6414
rect 31222 6466 31274 6478
rect 31222 6402 31274 6414
rect 1344 6298 34768 6332
rect 1344 6246 9530 6298
rect 9582 6246 9634 6298
rect 9686 6246 9738 6298
rect 9790 6246 17846 6298
rect 17898 6246 17950 6298
rect 18002 6246 18054 6298
rect 18106 6246 26162 6298
rect 26214 6246 26266 6298
rect 26318 6246 26370 6298
rect 26422 6246 34478 6298
rect 34530 6246 34582 6298
rect 34634 6246 34686 6298
rect 34738 6246 34768 6298
rect 1344 6212 34768 6246
rect 10670 6130 10722 6142
rect 10670 6066 10722 6078
rect 12014 6130 12066 6142
rect 15598 6130 15650 6142
rect 12014 6066 12066 6078
rect 14870 6074 14922 6086
rect 3110 6018 3162 6030
rect 7086 6018 7138 6030
rect 5226 5966 5238 6018
rect 5290 5966 5302 6018
rect 3110 5954 3162 5966
rect 2830 5906 2882 5918
rect 3378 5910 3390 5962
rect 3442 5910 3454 5962
rect 3602 5910 3614 5962
rect 3666 5910 3678 5962
rect 3826 5910 3838 5962
rect 3890 5910 3902 5962
rect 7086 5954 7138 5966
rect 8000 6018 8052 6030
rect 3950 5941 4002 5953
rect 3950 5877 4002 5889
rect 4734 5906 4786 5918
rect 2830 5842 2882 5854
rect 4734 5842 4786 5854
rect 4958 5906 5010 5918
rect 4958 5842 5010 5854
rect 6248 5906 6300 5918
rect 6526 5906 6578 5918
rect 7242 5910 7254 5962
rect 7306 5910 7318 5962
rect 8000 5954 8052 5966
rect 12910 6018 12962 6030
rect 12910 5954 12962 5966
rect 13302 6018 13354 6030
rect 15598 6066 15650 6078
rect 25286 6130 25338 6142
rect 14870 6010 14922 6022
rect 19518 6018 19570 6030
rect 16426 5966 16438 6018
rect 16490 5966 16502 6018
rect 13302 5954 13354 5966
rect 19518 5954 19570 5966
rect 19910 6018 19962 6030
rect 23874 6022 23886 6074
rect 23938 6022 23950 6074
rect 25286 6066 25338 6078
rect 25958 6130 26010 6142
rect 25958 6066 26010 6078
rect 19910 5954 19962 5966
rect 28814 6018 28866 6030
rect 32274 6022 32286 6074
rect 32338 6022 32350 6074
rect 33114 5966 33126 6018
rect 33178 5966 33190 6018
rect 6402 5854 6414 5906
rect 6466 5854 6478 5906
rect 6248 5842 6300 5854
rect 6526 5842 6578 5854
rect 7758 5906 7810 5918
rect 7758 5842 7810 5854
rect 11006 5906 11058 5918
rect 11678 5906 11730 5918
rect 11218 5854 11230 5906
rect 11282 5854 11294 5906
rect 11006 5842 11058 5854
rect 11678 5842 11730 5854
rect 12574 5906 12626 5918
rect 12574 5842 12626 5854
rect 12742 5906 12794 5918
rect 12742 5842 12794 5854
rect 13022 5906 13074 5918
rect 15934 5906 15986 5918
rect 15026 5854 15038 5906
rect 15090 5854 15102 5906
rect 13022 5842 13074 5854
rect 15934 5842 15986 5854
rect 16718 5906 16770 5918
rect 16718 5842 16770 5854
rect 16830 5906 16882 5918
rect 16830 5842 16882 5854
rect 17278 5906 17330 5918
rect 18162 5854 18174 5906
rect 18226 5854 18238 5906
rect 18902 5892 18914 5944
rect 18966 5892 18978 5944
rect 19182 5906 19234 5918
rect 19630 5906 19682 5918
rect 17278 5842 17330 5854
rect 19182 5842 19234 5854
rect 19350 5850 19402 5862
rect 5854 5794 5906 5806
rect 22306 5854 22318 5906
rect 22370 5854 22382 5906
rect 22642 5898 22654 5950
rect 22706 5898 22718 5950
rect 23426 5910 23438 5962
rect 23490 5910 23502 5962
rect 28814 5954 28866 5966
rect 23774 5906 23826 5918
rect 23202 5854 23214 5906
rect 23266 5854 23278 5906
rect 19630 5842 19682 5854
rect 23774 5842 23826 5854
rect 24222 5906 24274 5918
rect 26126 5906 26178 5918
rect 29486 5906 29538 5918
rect 25442 5854 25454 5906
rect 25506 5854 25518 5906
rect 26898 5854 26910 5906
rect 26962 5854 26974 5906
rect 24222 5842 24274 5854
rect 26126 5842 26178 5854
rect 29486 5842 29538 5854
rect 29822 5906 29874 5918
rect 30034 5910 30046 5962
rect 30098 5910 30110 5962
rect 31826 5910 31838 5962
rect 31890 5910 31902 5962
rect 32174 5906 32226 5918
rect 30370 5854 30382 5906
rect 30434 5854 30446 5906
rect 31602 5854 31614 5906
rect 31666 5854 31678 5906
rect 29822 5842 29874 5854
rect 32174 5842 32226 5854
rect 33406 5906 33458 5918
rect 33406 5842 33458 5854
rect 33630 5906 33682 5918
rect 33630 5842 33682 5854
rect 19350 5786 19402 5798
rect 30158 5794 30210 5806
rect 5854 5730 5906 5742
rect 18062 5738 18114 5750
rect 22754 5742 22766 5794
rect 22818 5742 22830 5794
rect 2494 5682 2546 5694
rect 2494 5618 2546 5630
rect 11398 5682 11450 5694
rect 11398 5618 11450 5630
rect 17614 5682 17666 5694
rect 30158 5730 30210 5742
rect 30998 5794 31050 5806
rect 30998 5730 31050 5742
rect 18062 5674 18114 5686
rect 24558 5682 24610 5694
rect 17614 5618 17666 5630
rect 24558 5618 24610 5630
rect 1344 5514 34608 5548
rect 1344 5462 5372 5514
rect 5424 5462 5476 5514
rect 5528 5462 5580 5514
rect 5632 5462 13688 5514
rect 13740 5462 13792 5514
rect 13844 5462 13896 5514
rect 13948 5462 22004 5514
rect 22056 5462 22108 5514
rect 22160 5462 22212 5514
rect 22264 5462 30320 5514
rect 30372 5462 30424 5514
rect 30476 5462 30528 5514
rect 30580 5462 34608 5514
rect 1344 5428 34608 5462
rect 2774 5346 2826 5358
rect 2774 5282 2826 5294
rect 3278 5346 3330 5358
rect 12462 5346 12514 5358
rect 3278 5282 3330 5294
rect 4286 5290 4338 5302
rect 10110 5290 10162 5302
rect 4946 5238 4958 5290
rect 5010 5238 5022 5290
rect 4286 5226 4338 5238
rect 6414 5234 6466 5246
rect 6414 5170 6466 5182
rect 7534 5234 7586 5246
rect 12462 5282 12514 5294
rect 18958 5346 19010 5358
rect 18958 5282 19010 5294
rect 21366 5346 21418 5358
rect 21366 5282 21418 5294
rect 26350 5346 26402 5358
rect 29194 5294 29206 5346
rect 29258 5294 29270 5346
rect 26350 5282 26402 5294
rect 10110 5226 10162 5238
rect 13638 5234 13690 5246
rect 18174 5234 18226 5246
rect 7534 5170 7586 5182
rect 11734 5178 11786 5190
rect 3614 5122 3666 5134
rect 6808 5122 6860 5134
rect 7086 5122 7138 5134
rect 2930 5070 2942 5122
rect 2994 5070 3006 5122
rect 3826 5070 3838 5122
rect 3890 5070 3902 5122
rect 4162 5070 4174 5122
rect 4226 5070 4238 5122
rect 4722 5070 4734 5122
rect 4786 5070 4798 5122
rect 4946 5070 4958 5122
rect 5010 5070 5022 5122
rect 6962 5070 6974 5122
rect 7026 5070 7038 5122
rect 3614 5058 3666 5070
rect 6808 5058 6860 5070
rect 7086 5058 7138 5070
rect 7926 5122 7978 5134
rect 8206 5122 8258 5134
rect 10988 5122 11040 5134
rect 8082 5070 8094 5122
rect 8146 5070 8158 5122
rect 10210 5070 10222 5122
rect 10274 5070 10286 5122
rect 10546 5070 10558 5122
rect 10610 5070 10622 5122
rect 7926 5058 7978 5070
rect 8206 5058 8258 5070
rect 10988 5058 11040 5070
rect 11230 5122 11282 5134
rect 14578 5182 14590 5234
rect 14642 5182 14654 5234
rect 23762 5182 23774 5234
rect 23826 5182 23838 5234
rect 27346 5182 27358 5234
rect 27410 5182 27422 5234
rect 34066 5182 34078 5234
rect 34130 5182 34142 5234
rect 13638 5170 13690 5182
rect 18174 5170 18226 5182
rect 11734 5114 11786 5126
rect 12126 5122 12178 5134
rect 11230 5058 11282 5070
rect 12126 5058 12178 5070
rect 13806 5122 13858 5134
rect 13806 5058 13858 5070
rect 16494 5122 16546 5134
rect 16494 5058 16546 5070
rect 17838 5122 17890 5134
rect 19350 5122 19402 5134
rect 19630 5122 19682 5134
rect 18498 5070 18510 5122
rect 18562 5070 18574 5122
rect 19506 5070 19518 5122
rect 19570 5070 19582 5122
rect 17838 5058 17890 5070
rect 18050 5014 18062 5066
rect 18114 5014 18126 5066
rect 19350 5058 19402 5070
rect 19630 5058 19682 5070
rect 20414 5122 20466 5134
rect 22430 5122 22482 5134
rect 21522 5070 21534 5122
rect 21586 5070 21598 5122
rect 21746 5070 21758 5122
rect 21810 5070 21822 5122
rect 22206 5083 22258 5095
rect 20414 5058 20466 5070
rect 22430 5058 22482 5070
rect 22990 5122 23042 5134
rect 22990 5058 23042 5070
rect 25678 5122 25730 5134
rect 25678 5058 25730 5070
rect 26686 5122 26738 5134
rect 28366 5122 28418 5134
rect 26898 5070 26910 5122
rect 26962 5070 26974 5122
rect 26686 5058 26738 5070
rect 27234 5055 27246 5107
rect 27298 5055 27310 5107
rect 27794 5070 27806 5122
rect 27858 5070 27870 5122
rect 28018 5043 28030 5095
rect 28082 5043 28094 5095
rect 28366 5058 28418 5070
rect 29486 5122 29538 5134
rect 29486 5058 29538 5070
rect 29598 5122 29650 5134
rect 30942 5122 30994 5134
rect 30370 5070 30382 5122
rect 30434 5070 30446 5122
rect 29598 5058 29650 5070
rect 22206 5019 22258 5031
rect 30594 5014 30606 5066
rect 30658 5014 30670 5066
rect 30942 5058 30994 5070
rect 31390 5122 31442 5134
rect 32162 5070 32174 5122
rect 32226 5070 32238 5122
rect 31390 5058 31442 5070
rect 11554 4902 11566 4954
rect 11618 4902 11630 4954
rect 20078 4898 20130 4910
rect 21858 4902 21870 4954
rect 21922 4902 21934 4954
rect 28354 4902 28366 4954
rect 28418 4902 28430 4954
rect 31042 4902 31054 4954
rect 31106 4902 31118 4954
rect 20078 4834 20130 4846
rect 1344 4730 34768 4764
rect 1344 4678 9530 4730
rect 9582 4678 9634 4730
rect 9686 4678 9738 4730
rect 9790 4678 17846 4730
rect 17898 4678 17950 4730
rect 18002 4678 18054 4730
rect 18106 4678 26162 4730
rect 26214 4678 26266 4730
rect 26318 4678 26370 4730
rect 26422 4678 34478 4730
rect 34530 4678 34582 4730
rect 34634 4678 34686 4730
rect 34738 4678 34768 4730
rect 1344 4644 34768 4678
rect 10446 4562 10498 4574
rect 10446 4498 10498 4510
rect 11118 4562 11170 4574
rect 11118 4498 11170 4510
rect 29766 4562 29818 4574
rect 4286 4450 4338 4462
rect 4286 4386 4338 4398
rect 7310 4450 7362 4462
rect 1598 4338 1650 4350
rect 4734 4338 4786 4350
rect 5598 4342 5610 4394
rect 5662 4342 5674 4394
rect 7310 4386 7362 4398
rect 16718 4450 16770 4462
rect 11936 4376 11988 4388
rect 16718 4386 16770 4398
rect 22318 4450 22370 4462
rect 23426 4454 23438 4506
rect 23490 4454 23502 4506
rect 29766 4498 29818 4510
rect 33294 4562 33346 4574
rect 33294 4498 33346 4510
rect 22318 4386 22370 4398
rect 29150 4450 29202 4462
rect 8430 4338 8482 4350
rect 2370 4286 2382 4338
rect 2434 4286 2446 4338
rect 7541 4286 7553 4338
rect 7605 4286 7617 4338
rect 1598 4274 1650 4286
rect 4734 4274 4786 4286
rect 8430 4274 8482 4286
rect 9662 4338 9714 4350
rect 9662 4274 9714 4286
rect 9998 4338 10050 4350
rect 9998 4274 10050 4286
rect 10782 4338 10834 4350
rect 10782 4274 10834 4286
rect 11454 4338 11506 4350
rect 11454 4274 11506 4286
rect 11678 4338 11730 4350
rect 11778 4286 11790 4338
rect 11842 4286 11854 4338
rect 11936 4312 11988 4324
rect 14030 4338 14082 4350
rect 17838 4338 17890 4350
rect 14802 4286 14814 4338
rect 14866 4286 14878 4338
rect 11678 4274 11730 4286
rect 14030 4274 14082 4286
rect 17838 4274 17890 4286
rect 18174 4338 18226 4350
rect 18174 4274 18226 4286
rect 19630 4338 19682 4350
rect 23314 4342 23326 4394
rect 23378 4342 23390 4394
rect 29150 4386 29202 4398
rect 23550 4338 23602 4350
rect 22978 4286 22990 4338
rect 23042 4286 23054 4338
rect 24210 4330 24222 4382
rect 24274 4330 24286 4382
rect 25118 4338 25170 4350
rect 24546 4286 24558 4338
rect 24610 4286 24622 4338
rect 19630 4274 19682 4286
rect 23550 4274 23602 4286
rect 25118 4274 25170 4286
rect 26350 4338 26402 4350
rect 26350 4274 26402 4286
rect 26462 4338 26514 4350
rect 32498 4313 32510 4365
rect 32562 4313 32574 4365
rect 32958 4338 33010 4350
rect 26462 4274 26514 4286
rect 32958 4274 33010 4286
rect 12350 4226 12402 4238
rect 26014 4226 26066 4238
rect 20402 4174 20414 4226
rect 20466 4174 20478 4226
rect 24098 4174 24110 4226
rect 24162 4174 24174 4226
rect 27234 4174 27246 4226
rect 27298 4174 27310 4226
rect 12350 4162 12402 4174
rect 26014 4162 26066 4174
rect 5854 4114 5906 4126
rect 5854 4050 5906 4062
rect 25454 4114 25506 4126
rect 25454 4050 25506 4062
rect 31502 4114 31554 4126
rect 31502 4050 31554 4062
rect 1344 3946 34608 3980
rect 1344 3894 5372 3946
rect 5424 3894 5476 3946
rect 5528 3894 5580 3946
rect 5632 3894 13688 3946
rect 13740 3894 13792 3946
rect 13844 3894 13896 3946
rect 13948 3894 22004 3946
rect 22056 3894 22108 3946
rect 22160 3894 22212 3946
rect 22264 3894 30320 3946
rect 30372 3894 30424 3946
rect 30476 3894 30528 3946
rect 30580 3894 34608 3946
rect 1344 3860 34608 3894
rect 11230 3778 11282 3790
rect 4398 3722 4450 3734
rect 11230 3714 11282 3726
rect 21086 3778 21138 3790
rect 33182 3778 33234 3790
rect 23482 3726 23494 3778
rect 23546 3726 23558 3778
rect 28634 3726 28646 3778
rect 28698 3726 28710 3778
rect 32554 3726 32566 3778
rect 32618 3726 32630 3778
rect 21086 3714 21138 3726
rect 33182 3714 33234 3726
rect 4398 3658 4450 3670
rect 5686 3666 5738 3678
rect 5686 3602 5738 3614
rect 22710 3666 22762 3678
rect 30662 3666 30714 3678
rect 26338 3614 26350 3666
rect 26402 3614 26414 3666
rect 30930 3614 30942 3666
rect 30994 3614 31006 3666
rect 22710 3602 22762 3614
rect 30662 3602 30714 3614
rect 10894 3554 10946 3566
rect 4498 3502 4510 3554
rect 4562 3502 4574 3554
rect 4834 3502 4846 3554
rect 4898 3502 4910 3554
rect 10894 3490 10946 3502
rect 18174 3554 18226 3566
rect 21422 3554 21474 3566
rect 18174 3490 18226 3502
rect 20066 3474 20078 3526
rect 20130 3474 20142 3526
rect 21422 3490 21474 3502
rect 23774 3554 23826 3566
rect 23774 3490 23826 3502
rect 23998 3554 24050 3566
rect 28926 3554 28978 3566
rect 23998 3490 24050 3502
rect 25442 3474 25454 3526
rect 25506 3474 25518 3526
rect 28926 3490 28978 3502
rect 29150 3554 29202 3566
rect 32062 3554 32114 3566
rect 29150 3490 29202 3502
rect 31042 3487 31054 3539
rect 31106 3487 31118 3539
rect 31266 3502 31278 3554
rect 31330 3502 31342 3554
rect 32062 3490 32114 3502
rect 32286 3554 32338 3566
rect 32286 3490 32338 3502
rect 32846 3554 32898 3566
rect 32846 3490 32898 3502
rect 6134 3442 6186 3454
rect 6134 3378 6186 3390
rect 10726 3442 10778 3454
rect 10726 3378 10778 3390
rect 1344 3162 34768 3196
rect 1344 3110 9530 3162
rect 9582 3110 9634 3162
rect 9686 3110 9738 3162
rect 9790 3110 17846 3162
rect 17898 3110 17950 3162
rect 18002 3110 18054 3162
rect 18106 3110 26162 3162
rect 26214 3110 26266 3162
rect 26318 3110 26370 3162
rect 26422 3110 34478 3162
rect 34530 3110 34582 3162
rect 34634 3110 34686 3162
rect 34738 3110 34768 3162
rect 1344 3076 34768 3110
<< via1 >>
rect 5372 32118 5424 32170
rect 5476 32118 5528 32170
rect 5580 32118 5632 32170
rect 13688 32118 13740 32170
rect 13792 32118 13844 32170
rect 13896 32118 13948 32170
rect 22004 32118 22056 32170
rect 22108 32118 22160 32170
rect 22212 32118 22264 32170
rect 30320 32118 30372 32170
rect 30424 32118 30476 32170
rect 30528 32118 30580 32170
rect 13134 31838 13186 31890
rect 19630 31838 19682 31890
rect 13470 31726 13522 31778
rect 16158 31726 16210 31778
rect 19182 31726 19234 31778
rect 13302 31670 13354 31722
rect 19462 31670 19514 31722
rect 15822 31502 15874 31554
rect 9530 31334 9582 31386
rect 9634 31334 9686 31386
rect 9738 31334 9790 31386
rect 17846 31334 17898 31386
rect 17950 31334 18002 31386
rect 18054 31334 18106 31386
rect 26162 31334 26214 31386
rect 26266 31334 26318 31386
rect 26370 31334 26422 31386
rect 34478 31334 34530 31386
rect 34582 31334 34634 31386
rect 34686 31334 34738 31386
rect 13134 30942 13186 30994
rect 13918 30942 13970 30994
rect 14030 30942 14082 30994
rect 14814 30942 14866 30994
rect 20526 30942 20578 30994
rect 21310 30942 21362 30994
rect 21870 30942 21922 30994
rect 25678 30942 25730 30994
rect 27246 30942 27298 30994
rect 11230 30830 11282 30882
rect 16718 30830 16770 30882
rect 18622 30830 18674 30882
rect 22654 30830 22706 30882
rect 24558 30830 24610 30882
rect 25342 30830 25394 30882
rect 27582 30718 27634 30770
rect 5372 30550 5424 30602
rect 5476 30550 5528 30602
rect 5580 30550 5632 30602
rect 13688 30550 13740 30602
rect 13792 30550 13844 30602
rect 13896 30550 13948 30602
rect 22004 30550 22056 30602
rect 22108 30550 22160 30602
rect 22212 30550 22264 30602
rect 30320 30550 30372 30602
rect 30424 30550 30476 30602
rect 30528 30550 30580 30602
rect 19966 30382 20018 30434
rect 17838 30326 17890 30378
rect 27918 30270 27970 30322
rect 9662 30158 9714 30210
rect 10446 30158 10498 30210
rect 13582 30158 13634 30210
rect 14702 30158 14754 30210
rect 15710 30158 15762 30210
rect 16382 30158 16434 30210
rect 13825 30102 13877 30154
rect 16046 30102 16098 30154
rect 16830 30158 16882 30210
rect 17054 30158 17106 30210
rect 17726 30158 17778 30210
rect 18062 30158 18114 30210
rect 18846 30158 18898 30210
rect 20302 30158 20354 30210
rect 19722 30102 19774 30154
rect 21646 30158 21698 30210
rect 22430 30158 22482 30210
rect 24670 30158 24722 30210
rect 24894 30158 24946 30210
rect 28702 30158 28754 30210
rect 29318 30158 29370 30210
rect 12350 30046 12402 30098
rect 17334 30046 17386 30098
rect 20638 30046 20690 30098
rect 16270 29990 16322 30042
rect 24334 30046 24386 30098
rect 25174 30046 25226 30098
rect 26014 30046 26066 30098
rect 12966 29934 13018 29986
rect 9530 29766 9582 29818
rect 9634 29766 9686 29818
rect 9738 29766 9790 29818
rect 17846 29766 17898 29818
rect 17950 29766 18002 29818
rect 18054 29766 18106 29818
rect 26162 29766 26214 29818
rect 26266 29766 26318 29818
rect 26370 29766 26422 29818
rect 34478 29766 34530 29818
rect 34582 29766 34634 29818
rect 34686 29766 34738 29818
rect 12798 29542 12850 29594
rect 16046 29542 16098 29594
rect 19630 29542 19682 29594
rect 23438 29542 23490 29594
rect 25790 29542 25842 29594
rect 27694 29542 27746 29594
rect 14646 29486 14698 29538
rect 20470 29486 20522 29538
rect 11790 29418 11842 29470
rect 12126 29374 12178 29426
rect 12686 29389 12738 29441
rect 12910 29374 12962 29426
rect 13358 29374 13410 29426
rect 13470 29374 13522 29426
rect 14254 29374 14306 29426
rect 14366 29374 14418 29426
rect 15934 29418 15986 29470
rect 16270 29374 16322 29426
rect 18174 29374 18226 29426
rect 18398 29418 18450 29470
rect 18958 29374 19010 29426
rect 19182 29401 19234 29453
rect 19518 29374 19570 29426
rect 19966 29374 20018 29426
rect 20190 29374 20242 29426
rect 20750 29374 20802 29426
rect 22654 29374 22706 29426
rect 22878 29418 22930 29470
rect 23326 29374 23378 29426
rect 23662 29401 23714 29453
rect 23998 29374 24050 29426
rect 25230 29374 25282 29426
rect 25566 29401 25618 29453
rect 25902 29374 25954 29426
rect 26910 29374 26962 29426
rect 27246 29401 27298 29453
rect 27582 29374 27634 29426
rect 11678 29262 11730 29314
rect 18510 29262 18562 29314
rect 22990 29262 23042 29314
rect 13750 29150 13802 29202
rect 21086 29150 21138 29202
rect 5372 28982 5424 29034
rect 5476 28982 5528 29034
rect 5580 28982 5632 29034
rect 13688 28982 13740 29034
rect 13792 28982 13844 29034
rect 13896 28982 13948 29034
rect 22004 28982 22056 29034
rect 22108 28982 22160 29034
rect 22212 28982 22264 29034
rect 30320 28982 30372 29034
rect 30424 28982 30476 29034
rect 30528 28982 30580 29034
rect 14198 28814 14250 28866
rect 15430 28814 15482 28866
rect 22990 28814 23042 28866
rect 25734 28814 25786 28866
rect 12350 28702 12402 28754
rect 12966 28702 13018 28754
rect 15038 28758 15090 28810
rect 18174 28702 18226 28754
rect 20078 28702 20130 28754
rect 23998 28702 24050 28754
rect 27134 28702 27186 28754
rect 9662 28590 9714 28642
rect 10446 28590 10498 28642
rect 13470 28590 13522 28642
rect 13638 28590 13690 28642
rect 13806 28590 13858 28642
rect 13918 28590 13970 28642
rect 14702 28590 14754 28642
rect 14926 28590 14978 28642
rect 15710 28590 15762 28642
rect 15822 28590 15874 28642
rect 17614 28590 17666 28642
rect 17838 28590 17890 28642
rect 20862 28590 20914 28642
rect 23326 28590 23378 28642
rect 23774 28590 23826 28642
rect 24110 28563 24162 28615
rect 24446 28590 24498 28642
rect 24782 28590 24834 28642
rect 25230 28590 25282 28642
rect 25454 28590 25506 28642
rect 26686 28590 26738 28642
rect 27022 28546 27074 28598
rect 27358 28590 27410 28642
rect 27582 28590 27634 28642
rect 17334 28478 17386 28530
rect 27862 28478 27914 28530
rect 9530 28198 9582 28250
rect 9634 28198 9686 28250
rect 9738 28198 9790 28250
rect 17846 28198 17898 28250
rect 17950 28198 18002 28250
rect 18054 28198 18106 28250
rect 26162 28198 26214 28250
rect 26266 28198 26318 28250
rect 26370 28198 26422 28250
rect 34478 28198 34530 28250
rect 34582 28198 34634 28250
rect 34686 28198 34738 28250
rect 11118 28030 11170 28082
rect 12350 27974 12402 28026
rect 27022 27974 27074 28026
rect 16718 27918 16770 27970
rect 28086 27918 28138 27970
rect 29206 27918 29258 27970
rect 8094 27806 8146 27858
rect 11454 27806 11506 27858
rect 12238 27806 12290 27858
rect 12686 27845 12738 27897
rect 12910 27806 12962 27858
rect 14030 27806 14082 27858
rect 21198 27806 21250 27858
rect 23774 27806 23826 27858
rect 25510 27862 25562 27914
rect 23886 27806 23938 27858
rect 25230 27806 25282 27858
rect 26798 27806 26850 27858
rect 27246 27845 27298 27897
rect 27470 27806 27522 27858
rect 28366 27806 28418 27858
rect 28478 27806 28530 27858
rect 28702 27806 28754 27858
rect 28926 27806 28978 27858
rect 14814 27694 14866 27746
rect 25678 27694 25730 27746
rect 8430 27582 8482 27634
rect 21534 27582 21586 27634
rect 23494 27582 23546 27634
rect 5372 27414 5424 27466
rect 5476 27414 5528 27466
rect 5580 27414 5632 27466
rect 13688 27414 13740 27466
rect 13792 27414 13844 27466
rect 13896 27414 13948 27466
rect 22004 27414 22056 27466
rect 22108 27414 22160 27466
rect 22212 27414 22264 27466
rect 30320 27414 30372 27466
rect 30424 27414 30476 27466
rect 30528 27414 30580 27466
rect 14478 27190 14530 27242
rect 8318 27134 8370 27186
rect 14814 27134 14866 27186
rect 17614 27134 17666 27186
rect 21982 27134 22034 27186
rect 23886 27134 23938 27186
rect 27806 27134 27858 27186
rect 7310 27022 7362 27074
rect 7534 27022 7586 27074
rect 14030 27022 14082 27074
rect 14366 27022 14418 27074
rect 14926 27007 14978 27059
rect 15262 27022 15314 27074
rect 16718 27022 16770 27074
rect 16942 27022 16994 27074
rect 17166 27022 17218 27074
rect 17502 27007 17554 27059
rect 20190 27022 20242 27074
rect 20414 27022 20466 27074
rect 21198 27022 21250 27074
rect 25118 27022 25170 27074
rect 25902 27022 25954 27074
rect 6974 26910 7026 26962
rect 10222 26910 10274 26962
rect 16438 26910 16490 26962
rect 20694 26910 20746 26962
rect 5798 26798 5850 26850
rect 10838 26798 10890 26850
rect 9530 26630 9582 26682
rect 9634 26630 9686 26682
rect 9738 26630 9790 26682
rect 17846 26630 17898 26682
rect 17950 26630 18002 26682
rect 18054 26630 18106 26682
rect 26162 26630 26214 26682
rect 26266 26630 26318 26682
rect 26370 26630 26422 26682
rect 34478 26630 34530 26682
rect 34582 26630 34634 26682
rect 34686 26630 34738 26682
rect 23214 26462 23266 26514
rect 26574 26462 26626 26514
rect 21254 26350 21306 26402
rect 2270 26238 2322 26290
rect 5294 26238 5346 26290
rect 6078 26238 6130 26290
rect 8766 26238 8818 26290
rect 8878 26238 8930 26290
rect 9662 26253 9714 26305
rect 9998 26238 10050 26290
rect 11566 26238 11618 26290
rect 12574 26238 12626 26290
rect 12686 26238 12738 26290
rect 17278 26238 17330 26290
rect 20862 26238 20914 26290
rect 20974 26238 21026 26290
rect 22878 26238 22930 26290
rect 23886 26253 23938 26305
rect 24110 26238 24162 26290
rect 26910 26238 26962 26290
rect 27582 26253 27634 26305
rect 27806 26238 27858 26290
rect 28590 26282 28642 26334
rect 28926 26238 28978 26290
rect 29262 26238 29314 26290
rect 29374 26238 29426 26290
rect 3054 26126 3106 26178
rect 4958 26126 5010 26178
rect 7982 26126 8034 26178
rect 9550 26126 9602 26178
rect 10502 26126 10554 26178
rect 11958 26126 12010 26178
rect 13190 26126 13242 26178
rect 15990 26126 16042 26178
rect 16438 26126 16490 26178
rect 18062 26126 18114 26178
rect 19966 26126 20018 26178
rect 23774 26126 23826 26178
rect 27470 26126 27522 26178
rect 28478 26126 28530 26178
rect 8486 26014 8538 26066
rect 11230 26014 11282 26066
rect 12294 26014 12346 26066
rect 29654 26014 29706 26066
rect 5372 25846 5424 25898
rect 5476 25846 5528 25898
rect 5580 25846 5632 25898
rect 13688 25846 13740 25898
rect 13792 25846 13844 25898
rect 13896 25846 13948 25898
rect 22004 25846 22056 25898
rect 22108 25846 22160 25898
rect 22212 25846 22264 25898
rect 30320 25846 30372 25898
rect 30424 25846 30476 25898
rect 30528 25846 30580 25898
rect 4846 25678 4898 25730
rect 7814 25678 7866 25730
rect 17502 25678 17554 25730
rect 19182 25622 19234 25674
rect 5798 25566 5850 25618
rect 10894 25566 10946 25618
rect 12798 25566 12850 25618
rect 15598 25566 15650 25618
rect 20414 25566 20466 25618
rect 28142 25566 28194 25618
rect 1598 25454 1650 25506
rect 2382 25454 2434 25506
rect 5182 25454 5234 25506
rect 6526 25454 6578 25506
rect 6750 25454 6802 25506
rect 7310 25454 7362 25506
rect 7422 25454 7474 25506
rect 8094 25454 8146 25506
rect 8542 25454 8594 25506
rect 8766 25454 8818 25506
rect 10110 25454 10162 25506
rect 13358 25454 13410 25506
rect 14478 25454 14530 25506
rect 8374 25398 8426 25450
rect 14590 25454 14642 25506
rect 15262 25454 15314 25506
rect 16046 25398 16098 25450
rect 16158 25426 16210 25478
rect 16886 25454 16938 25506
rect 16382 25398 16434 25450
rect 16606 25398 16658 25450
rect 17166 25454 17218 25506
rect 18958 25454 19010 25506
rect 19294 25454 19346 25506
rect 19742 25398 19794 25450
rect 19854 25416 19906 25468
rect 4286 25342 4338 25394
rect 6246 25342 6298 25394
rect 7030 25342 7082 25394
rect 8206 25342 8258 25394
rect 20582 25398 20634 25450
rect 23998 25454 24050 25506
rect 24110 25454 24162 25506
rect 24446 25454 24498 25506
rect 24558 25454 24610 25506
rect 27358 25454 27410 25506
rect 27694 25454 27746 25506
rect 28366 25454 28418 25506
rect 31166 25454 31218 25506
rect 31950 25454 32002 25506
rect 28030 25398 28082 25450
rect 32342 25454 32394 25506
rect 23718 25342 23770 25394
rect 24838 25342 24890 25394
rect 29262 25342 29314 25394
rect 9830 25230 9882 25282
rect 13526 25286 13578 25338
rect 14142 25230 14194 25282
rect 14926 25230 14978 25282
rect 23382 25230 23434 25282
rect 9530 25062 9582 25114
rect 9634 25062 9686 25114
rect 9738 25062 9790 25114
rect 17846 25062 17898 25114
rect 17950 25062 18002 25114
rect 18054 25062 18106 25114
rect 26162 25062 26214 25114
rect 26266 25062 26318 25114
rect 26370 25062 26422 25114
rect 34478 25062 34530 25114
rect 34582 25062 34634 25114
rect 34686 25062 34738 25114
rect 2718 24894 2770 24946
rect 17614 24894 17666 24946
rect 29710 24894 29762 24946
rect 24446 24838 24498 24890
rect 29038 24838 29090 24890
rect 12742 24782 12794 24834
rect 16102 24782 16154 24834
rect 19070 24782 19122 24834
rect 27862 24782 27914 24834
rect 3054 24670 3106 24722
rect 4398 24670 4450 24722
rect 4510 24670 4562 24722
rect 5182 24670 5234 24722
rect 5294 24670 5346 24722
rect 6638 24670 6690 24722
rect 6862 24670 6914 24722
rect 7702 24726 7754 24778
rect 7534 24670 7586 24722
rect 7870 24670 7922 24722
rect 7982 24670 8034 24722
rect 8262 24670 8314 24722
rect 11902 24697 11954 24749
rect 12238 24670 12290 24722
rect 12462 24670 12514 24722
rect 13246 24697 13298 24749
rect 16382 24670 16434 24722
rect 16494 24670 16546 24722
rect 17278 24670 17330 24722
rect 18398 24670 18450 24722
rect 20974 24670 21026 24722
rect 21758 24670 21810 24722
rect 22094 24670 22146 24722
rect 22430 24670 22482 24722
rect 22990 24714 23042 24766
rect 23326 24670 23378 24722
rect 23662 24670 23714 24722
rect 23998 24697 24050 24749
rect 24334 24670 24386 24722
rect 25118 24670 25170 24722
rect 27358 24670 27410 24722
rect 28590 24726 28642 24778
rect 27582 24670 27634 24722
rect 28254 24670 28306 24722
rect 28926 24670 28978 24722
rect 29374 24670 29426 24722
rect 22878 24558 22930 24610
rect 26742 24558 26794 24610
rect 4118 24446 4170 24498
rect 4902 24446 4954 24498
rect 7142 24446 7194 24498
rect 10334 24446 10386 24498
rect 14254 24446 14306 24498
rect 18566 24446 18618 24498
rect 21982 24502 22034 24554
rect 27190 24558 27242 24610
rect 25454 24446 25506 24498
rect 5372 24278 5424 24330
rect 5476 24278 5528 24330
rect 5580 24278 5632 24330
rect 13688 24278 13740 24330
rect 13792 24278 13844 24330
rect 13896 24278 13948 24330
rect 22004 24278 22056 24330
rect 22108 24278 22160 24330
rect 22212 24278 22264 24330
rect 30320 24278 30372 24330
rect 30424 24278 30476 24330
rect 30528 24278 30580 24330
rect 4342 24110 4394 24162
rect 6582 24110 6634 24162
rect 12798 24110 12850 24162
rect 16326 24110 16378 24162
rect 20694 24110 20746 24162
rect 3838 23886 3890 23938
rect 3950 23886 4002 23938
rect 4622 23886 4674 23938
rect 4902 23942 4954 23994
rect 11678 23998 11730 24050
rect 5070 23886 5122 23938
rect 5798 23886 5850 23938
rect 6078 23886 6130 23938
rect 6302 23886 6354 23938
rect 6862 23886 6914 23938
rect 7142 23942 7194 23994
rect 7310 23886 7362 23938
rect 7870 23886 7922 23938
rect 8206 23859 8258 23911
rect 8542 23886 8594 23938
rect 9326 23886 9378 23938
rect 9550 23886 9602 23938
rect 9830 23886 9882 23938
rect 10110 23886 10162 23938
rect 11006 23942 11058 23994
rect 11846 23942 11898 23994
rect 24334 23998 24386 24050
rect 26238 23998 26290 24050
rect 10222 23886 10274 23938
rect 11230 23858 11282 23910
rect 12126 23886 12178 23938
rect 12238 23886 12290 23938
rect 12404 23886 12456 23938
rect 13806 23858 13858 23910
rect 16606 23886 16658 23938
rect 16718 23886 16770 23938
rect 16942 23886 16994 23938
rect 18174 23886 18226 23938
rect 18790 23942 18842 23994
rect 19630 23942 19682 23994
rect 19518 23848 19570 23900
rect 19966 23886 20018 23938
rect 20134 23942 20186 23994
rect 20414 23886 20466 23938
rect 22654 23886 22706 23938
rect 23550 23886 23602 23938
rect 27022 23871 27074 23923
rect 27246 23886 27298 23938
rect 27694 23886 27746 23938
rect 28366 23886 28418 23938
rect 3558 23774 3610 23826
rect 4734 23774 4786 23826
rect 6974 23774 7026 23826
rect 9046 23774 9098 23826
rect 17838 23774 17890 23826
rect 8206 23718 8258 23770
rect 18958 23774 19010 23826
rect 27974 23830 28026 23882
rect 29038 23886 29090 23938
rect 20302 23774 20354 23826
rect 17278 23662 17330 23714
rect 27246 23718 27298 23770
rect 28478 23718 28530 23770
rect 22990 23662 23042 23714
rect 29374 23662 29426 23714
rect 9530 23494 9582 23546
rect 9634 23494 9686 23546
rect 9738 23494 9790 23546
rect 17846 23494 17898 23546
rect 17950 23494 18002 23546
rect 18054 23494 18106 23546
rect 26162 23494 26214 23546
rect 26266 23494 26318 23546
rect 26370 23494 26422 23546
rect 34478 23494 34530 23546
rect 34582 23494 34634 23546
rect 34686 23494 34738 23546
rect 20134 23326 20186 23378
rect 20638 23326 20690 23378
rect 26182 23326 26234 23378
rect 29878 23326 29930 23378
rect 4286 23214 4338 23266
rect 8318 23214 8370 23266
rect 1598 23102 1650 23154
rect 5610 23158 5662 23210
rect 10110 23214 10162 23266
rect 13358 23214 13410 23266
rect 26798 23214 26850 23266
rect 4734 23102 4786 23154
rect 6302 23102 6354 23154
rect 6638 23146 6690 23198
rect 8206 23102 8258 23154
rect 8486 23046 8538 23098
rect 8654 23102 8706 23154
rect 12798 23102 12850 23154
rect 13022 23102 13074 23154
rect 2382 22990 2434 23042
rect 6750 22990 6802 23042
rect 13190 23046 13242 23098
rect 13470 23102 13522 23154
rect 14030 23102 14082 23154
rect 14814 23102 14866 23154
rect 18174 23102 18226 23154
rect 18510 23140 18562 23192
rect 19294 23102 19346 23154
rect 19630 23102 19682 23154
rect 20302 23102 20354 23154
rect 22206 23129 22258 23181
rect 12014 22990 12066 23042
rect 17782 23046 17834 23098
rect 25566 23102 25618 23154
rect 25790 23102 25842 23154
rect 28702 23102 28754 23154
rect 29486 23102 29538 23154
rect 30942 23102 30994 23154
rect 16718 22990 16770 23042
rect 17950 22990 18002 23042
rect 5854 22878 5906 22930
rect 7926 22878 7978 22930
rect 13750 22878 13802 22930
rect 19182 22934 19234 22986
rect 21926 22990 21978 23042
rect 23214 22878 23266 22930
rect 25286 22878 25338 22930
rect 30606 22878 30658 22930
rect 5372 22710 5424 22762
rect 5476 22710 5528 22762
rect 5580 22710 5632 22762
rect 13688 22710 13740 22762
rect 13792 22710 13844 22762
rect 13896 22710 13948 22762
rect 22004 22710 22056 22762
rect 22108 22710 22160 22762
rect 22212 22710 22264 22762
rect 30320 22710 30372 22762
rect 30424 22710 30476 22762
rect 30528 22710 30580 22762
rect 2718 22542 2770 22594
rect 9886 22542 9938 22594
rect 12070 22542 12122 22594
rect 14366 22542 14418 22594
rect 5014 22430 5066 22482
rect 9270 22430 9322 22482
rect 12798 22430 12850 22482
rect 18510 22430 18562 22482
rect 22878 22486 22930 22538
rect 32118 22430 32170 22482
rect 3054 22318 3106 22370
rect 3726 22318 3778 22370
rect 4062 22318 4114 22370
rect 4174 22318 4226 22370
rect 3894 22262 3946 22314
rect 4454 22318 4506 22370
rect 7534 22280 7586 22332
rect 7870 22318 7922 22370
rect 8094 22318 8146 22370
rect 8262 22262 8314 22314
rect 8542 22318 8594 22370
rect 8710 22318 8762 22370
rect 8990 22318 9042 22370
rect 9550 22318 9602 22370
rect 11174 22302 11226 22354
rect 11398 22283 11450 22335
rect 12462 22318 12514 22370
rect 11566 22262 11618 22314
rect 11790 22262 11842 22314
rect 13806 22318 13858 22370
rect 14030 22318 14082 22370
rect 14702 22318 14754 22370
rect 17166 22318 17218 22370
rect 17614 22279 17666 22331
rect 17838 22318 17890 22370
rect 19070 22318 19122 22370
rect 19182 22318 19234 22370
rect 22430 22318 22482 22370
rect 22766 22318 22818 22370
rect 23102 22318 23154 22370
rect 23886 22318 23938 22370
rect 18904 22262 18956 22314
rect 29486 22290 29538 22342
rect 8878 22206 8930 22258
rect 13526 22206 13578 22258
rect 25790 22206 25842 22258
rect 10950 22094 11002 22146
rect 17278 22150 17330 22202
rect 15990 22094 16042 22146
rect 9530 21926 9582 21978
rect 9634 21926 9686 21978
rect 9738 21926 9790 21978
rect 17846 21926 17898 21978
rect 17950 21926 18002 21978
rect 18054 21926 18106 21978
rect 26162 21926 26214 21978
rect 26266 21926 26318 21978
rect 26370 21926 26422 21978
rect 34478 21926 34530 21978
rect 34582 21926 34634 21978
rect 34686 21926 34738 21978
rect 11790 21758 11842 21810
rect 18062 21758 18114 21810
rect 18566 21758 18618 21810
rect 21870 21758 21922 21810
rect 4230 21646 4282 21698
rect 4510 21534 4562 21586
rect 4734 21534 4786 21586
rect 4846 21534 4898 21586
rect 8318 21534 8370 21586
rect 8654 21534 8706 21586
rect 12126 21534 12178 21586
rect 13134 21534 13186 21586
rect 17726 21534 17778 21586
rect 18734 21534 18786 21586
rect 21422 21534 21474 21586
rect 21534 21534 21586 21586
rect 23158 21590 23210 21642
rect 23326 21646 23378 21698
rect 33238 21646 33290 21698
rect 23550 21534 23602 21586
rect 23774 21562 23826 21614
rect 29374 21534 29426 21586
rect 29486 21534 29538 21586
rect 32622 21534 32674 21586
rect 9046 21422 9098 21474
rect 22934 21422 22986 21474
rect 29934 21422 29986 21474
rect 31838 21422 31890 21474
rect 5014 21310 5066 21362
rect 13302 21310 13354 21362
rect 21086 21310 21138 21362
rect 29094 21310 29146 21362
rect 5372 21142 5424 21194
rect 5476 21142 5528 21194
rect 5580 21142 5632 21194
rect 13688 21142 13740 21194
rect 13792 21142 13844 21194
rect 13896 21142 13948 21194
rect 22004 21142 22056 21194
rect 22108 21142 22160 21194
rect 22212 21142 22264 21194
rect 30320 21142 30372 21194
rect 30424 21142 30476 21194
rect 30528 21142 30580 21194
rect 6358 20974 6410 21026
rect 32342 20974 32394 21026
rect 7646 20918 7698 20970
rect 3670 20862 3722 20914
rect 12686 20862 12738 20914
rect 15038 20862 15090 20914
rect 3950 20750 4002 20802
rect 4062 20750 4114 20802
rect 5630 20750 5682 20802
rect 5966 20750 6018 20802
rect 6078 20750 6130 20802
rect 7198 20750 7250 20802
rect 7534 20750 7586 20802
rect 11790 20750 11842 20802
rect 5798 20694 5850 20746
rect 12014 20750 12066 20802
rect 12238 20750 12290 20802
rect 14030 20750 14082 20802
rect 12518 20694 12570 20746
rect 14422 20720 14474 20772
rect 15150 20706 15202 20758
rect 15486 20750 15538 20802
rect 16158 20750 16210 20802
rect 20078 20750 20130 20802
rect 20302 20750 20354 20802
rect 20414 20750 20466 20802
rect 21366 20750 21418 20802
rect 21646 20750 21698 20802
rect 21758 20750 21810 20802
rect 22094 20750 22146 20802
rect 21926 20694 21978 20746
rect 22430 20750 22482 20802
rect 22598 20750 22650 20802
rect 22878 20750 22930 20802
rect 23438 20750 23490 20802
rect 24222 20750 24274 20802
rect 26126 20750 26178 20802
rect 26462 20750 26514 20802
rect 26686 20750 26738 20802
rect 27750 20750 27802 20802
rect 28478 20750 28530 20802
rect 29150 20722 29202 20774
rect 31390 20750 31442 20802
rect 31838 20750 31890 20802
rect 32062 20750 32114 20802
rect 11510 20638 11562 20690
rect 20694 20638 20746 20690
rect 22766 20638 22818 20690
rect 14366 20582 14418 20634
rect 23158 20638 23210 20690
rect 26966 20638 27018 20690
rect 15990 20526 16042 20578
rect 19742 20526 19794 20578
rect 28142 20526 28194 20578
rect 9530 20358 9582 20410
rect 9634 20358 9686 20410
rect 9738 20358 9790 20410
rect 17846 20358 17898 20410
rect 17950 20358 18002 20410
rect 18054 20358 18106 20410
rect 26162 20358 26214 20410
rect 26266 20358 26318 20410
rect 26370 20358 26422 20410
rect 34478 20358 34530 20410
rect 34582 20358 34634 20410
rect 34686 20358 34738 20410
rect 23886 20190 23938 20242
rect 4454 20078 4506 20130
rect 22374 20078 22426 20130
rect 30830 20078 30882 20130
rect 3054 19966 3106 20018
rect 3222 19910 3274 19962
rect 3726 19966 3778 20018
rect 3968 19966 4020 20018
rect 4734 19966 4786 20018
rect 5518 20022 5570 20074
rect 4846 19966 4898 20018
rect 5182 19966 5234 20018
rect 5854 19966 5906 20018
rect 6862 19966 6914 20018
rect 7310 20005 7362 20057
rect 7534 19966 7586 20018
rect 7870 19966 7922 20018
rect 8318 19966 8370 20018
rect 8542 19966 8594 20018
rect 8822 19966 8874 20018
rect 9438 19966 9490 20018
rect 12518 20022 12570 20074
rect 12910 19966 12962 20018
rect 13134 19994 13186 20046
rect 13862 19966 13914 20018
rect 14030 19966 14082 20018
rect 14814 19966 14866 20018
rect 18174 19966 18226 20018
rect 18398 19966 18450 20018
rect 18846 19966 18898 20018
rect 19630 19966 19682 20018
rect 21870 19966 21922 20018
rect 22094 19966 22146 20018
rect 23550 19966 23602 20018
rect 26910 19966 26962 20018
rect 27022 19966 27074 20018
rect 27806 19966 27858 20018
rect 30270 20004 30322 20056
rect 30606 19966 30658 20018
rect 31950 19981 32002 20033
rect 32286 19966 32338 20018
rect 32958 19966 33010 20018
rect 30998 19910 31050 19962
rect 5518 19854 5570 19906
rect 6974 19854 7026 19906
rect 10222 19854 10274 19906
rect 12126 19854 12178 19906
rect 12686 19854 12738 19906
rect 16718 19854 16770 19906
rect 21534 19854 21586 19906
rect 29710 19854 29762 19906
rect 31838 19854 31890 19906
rect 17894 19742 17946 19794
rect 26574 19742 26626 19794
rect 33294 19742 33346 19794
rect 5372 19574 5424 19626
rect 5476 19574 5528 19626
rect 5580 19574 5632 19626
rect 13688 19574 13740 19626
rect 13792 19574 13844 19626
rect 13896 19574 13948 19626
rect 22004 19574 22056 19626
rect 22108 19574 22160 19626
rect 22212 19574 22264 19626
rect 30320 19574 30372 19626
rect 30424 19574 30476 19626
rect 30528 19574 30580 19626
rect 2942 19350 2994 19402
rect 7590 19406 7642 19458
rect 3838 19294 3890 19346
rect 4958 19350 5010 19402
rect 5854 19350 5906 19402
rect 7982 19350 8034 19402
rect 9214 19350 9266 19402
rect 10670 19406 10722 19458
rect 15280 19406 15332 19458
rect 2606 19182 2658 19234
rect 2830 19182 2882 19234
rect 3502 19182 3554 19234
rect 4174 19182 4226 19234
rect 4510 19182 4562 19234
rect 4846 19182 4898 19234
rect 5742 19182 5794 19234
rect 3838 19126 3890 19178
rect 6418 19144 6470 19196
rect 6862 19182 6914 19234
rect 7030 19182 7082 19234
rect 7198 19182 7250 19234
rect 7310 19182 7362 19234
rect 8094 19182 8146 19234
rect 8430 19182 8482 19234
rect 8766 19182 8818 19234
rect 9102 19182 9154 19234
rect 11006 19182 11058 19234
rect 11286 19182 11338 19234
rect 11566 19182 11618 19234
rect 12126 19238 12178 19290
rect 11790 19182 11842 19234
rect 12238 19144 12290 19196
rect 12966 19182 13018 19234
rect 13526 19182 13578 19234
rect 13806 19182 13858 19234
rect 13918 19182 13970 19234
rect 14366 19182 14418 19234
rect 14534 19238 14586 19290
rect 15038 19182 15090 19234
rect 16158 19182 16210 19234
rect 16326 19238 16378 19290
rect 17614 19294 17666 19346
rect 21982 19294 22034 19346
rect 25902 19294 25954 19346
rect 29150 19294 29202 19346
rect 31222 19294 31274 19346
rect 33518 19294 33570 19346
rect 16494 19182 16546 19234
rect 16606 19182 16658 19234
rect 16886 19182 16938 19234
rect 17278 19182 17330 19234
rect 17950 19182 18002 19234
rect 17726 19126 17778 19178
rect 18286 19182 18338 19234
rect 19406 19167 19458 19219
rect 19742 19182 19794 19234
rect 19966 19182 20018 19234
rect 21534 19182 21586 19234
rect 23886 19182 23938 19234
rect 24670 19182 24722 19234
rect 25118 19182 25170 19234
rect 29598 19182 29650 19234
rect 34302 19182 34354 19234
rect 12798 19070 12850 19122
rect 29318 19126 29370 19178
rect 19630 19014 19682 19066
rect 20302 18958 20354 19010
rect 21366 19014 21418 19066
rect 27806 19070 27858 19122
rect 31614 19070 31666 19122
rect 30102 18958 30154 19010
rect 9530 18790 9582 18842
rect 9634 18790 9686 18842
rect 9738 18790 9790 18842
rect 17846 18790 17898 18842
rect 17950 18790 18002 18842
rect 18054 18790 18106 18842
rect 26162 18790 26214 18842
rect 26266 18790 26318 18842
rect 26370 18790 26422 18842
rect 34478 18790 34530 18842
rect 34582 18790 34634 18842
rect 34686 18790 34738 18842
rect 8542 18566 8594 18618
rect 4902 18510 4954 18562
rect 6694 18510 6746 18562
rect 7086 18510 7138 18562
rect 14048 18510 14100 18562
rect 3278 18398 3330 18450
rect 3614 18398 3666 18450
rect 4062 18398 4114 18450
rect 4398 18398 4450 18450
rect 5182 18398 5234 18450
rect 5294 18398 5346 18450
rect 6302 18398 6354 18450
rect 7254 18454 7306 18506
rect 14814 18510 14866 18562
rect 27134 18566 27186 18618
rect 28926 18566 28978 18618
rect 32174 18566 32226 18618
rect 15934 18510 15986 18562
rect 6414 18398 6466 18450
rect 7758 18398 7810 18450
rect 8430 18398 8482 18450
rect 8766 18413 8818 18465
rect 12238 18398 12290 18450
rect 12462 18398 12514 18450
rect 13134 18398 13186 18450
rect 3502 18286 3554 18338
rect 8000 18286 8052 18338
rect 13302 18342 13354 18394
rect 13806 18398 13858 18450
rect 14478 18398 14530 18450
rect 14646 18342 14698 18394
rect 14926 18398 14978 18450
rect 15206 18398 15258 18450
rect 15598 18398 15650 18450
rect 15766 18342 15818 18394
rect 16046 18398 16098 18450
rect 17502 18398 17554 18450
rect 17726 18398 17778 18450
rect 18174 18425 18226 18477
rect 20974 18398 21026 18450
rect 21086 18398 21138 18450
rect 21232 18435 21284 18487
rect 22038 18398 22090 18450
rect 22206 18398 22258 18450
rect 22430 18398 22482 18450
rect 22766 18436 22818 18488
rect 27134 18398 27186 18450
rect 27470 18437 27522 18489
rect 27694 18398 27746 18450
rect 28478 18398 28530 18450
rect 28814 18425 28866 18477
rect 29038 18398 29090 18450
rect 30046 18398 30098 18450
rect 30158 18398 30210 18450
rect 30718 18398 30770 18450
rect 30942 18413 30994 18465
rect 31838 18454 31890 18506
rect 31390 18398 31442 18450
rect 32062 18398 32114 18450
rect 33294 18398 33346 18450
rect 12742 18174 12794 18226
rect 16326 18174 16378 18226
rect 17838 18230 17890 18282
rect 21646 18286 21698 18338
rect 31054 18286 31106 18338
rect 19518 18174 19570 18226
rect 29766 18174 29818 18226
rect 33126 18174 33178 18226
rect 5372 18006 5424 18058
rect 5476 18006 5528 18058
rect 5580 18006 5632 18058
rect 13688 18006 13740 18058
rect 13792 18006 13844 18058
rect 13896 18006 13948 18058
rect 22004 18006 22056 18058
rect 22108 18006 22160 18058
rect 22212 18006 22264 18058
rect 30320 18006 30372 18058
rect 30424 18006 30476 18058
rect 30528 18006 30580 18058
rect 3166 17838 3218 17890
rect 3782 17838 3834 17890
rect 4734 17838 4786 17890
rect 6078 17782 6130 17834
rect 7422 17782 7474 17834
rect 12144 17838 12196 17890
rect 19350 17838 19402 17890
rect 12630 17782 12682 17834
rect 18622 17782 18674 17834
rect 20638 17838 20690 17890
rect 3502 17614 3554 17666
rect 4062 17614 4114 17666
rect 4286 17614 4338 17666
rect 4398 17614 4450 17666
rect 5742 17614 5794 17666
rect 5966 17614 6018 17666
rect 6974 17614 7026 17666
rect 7310 17614 7362 17666
rect 7646 17614 7698 17666
rect 10894 17614 10946 17666
rect 11230 17614 11282 17666
rect 11902 17614 11954 17666
rect 12798 17614 12850 17666
rect 13582 17614 13634 17666
rect 13750 17670 13802 17722
rect 15822 17726 15874 17778
rect 22094 17726 22146 17778
rect 27806 17726 27858 17778
rect 30830 17726 30882 17778
rect 31614 17726 31666 17778
rect 11398 17558 11450 17610
rect 14254 17614 14306 17666
rect 15262 17614 15314 17666
rect 15486 17614 15538 17666
rect 16158 17614 16210 17666
rect 17054 17614 17106 17666
rect 17390 17614 17442 17666
rect 18510 17614 18562 17666
rect 18846 17614 18898 17666
rect 19630 17614 19682 17666
rect 20078 17614 20130 17666
rect 19910 17558 19962 17610
rect 20302 17614 20354 17666
rect 22654 17614 22706 17666
rect 22766 17614 22818 17666
rect 23326 17614 23378 17666
rect 22486 17558 22538 17610
rect 26686 17558 26738 17610
rect 27134 17558 27186 17610
rect 27582 17577 27634 17629
rect 27780 17574 27832 17626
rect 28478 17614 28530 17666
rect 29486 17614 29538 17666
rect 29598 17614 29650 17666
rect 30158 17614 30210 17666
rect 30494 17614 30546 17666
rect 30718 17575 30770 17627
rect 31166 17614 31218 17666
rect 33518 17614 33570 17666
rect 34302 17614 34354 17666
rect 14496 17502 14548 17554
rect 14982 17502 15034 17554
rect 19742 17502 19794 17554
rect 29206 17502 29258 17554
rect 7814 17390 7866 17442
rect 10558 17390 10610 17442
rect 17894 17390 17946 17442
rect 23158 17446 23210 17498
rect 28310 17390 28362 17442
rect 9530 17222 9582 17274
rect 9634 17222 9686 17274
rect 9738 17222 9790 17274
rect 17846 17222 17898 17274
rect 17950 17222 18002 17274
rect 18054 17222 18106 17274
rect 26162 17222 26214 17274
rect 26266 17222 26318 17274
rect 26370 17222 26422 17274
rect 34478 17222 34530 17274
rect 34582 17222 34634 17274
rect 34686 17222 34738 17274
rect 4958 17054 5010 17106
rect 8710 17054 8762 17106
rect 17838 17054 17890 17106
rect 8094 16942 8146 16994
rect 12126 16942 12178 16994
rect 12686 16942 12738 16994
rect 4174 16830 4226 16882
rect 4510 16830 4562 16882
rect 4622 16830 4674 16882
rect 5406 16830 5458 16882
rect 9438 16830 9490 16882
rect 10222 16830 10274 16882
rect 12929 16830 12981 16882
rect 13806 16830 13858 16882
rect 14590 16830 14642 16882
rect 14814 16830 14866 16882
rect 15094 16830 15146 16882
rect 15374 16830 15426 16882
rect 18174 16830 18226 16882
rect 18398 16830 18450 16882
rect 18510 16830 18562 16882
rect 18696 16868 18748 16920
rect 20190 16886 20242 16938
rect 19462 16830 19514 16882
rect 19854 16830 19906 16882
rect 20974 16868 21026 16920
rect 21702 16886 21754 16938
rect 23102 16942 23154 16994
rect 23606 16998 23658 17050
rect 28814 16998 28866 17050
rect 29598 16998 29650 17050
rect 32062 16998 32114 17050
rect 21310 16830 21362 16882
rect 28590 16886 28642 16938
rect 29766 16886 29818 16938
rect 31726 16886 31778 16938
rect 21982 16830 22034 16882
rect 22858 16830 22910 16882
rect 23438 16830 23490 16882
rect 28030 16830 28082 16882
rect 28366 16830 28418 16882
rect 28926 16830 28978 16882
rect 29486 16830 29538 16882
rect 30158 16830 30210 16882
rect 31054 16830 31106 16882
rect 31278 16830 31330 16882
rect 31950 16830 32002 16882
rect 32958 16830 33010 16882
rect 33182 16830 33234 16882
rect 6190 16718 6242 16770
rect 19070 16718 19122 16770
rect 19630 16718 19682 16770
rect 21534 16718 21586 16770
rect 25342 16718 25394 16770
rect 27246 16718 27298 16770
rect 15710 16606 15762 16658
rect 30886 16606 30938 16658
rect 33462 16606 33514 16658
rect 5372 16438 5424 16490
rect 5476 16438 5528 16490
rect 5580 16438 5632 16490
rect 13688 16438 13740 16490
rect 13792 16438 13844 16490
rect 13896 16438 13948 16490
rect 22004 16438 22056 16490
rect 22108 16438 22160 16490
rect 22212 16438 22264 16490
rect 30320 16438 30372 16490
rect 30424 16438 30476 16490
rect 30528 16438 30580 16490
rect 19854 16270 19906 16322
rect 26294 16270 26346 16322
rect 32846 16270 32898 16322
rect 33462 16270 33514 16322
rect 4510 16158 4562 16210
rect 10558 16158 10610 16210
rect 14254 16158 14306 16210
rect 16158 16158 16210 16210
rect 19294 16158 19346 16210
rect 22318 16158 22370 16210
rect 24222 16158 24274 16210
rect 27358 16158 27410 16210
rect 29318 16158 29370 16210
rect 31222 16158 31274 16210
rect 32286 16158 32338 16210
rect 1822 16046 1874 16098
rect 2606 16046 2658 16098
rect 5126 16046 5178 16098
rect 7870 16046 7922 16098
rect 8654 16046 8706 16098
rect 16942 16046 16994 16098
rect 18846 16046 18898 16098
rect 19126 16016 19178 16068
rect 19518 16046 19570 16098
rect 21534 16046 21586 16098
rect 26126 16046 26178 16098
rect 26910 16018 26962 16070
rect 27134 16046 27186 16098
rect 27526 15990 27578 16042
rect 27806 16046 27858 16098
rect 27974 16046 28026 16098
rect 31614 16102 31666 16154
rect 32454 16102 32506 16154
rect 28254 16046 28306 16098
rect 31838 16018 31890 16070
rect 28142 15934 28194 15986
rect 28534 15934 28586 15986
rect 11174 15822 11226 15874
rect 12518 15822 12570 15874
rect 24838 15822 24890 15874
rect 9530 15654 9582 15706
rect 9634 15654 9686 15706
rect 9738 15654 9790 15706
rect 17846 15654 17898 15706
rect 17950 15654 18002 15706
rect 18054 15654 18106 15706
rect 26162 15654 26214 15706
rect 26266 15654 26318 15706
rect 26370 15654 26422 15706
rect 34478 15654 34530 15706
rect 34582 15654 34634 15706
rect 34686 15654 34738 15706
rect 4902 15486 4954 15538
rect 12518 15486 12570 15538
rect 17838 15486 17890 15538
rect 4286 15374 4338 15426
rect 6302 15374 6354 15426
rect 14814 15374 14866 15426
rect 1598 15262 1650 15314
rect 8990 15262 9042 15314
rect 9774 15262 9826 15314
rect 12014 15289 12066 15341
rect 14646 15318 14698 15370
rect 15206 15374 15258 15426
rect 18342 15430 18394 15482
rect 28926 15486 28978 15538
rect 30494 15486 30546 15538
rect 21758 15374 21810 15426
rect 14478 15262 14530 15314
rect 14926 15262 14978 15314
rect 16382 15262 16434 15314
rect 28198 15318 28250 15370
rect 17502 15262 17554 15314
rect 18510 15262 18562 15314
rect 19070 15262 19122 15314
rect 19854 15262 19906 15314
rect 27246 15262 27298 15314
rect 27582 15262 27634 15314
rect 28478 15262 28530 15314
rect 29262 15262 29314 15314
rect 30158 15262 30210 15314
rect 31614 15262 31666 15314
rect 31726 15262 31778 15314
rect 2382 15150 2434 15202
rect 8206 15150 8258 15202
rect 16718 15150 16770 15202
rect 22374 15150 22426 15202
rect 28030 15150 28082 15202
rect 27358 15094 27410 15146
rect 32006 15038 32058 15090
rect 5372 14870 5424 14922
rect 5476 14870 5528 14922
rect 5580 14870 5632 14922
rect 13688 14870 13740 14922
rect 13792 14870 13844 14922
rect 13896 14870 13948 14922
rect 22004 14870 22056 14922
rect 22108 14870 22160 14922
rect 22212 14870 22264 14922
rect 30320 14870 30372 14922
rect 30424 14870 30476 14922
rect 30528 14870 30580 14922
rect 3054 14702 3106 14754
rect 6750 14702 6802 14754
rect 7310 14702 7362 14754
rect 31166 14590 31218 14642
rect 3390 14478 3442 14530
rect 6414 14478 6466 14530
rect 7646 14478 7698 14530
rect 7870 14478 7922 14530
rect 11454 14478 11506 14530
rect 12238 14478 12290 14530
rect 17838 14478 17890 14530
rect 26033 14478 26085 14530
rect 26910 14478 26962 14530
rect 27694 14478 27746 14530
rect 28030 14451 28082 14503
rect 28366 14478 28418 14530
rect 29150 14478 29202 14530
rect 29262 14478 29314 14530
rect 29542 14478 29594 14530
rect 30438 14478 30490 14530
rect 30718 14478 30770 14530
rect 31054 14434 31106 14486
rect 33518 14478 33570 14530
rect 34302 14478 34354 14530
rect 9550 14366 9602 14418
rect 25790 14366 25842 14418
rect 31614 14366 31666 14418
rect 14646 14254 14698 14306
rect 28254 14310 28306 14362
rect 18174 14254 18226 14306
rect 9530 14086 9582 14138
rect 9634 14086 9686 14138
rect 9738 14086 9790 14138
rect 17846 14086 17898 14138
rect 17950 14086 18002 14138
rect 18054 14086 18106 14138
rect 26162 14086 26214 14138
rect 26266 14086 26318 14138
rect 26370 14086 26422 14138
rect 34478 14086 34530 14138
rect 34582 14086 34634 14138
rect 34686 14086 34738 14138
rect 9046 13918 9098 13970
rect 9718 13918 9770 13970
rect 15150 13918 15202 13970
rect 22934 13918 22986 13970
rect 29878 13918 29930 13970
rect 30326 13918 30378 13970
rect 33294 13918 33346 13970
rect 31054 13862 31106 13914
rect 17838 13806 17890 13858
rect 2942 13694 2994 13746
rect 3614 13750 3666 13802
rect 3054 13694 3106 13746
rect 3838 13694 3890 13746
rect 4062 13582 4114 13634
rect 4230 13638 4282 13690
rect 4846 13694 4898 13746
rect 5182 13732 5234 13784
rect 11790 13694 11842 13746
rect 4454 13638 4506 13690
rect 14814 13694 14866 13746
rect 16382 13694 16434 13746
rect 16494 13694 16546 13746
rect 16662 13694 16714 13746
rect 16830 13694 16882 13746
rect 17726 13694 17778 13746
rect 18006 13694 18058 13746
rect 18174 13694 18226 13746
rect 18846 13694 18898 13746
rect 18958 13694 19010 13746
rect 21086 13694 21138 13746
rect 21310 13694 21362 13746
rect 21590 13694 21642 13746
rect 21870 13694 21922 13746
rect 23214 13694 23266 13746
rect 23550 13694 23602 13746
rect 25342 13738 25394 13790
rect 25678 13694 25730 13746
rect 26126 13694 26178 13746
rect 26462 13694 26514 13746
rect 26574 13694 26626 13746
rect 30942 13694 30994 13746
rect 31222 13723 31274 13775
rect 31950 13750 32002 13802
rect 31726 13694 31778 13746
rect 32286 13694 32338 13746
rect 32958 13694 33010 13746
rect 4622 13582 4674 13634
rect 12574 13582 12626 13634
rect 14478 13582 14530 13634
rect 24166 13582 24218 13634
rect 25230 13582 25282 13634
rect 27358 13582 27410 13634
rect 29262 13582 29314 13634
rect 31950 13582 32002 13634
rect 2662 13470 2714 13522
rect 16102 13470 16154 13522
rect 23326 13526 23378 13578
rect 17446 13470 17498 13522
rect 18566 13470 18618 13522
rect 22206 13470 22258 13522
rect 5372 13302 5424 13354
rect 5476 13302 5528 13354
rect 5580 13302 5632 13354
rect 13688 13302 13740 13354
rect 13792 13302 13844 13354
rect 13896 13302 13948 13354
rect 22004 13302 22056 13354
rect 22108 13302 22160 13354
rect 22212 13302 22264 13354
rect 30320 13302 30372 13354
rect 30424 13302 30476 13354
rect 30528 13302 30580 13354
rect 2718 13078 2770 13130
rect 3614 13022 3666 13074
rect 4622 13078 4674 13130
rect 6470 13134 6522 13186
rect 7646 13078 7698 13130
rect 5630 13022 5682 13074
rect 9774 13022 9826 13074
rect 11006 13078 11058 13130
rect 22654 13134 22706 13186
rect 26966 13134 27018 13186
rect 27694 13134 27746 13186
rect 29374 13134 29426 13186
rect 15822 13022 15874 13074
rect 17502 13022 17554 13074
rect 23886 13022 23938 13074
rect 25790 13022 25842 13074
rect 33070 13022 33122 13074
rect 2382 12910 2434 12962
rect 2606 12910 2658 12962
rect 3054 12910 3106 12962
rect 3390 12910 3442 12962
rect 3838 12910 3890 12962
rect 4286 12910 4338 12962
rect 4734 12910 4786 12962
rect 5070 12910 5122 12962
rect 5742 12895 5794 12947
rect 5966 12910 6018 12962
rect 6750 12854 6802 12906
rect 6974 12882 7026 12934
rect 7198 12854 7250 12906
rect 7366 12875 7418 12927
rect 7758 12910 7810 12962
rect 8434 12872 8486 12924
rect 10166 12910 10218 12962
rect 10334 12910 10386 12962
rect 10446 12910 10498 12962
rect 11118 12910 11170 12962
rect 11342 12910 11394 12962
rect 12014 12910 12066 12962
rect 13358 12910 13410 12962
rect 14366 12910 14418 12962
rect 15038 12910 15090 12962
rect 15598 12910 15650 12962
rect 15934 12883 15986 12935
rect 16270 12910 16322 12962
rect 16606 12910 16658 12962
rect 18062 12910 18114 12962
rect 18174 12910 18226 12962
rect 17894 12854 17946 12906
rect 18510 12910 18562 12962
rect 18846 12910 18898 12962
rect 18958 12910 19010 12962
rect 19518 12910 19570 12962
rect 21534 12910 21586 12962
rect 22410 12910 22462 12962
rect 23102 12910 23154 12962
rect 18678 12854 18730 12906
rect 26462 12910 26514 12962
rect 26686 12910 26738 12962
rect 28030 12910 28082 12962
rect 28702 12910 28754 12962
rect 29038 12910 29090 12962
rect 29934 12910 29986 12962
rect 30270 12910 30322 12962
rect 30382 12910 30434 12962
rect 31166 12910 31218 12962
rect 33630 12895 33682 12947
rect 33854 12910 33906 12962
rect 13694 12686 13746 12738
rect 14198 12686 14250 12738
rect 14870 12686 14922 12738
rect 15206 12742 15258 12794
rect 19238 12798 19290 12850
rect 19686 12742 19738 12794
rect 28366 12686 28418 12738
rect 33630 12742 33682 12794
rect 9530 12518 9582 12570
rect 9634 12518 9686 12570
rect 9738 12518 9790 12570
rect 17846 12518 17898 12570
rect 17950 12518 18002 12570
rect 18054 12518 18106 12570
rect 26162 12518 26214 12570
rect 26266 12518 26318 12570
rect 26370 12518 26422 12570
rect 34478 12518 34530 12570
rect 34582 12518 34634 12570
rect 34686 12518 34738 12570
rect 15318 12350 15370 12402
rect 2830 12238 2882 12290
rect 6974 12238 7026 12290
rect 2662 12126 2714 12178
rect 3054 12126 3106 12178
rect 3278 12154 3330 12206
rect 4006 12182 4058 12234
rect 3838 12126 3890 12178
rect 6302 12182 6354 12234
rect 6526 12182 6578 12234
rect 8766 12238 8818 12290
rect 10782 12238 10834 12290
rect 17502 12294 17554 12346
rect 31278 12294 31330 12346
rect 16494 12238 16546 12290
rect 4510 12126 4562 12178
rect 5294 12126 5346 12178
rect 5518 12126 5570 12178
rect 7534 12159 7586 12211
rect 7982 12162 8034 12214
rect 8318 12159 8370 12211
rect 8628 12159 8680 12211
rect 10334 12154 10386 12206
rect 10558 12126 10610 12178
rect 10950 12126 11002 12178
rect 11756 12163 11808 12215
rect 11902 12126 11954 12178
rect 12014 12126 12066 12178
rect 12462 12153 12514 12205
rect 16662 12182 16714 12234
rect 14590 12126 14642 12178
rect 16382 12126 16434 12178
rect 4752 12014 4804 12066
rect 7142 12070 7194 12122
rect 17726 12182 17778 12234
rect 24222 12182 24274 12234
rect 16830 12126 16882 12178
rect 17390 12126 17442 12178
rect 18062 12126 18114 12178
rect 18622 12126 18674 12178
rect 18958 12126 19010 12178
rect 21870 12126 21922 12178
rect 22654 12126 22706 12178
rect 22878 12126 22930 12178
rect 23774 12126 23826 12178
rect 24446 12126 24498 12178
rect 25454 12153 25506 12205
rect 28030 12153 28082 12205
rect 31614 12182 31666 12234
rect 30270 12126 30322 12178
rect 31166 12126 31218 12178
rect 31838 12126 31890 12178
rect 5182 11958 5234 12010
rect 11342 12014 11394 12066
rect 19966 12014 20018 12066
rect 23886 12014 23938 12066
rect 18734 11958 18786 12010
rect 16102 11902 16154 11954
rect 26238 11902 26290 11954
rect 5372 11734 5424 11786
rect 5476 11734 5528 11786
rect 5580 11734 5632 11786
rect 13688 11734 13740 11786
rect 13792 11734 13844 11786
rect 13896 11734 13948 11786
rect 22004 11734 22056 11786
rect 22108 11734 22160 11786
rect 22212 11734 22264 11786
rect 30320 11734 30372 11786
rect 30424 11734 30476 11786
rect 30528 11734 30580 11786
rect 3558 11566 3610 11618
rect 11902 11566 11954 11618
rect 12574 11566 12626 11618
rect 14982 11566 15034 11618
rect 16046 11510 16098 11562
rect 18734 11566 18786 11618
rect 32006 11566 32058 11618
rect 24334 11454 24386 11506
rect 25342 11454 25394 11506
rect 29318 11454 29370 11506
rect 3838 11342 3890 11394
rect 4118 11398 4170 11450
rect 29766 11454 29818 11506
rect 30214 11454 30266 11506
rect 32734 11454 32786 11506
rect 4286 11342 4338 11394
rect 6974 11307 7026 11359
rect 7086 11286 7138 11338
rect 7310 11314 7362 11366
rect 9102 11342 9154 11394
rect 7534 11286 7586 11338
rect 9326 11303 9378 11355
rect 9662 11342 9714 11394
rect 10558 11342 10610 11394
rect 11230 11342 11282 11394
rect 11454 11342 11506 11394
rect 12238 11342 12290 11394
rect 12910 11342 12962 11394
rect 13694 11342 13746 11394
rect 14478 11342 14530 11394
rect 15262 11342 15314 11394
rect 15542 11342 15594 11394
rect 15710 11342 15762 11394
rect 16102 11342 16154 11394
rect 16898 11304 16950 11356
rect 17670 11342 17722 11394
rect 17950 11342 18002 11394
rect 18062 11342 18114 11394
rect 19070 11342 19122 11394
rect 22430 11342 22482 11394
rect 25118 11342 25170 11394
rect 3950 11230 4002 11282
rect 25454 11298 25506 11350
rect 25790 11342 25842 11394
rect 26742 11342 26794 11394
rect 27470 11342 27522 11394
rect 27582 11342 27634 11394
rect 32286 11342 32338 11394
rect 32398 11342 32450 11394
rect 33182 11342 33234 11394
rect 32902 11286 32954 11338
rect 7814 11230 7866 11282
rect 10950 11230 11002 11282
rect 15374 11230 15426 11282
rect 9214 11174 9266 11226
rect 3222 11118 3274 11170
rect 10222 11118 10274 11170
rect 13526 11118 13578 11170
rect 14142 11118 14194 11170
rect 22038 11118 22090 11170
rect 26294 11118 26346 11170
rect 27134 11118 27186 11170
rect 9530 10950 9582 11002
rect 9634 10950 9686 11002
rect 9738 10950 9790 11002
rect 17846 10950 17898 11002
rect 17950 10950 18002 11002
rect 18054 10950 18106 11002
rect 26162 10950 26214 11002
rect 26266 10950 26318 11002
rect 26370 10950 26422 11002
rect 34478 10950 34530 11002
rect 34582 10950 34634 11002
rect 34686 10950 34738 11002
rect 15374 10782 15426 10834
rect 15822 10782 15874 10834
rect 24726 10782 24778 10834
rect 4734 10670 4786 10722
rect 7590 10670 7642 10722
rect 31950 10726 32002 10778
rect 33462 10670 33514 10722
rect 3054 10558 3106 10610
rect 3614 10558 3666 10610
rect 3838 10558 3890 10610
rect 4510 10558 4562 10610
rect 4872 10591 4924 10643
rect 5182 10614 5234 10666
rect 5630 10591 5682 10643
rect 5854 10614 5906 10666
rect 8150 10614 8202 10666
rect 7870 10558 7922 10610
rect 7982 10558 8034 10610
rect 8318 10558 8370 10610
rect 10110 10558 10162 10610
rect 12014 10558 12066 10610
rect 12798 10602 12850 10654
rect 13134 10558 13186 10610
rect 13918 10558 13970 10610
rect 14702 10558 14754 10610
rect 14814 10558 14866 10610
rect 21310 10558 21362 10610
rect 23121 10558 23173 10610
rect 23998 10558 24050 10610
rect 25342 10573 25394 10625
rect 25678 10558 25730 10610
rect 25902 10558 25954 10610
rect 26686 10558 26738 10610
rect 29262 10558 29314 10610
rect 29598 10558 29650 10610
rect 29822 10597 29874 10649
rect 30270 10558 30322 10610
rect 30942 10573 30994 10625
rect 32062 10614 32114 10666
rect 31278 10558 31330 10610
rect 31726 10558 31778 10610
rect 32286 10558 32338 10610
rect 32958 10558 33010 10610
rect 33182 10558 33234 10610
rect 12686 10446 12738 10498
rect 25230 10446 25282 10498
rect 28590 10446 28642 10498
rect 29934 10446 29986 10498
rect 30830 10446 30882 10498
rect 2718 10334 2770 10386
rect 3334 10334 3386 10386
rect 4174 10334 4226 10386
rect 9774 10334 9826 10386
rect 12182 10390 12234 10442
rect 13582 10334 13634 10386
rect 14422 10334 14474 10386
rect 20974 10334 21026 10386
rect 22878 10334 22930 10386
rect 5372 10166 5424 10218
rect 5476 10166 5528 10218
rect 5580 10166 5632 10218
rect 13688 10166 13740 10218
rect 13792 10166 13844 10218
rect 13896 10166 13948 10218
rect 22004 10166 22056 10218
rect 22108 10166 22160 10218
rect 22212 10166 22264 10218
rect 30320 10166 30372 10218
rect 30424 10166 30476 10218
rect 30528 10166 30580 10218
rect 3110 9998 3162 10050
rect 8038 9998 8090 10050
rect 4734 9942 4786 9994
rect 5742 9942 5794 9994
rect 10558 9942 10610 9994
rect 27302 9998 27354 10050
rect 13582 9886 13634 9938
rect 14422 9886 14474 9938
rect 16046 9886 16098 9938
rect 17838 9886 17890 9938
rect 19742 9886 19794 9938
rect 23942 9886 23994 9938
rect 25678 9886 25730 9938
rect 30382 9886 30434 9938
rect 34078 9886 34130 9938
rect 3390 9718 3442 9770
rect 3558 9739 3610 9791
rect 3838 9746 3890 9798
rect 4006 9758 4058 9810
rect 4286 9774 4338 9826
rect 4622 9774 4674 9826
rect 5742 9774 5794 9826
rect 5966 9774 6018 9826
rect 7086 9774 7138 9826
rect 7310 9774 7362 9826
rect 8318 9774 8370 9826
rect 8430 9774 8482 9826
rect 10670 9774 10722 9826
rect 10894 9774 10946 9826
rect 11398 9774 11450 9826
rect 11678 9774 11730 9826
rect 11790 9774 11842 9826
rect 12462 9774 12514 9826
rect 12686 9774 12738 9826
rect 15710 9774 15762 9826
rect 15934 9735 15986 9787
rect 16382 9774 16434 9826
rect 17054 9774 17106 9826
rect 21870 9730 21922 9782
rect 22206 9774 22258 9826
rect 22766 9774 22818 9826
rect 23102 9747 23154 9799
rect 23326 9774 23378 9826
rect 24782 9774 24834 9826
rect 25566 9774 25618 9826
rect 26014 9735 26066 9787
rect 26238 9774 26290 9826
rect 26574 9774 26626 9826
rect 27470 9774 27522 9826
rect 27806 9774 27858 9826
rect 28366 9774 28418 9826
rect 27974 9718 28026 9770
rect 29374 9774 29426 9826
rect 29598 9735 29650 9787
rect 29934 9774 29986 9826
rect 30494 9730 30546 9782
rect 30718 9774 30770 9826
rect 31390 9774 31442 9826
rect 32174 9774 32226 9826
rect 7590 9662 7642 9714
rect 12182 9662 12234 9714
rect 21982 9606 22034 9658
rect 22654 9606 22706 9658
rect 2774 9550 2826 9602
rect 28478 9606 28530 9658
rect 29262 9606 29314 9658
rect 25118 9550 25170 9602
rect 9530 9382 9582 9434
rect 9634 9382 9686 9434
rect 9738 9382 9790 9434
rect 17846 9382 17898 9434
rect 17950 9382 18002 9434
rect 18054 9382 18106 9434
rect 26162 9382 26214 9434
rect 26266 9382 26318 9434
rect 26370 9382 26422 9434
rect 34478 9382 34530 9434
rect 34582 9382 34634 9434
rect 34686 9382 34738 9434
rect 33294 9214 33346 9266
rect 3054 9018 3106 9070
rect 3670 9046 3722 9098
rect 3278 8990 3330 9042
rect 4174 9005 4226 9057
rect 6078 9046 6130 9098
rect 4510 8990 4562 9042
rect 6302 8990 6354 9042
rect 6526 8990 6578 9042
rect 6694 9046 6746 9098
rect 23046 9102 23098 9154
rect 7310 9028 7362 9080
rect 8038 9046 8090 9098
rect 7646 8990 7698 9042
rect 8430 8990 8482 9042
rect 8654 8990 8706 9042
rect 11118 8990 11170 9042
rect 12462 8990 12514 9042
rect 12686 8990 12738 9042
rect 13436 9027 13488 9079
rect 13582 8990 13634 9042
rect 13694 8990 13746 9042
rect 14198 8990 14250 9042
rect 15598 9046 15650 9098
rect 14366 8990 14418 9042
rect 15150 8990 15202 9042
rect 15822 8990 15874 9042
rect 19518 8990 19570 9042
rect 20302 8990 20354 9042
rect 22654 8990 22706 9042
rect 22766 8990 22818 9042
rect 25342 8990 25394 9042
rect 25566 9005 25618 9057
rect 28030 8990 28082 9042
rect 28254 9005 28306 9057
rect 28926 9018 28978 9070
rect 29150 8990 29202 9042
rect 3502 8878 3554 8930
rect 4062 8878 4114 8930
rect 7870 8878 7922 8930
rect 8318 8822 8370 8874
rect 13022 8878 13074 8930
rect 15262 8878 15314 8930
rect 22206 8878 22258 8930
rect 23606 8878 23658 8930
rect 25678 8878 25730 8930
rect 28366 8878 28418 8930
rect 29374 8878 29426 8930
rect 29542 8934 29594 8986
rect 29710 8990 29762 9042
rect 32958 8990 33010 9042
rect 30494 8878 30546 8930
rect 32398 8878 32450 8930
rect 11286 8766 11338 8818
rect 12182 8766 12234 8818
rect 14702 8766 14754 8818
rect 5372 8598 5424 8650
rect 5476 8598 5528 8650
rect 5580 8598 5632 8650
rect 13688 8598 13740 8650
rect 13792 8598 13844 8650
rect 13896 8598 13948 8650
rect 22004 8598 22056 8650
rect 22108 8598 22160 8650
rect 22212 8598 22264 8650
rect 30320 8598 30372 8650
rect 30424 8598 30476 8650
rect 30528 8598 30580 8650
rect 29542 8430 29594 8482
rect 31894 8430 31946 8482
rect 4174 8374 4226 8426
rect 3894 8262 3946 8314
rect 7086 8318 7138 8370
rect 9550 8318 9602 8370
rect 13918 8318 13970 8370
rect 15150 8318 15202 8370
rect 18958 8318 19010 8370
rect 21310 8318 21362 8370
rect 22766 8318 22818 8370
rect 28478 8318 28530 8370
rect 30102 8318 30154 8370
rect 3054 8150 3106 8202
rect 3278 8178 3330 8230
rect 4286 8206 4338 8258
rect 4510 8206 4562 8258
rect 7422 8206 7474 8258
rect 7870 8206 7922 8258
rect 8206 8206 8258 8258
rect 8430 8206 8482 8258
rect 8654 8206 8706 8258
rect 9102 8206 9154 8258
rect 9438 8206 9490 8258
rect 10110 8206 10162 8258
rect 9774 8150 9826 8202
rect 11566 8206 11618 8258
rect 13582 8206 13634 8258
rect 11118 8150 11170 8202
rect 12126 8150 12178 8202
rect 12574 8150 12626 8202
rect 13806 8162 13858 8214
rect 15486 8150 15538 8202
rect 15598 8206 15650 8258
rect 15934 8206 15986 8258
rect 16270 8206 16322 8258
rect 17054 8206 17106 8258
rect 21422 8162 21474 8214
rect 21758 8206 21810 8258
rect 22430 8206 22482 8258
rect 23102 8206 23154 8258
rect 22766 8150 22818 8202
rect 23438 8206 23490 8258
rect 24110 8162 24162 8214
rect 24334 8206 24386 8258
rect 27918 8206 27970 8258
rect 28142 8206 28194 8258
rect 29038 8206 29090 8258
rect 29262 8206 29314 8258
rect 32062 8206 32114 8258
rect 3726 8094 3778 8146
rect 24222 8038 24274 8090
rect 27582 7982 27634 8034
rect 31222 7982 31274 8034
rect 9530 7814 9582 7866
rect 9634 7814 9686 7866
rect 9738 7814 9790 7866
rect 17846 7814 17898 7866
rect 17950 7814 18002 7866
rect 18054 7814 18106 7866
rect 26162 7814 26214 7866
rect 26266 7814 26318 7866
rect 26370 7814 26422 7866
rect 34478 7814 34530 7866
rect 34582 7814 34634 7866
rect 34686 7814 34738 7866
rect 4510 7646 4562 7698
rect 4734 7646 4786 7698
rect 11566 7590 11618 7642
rect 7366 7534 7418 7586
rect 14870 7534 14922 7586
rect 3166 7422 3218 7474
rect 3726 7422 3778 7474
rect 4286 7422 4338 7474
rect 4622 7422 4674 7474
rect 7646 7422 7698 7474
rect 7870 7422 7922 7474
rect 10392 7422 10444 7474
rect 10558 7422 10610 7474
rect 10670 7422 10722 7474
rect 11454 7422 11506 7474
rect 11678 7461 11730 7513
rect 12014 7422 12066 7474
rect 12462 7422 12514 7474
rect 12630 7422 12682 7474
rect 12798 7422 12850 7474
rect 12910 7422 12962 7474
rect 14030 7457 14082 7509
rect 14198 7457 14250 7509
rect 14366 7450 14418 7502
rect 14590 7478 14642 7530
rect 22094 7534 22146 7586
rect 23214 7534 23266 7586
rect 29766 7534 29818 7586
rect 15766 7422 15818 7474
rect 15934 7422 15986 7474
rect 16046 7422 16098 7474
rect 23046 7478 23098 7530
rect 19406 7422 19458 7474
rect 20190 7422 20242 7474
rect 22878 7422 22930 7474
rect 23326 7422 23378 7474
rect 23606 7422 23658 7474
rect 24110 7422 24162 7474
rect 24446 7422 24498 7474
rect 26910 7422 26962 7474
rect 27302 7451 27354 7503
rect 29262 7422 29314 7474
rect 29486 7422 29538 7474
rect 31614 7422 31666 7474
rect 31950 7437 32002 7489
rect 32958 7422 33010 7474
rect 9998 7310 10050 7362
rect 2942 7254 2994 7306
rect 27358 7310 27410 7362
rect 32062 7310 32114 7362
rect 13190 7198 13242 7250
rect 15374 7198 15426 7250
rect 23998 7254 24050 7306
rect 33294 7198 33346 7250
rect 5372 7030 5424 7082
rect 5476 7030 5528 7082
rect 5580 7030 5632 7082
rect 13688 7030 13740 7082
rect 13792 7030 13844 7082
rect 13896 7030 13948 7082
rect 22004 7030 22056 7082
rect 22108 7030 22160 7082
rect 22212 7030 22264 7082
rect 30320 7030 30372 7082
rect 30424 7030 30476 7082
rect 30528 7030 30580 7082
rect 5854 6862 5906 6914
rect 8654 6862 8706 6914
rect 11174 6862 11226 6914
rect 13862 6862 13914 6914
rect 15710 6862 15762 6914
rect 22206 6862 22258 6914
rect 17390 6806 17442 6858
rect 23886 6750 23938 6802
rect 25790 6750 25842 6802
rect 28030 6750 28082 6802
rect 32174 6750 32226 6802
rect 2774 6638 2826 6690
rect 3110 6638 3162 6690
rect 5070 6694 5122 6746
rect 3390 6610 3442 6662
rect 3614 6582 3666 6634
rect 3838 6582 3890 6634
rect 3950 6582 4002 6634
rect 4230 6638 4282 6690
rect 4958 6600 5010 6652
rect 5518 6638 5570 6690
rect 7870 6638 7922 6690
rect 8094 6638 8146 6690
rect 4398 6526 4450 6578
rect 7534 6582 7586 6634
rect 8262 6582 8314 6634
rect 8990 6638 9042 6690
rect 11454 6638 11506 6690
rect 11902 6638 11954 6690
rect 11734 6582 11786 6634
rect 13358 6638 13410 6690
rect 13582 6638 13634 6690
rect 14366 6638 14418 6690
rect 14590 6638 14642 6690
rect 15374 6638 15426 6690
rect 16606 6638 16658 6690
rect 17054 6638 17106 6690
rect 17278 6638 17330 6690
rect 17614 6638 17666 6690
rect 18006 6638 18058 6690
rect 18398 6638 18450 6690
rect 11566 6526 11618 6578
rect 14870 6526 14922 6578
rect 16270 6526 16322 6578
rect 18174 6526 18226 6578
rect 18734 6582 18786 6634
rect 22542 6638 22594 6690
rect 22934 6638 22986 6690
rect 23102 6638 23154 6690
rect 26406 6638 26458 6690
rect 28142 6594 28194 6646
rect 28478 6638 28530 6690
rect 29486 6638 29538 6690
rect 30362 6638 30414 6690
rect 31390 6638 31442 6690
rect 34078 6638 34130 6690
rect 29038 6526 29090 6578
rect 29262 6526 29314 6578
rect 30606 6526 30658 6578
rect 12350 6414 12402 6466
rect 12742 6414 12794 6466
rect 16886 6414 16938 6466
rect 31222 6414 31274 6466
rect 9530 6246 9582 6298
rect 9634 6246 9686 6298
rect 9738 6246 9790 6298
rect 17846 6246 17898 6298
rect 17950 6246 18002 6298
rect 18054 6246 18106 6298
rect 26162 6246 26214 6298
rect 26266 6246 26318 6298
rect 26370 6246 26422 6298
rect 34478 6246 34530 6298
rect 34582 6246 34634 6298
rect 34686 6246 34738 6298
rect 10670 6078 10722 6130
rect 12014 6078 12066 6130
rect 3110 5966 3162 6018
rect 5238 5966 5290 6018
rect 7086 5966 7138 6018
rect 3390 5910 3442 5962
rect 3614 5910 3666 5962
rect 3838 5910 3890 5962
rect 8000 5966 8052 6018
rect 2830 5854 2882 5906
rect 3950 5889 4002 5941
rect 4734 5854 4786 5906
rect 4958 5854 5010 5906
rect 7254 5910 7306 5962
rect 12910 5966 12962 6018
rect 13302 5966 13354 6018
rect 14870 6022 14922 6074
rect 15598 6078 15650 6130
rect 25286 6078 25338 6130
rect 16438 5966 16490 6018
rect 19518 5966 19570 6018
rect 23886 6022 23938 6074
rect 25958 6078 26010 6130
rect 19910 5966 19962 6018
rect 32286 6022 32338 6074
rect 28814 5966 28866 6018
rect 33126 5966 33178 6018
rect 6248 5854 6300 5906
rect 6414 5854 6466 5906
rect 6526 5854 6578 5906
rect 7758 5854 7810 5906
rect 11006 5854 11058 5906
rect 11230 5854 11282 5906
rect 11678 5854 11730 5906
rect 12574 5854 12626 5906
rect 12742 5854 12794 5906
rect 13022 5854 13074 5906
rect 15038 5854 15090 5906
rect 15934 5854 15986 5906
rect 16718 5854 16770 5906
rect 16830 5854 16882 5906
rect 17278 5854 17330 5906
rect 18174 5854 18226 5906
rect 18914 5892 18966 5944
rect 19182 5854 19234 5906
rect 5854 5742 5906 5794
rect 19350 5798 19402 5850
rect 19630 5854 19682 5906
rect 22318 5854 22370 5906
rect 22654 5898 22706 5950
rect 23438 5910 23490 5962
rect 23214 5854 23266 5906
rect 23774 5854 23826 5906
rect 24222 5854 24274 5906
rect 25454 5854 25506 5906
rect 26126 5854 26178 5906
rect 26910 5854 26962 5906
rect 29486 5854 29538 5906
rect 30046 5910 30098 5962
rect 31838 5910 31890 5962
rect 29822 5854 29874 5906
rect 30382 5854 30434 5906
rect 31614 5854 31666 5906
rect 32174 5854 32226 5906
rect 33406 5854 33458 5906
rect 33630 5854 33682 5906
rect 22766 5742 22818 5794
rect 30158 5742 30210 5794
rect 2494 5630 2546 5682
rect 11398 5630 11450 5682
rect 17614 5630 17666 5682
rect 18062 5686 18114 5738
rect 30998 5742 31050 5794
rect 24558 5630 24610 5682
rect 5372 5462 5424 5514
rect 5476 5462 5528 5514
rect 5580 5462 5632 5514
rect 13688 5462 13740 5514
rect 13792 5462 13844 5514
rect 13896 5462 13948 5514
rect 22004 5462 22056 5514
rect 22108 5462 22160 5514
rect 22212 5462 22264 5514
rect 30320 5462 30372 5514
rect 30424 5462 30476 5514
rect 30528 5462 30580 5514
rect 2774 5294 2826 5346
rect 3278 5294 3330 5346
rect 4286 5238 4338 5290
rect 4958 5238 5010 5290
rect 6414 5182 6466 5234
rect 7534 5182 7586 5234
rect 10110 5238 10162 5290
rect 12462 5294 12514 5346
rect 18958 5294 19010 5346
rect 21366 5294 21418 5346
rect 26350 5294 26402 5346
rect 29206 5294 29258 5346
rect 2942 5070 2994 5122
rect 3614 5070 3666 5122
rect 3838 5070 3890 5122
rect 4174 5070 4226 5122
rect 4734 5070 4786 5122
rect 4958 5070 5010 5122
rect 6808 5070 6860 5122
rect 6974 5070 7026 5122
rect 7086 5070 7138 5122
rect 7926 5070 7978 5122
rect 8094 5070 8146 5122
rect 8206 5070 8258 5122
rect 10222 5070 10274 5122
rect 10558 5070 10610 5122
rect 10988 5070 11040 5122
rect 11230 5070 11282 5122
rect 11734 5126 11786 5178
rect 13638 5182 13690 5234
rect 14590 5182 14642 5234
rect 18174 5182 18226 5234
rect 23774 5182 23826 5234
rect 27358 5182 27410 5234
rect 34078 5182 34130 5234
rect 12126 5070 12178 5122
rect 13806 5070 13858 5122
rect 16494 5070 16546 5122
rect 17838 5070 17890 5122
rect 18510 5070 18562 5122
rect 19350 5070 19402 5122
rect 19518 5070 19570 5122
rect 19630 5070 19682 5122
rect 18062 5014 18114 5066
rect 20414 5070 20466 5122
rect 21534 5070 21586 5122
rect 21758 5070 21810 5122
rect 22206 5031 22258 5083
rect 22430 5070 22482 5122
rect 22990 5070 23042 5122
rect 25678 5070 25730 5122
rect 26686 5070 26738 5122
rect 26910 5070 26962 5122
rect 27246 5055 27298 5107
rect 27806 5070 27858 5122
rect 28030 5043 28082 5095
rect 28366 5070 28418 5122
rect 29486 5070 29538 5122
rect 29598 5070 29650 5122
rect 30382 5070 30434 5122
rect 30942 5070 30994 5122
rect 30606 5014 30658 5066
rect 31390 5070 31442 5122
rect 32174 5070 32226 5122
rect 11566 4902 11618 4954
rect 21870 4902 21922 4954
rect 28366 4902 28418 4954
rect 31054 4902 31106 4954
rect 20078 4846 20130 4898
rect 9530 4678 9582 4730
rect 9634 4678 9686 4730
rect 9738 4678 9790 4730
rect 17846 4678 17898 4730
rect 17950 4678 18002 4730
rect 18054 4678 18106 4730
rect 26162 4678 26214 4730
rect 26266 4678 26318 4730
rect 26370 4678 26422 4730
rect 34478 4678 34530 4730
rect 34582 4678 34634 4730
rect 34686 4678 34738 4730
rect 10446 4510 10498 4562
rect 11118 4510 11170 4562
rect 29766 4510 29818 4562
rect 4286 4398 4338 4450
rect 7310 4398 7362 4450
rect 5610 4342 5662 4394
rect 16718 4398 16770 4450
rect 23438 4454 23490 4506
rect 33294 4510 33346 4562
rect 22318 4398 22370 4450
rect 29150 4398 29202 4450
rect 1598 4286 1650 4338
rect 2382 4286 2434 4338
rect 4734 4286 4786 4338
rect 7553 4286 7605 4338
rect 8430 4286 8482 4338
rect 9662 4286 9714 4338
rect 9998 4286 10050 4338
rect 10782 4286 10834 4338
rect 11454 4286 11506 4338
rect 11678 4286 11730 4338
rect 11790 4286 11842 4338
rect 11936 4324 11988 4376
rect 14030 4286 14082 4338
rect 14814 4286 14866 4338
rect 17838 4286 17890 4338
rect 18174 4286 18226 4338
rect 23326 4342 23378 4394
rect 19630 4286 19682 4338
rect 22990 4286 23042 4338
rect 23550 4286 23602 4338
rect 24222 4330 24274 4382
rect 24558 4286 24610 4338
rect 25118 4286 25170 4338
rect 26350 4286 26402 4338
rect 26462 4286 26514 4338
rect 32510 4313 32562 4365
rect 32958 4286 33010 4338
rect 12350 4174 12402 4226
rect 20414 4174 20466 4226
rect 24110 4174 24162 4226
rect 26014 4174 26066 4226
rect 27246 4174 27298 4226
rect 5854 4062 5906 4114
rect 25454 4062 25506 4114
rect 31502 4062 31554 4114
rect 5372 3894 5424 3946
rect 5476 3894 5528 3946
rect 5580 3894 5632 3946
rect 13688 3894 13740 3946
rect 13792 3894 13844 3946
rect 13896 3894 13948 3946
rect 22004 3894 22056 3946
rect 22108 3894 22160 3946
rect 22212 3894 22264 3946
rect 30320 3894 30372 3946
rect 30424 3894 30476 3946
rect 30528 3894 30580 3946
rect 4398 3670 4450 3722
rect 11230 3726 11282 3778
rect 21086 3726 21138 3778
rect 23494 3726 23546 3778
rect 28646 3726 28698 3778
rect 32566 3726 32618 3778
rect 33182 3726 33234 3778
rect 5686 3614 5738 3666
rect 22710 3614 22762 3666
rect 26350 3614 26402 3666
rect 30662 3614 30714 3666
rect 30942 3614 30994 3666
rect 4510 3502 4562 3554
rect 4846 3502 4898 3554
rect 10894 3502 10946 3554
rect 18174 3502 18226 3554
rect 20078 3474 20130 3526
rect 21422 3502 21474 3554
rect 23774 3502 23826 3554
rect 23998 3502 24050 3554
rect 25454 3474 25506 3526
rect 28926 3502 28978 3554
rect 29150 3502 29202 3554
rect 31054 3487 31106 3539
rect 31278 3502 31330 3554
rect 32062 3502 32114 3554
rect 32286 3502 32338 3554
rect 32846 3502 32898 3554
rect 6134 3390 6186 3442
rect 10726 3390 10778 3442
rect 9530 3110 9582 3162
rect 9634 3110 9686 3162
rect 9738 3110 9790 3162
rect 17846 3110 17898 3162
rect 17950 3110 18002 3162
rect 18054 3110 18106 3162
rect 26162 3110 26214 3162
rect 26266 3110 26318 3162
rect 26370 3110 26422 3162
rect 34478 3110 34530 3162
rect 34582 3110 34634 3162
rect 34686 3110 34738 3162
<< metal2 >>
rect 5370 32172 5634 32182
rect 5426 32116 5474 32172
rect 5530 32116 5578 32172
rect 5370 32106 5634 32116
rect 13686 32172 13950 32182
rect 13742 32116 13790 32172
rect 13846 32116 13894 32172
rect 13686 32106 13950 32116
rect 22002 32172 22266 32182
rect 22058 32116 22106 32172
rect 22162 32116 22210 32172
rect 22002 32106 22266 32116
rect 30318 32172 30582 32182
rect 30374 32116 30422 32172
rect 30478 32116 30526 32172
rect 30318 32106 30582 32116
rect 13132 31890 13188 31902
rect 13132 31838 13134 31890
rect 13186 31838 13188 31890
rect 9528 31388 9792 31398
rect 9584 31332 9632 31388
rect 9688 31332 9736 31388
rect 9528 31322 9792 31332
rect 13132 30994 13188 31838
rect 19628 31892 19684 31902
rect 19628 31798 19684 31836
rect 20524 31892 20580 31902
rect 13468 31778 13524 31790
rect 13300 31722 13356 31734
rect 13300 31670 13302 31722
rect 13354 31670 13356 31722
rect 13300 31668 13356 31670
rect 13468 31726 13470 31778
rect 13522 31726 13524 31778
rect 13300 31612 13412 31668
rect 13132 30942 13134 30994
rect 13186 30942 13188 30994
rect 13132 30930 13188 30942
rect 11228 30884 11284 30894
rect 11228 30882 11620 30884
rect 11228 30830 11230 30882
rect 11282 30830 11620 30882
rect 11228 30828 11620 30830
rect 11228 30818 11284 30828
rect 5370 30604 5634 30614
rect 5426 30548 5474 30604
rect 5530 30548 5578 30604
rect 5370 30538 5634 30548
rect 9660 30210 9716 30222
rect 9660 30158 9662 30210
rect 9714 30158 9716 30210
rect 9660 29988 9716 30158
rect 10444 30212 10500 30222
rect 10444 30118 10500 30156
rect 11564 30100 11620 30828
rect 11564 30034 11620 30044
rect 11676 30212 11732 30222
rect 13356 30212 13412 31612
rect 13468 30436 13524 31726
rect 16156 31780 16212 31790
rect 16156 31778 16324 31780
rect 16156 31726 16158 31778
rect 16210 31726 16324 31778
rect 16156 31724 16324 31726
rect 16156 31714 16212 31724
rect 14812 31556 14868 31566
rect 13916 30996 13972 31006
rect 14028 30996 14084 31006
rect 13916 30994 14084 30996
rect 13916 30942 13918 30994
rect 13970 30942 14030 30994
rect 14082 30942 14084 30994
rect 13916 30940 14084 30942
rect 13916 30930 13972 30940
rect 13686 30604 13950 30614
rect 13742 30548 13790 30604
rect 13846 30548 13894 30604
rect 13686 30538 13950 30548
rect 13468 30380 13748 30436
rect 13580 30212 13636 30222
rect 13356 30210 13636 30212
rect 13356 30158 13582 30210
rect 13634 30158 13636 30210
rect 13356 30156 13636 30158
rect 9660 29932 9940 29988
rect 9528 29820 9792 29830
rect 9584 29764 9632 29820
rect 9688 29764 9736 29820
rect 9528 29754 9792 29764
rect 5370 29036 5634 29046
rect 5426 28980 5474 29036
rect 5530 28980 5578 29036
rect 5370 28970 5634 28980
rect 9660 28644 9716 28654
rect 9884 28644 9940 29932
rect 11676 29314 11732 30156
rect 13580 30146 13636 30156
rect 12348 30098 12404 30110
rect 12348 30046 12350 30098
rect 12402 30046 12404 30098
rect 11788 29988 11844 29998
rect 11788 29470 11844 29932
rect 11788 29418 11790 29470
rect 11842 29418 11844 29470
rect 11788 29406 11844 29418
rect 12124 29426 12180 29438
rect 11676 29262 11678 29314
rect 11730 29262 11732 29314
rect 11676 29250 11732 29262
rect 12124 29374 12126 29426
rect 12178 29374 12180 29426
rect 12124 29316 12180 29374
rect 12124 29250 12180 29260
rect 12348 29316 12404 30046
rect 12964 29988 13020 29998
rect 13692 29988 13748 30380
rect 12964 29986 13076 29988
rect 12964 29934 12966 29986
rect 13018 29934 13076 29986
rect 12964 29922 13076 29934
rect 13692 29922 13748 29932
rect 13823 30154 13879 30166
rect 13823 30102 13825 30154
rect 13877 30102 13879 30154
rect 12796 29594 12852 29606
rect 12796 29542 12798 29594
rect 12850 29542 12852 29594
rect 12348 29250 12404 29260
rect 12684 29441 12740 29453
rect 12684 29428 12686 29441
rect 12738 29428 12740 29441
rect 12348 28756 12404 28766
rect 12684 28756 12740 29372
rect 12348 28754 12740 28756
rect 12348 28702 12350 28754
rect 12402 28702 12740 28754
rect 12348 28700 12740 28702
rect 12348 28690 12404 28700
rect 9660 28642 9940 28644
rect 9660 28590 9662 28642
rect 9714 28590 9940 28642
rect 9660 28588 9940 28590
rect 9660 28578 9716 28588
rect 9528 28252 9792 28262
rect 9584 28196 9632 28252
rect 9688 28196 9736 28252
rect 9528 28186 9792 28196
rect 8092 27858 8148 27870
rect 8092 27806 8094 27858
rect 8146 27806 8148 27858
rect 5370 27468 5634 27478
rect 5426 27412 5474 27468
rect 5530 27412 5578 27468
rect 5370 27402 5634 27412
rect 7308 27076 7364 27086
rect 7308 27074 7476 27076
rect 7308 27022 7310 27074
rect 7362 27022 7476 27074
rect 7308 27020 7476 27022
rect 7308 27010 7364 27020
rect 6076 26964 6132 26974
rect 5796 26852 5852 26862
rect 2268 26290 2324 26302
rect 2268 26238 2270 26290
rect 2322 26238 2324 26290
rect 1596 25506 1652 25518
rect 1596 25454 1598 25506
rect 1650 25454 1652 25506
rect 1596 25284 1652 25454
rect 1596 23154 1652 25228
rect 2268 25284 2324 26238
rect 4620 26292 4676 26302
rect 3052 26180 3108 26190
rect 3052 26086 3108 26124
rect 2380 25508 2436 25518
rect 2380 25506 2660 25508
rect 2380 25454 2382 25506
rect 2434 25454 2660 25506
rect 2380 25452 2660 25454
rect 2380 25442 2436 25452
rect 2268 25218 2324 25228
rect 2604 24948 2660 25452
rect 4284 25394 4340 25406
rect 4284 25342 4286 25394
rect 4338 25342 4340 25394
rect 2716 24948 2772 24958
rect 2604 24946 2772 24948
rect 2604 24894 2718 24946
rect 2770 24894 2772 24946
rect 2604 24892 2772 24894
rect 2716 24882 2772 24892
rect 3052 24722 3108 24734
rect 4284 24724 4340 25342
rect 4620 25284 4676 26236
rect 5292 26292 5348 26302
rect 5292 26198 5348 26236
rect 5796 26292 5852 26796
rect 4844 26180 4900 26190
rect 4844 25730 4900 26124
rect 4844 25678 4846 25730
rect 4898 25678 4900 25730
rect 4844 25666 4900 25678
rect 4956 26178 5012 26190
rect 4956 26126 4958 26178
rect 5010 26126 5012 26178
rect 3052 24670 3054 24722
rect 3106 24670 3108 24722
rect 3052 24164 3108 24670
rect 3052 24098 3108 24108
rect 3948 24668 4340 24724
rect 4396 24836 4452 24846
rect 4396 24722 4452 24780
rect 4396 24670 4398 24722
rect 4450 24670 4452 24722
rect 3836 23938 3892 23950
rect 3836 23886 3838 23938
rect 3890 23886 3892 23938
rect 3556 23828 3612 23838
rect 1596 23102 1598 23154
rect 1650 23102 1652 23154
rect 1596 23090 1652 23102
rect 3500 23826 3612 23828
rect 3500 23774 3558 23826
rect 3610 23774 3612 23826
rect 3500 23762 3612 23774
rect 2380 23044 2436 23054
rect 2380 23042 2660 23044
rect 2380 22990 2382 23042
rect 2434 22990 2660 23042
rect 2380 22988 2660 22990
rect 2380 22978 2436 22988
rect 2604 22596 2660 22988
rect 2716 22596 2772 22606
rect 2604 22594 2772 22596
rect 2604 22542 2718 22594
rect 2770 22542 2772 22594
rect 2604 22540 2772 22542
rect 2716 22530 2772 22540
rect 3388 22484 3444 22494
rect 3500 22484 3556 23762
rect 3444 22428 3556 22484
rect 3612 23492 3668 23502
rect 3388 22418 3444 22428
rect 3052 22372 3108 22382
rect 3052 22278 3108 22316
rect 3612 21588 3668 23436
rect 3836 23492 3892 23886
rect 3948 23938 4004 24668
rect 4396 24658 4452 24670
rect 4508 24722 4564 24734
rect 4508 24670 4510 24722
rect 4562 24670 4564 24722
rect 4116 24500 4172 24510
rect 3948 23886 3950 23938
rect 4002 23886 4004 23938
rect 3948 23604 4004 23886
rect 3948 23538 4004 23548
rect 4060 24498 4172 24500
rect 4060 24446 4118 24498
rect 4170 24446 4172 24498
rect 4060 24434 4172 24446
rect 3836 23426 3892 23436
rect 4060 23268 4116 24434
rect 4508 24388 4564 24670
rect 4228 24332 4564 24388
rect 4228 24276 4284 24332
rect 3724 23212 4116 23268
rect 4172 24220 4284 24276
rect 4172 23268 4228 24220
rect 4340 24164 4396 24174
rect 4620 24164 4676 25228
rect 4956 24724 5012 26126
rect 5370 25900 5634 25910
rect 5426 25844 5474 25900
rect 5530 25844 5578 25900
rect 5370 25834 5634 25844
rect 5796 25618 5852 26236
rect 6076 26290 6132 26908
rect 6972 26964 7028 26974
rect 6972 26870 7028 26908
rect 6076 26238 6078 26290
rect 6130 26238 6132 26290
rect 6076 26226 6132 26238
rect 6748 25844 6804 25854
rect 5796 25566 5798 25618
rect 5850 25566 5852 25618
rect 5796 25554 5852 25566
rect 6524 25620 6580 25630
rect 5180 25506 5236 25518
rect 5180 25454 5182 25506
rect 5234 25454 5236 25506
rect 5068 25060 5124 25070
rect 5068 24836 5124 25004
rect 5180 24948 5236 25454
rect 6524 25506 6580 25564
rect 6524 25454 6526 25506
rect 6578 25454 6580 25506
rect 6524 25442 6580 25454
rect 6748 25506 6804 25788
rect 7420 25732 7476 27020
rect 7420 25666 7476 25676
rect 7532 27074 7588 27086
rect 7532 27022 7534 27074
rect 7586 27022 7588 27074
rect 7532 26852 7588 27022
rect 6748 25454 6750 25506
rect 6802 25454 6804 25506
rect 6748 25442 6804 25454
rect 6860 25620 6916 25630
rect 5180 24882 5236 24892
rect 6244 25394 6300 25406
rect 6244 25342 6246 25394
rect 6298 25342 6300 25394
rect 5068 24724 5124 24780
rect 6244 24836 6300 25342
rect 6748 25172 6804 25182
rect 6244 24770 6300 24780
rect 6524 24948 6580 24958
rect 5180 24724 5236 24734
rect 5068 24722 5236 24724
rect 5068 24670 5182 24722
rect 5234 24670 5236 24722
rect 5068 24668 5236 24670
rect 4956 24658 5012 24668
rect 5180 24658 5236 24668
rect 5292 24722 5348 24734
rect 5292 24670 5294 24722
rect 5346 24670 5348 24722
rect 4900 24500 4956 24510
rect 5292 24500 5348 24670
rect 4900 24498 5124 24500
rect 4900 24446 4902 24498
rect 4954 24446 5124 24498
rect 4900 24444 5124 24446
rect 4900 24434 4956 24444
rect 4340 24070 4396 24108
rect 4508 24108 4676 24164
rect 4396 23828 4452 23838
rect 4284 23268 4340 23278
rect 4172 23212 4284 23268
rect 3724 22370 3780 23212
rect 4284 23174 4340 23212
rect 4172 23044 4228 23054
rect 3724 22318 3726 22370
rect 3778 22318 3780 22370
rect 4060 22484 4116 22494
rect 4060 22370 4116 22428
rect 3724 22306 3780 22318
rect 3892 22314 3948 22326
rect 3892 22262 3894 22314
rect 3946 22262 3948 22314
rect 4060 22318 4062 22370
rect 4114 22318 4116 22370
rect 4060 22306 4116 22318
rect 4172 22370 4228 22988
rect 4396 22596 4452 23772
rect 4508 22708 4564 24108
rect 4900 24052 4956 24062
rect 4900 23994 4956 23996
rect 4620 23940 4676 23950
rect 4620 23846 4676 23884
rect 4900 23942 4902 23994
rect 4954 23942 4956 23994
rect 4732 23828 4788 23838
rect 4732 23734 4788 23772
rect 4732 23604 4788 23614
rect 4732 23154 4788 23548
rect 4900 23492 4956 23942
rect 5068 23938 5124 24444
rect 5068 23886 5070 23938
rect 5122 23886 5124 23938
rect 5068 23874 5124 23886
rect 5180 24444 5348 24500
rect 6300 24612 6356 24622
rect 5180 23604 5236 24444
rect 5370 24332 5634 24342
rect 5426 24276 5474 24332
rect 5530 24276 5578 24332
rect 5370 24266 5634 24276
rect 5796 23940 5852 23950
rect 5796 23846 5852 23884
rect 6076 23938 6132 23950
rect 6076 23886 6078 23938
rect 6130 23886 6132 23938
rect 6076 23716 6132 23886
rect 6300 23938 6356 24556
rect 6524 24174 6580 24892
rect 6636 24724 6692 24734
rect 6636 24630 6692 24668
rect 6524 24162 6636 24174
rect 6524 24110 6582 24162
rect 6634 24110 6636 24162
rect 6524 24108 6636 24110
rect 6580 24098 6636 24108
rect 6300 23886 6302 23938
rect 6354 23886 6356 23938
rect 6300 23828 6356 23886
rect 6300 23762 6356 23772
rect 6748 23716 6804 25116
rect 6860 24722 6916 25564
rect 7308 25506 7364 25518
rect 7308 25454 7310 25506
rect 7362 25454 7364 25506
rect 7028 25396 7084 25406
rect 7028 25394 7252 25396
rect 7028 25342 7030 25394
rect 7082 25342 7252 25394
rect 7028 25340 7252 25342
rect 7028 25330 7084 25340
rect 7196 25060 7252 25340
rect 7308 25284 7364 25454
rect 7420 25506 7476 25518
rect 7420 25454 7422 25506
rect 7474 25454 7476 25506
rect 7420 25284 7476 25454
rect 7532 25508 7588 26796
rect 7980 26292 8036 26302
rect 7980 26178 8036 26236
rect 7980 26126 7982 26178
rect 8034 26126 8036 26178
rect 7980 26068 8036 26126
rect 7532 25442 7588 25452
rect 7644 26012 8036 26068
rect 7644 25284 7700 26012
rect 7812 25732 7868 25742
rect 8092 25732 8148 27806
rect 8428 27636 8484 27646
rect 8316 27634 8484 27636
rect 8316 27582 8430 27634
rect 8482 27582 8484 27634
rect 8316 27580 8484 27582
rect 8316 27186 8372 27580
rect 8428 27570 8484 27580
rect 8316 27134 8318 27186
rect 8370 27134 8372 27186
rect 8316 27122 8372 27134
rect 9528 26684 9792 26694
rect 9584 26628 9632 26684
rect 9688 26628 9736 26684
rect 9528 26618 9792 26628
rect 9884 26516 9940 28588
rect 10444 28644 10500 28654
rect 12796 28644 12852 29542
rect 12908 29426 12964 29438
rect 12908 29374 12910 29426
rect 12962 29374 12964 29426
rect 12908 29316 12964 29374
rect 12908 29250 12964 29260
rect 13020 28766 13076 29922
rect 13823 29540 13879 30102
rect 13804 29484 13879 29540
rect 13356 29426 13412 29438
rect 13356 29374 13358 29426
rect 13410 29374 13412 29426
rect 13356 29316 13412 29374
rect 12964 28756 13076 28766
rect 13244 29204 13300 29214
rect 12964 28754 13188 28756
rect 12964 28702 12966 28754
rect 13018 28702 13188 28754
rect 12964 28700 13188 28702
rect 12964 28690 13020 28700
rect 10444 28642 10724 28644
rect 10444 28590 10446 28642
rect 10498 28590 10724 28642
rect 10444 28588 10724 28590
rect 10444 28578 10500 28588
rect 10668 28196 10724 28588
rect 12684 28588 12852 28644
rect 10668 28140 11172 28196
rect 11116 28082 11172 28140
rect 11116 28030 11118 28082
rect 11170 28030 11172 28082
rect 11116 28018 11172 28030
rect 12348 28026 12404 28038
rect 12348 27974 12350 28026
rect 12402 27974 12404 28026
rect 11452 27860 11508 27870
rect 11452 27766 11508 27804
rect 12236 27858 12292 27870
rect 12236 27806 12238 27858
rect 12290 27806 12292 27858
rect 9772 26460 9940 26516
rect 10220 26962 10276 26974
rect 10220 26910 10222 26962
rect 10274 26910 10276 26962
rect 9660 26305 9716 26330
rect 8764 26290 8820 26302
rect 8764 26238 8766 26290
rect 8818 26238 8820 26290
rect 7812 25638 7868 25676
rect 7980 25676 8148 25732
rect 8204 26068 8260 26078
rect 7420 25228 7700 25284
rect 7980 25284 8036 25676
rect 8204 25620 8260 26012
rect 8092 25564 8260 25620
rect 8484 26066 8540 26078
rect 8484 26014 8486 26066
rect 8538 26014 8540 26066
rect 8092 25506 8148 25564
rect 8092 25454 8094 25506
rect 8146 25454 8148 25506
rect 8484 25518 8540 26014
rect 8652 25844 8708 25854
rect 8484 25506 8596 25518
rect 8092 25442 8148 25454
rect 8372 25450 8428 25462
rect 8484 25454 8542 25506
rect 8594 25454 8596 25506
rect 8484 25452 8596 25454
rect 8204 25394 8260 25406
rect 8204 25342 8206 25394
rect 8258 25342 8260 25394
rect 8204 25284 8260 25342
rect 7308 25218 7364 25228
rect 7980 25218 8036 25228
rect 8092 25228 8260 25284
rect 8372 25398 8374 25450
rect 8426 25398 8428 25450
rect 8540 25442 8596 25452
rect 8372 25284 8428 25398
rect 7196 25004 8036 25060
rect 6860 24670 6862 24722
rect 6914 24670 6916 24722
rect 6860 24658 6916 24670
rect 7532 24836 7588 24846
rect 7532 24722 7588 24780
rect 7532 24670 7534 24722
rect 7586 24670 7588 24722
rect 7700 24836 7756 24846
rect 7700 24778 7756 24780
rect 7700 24726 7702 24778
rect 7754 24726 7756 24778
rect 7700 24714 7756 24726
rect 7868 24722 7924 24734
rect 7532 24658 7588 24670
rect 7868 24670 7870 24722
rect 7922 24670 7924 24722
rect 7140 24500 7196 24510
rect 7140 24498 7364 24500
rect 7140 24446 7142 24498
rect 7194 24446 7364 24498
rect 7140 24444 7364 24446
rect 7140 24434 7196 24444
rect 7140 24276 7196 24286
rect 7140 24052 7196 24220
rect 7140 23994 7196 23996
rect 6860 23940 6916 23950
rect 7140 23942 7142 23994
rect 7194 23942 7196 23994
rect 7140 23930 7196 23942
rect 7308 23938 7364 24444
rect 7868 24276 7924 24670
rect 7980 24722 8036 25004
rect 7980 24670 7982 24722
rect 8034 24670 8036 24722
rect 7980 24658 8036 24670
rect 6860 23846 6916 23884
rect 7308 23886 7310 23938
rect 7362 23886 7364 23938
rect 7308 23874 7364 23886
rect 7532 24220 7924 24276
rect 6972 23826 7028 23838
rect 6972 23774 6974 23826
rect 7026 23774 7028 23826
rect 6860 23716 6916 23726
rect 6748 23660 6860 23716
rect 6076 23650 6132 23660
rect 5180 23538 5236 23548
rect 6300 23604 6356 23614
rect 4732 23102 4734 23154
rect 4786 23102 4788 23154
rect 4732 23090 4788 23102
rect 4844 23436 4956 23492
rect 4844 23156 4900 23436
rect 5608 23268 5664 23278
rect 5608 23210 5664 23212
rect 5608 23158 5610 23210
rect 5662 23158 5664 23210
rect 5608 23146 5664 23158
rect 6300 23154 6356 23548
rect 6636 23268 6692 23278
rect 6636 23198 6692 23212
rect 4844 23090 4900 23100
rect 6300 23102 6302 23154
rect 6354 23102 6356 23154
rect 6300 23090 6356 23102
rect 6412 23156 6468 23166
rect 6636 23146 6638 23198
rect 6690 23146 6692 23198
rect 6636 23134 6692 23146
rect 5852 22932 5908 22942
rect 5852 22838 5908 22876
rect 5370 22764 5634 22774
rect 5426 22708 5474 22764
rect 5530 22708 5578 22764
rect 4508 22652 5068 22708
rect 5370 22698 5634 22708
rect 4172 22318 4174 22370
rect 4226 22318 4228 22370
rect 4172 22306 4228 22318
rect 4284 22540 4452 22596
rect 3892 21700 3948 22262
rect 4284 21710 4340 22540
rect 5012 22482 5068 22652
rect 5012 22430 5014 22482
rect 5066 22430 5068 22482
rect 5012 22418 5068 22430
rect 4452 22372 4508 22382
rect 4452 22278 4508 22316
rect 3612 21522 3668 21532
rect 3836 21644 3948 21700
rect 4228 21698 4340 21710
rect 4228 21646 4230 21698
rect 4282 21646 4340 21698
rect 4228 21644 4340 21646
rect 3668 20916 3724 20926
rect 3668 20822 3724 20860
rect 2828 20132 2884 20142
rect 2604 19234 2660 19246
rect 2604 19182 2606 19234
rect 2658 19182 2660 19234
rect 2604 18452 2660 19182
rect 2828 19234 2884 20076
rect 3612 20132 3668 20142
rect 3052 20020 3108 20030
rect 2940 20018 3108 20020
rect 2940 19966 3054 20018
rect 3106 19966 3108 20018
rect 2940 19964 3108 19966
rect 2940 19402 2996 19964
rect 3052 19954 3108 19964
rect 3220 19962 3276 19974
rect 3220 19910 3222 19962
rect 3274 19910 3276 19962
rect 3220 19460 3276 19910
rect 3220 19404 3332 19460
rect 2940 19350 2942 19402
rect 2994 19350 2996 19402
rect 2940 19338 2996 19350
rect 2828 19182 2830 19234
rect 2882 19182 2884 19234
rect 2828 19170 2884 19182
rect 3276 19236 3332 19404
rect 3500 19236 3556 19246
rect 3276 19234 3556 19236
rect 3276 19182 3502 19234
rect 3554 19182 3556 19234
rect 3276 19180 3556 19182
rect 2604 18386 2660 18396
rect 3276 18900 3332 18910
rect 3276 18450 3332 18844
rect 3276 18398 3278 18450
rect 3330 18398 3332 18450
rect 3276 18386 3332 18398
rect 3388 18340 3444 18350
rect 3164 17892 3220 17902
rect 3388 17892 3444 18284
rect 3500 18338 3556 19180
rect 3612 19012 3668 20076
rect 3724 20018 3780 20030
rect 3724 19966 3726 20018
rect 3778 19966 3780 20018
rect 3724 19908 3780 19966
rect 3724 19842 3780 19852
rect 3836 19346 3892 21644
rect 4228 21634 4284 21644
rect 4060 21588 4116 21598
rect 4508 21588 4564 21598
rect 3948 20802 4004 20814
rect 3948 20750 3950 20802
rect 4002 20750 4004 20802
rect 3948 20692 4004 20750
rect 4060 20802 4116 21532
rect 4396 21586 4564 21588
rect 4396 21534 4510 21586
rect 4562 21534 4564 21586
rect 4396 21532 4564 21534
rect 4060 20750 4062 20802
rect 4114 20750 4116 20802
rect 4060 20738 4116 20750
rect 4172 20916 4228 20926
rect 3948 20626 4004 20636
rect 3966 20020 4022 20030
rect 3966 19926 4022 19964
rect 3836 19294 3838 19346
rect 3890 19294 3892 19346
rect 3836 19282 3892 19294
rect 4172 19234 4228 20860
rect 4396 20356 4452 21532
rect 4508 21522 4564 21532
rect 4732 21586 4788 21598
rect 4732 21534 4734 21586
rect 4786 21534 4788 21586
rect 4732 21364 4788 21534
rect 4844 21588 4900 21598
rect 4844 21494 4900 21532
rect 5012 21364 5068 21374
rect 4732 21362 5068 21364
rect 4732 21310 5014 21362
rect 5066 21310 5068 21362
rect 4732 21308 5068 21310
rect 5012 21028 5068 21308
rect 5370 21196 5634 21206
rect 5426 21140 5474 21196
rect 5530 21140 5578 21196
rect 5370 21130 5634 21140
rect 6412 21038 6468 23100
rect 6748 23044 6804 23054
rect 6748 22950 6804 22988
rect 5012 20962 5068 20972
rect 5628 21028 5684 21038
rect 5628 20802 5684 20972
rect 6356 21026 6468 21038
rect 6356 20974 6358 21026
rect 6410 20974 6468 21026
rect 6356 20972 6468 20974
rect 6860 22596 6916 23660
rect 6356 20962 6412 20972
rect 5628 20750 5630 20802
rect 5682 20750 5684 20802
rect 5964 20804 6020 20814
rect 5628 20738 5684 20750
rect 5796 20746 5852 20758
rect 5796 20694 5798 20746
rect 5850 20694 5852 20746
rect 5964 20710 6020 20748
rect 6076 20802 6132 20814
rect 6076 20750 6078 20802
rect 6130 20750 6132 20802
rect 4284 20300 4452 20356
rect 4508 20356 4564 20366
rect 4284 20020 4340 20300
rect 4508 20142 4564 20300
rect 5796 20356 5852 20694
rect 5796 20290 5852 20300
rect 6076 20188 6132 20750
rect 4452 20130 4564 20142
rect 4452 20078 4454 20130
rect 4506 20078 4564 20130
rect 4452 20076 4564 20078
rect 5516 20132 5572 20142
rect 4452 20066 4508 20076
rect 5516 20074 5572 20076
rect 4284 19954 4340 19964
rect 4732 20020 4788 20030
rect 4732 19926 4788 19964
rect 4844 20020 4900 20030
rect 5180 20020 5236 20030
rect 4844 20018 5236 20020
rect 4844 19966 4846 20018
rect 4898 19966 5182 20018
rect 5234 19966 5236 20018
rect 5516 20022 5518 20074
rect 5570 20022 5572 20074
rect 5516 20010 5572 20022
rect 5628 20132 6132 20188
rect 4844 19964 5236 19966
rect 3836 19178 3892 19190
rect 3836 19126 3838 19178
rect 3890 19126 3892 19178
rect 4172 19182 4174 19234
rect 4226 19182 4228 19234
rect 4172 19170 4228 19182
rect 4508 19908 4564 19918
rect 4508 19234 4564 19852
rect 4844 19236 4900 19964
rect 5180 19954 5236 19964
rect 5516 19908 5572 19918
rect 5628 19908 5684 20132
rect 5516 19906 5684 19908
rect 5516 19854 5518 19906
rect 5570 19854 5684 19906
rect 5516 19852 5684 19854
rect 5852 20020 5908 20030
rect 5516 19842 5572 19852
rect 5370 19628 5634 19638
rect 5426 19572 5474 19628
rect 5530 19572 5578 19628
rect 5370 19562 5634 19572
rect 4508 19182 4510 19234
rect 4562 19182 4564 19234
rect 3612 18956 3780 19012
rect 3500 18286 3502 18338
rect 3554 18286 3556 18338
rect 3500 18274 3556 18286
rect 3612 18450 3668 18462
rect 3612 18398 3614 18450
rect 3666 18398 3668 18450
rect 3164 17890 3444 17892
rect 3164 17838 3166 17890
rect 3218 17838 3444 17890
rect 3164 17836 3444 17838
rect 3612 17892 3668 18398
rect 3724 17902 3780 18956
rect 3836 18788 3892 19126
rect 3836 18722 3892 18732
rect 3948 18900 4004 18910
rect 3724 17890 3836 17902
rect 3724 17838 3782 17890
rect 3834 17838 3836 17890
rect 3724 17836 3836 17838
rect 3164 17826 3220 17836
rect 3612 17826 3668 17836
rect 3780 17826 3836 17836
rect 3500 17668 3556 17678
rect 3500 17666 3668 17668
rect 3500 17614 3502 17666
rect 3554 17614 3668 17666
rect 3500 17612 3668 17614
rect 3500 17602 3556 17612
rect 3612 17108 3668 17612
rect 3948 17332 4004 18844
rect 4060 18452 4116 18462
rect 4396 18452 4452 18462
rect 4060 18228 4116 18396
rect 4060 18162 4116 18172
rect 4172 18450 4452 18452
rect 4172 18398 4398 18450
rect 4450 18398 4452 18450
rect 4172 18396 4452 18398
rect 4060 17892 4116 17902
rect 4060 17666 4116 17836
rect 4060 17614 4062 17666
rect 4114 17614 4116 17666
rect 4060 17602 4116 17614
rect 4172 17556 4228 18396
rect 4396 18386 4452 18396
rect 4508 18340 4564 19182
rect 4508 18274 4564 18284
rect 4732 19234 4900 19236
rect 4732 19182 4846 19234
rect 4898 19182 4900 19234
rect 4732 19180 4900 19182
rect 4396 17892 4452 17902
rect 4284 17668 4340 17678
rect 4284 17574 4340 17612
rect 4396 17668 4452 17836
rect 4732 17892 4788 19180
rect 4844 19170 4900 19180
rect 4956 19402 5012 19414
rect 4956 19350 4958 19402
rect 5010 19350 5012 19402
rect 4956 19236 5012 19350
rect 5852 19402 5908 19964
rect 6860 20018 6916 22540
rect 6860 19966 6862 20018
rect 6914 19966 6916 20018
rect 6860 19954 6916 19966
rect 6972 19906 7028 23774
rect 7532 23156 7588 24220
rect 7868 23938 7924 23950
rect 7868 23886 7870 23938
rect 7922 23886 7924 23938
rect 7868 23828 7924 23886
rect 7868 23762 7924 23772
rect 8092 23156 8148 25228
rect 8372 24846 8428 25228
rect 8372 24836 8484 24846
rect 8372 24780 8428 24836
rect 8428 24770 8484 24780
rect 8260 24724 8316 24734
rect 8260 24630 8316 24668
rect 8316 24164 8372 24174
rect 8204 24052 8260 24062
rect 8204 23911 8260 23996
rect 8204 23859 8206 23911
rect 8258 23859 8260 23911
rect 8204 23847 8260 23859
rect 7532 23090 7588 23100
rect 7644 23100 8148 23156
rect 8204 23770 8260 23782
rect 8204 23718 8206 23770
rect 8258 23718 8260 23770
rect 8204 23154 8260 23718
rect 8316 23266 8372 24108
rect 8540 23940 8596 23950
rect 8652 23940 8708 25788
rect 8764 25732 8820 26238
rect 8876 26292 8932 26302
rect 8876 26198 8932 26236
rect 9660 26292 9662 26305
rect 9714 26292 9716 26305
rect 9660 26226 9716 26236
rect 9548 26180 9604 26190
rect 8764 25666 8820 25676
rect 9324 26178 9604 26180
rect 9324 26126 9550 26178
rect 9602 26126 9604 26178
rect 9324 26124 9604 26126
rect 8764 25508 8820 25518
rect 8764 25414 8820 25452
rect 8540 23938 8708 23940
rect 8540 23886 8542 23938
rect 8594 23886 8708 23938
rect 8540 23884 8708 23886
rect 9212 24276 9268 24286
rect 8540 23716 8596 23884
rect 8540 23650 8596 23660
rect 8876 23828 8932 23838
rect 9044 23828 9100 23838
rect 8316 23214 8318 23266
rect 8370 23214 8372 23266
rect 8316 23202 8372 23214
rect 8204 23102 8206 23154
rect 8258 23102 8260 23154
rect 8652 23154 8708 23166
rect 7532 22932 7588 22942
rect 7532 22332 7588 22876
rect 7532 22280 7534 22332
rect 7586 22280 7588 22332
rect 7532 22268 7588 22280
rect 7644 20970 7700 23100
rect 8204 23090 8260 23102
rect 8484 23098 8540 23110
rect 8484 23046 8486 23098
rect 8538 23046 8540 23098
rect 8484 23044 8540 23046
rect 8484 22978 8540 22988
rect 8652 23102 8654 23154
rect 8706 23102 8708 23154
rect 7924 22932 7980 22942
rect 7924 22838 7980 22876
rect 8428 22820 8484 22830
rect 7868 22484 7924 22494
rect 7868 22370 7924 22428
rect 7868 22318 7870 22370
rect 7922 22318 7924 22370
rect 7868 22306 7924 22318
rect 8092 22372 8148 22382
rect 8092 22278 8148 22316
rect 8260 22314 8316 22326
rect 8260 22262 8262 22314
rect 8314 22262 8316 22314
rect 8260 22260 8316 22262
rect 8428 22260 8484 22764
rect 8652 22708 8708 23102
rect 8652 22642 8708 22652
rect 8876 22484 8932 23772
rect 8988 23826 9100 23828
rect 8988 23774 9046 23826
rect 9098 23774 9100 23826
rect 8988 23762 9100 23774
rect 8988 22820 9044 23762
rect 8988 22754 9044 22764
rect 9212 22494 9268 24220
rect 9324 24164 9380 26124
rect 9548 26114 9604 26124
rect 9772 25518 9828 26460
rect 9996 26290 10052 26302
rect 9996 26238 9998 26290
rect 10050 26238 10052 26290
rect 9772 25508 9884 25518
rect 9772 25452 9828 25508
rect 9828 25284 9884 25452
rect 9996 25508 10052 26238
rect 10220 25844 10276 26910
rect 10836 26852 10892 26862
rect 10836 26850 10948 26852
rect 10836 26798 10838 26850
rect 10890 26798 10948 26850
rect 10836 26786 10948 26798
rect 10500 26180 10556 26190
rect 10220 25778 10276 25788
rect 10444 26124 10500 26180
rect 10444 26086 10556 26124
rect 10892 26180 10948 26786
rect 10892 26114 10948 26124
rect 11564 26290 11620 26302
rect 11564 26238 11566 26290
rect 11618 26238 11620 26290
rect 9996 25442 10052 25452
rect 10108 25508 10164 25518
rect 10444 25508 10500 26086
rect 11228 26068 11284 26078
rect 11004 26066 11284 26068
rect 11004 26014 11230 26066
rect 11282 26014 11284 26066
rect 11004 26012 11284 26014
rect 10892 25620 10948 25630
rect 11004 25620 11060 26012
rect 11228 26002 11284 26012
rect 11564 25844 11620 26238
rect 12124 26292 12180 26302
rect 12236 26292 12292 27806
rect 12348 27860 12404 27974
rect 12348 27794 12404 27804
rect 12684 27897 12740 28588
rect 12684 27845 12686 27897
rect 12738 27845 12740 27897
rect 12684 27076 12740 27845
rect 12908 27860 12964 27870
rect 12908 27766 12964 27804
rect 12684 27010 12740 27020
rect 12236 26236 12516 26292
rect 11956 26180 12012 26190
rect 11956 26178 12068 26180
rect 11956 26126 11958 26178
rect 12010 26126 12068 26178
rect 11956 26114 12068 26126
rect 10892 25618 11060 25620
rect 10892 25566 10894 25618
rect 10946 25566 11060 25618
rect 10892 25564 11060 25566
rect 11116 25788 11620 25844
rect 10892 25554 10948 25564
rect 10108 25506 10500 25508
rect 10108 25454 10110 25506
rect 10162 25454 10500 25506
rect 10108 25452 10500 25454
rect 10108 25284 10164 25452
rect 9828 25282 10164 25284
rect 9828 25230 9830 25282
rect 9882 25230 10164 25282
rect 9828 25228 10164 25230
rect 9828 25218 9884 25228
rect 9528 25116 9792 25126
rect 9584 25060 9632 25116
rect 9688 25060 9736 25116
rect 9528 25050 9792 25060
rect 10108 24500 10164 25228
rect 11004 25396 11060 25406
rect 10332 24500 10388 24510
rect 10108 24498 10388 24500
rect 10108 24446 10334 24498
rect 10386 24446 10388 24498
rect 10108 24444 10388 24446
rect 9324 24098 9380 24108
rect 10220 24052 10276 24062
rect 9324 23938 9380 23950
rect 9324 23886 9326 23938
rect 9378 23886 9380 23938
rect 9324 22932 9380 23886
rect 9548 23938 9604 23950
rect 9548 23886 9550 23938
rect 9602 23886 9604 23938
rect 9548 23828 9604 23886
rect 9828 23940 9884 23950
rect 9828 23846 9884 23884
rect 10108 23938 10164 23950
rect 10108 23886 10110 23938
rect 10162 23886 10164 23938
rect 9548 23762 9604 23772
rect 9528 23548 9792 23558
rect 9584 23492 9632 23548
rect 9688 23492 9736 23548
rect 10108 23492 10164 23886
rect 9528 23482 9792 23492
rect 9324 22708 9380 22876
rect 9996 23436 10164 23492
rect 10220 23938 10276 23996
rect 10220 23886 10222 23938
rect 10274 23886 10276 23938
rect 9324 22652 9604 22708
rect 9212 22482 9324 22494
rect 9212 22430 9270 22482
rect 9322 22430 9324 22482
rect 9212 22428 9324 22430
rect 8876 22418 8932 22428
rect 9268 22418 9324 22428
rect 8540 22372 8596 22382
rect 8540 22278 8596 22316
rect 8708 22372 8764 22382
rect 8708 22370 8820 22372
rect 8708 22318 8710 22370
rect 8762 22318 8820 22370
rect 8708 22306 8820 22318
rect 8260 22204 8484 22260
rect 8316 21588 8372 21598
rect 8316 21494 8372 21532
rect 8428 21476 8484 22204
rect 8652 22148 8708 22158
rect 8652 21586 8708 22092
rect 8652 21534 8654 21586
rect 8706 21534 8708 21586
rect 8652 21522 8708 21534
rect 8764 21588 8820 22306
rect 8988 22370 9044 22382
rect 8988 22318 8990 22370
rect 9042 22318 9044 22370
rect 8764 21522 8820 21532
rect 8876 22260 8932 22270
rect 8428 21410 8484 21420
rect 7196 20916 7252 20926
rect 7644 20918 7646 20970
rect 7698 20918 7700 20970
rect 7644 20906 7700 20918
rect 8876 20916 8932 22204
rect 8988 21700 9044 22318
rect 9548 22370 9604 22652
rect 9884 22596 9940 22606
rect 9996 22596 10052 23436
rect 10108 23268 10164 23278
rect 10220 23268 10276 23886
rect 10108 23266 10276 23268
rect 10108 23214 10110 23266
rect 10162 23214 10276 23266
rect 10108 23212 10276 23214
rect 10108 23202 10164 23212
rect 9940 22540 10052 22596
rect 9884 22502 9940 22540
rect 9548 22318 9550 22370
rect 9602 22318 9604 22370
rect 9548 22148 9604 22318
rect 9548 22082 9604 22092
rect 9528 21980 9792 21990
rect 9584 21924 9632 21980
rect 9688 21924 9736 21980
rect 9528 21914 9792 21924
rect 8988 21644 9268 21700
rect 9044 21476 9100 21486
rect 9044 21382 9100 21420
rect 8876 20860 9044 20916
rect 7196 20802 7252 20860
rect 7196 20750 7198 20802
rect 7250 20750 7252 20802
rect 7196 20738 7252 20750
rect 7532 20804 7588 20814
rect 7532 20802 7700 20804
rect 7532 20750 7534 20802
rect 7586 20750 7700 20802
rect 7532 20748 7700 20750
rect 7532 20738 7588 20748
rect 6972 19854 6974 19906
rect 7026 19854 7028 19906
rect 6972 19842 7028 19854
rect 7084 20132 7140 20142
rect 5852 19350 5854 19402
rect 5906 19350 5908 19402
rect 5852 19338 5908 19350
rect 7084 19256 7140 20076
rect 7308 20057 7364 20069
rect 7308 20005 7310 20057
rect 7362 20005 7364 20057
rect 4956 19170 5012 19180
rect 5740 19234 5796 19246
rect 6860 19236 6916 19246
rect 5740 19182 5742 19234
rect 5794 19182 5796 19234
rect 6748 19234 6916 19236
rect 4900 18788 4956 18798
rect 4900 18562 4956 18732
rect 4900 18510 4902 18562
rect 4954 18510 4956 18562
rect 4900 18498 4956 18510
rect 5180 18450 5236 18462
rect 5180 18398 5182 18450
rect 5234 18398 5236 18450
rect 5180 17892 5236 18398
rect 5292 18450 5348 18462
rect 5292 18398 5294 18450
rect 5346 18398 5348 18450
rect 5292 18340 5348 18398
rect 5292 18274 5348 18284
rect 5740 18340 5796 19182
rect 6416 19196 6472 19208
rect 6416 19144 6418 19196
rect 6470 19144 6472 19196
rect 6416 18900 6472 19144
rect 6416 18834 6472 18844
rect 6748 19182 6862 19234
rect 6914 19182 6916 19234
rect 6748 19180 6916 19182
rect 6412 18676 6468 18686
rect 6300 18564 6356 18574
rect 6300 18452 6356 18508
rect 5740 18274 5796 18284
rect 6076 18450 6356 18452
rect 6076 18398 6302 18450
rect 6354 18398 6356 18450
rect 6076 18396 6356 18398
rect 5370 18060 5634 18070
rect 5426 18004 5474 18060
rect 5530 18004 5578 18060
rect 5370 17994 5634 18004
rect 4732 17890 5236 17892
rect 4732 17838 4734 17890
rect 4786 17838 5236 17890
rect 4732 17836 5236 17838
rect 5964 17892 6020 17902
rect 4732 17826 4788 17836
rect 5740 17668 5796 17678
rect 4396 17666 4788 17668
rect 4396 17614 4398 17666
rect 4450 17614 4788 17666
rect 4396 17612 4788 17614
rect 4396 17602 4452 17612
rect 4172 17490 4228 17500
rect 3948 17266 4004 17276
rect 3612 17052 4676 17108
rect 4172 16884 4228 16894
rect 4172 16790 4228 16828
rect 1820 16100 1876 16110
rect 2604 16100 2660 16110
rect 1596 15316 1652 15326
rect 1820 15316 1876 16044
rect 1596 15314 1876 15316
rect 1596 15262 1598 15314
rect 1650 15262 1876 15314
rect 1596 15260 1876 15262
rect 2268 16098 2660 16100
rect 2268 16046 2606 16098
rect 2658 16046 2660 16098
rect 2268 16044 2660 16046
rect 1596 15250 1652 15260
rect 2268 13524 2324 16044
rect 2604 16034 2660 16044
rect 4284 15426 4340 17052
rect 4508 16884 4564 16894
rect 4508 16790 4564 16828
rect 4620 16882 4676 17052
rect 4620 16830 4622 16882
rect 4674 16830 4676 16882
rect 4620 16818 4676 16830
rect 4508 16212 4564 16222
rect 4732 16212 4788 17612
rect 5740 17574 5796 17612
rect 5964 17666 6020 17836
rect 6076 17834 6132 18396
rect 6300 18386 6356 18396
rect 6412 18450 6468 18620
rect 6748 18574 6804 19180
rect 6860 19170 6916 19180
rect 7028 19234 7140 19256
rect 7028 19182 7030 19234
rect 7082 19182 7140 19234
rect 7028 19170 7140 19182
rect 7084 18900 7140 19170
rect 6692 18562 6804 18574
rect 6692 18510 6694 18562
rect 6746 18510 6804 18562
rect 6692 18508 6804 18510
rect 6972 18844 7140 18900
rect 7196 19348 7252 19358
rect 7196 19234 7252 19292
rect 7196 19182 7198 19234
rect 7250 19182 7252 19234
rect 6692 18498 6748 18508
rect 6412 18398 6414 18450
rect 6466 18398 6468 18450
rect 6412 18386 6468 18398
rect 6972 18116 7028 18844
rect 7196 18788 7252 19182
rect 7308 19236 7364 20005
rect 7532 20020 7588 20030
rect 7532 19926 7588 19964
rect 7644 19470 7700 20748
rect 7868 20020 7924 20030
rect 7868 20018 8036 20020
rect 7868 19966 7870 20018
rect 7922 19966 8036 20018
rect 7868 19964 8036 19966
rect 7868 19954 7924 19964
rect 7588 19458 7700 19470
rect 7588 19406 7590 19458
rect 7642 19406 7700 19458
rect 7588 19404 7700 19406
rect 7588 19394 7644 19404
rect 7980 19402 8036 19964
rect 7980 19350 7982 19402
rect 8034 19350 8036 19402
rect 7980 19338 8036 19350
rect 8316 20018 8372 20030
rect 8316 19966 8318 20018
rect 8370 19966 8372 20018
rect 8092 19236 8148 19246
rect 7308 19142 7364 19180
rect 7420 19234 8148 19236
rect 7420 19182 8094 19234
rect 8146 19182 8148 19234
rect 7420 19180 8148 19182
rect 7196 18722 7252 18732
rect 7084 18564 7140 18574
rect 7420 18564 7476 19180
rect 8092 19170 8148 19180
rect 7084 18470 7140 18508
rect 7252 18508 7476 18564
rect 7252 18506 7308 18508
rect 7252 18454 7254 18506
rect 7306 18454 7308 18506
rect 7252 18442 7308 18454
rect 6972 18060 7252 18116
rect 6076 17782 6078 17834
rect 6130 17782 6132 17834
rect 6076 17770 6132 17782
rect 5964 17614 5966 17666
rect 6018 17614 6020 17666
rect 5964 17602 6020 17614
rect 6300 17668 6356 17678
rect 4956 17556 5012 17566
rect 4956 17106 5012 17500
rect 4956 17054 4958 17106
rect 5010 17054 5012 17106
rect 4956 17042 5012 17054
rect 5404 16882 5460 16894
rect 5404 16830 5406 16882
rect 5458 16830 5460 16882
rect 5404 16660 5460 16830
rect 6300 16884 6356 17612
rect 6972 17666 7028 17678
rect 6972 17614 6974 17666
rect 7026 17614 7028 17666
rect 6972 17556 7028 17614
rect 7196 17668 7252 18060
rect 7420 17834 7476 18508
rect 7756 18452 7812 18462
rect 7420 17782 7422 17834
rect 7474 17782 7476 17834
rect 7420 17770 7476 17782
rect 7644 18228 7700 18238
rect 7644 17780 7700 18172
rect 7308 17668 7364 17678
rect 7196 17666 7364 17668
rect 7196 17614 7310 17666
rect 7362 17614 7364 17666
rect 7196 17612 7364 17614
rect 6972 17490 7028 17500
rect 7308 17444 7364 17612
rect 7644 17666 7700 17724
rect 7644 17614 7646 17666
rect 7698 17614 7700 17666
rect 7644 17602 7700 17614
rect 7756 17668 7812 18396
rect 7998 18340 8054 18350
rect 7998 18246 8054 18284
rect 7756 17602 7812 17612
rect 8092 17780 8148 17790
rect 7308 17378 7364 17388
rect 7812 17444 7868 17454
rect 7812 17350 7868 17388
rect 8092 16994 8148 17724
rect 8316 17780 8372 19966
rect 8540 20018 8596 20030
rect 8540 19966 8542 20018
rect 8594 19966 8596 20018
rect 8540 19348 8596 19966
rect 8820 20020 8876 20030
rect 8820 19926 8876 19964
rect 8540 19282 8596 19292
rect 8428 19234 8484 19246
rect 8428 19182 8430 19234
rect 8482 19182 8484 19234
rect 8428 19124 8484 19182
rect 8764 19234 8820 19246
rect 8764 19182 8766 19234
rect 8818 19182 8820 19234
rect 8764 19124 8820 19182
rect 8428 19068 8820 19124
rect 8428 18900 8484 19068
rect 8428 18834 8484 18844
rect 8540 18676 8596 18686
rect 8540 18618 8596 18620
rect 8540 18566 8542 18618
rect 8594 18566 8596 18618
rect 8540 18554 8596 18566
rect 8764 18465 8820 18477
rect 8428 18452 8484 18462
rect 8428 18358 8484 18396
rect 8764 18413 8766 18465
rect 8818 18413 8820 18465
rect 8316 17714 8372 17724
rect 8764 17444 8820 18413
rect 8988 18340 9044 20860
rect 9212 20804 9268 21644
rect 9212 19402 9268 20748
rect 9528 20412 9792 20422
rect 9584 20356 9632 20412
rect 9688 20356 9736 20412
rect 9528 20346 9792 20356
rect 9436 20020 9492 20030
rect 9436 19926 9492 19964
rect 10332 20020 10388 24444
rect 10892 24052 10948 24062
rect 10892 22372 10948 23996
rect 11004 23994 11060 25340
rect 11116 24948 11172 25788
rect 11116 24882 11172 24892
rect 12012 24836 12068 26114
rect 11900 24780 12012 24836
rect 11900 24749 11956 24780
rect 11004 23942 11006 23994
rect 11058 23942 11060 23994
rect 11676 24724 11732 24734
rect 11900 24697 11902 24749
rect 11954 24697 11956 24749
rect 12012 24742 12068 24780
rect 11900 24685 11956 24697
rect 11676 24050 11732 24668
rect 11676 23998 11678 24050
rect 11730 23998 11732 24050
rect 11676 23986 11732 23998
rect 11844 24052 11900 24062
rect 11844 23994 11900 23996
rect 11004 23930 11060 23942
rect 11228 23940 11284 23950
rect 11228 23858 11230 23884
rect 11282 23858 11284 23884
rect 11228 23846 11284 23858
rect 11564 23940 11620 23950
rect 11844 23942 11846 23994
rect 11898 23942 11900 23994
rect 11844 23930 11900 23942
rect 12124 23938 12180 26236
rect 12292 26068 12348 26078
rect 12292 25974 12348 26012
rect 12460 24948 12516 26236
rect 12572 26290 12628 26302
rect 12572 26238 12574 26290
rect 12626 26238 12628 26290
rect 12572 25620 12628 26238
rect 12684 26292 12740 26302
rect 12684 26198 12740 26236
rect 13132 26190 13188 28700
rect 13244 27860 13300 29148
rect 13356 28644 13412 29260
rect 13468 29428 13524 29438
rect 13468 28868 13524 29372
rect 13804 29242 13860 29484
rect 13748 29204 13860 29242
rect 13804 29148 13860 29204
rect 13748 29138 13804 29148
rect 13686 29036 13950 29046
rect 13742 28980 13790 29036
rect 13846 28980 13894 29036
rect 13686 28970 13950 28980
rect 13916 28868 13972 28878
rect 13468 28812 13860 28868
rect 13356 28578 13412 28588
rect 13468 28642 13524 28654
rect 13468 28590 13470 28642
rect 13522 28590 13524 28642
rect 13468 28532 13524 28590
rect 13636 28644 13692 28654
rect 13636 28550 13692 28588
rect 13804 28642 13860 28812
rect 13804 28590 13806 28642
rect 13858 28590 13860 28642
rect 13804 28578 13860 28590
rect 13916 28642 13972 28812
rect 13916 28590 13918 28642
rect 13970 28590 13972 28642
rect 13916 28578 13972 28590
rect 13468 28466 13524 28476
rect 13244 27794 13300 27804
rect 14028 27860 14084 30940
rect 14812 30994 14868 31500
rect 15820 31556 15876 31566
rect 15820 31462 15876 31500
rect 14812 30942 14814 30994
rect 14866 30942 14868 30994
rect 14812 30930 14868 30942
rect 14700 30210 14756 30222
rect 14700 30158 14702 30210
rect 14754 30158 14756 30210
rect 14700 30100 14756 30158
rect 15708 30210 15764 30222
rect 15708 30158 15710 30210
rect 15762 30158 15764 30210
rect 14756 30044 14868 30100
rect 14700 30034 14756 30044
rect 14644 29540 14700 29550
rect 14644 29446 14700 29484
rect 14252 29428 14308 29438
rect 14252 29334 14308 29372
rect 14364 29426 14420 29438
rect 14364 29374 14366 29426
rect 14418 29374 14420 29426
rect 14364 29204 14420 29374
rect 14364 29138 14420 29148
rect 14812 29204 14868 30044
rect 15708 29988 15764 30158
rect 15708 29922 15764 29932
rect 16044 30154 16100 30166
rect 16044 30102 16046 30154
rect 16098 30102 16100 30154
rect 16044 29594 16100 30102
rect 16268 30042 16324 31724
rect 19180 31778 19236 31790
rect 19180 31726 19182 31778
rect 19234 31726 19236 31778
rect 17844 31388 18108 31398
rect 17900 31332 17948 31388
rect 18004 31332 18052 31388
rect 17844 31322 18108 31332
rect 19180 31108 19236 31726
rect 19460 31722 19516 31734
rect 19460 31670 19462 31722
rect 19514 31670 19516 31722
rect 19460 31668 19516 31670
rect 18508 31052 19236 31108
rect 19404 31612 19516 31668
rect 16716 30882 16772 30894
rect 16716 30830 16718 30882
rect 16770 30830 16772 30882
rect 16268 29990 16270 30042
rect 16322 29990 16324 30042
rect 16268 29978 16324 29990
rect 16380 30210 16436 30222
rect 16380 30158 16382 30210
rect 16434 30158 16436 30210
rect 15932 29540 15988 29550
rect 16044 29542 16046 29594
rect 16098 29542 16100 29594
rect 16380 29652 16436 30158
rect 16716 30212 16772 30830
rect 17836 30378 17892 30390
rect 17836 30326 17838 30378
rect 17890 30326 17892 30378
rect 16828 30212 16884 30222
rect 16716 30156 16828 30212
rect 16380 29586 16436 29596
rect 16044 29530 16100 29542
rect 15932 29470 15988 29484
rect 14812 29138 14868 29148
rect 15428 29428 15484 29438
rect 14196 28924 14980 28980
rect 14196 28866 14252 28924
rect 14196 28814 14198 28866
rect 14250 28814 14252 28866
rect 14196 28802 14252 28814
rect 14364 28756 14420 28766
rect 14028 27858 14308 27860
rect 14028 27806 14030 27858
rect 14082 27806 14308 27858
rect 14028 27804 14308 27806
rect 14028 27794 14084 27804
rect 13686 27468 13950 27478
rect 13742 27412 13790 27468
rect 13846 27412 13894 27468
rect 13686 27402 13950 27412
rect 14028 27076 14084 27086
rect 14028 26982 14084 27020
rect 14252 26292 14308 27804
rect 14364 27074 14420 28700
rect 14700 28642 14756 28654
rect 14700 28590 14702 28642
rect 14754 28590 14756 28642
rect 14364 27022 14366 27074
rect 14418 27022 14420 27074
rect 14364 27010 14420 27022
rect 14476 27242 14532 27254
rect 14476 27190 14478 27242
rect 14530 27190 14532 27242
rect 14476 27076 14532 27190
rect 14476 27010 14532 27020
rect 13132 26180 13244 26190
rect 13132 26124 13188 26180
rect 13188 26086 13244 26124
rect 13686 25900 13950 25910
rect 13742 25844 13790 25900
rect 13846 25844 13894 25900
rect 13686 25834 13950 25844
rect 12796 25620 12852 25630
rect 13692 25620 13748 25630
rect 12572 25618 13412 25620
rect 12572 25566 12798 25618
rect 12850 25566 13412 25618
rect 12572 25564 13412 25566
rect 12796 25554 12852 25564
rect 13356 25506 13412 25564
rect 13356 25454 13358 25506
rect 13410 25454 13412 25506
rect 13356 25442 13412 25454
rect 13524 25508 13580 25518
rect 12348 24892 12516 24948
rect 12572 25396 12628 25406
rect 12236 24722 12292 24734
rect 12236 24670 12238 24722
rect 12290 24670 12292 24722
rect 12236 24276 12292 24670
rect 12236 24210 12292 24220
rect 12348 24052 12404 24892
rect 12460 24724 12516 24734
rect 12460 24630 12516 24668
rect 12572 24164 12628 25340
rect 13524 25338 13580 25452
rect 13524 25286 13526 25338
rect 13578 25286 13580 25338
rect 13524 25274 13580 25286
rect 13468 25172 13524 25182
rect 12740 24948 12796 24958
rect 12740 24834 12796 24892
rect 12740 24782 12742 24834
rect 12794 24782 12796 24834
rect 12740 24770 12796 24782
rect 12908 24836 12964 24846
rect 12796 24164 12852 24174
rect 12572 24162 12852 24164
rect 12572 24110 12798 24162
rect 12850 24110 12852 24162
rect 12572 24108 12852 24110
rect 12796 24098 12852 24108
rect 12348 23950 12404 23996
rect 11564 23380 11620 23884
rect 12124 23886 12126 23938
rect 12178 23886 12180 23938
rect 11564 23324 11844 23380
rect 11788 22820 11844 23324
rect 12012 23044 12068 23054
rect 11452 22764 11844 22820
rect 11900 23042 12068 23044
rect 11900 22990 12014 23042
rect 12066 22990 12068 23042
rect 11900 22988 12068 22990
rect 11452 22372 11508 22764
rect 10892 22354 11228 22372
rect 10892 22316 11174 22354
rect 11172 22302 11174 22316
rect 11226 22302 11228 22354
rect 11172 22290 11228 22302
rect 11396 22335 11508 22372
rect 11396 22283 11398 22335
rect 11450 22316 11508 22335
rect 11450 22283 11452 22316
rect 11396 22271 11452 22283
rect 11564 22314 11620 22326
rect 11564 22262 11566 22314
rect 11618 22262 11620 22314
rect 10948 22148 11004 22158
rect 10948 22054 11004 22092
rect 11564 22148 11620 22262
rect 11788 22314 11844 22326
rect 11788 22262 11790 22314
rect 11842 22262 11844 22314
rect 11788 22260 11844 22262
rect 11788 22194 11844 22204
rect 11564 21476 11620 22092
rect 11788 21812 11844 21822
rect 11900 21812 11956 22988
rect 12012 22978 12068 22988
rect 12124 22820 12180 23886
rect 12236 23940 12292 23950
rect 12348 23938 12458 23950
rect 12348 23886 12404 23938
rect 12456 23886 12458 23938
rect 12348 23884 12458 23886
rect 12236 23846 12292 23884
rect 12402 23380 12458 23884
rect 12402 23314 12458 23324
rect 12684 23380 12740 23390
rect 12124 22764 12292 22820
rect 12068 22596 12124 22606
rect 12068 22502 12124 22540
rect 12236 22484 12292 22764
rect 12236 22418 12292 22428
rect 12460 22708 12516 22718
rect 12460 22370 12516 22652
rect 12460 22318 12462 22370
rect 12514 22318 12516 22370
rect 12460 22306 12516 22318
rect 11788 21810 11956 21812
rect 11788 21758 11790 21810
rect 11842 21758 11956 21810
rect 11788 21756 11956 21758
rect 12124 22260 12180 22270
rect 11788 21746 11844 21756
rect 12124 21586 12180 22204
rect 12124 21534 12126 21586
rect 12178 21534 12180 21586
rect 12124 21522 12180 21534
rect 11564 21410 11620 21420
rect 12684 21364 12740 23324
rect 12796 23156 12852 23166
rect 12796 23062 12852 23100
rect 12796 22484 12852 22494
rect 12796 21588 12852 22428
rect 12796 21522 12852 21532
rect 12684 21308 12852 21364
rect 11900 20972 12180 21028
rect 11788 20804 11844 20814
rect 11788 20710 11844 20748
rect 11508 20692 11564 20702
rect 11508 20690 11732 20692
rect 11508 20638 11510 20690
rect 11562 20638 11732 20690
rect 11508 20636 11732 20638
rect 11508 20626 11564 20636
rect 10332 19954 10388 19964
rect 10220 19906 10276 19918
rect 10220 19854 10222 19906
rect 10274 19854 10276 19906
rect 10220 19572 10276 19854
rect 11564 19908 11620 19918
rect 10220 19516 10724 19572
rect 9212 19350 9214 19402
rect 9266 19350 9268 19402
rect 10668 19458 10724 19516
rect 10668 19406 10670 19458
rect 10722 19406 10724 19458
rect 10668 19394 10724 19406
rect 9212 19338 9268 19350
rect 9100 19234 9156 19246
rect 9100 19182 9102 19234
rect 9154 19182 9156 19234
rect 9100 18676 9156 19182
rect 11004 19236 11060 19246
rect 11284 19236 11340 19246
rect 11004 19234 11340 19236
rect 11004 19182 11006 19234
rect 11058 19182 11286 19234
rect 11338 19182 11340 19234
rect 11004 19180 11340 19182
rect 11004 19170 11060 19180
rect 11284 19170 11340 19180
rect 11564 19234 11620 19852
rect 11564 19182 11566 19234
rect 11618 19182 11620 19234
rect 11564 19170 11620 19182
rect 11676 19236 11732 20636
rect 11900 19348 11956 20972
rect 12012 20802 12068 20814
rect 12012 20750 12014 20802
rect 12066 20750 12068 20802
rect 12012 19908 12068 20750
rect 12124 20804 12180 20972
rect 12684 20914 12740 20926
rect 12684 20862 12686 20914
rect 12738 20862 12740 20914
rect 12236 20804 12292 20814
rect 12124 20802 12292 20804
rect 12124 20750 12238 20802
rect 12290 20750 12292 20802
rect 12124 20748 12292 20750
rect 12236 20738 12292 20748
rect 12348 20746 12572 20760
rect 12348 20704 12518 20746
rect 12124 19908 12180 19918
rect 12348 19908 12404 20704
rect 12516 20694 12518 20704
rect 12570 20694 12572 20746
rect 12516 20682 12572 20694
rect 12516 20468 12572 20478
rect 12516 20074 12572 20412
rect 12516 20022 12518 20074
rect 12570 20022 12572 20074
rect 12684 20132 12740 20862
rect 12796 20468 12852 21308
rect 12796 20402 12852 20412
rect 12908 20244 12964 24780
rect 13244 24836 13300 24846
rect 13244 24749 13300 24780
rect 13244 24697 13246 24749
rect 13298 24697 13300 24749
rect 13244 24685 13300 24697
rect 13468 24388 13524 25116
rect 13692 25060 13748 25564
rect 14140 25282 14196 25294
rect 14140 25230 14142 25282
rect 14194 25230 14196 25282
rect 14140 25172 14196 25230
rect 14140 25106 14196 25116
rect 13692 24994 13748 25004
rect 14252 24500 14308 26236
rect 14700 25620 14756 28590
rect 14924 28642 14980 28924
rect 15428 28866 15484 29372
rect 15932 29418 15934 29470
rect 15986 29418 15988 29470
rect 14924 28590 14926 28642
rect 14978 28590 14980 28642
rect 14924 28578 14980 28590
rect 15036 28810 15092 28822
rect 15036 28758 15038 28810
rect 15090 28758 15092 28810
rect 15036 27972 15092 28758
rect 15428 28814 15430 28866
rect 15482 28814 15484 28866
rect 15428 28756 15484 28814
rect 15428 28690 15484 28700
rect 15708 28868 15764 28878
rect 15708 28642 15764 28812
rect 15708 28590 15710 28642
rect 15762 28590 15764 28642
rect 15708 28578 15764 28590
rect 15820 28644 15876 28654
rect 15820 28550 15876 28588
rect 14924 27916 15092 27972
rect 14812 27746 14868 27758
rect 14812 27694 14814 27746
rect 14866 27694 14868 27746
rect 14812 27186 14868 27694
rect 14812 27134 14814 27186
rect 14866 27134 14868 27186
rect 14812 27122 14868 27134
rect 14924 27059 14980 27916
rect 15932 27524 15988 29418
rect 16268 29428 16324 29438
rect 16268 29334 16324 29372
rect 16828 29428 16884 30156
rect 17052 30210 17108 30222
rect 17052 30158 17054 30210
rect 17106 30158 17108 30210
rect 17052 29540 17108 30158
rect 17724 30212 17780 30222
rect 17724 30118 17780 30156
rect 17332 30098 17388 30110
rect 17332 30046 17334 30098
rect 17386 30046 17388 30098
rect 17332 29652 17388 30046
rect 17836 29988 17892 30326
rect 18060 30212 18116 30222
rect 18060 30118 18116 30156
rect 17332 29586 17388 29596
rect 17612 29932 17892 29988
rect 18508 29988 18564 31052
rect 18620 30882 18676 30894
rect 18620 30830 18622 30882
rect 18674 30830 18676 30882
rect 18620 30212 18676 30830
rect 19404 30660 19460 31612
rect 20524 30994 20580 31836
rect 26160 31388 26424 31398
rect 26216 31332 26264 31388
rect 26320 31332 26368 31388
rect 26160 31322 26424 31332
rect 34476 31388 34740 31398
rect 34532 31332 34580 31388
rect 34636 31332 34684 31388
rect 34476 31322 34740 31332
rect 20524 30942 20526 30994
rect 20578 30942 20580 30994
rect 20524 30930 20580 30942
rect 21308 30994 21364 31006
rect 21308 30942 21310 30994
rect 21362 30942 21364 30994
rect 19404 30604 20020 30660
rect 19964 30434 20020 30604
rect 19964 30382 19966 30434
rect 20018 30382 20020 30434
rect 19964 30370 20020 30382
rect 20860 30324 20916 30334
rect 18844 30212 18900 30222
rect 18676 30210 18900 30212
rect 18676 30158 18846 30210
rect 18898 30158 18900 30210
rect 18676 30156 18900 30158
rect 18620 30118 18676 30156
rect 18844 30146 18900 30156
rect 18956 30212 19012 30222
rect 20300 30212 20356 30222
rect 17052 29474 17108 29484
rect 16828 29362 16884 29372
rect 16716 28644 16772 28654
rect 16716 27970 16772 28588
rect 17612 28642 17668 29932
rect 18508 29922 18564 29932
rect 17844 29820 18108 29830
rect 17900 29764 17948 29820
rect 18004 29764 18052 29820
rect 17844 29754 18108 29764
rect 18396 29652 18452 29662
rect 18396 29470 18452 29596
rect 18172 29426 18228 29438
rect 18172 29374 18174 29426
rect 18226 29374 18228 29426
rect 18396 29418 18398 29470
rect 18450 29418 18452 29470
rect 18396 29406 18452 29418
rect 18956 29426 19012 30156
rect 19720 30154 19776 30166
rect 19720 30102 19722 30154
rect 19774 30102 19776 30154
rect 20300 30118 20356 30156
rect 19720 29764 19776 30102
rect 20636 30100 20692 30110
rect 20636 30006 20692 30044
rect 19720 29708 19796 29764
rect 19628 29594 19684 29606
rect 19516 29540 19572 29550
rect 18172 29204 18228 29374
rect 18956 29374 18958 29426
rect 19010 29374 19012 29426
rect 18508 29316 18564 29326
rect 18508 29222 18564 29260
rect 18172 28756 18228 29148
rect 17612 28590 17614 28642
rect 17666 28590 17668 28642
rect 17612 28578 17668 28590
rect 17836 28754 18228 28756
rect 17836 28702 18174 28754
rect 18226 28702 18228 28754
rect 17836 28700 18228 28702
rect 17836 28642 17892 28700
rect 18172 28690 18228 28700
rect 17836 28590 17838 28642
rect 17890 28590 17892 28642
rect 17836 28578 17892 28590
rect 17332 28532 17388 28542
rect 16716 27918 16718 27970
rect 16770 27918 16772 27970
rect 16716 27906 16772 27918
rect 17164 28530 17388 28532
rect 17164 28478 17334 28530
rect 17386 28478 17388 28530
rect 17164 28476 17388 28478
rect 14924 27007 14926 27059
rect 14978 27007 14980 27059
rect 15260 27468 15988 27524
rect 15260 27074 15316 27468
rect 15260 27022 15262 27074
rect 15314 27022 15316 27074
rect 15260 27010 15316 27022
rect 16716 27076 16772 27086
rect 14924 26995 14980 27007
rect 16716 26982 16772 27020
rect 16940 27076 16996 27086
rect 17164 27076 17220 28476
rect 17332 28466 17388 28476
rect 18956 28420 19012 29374
rect 19180 29453 19236 29465
rect 19180 29401 19182 29453
rect 19234 29401 19236 29453
rect 19180 29316 19236 29401
rect 19516 29426 19572 29484
rect 19516 29374 19518 29426
rect 19570 29374 19572 29426
rect 19516 29362 19572 29374
rect 19628 29542 19630 29594
rect 19682 29542 19684 29594
rect 19628 29428 19684 29542
rect 19740 29540 19796 29708
rect 19740 29474 19796 29484
rect 20188 29652 20244 29662
rect 19628 29362 19684 29372
rect 19964 29426 20020 29438
rect 19964 29374 19966 29426
rect 20018 29374 20020 29426
rect 19180 29250 19236 29260
rect 19964 29204 20020 29374
rect 20188 29426 20244 29596
rect 20468 29540 20524 29550
rect 20468 29446 20524 29484
rect 20188 29374 20190 29426
rect 20242 29374 20244 29426
rect 20188 29362 20244 29374
rect 20748 29428 20804 29438
rect 20748 29334 20804 29372
rect 19964 29138 20020 29148
rect 20076 28756 20132 28766
rect 20076 28662 20132 28700
rect 20860 28642 20916 30268
rect 21308 30324 21364 30942
rect 21868 30994 21924 31006
rect 21868 30942 21870 30994
rect 21922 30942 21924 30994
rect 21308 30258 21364 30268
rect 21644 30324 21700 30334
rect 21868 30324 21924 30942
rect 25676 30996 25732 31006
rect 25676 30994 25844 30996
rect 25676 30942 25678 30994
rect 25730 30942 25844 30994
rect 25676 30940 25844 30942
rect 25676 30930 25732 30940
rect 22652 30884 22708 30894
rect 22652 30790 22708 30828
rect 24556 30882 24612 30894
rect 24556 30830 24558 30882
rect 24610 30830 24612 30882
rect 22002 30604 22266 30614
rect 22058 30548 22106 30604
rect 22162 30548 22210 30604
rect 22002 30538 22266 30548
rect 21700 30268 21924 30324
rect 21644 30210 21700 30268
rect 21644 30158 21646 30210
rect 21698 30158 21700 30210
rect 21644 30146 21700 30158
rect 22428 30210 22484 30222
rect 22428 30158 22430 30210
rect 22482 30158 22484 30210
rect 21084 29202 21140 29214
rect 21084 29150 21086 29202
rect 21138 29150 21140 29202
rect 21084 28756 21140 29150
rect 22002 29036 22266 29046
rect 22058 28980 22106 29036
rect 22162 28980 22210 29036
rect 22002 28970 22266 28980
rect 22428 28868 22484 30158
rect 24332 30212 24388 30222
rect 23996 30100 24052 30110
rect 22876 29988 22932 29998
rect 22876 29470 22932 29932
rect 23436 29594 23492 29606
rect 22652 29428 22708 29438
rect 22876 29418 22878 29470
rect 22930 29418 22932 29470
rect 23324 29540 23380 29550
rect 23324 29428 23380 29484
rect 22876 29406 22932 29418
rect 23212 29426 23380 29428
rect 22652 29334 22708 29372
rect 23212 29374 23326 29426
rect 23378 29374 23380 29426
rect 23212 29372 23380 29374
rect 22988 29316 23044 29326
rect 22988 29222 23044 29260
rect 22988 28868 23044 28878
rect 22428 28866 23044 28868
rect 22428 28814 22990 28866
rect 23042 28814 23044 28866
rect 22428 28812 23044 28814
rect 22988 28802 23044 28812
rect 21084 28690 21140 28700
rect 20860 28590 20862 28642
rect 20914 28590 20916 28642
rect 18956 28364 19236 28420
rect 17844 28252 18108 28262
rect 17900 28196 17948 28252
rect 18004 28196 18052 28252
rect 17844 28186 18108 28196
rect 17612 27186 17668 27198
rect 17612 27134 17614 27186
rect 17666 27134 17668 27186
rect 16940 27074 17220 27076
rect 16940 27022 16942 27074
rect 16994 27022 17166 27074
rect 17218 27022 17220 27074
rect 16940 27020 17220 27022
rect 16940 27010 16996 27020
rect 17164 27010 17220 27020
rect 17500 27076 17556 27086
rect 17500 27007 17502 27020
rect 17554 27007 17556 27020
rect 17500 26982 17556 27007
rect 16436 26964 16492 26974
rect 16268 26962 16492 26964
rect 16268 26910 16438 26962
rect 16490 26910 16492 26962
rect 16268 26908 16492 26910
rect 15988 26180 16044 26190
rect 15820 26178 16044 26180
rect 15820 26126 15990 26178
rect 16042 26126 16044 26178
rect 15820 26124 16044 26126
rect 14700 25554 14756 25564
rect 15260 25732 15316 25742
rect 14476 25508 14532 25518
rect 14476 25284 14532 25452
rect 14588 25506 14644 25518
rect 14588 25454 14590 25506
rect 14642 25454 14644 25506
rect 14588 25396 14644 25454
rect 14588 25330 14644 25340
rect 15260 25506 15316 25676
rect 15596 25620 15652 25630
rect 15596 25526 15652 25564
rect 15260 25454 15262 25506
rect 15314 25454 15316 25506
rect 15260 25396 15316 25454
rect 15260 25330 15316 25340
rect 15708 25508 15764 25518
rect 14476 25218 14532 25228
rect 14924 25282 14980 25294
rect 14924 25230 14926 25282
rect 14978 25230 14980 25282
rect 14140 24498 14308 24500
rect 14140 24446 14254 24498
rect 14306 24446 14308 24498
rect 14140 24444 14308 24446
rect 13468 24322 13524 24332
rect 13686 24332 13950 24342
rect 13742 24276 13790 24332
rect 13846 24276 13894 24332
rect 13686 24266 13950 24276
rect 13804 23910 13860 23922
rect 13804 23858 13806 23910
rect 13858 23858 13860 23910
rect 13468 23716 13524 23726
rect 13356 23604 13412 23614
rect 13356 23266 13412 23548
rect 13356 23214 13358 23266
rect 13410 23214 13412 23266
rect 13356 23202 13412 23214
rect 13020 23154 13076 23166
rect 13020 23102 13022 23154
rect 13074 23102 13076 23154
rect 13468 23154 13524 23660
rect 13020 22596 13076 23102
rect 13020 22530 13076 22540
rect 13188 23098 13244 23110
rect 13188 23046 13190 23098
rect 13242 23046 13244 23098
rect 13468 23102 13470 23154
rect 13522 23102 13524 23154
rect 13468 23090 13524 23102
rect 13804 23156 13860 23858
rect 14028 23156 14084 23166
rect 14140 23156 14196 24444
rect 14252 24434 14308 24444
rect 13860 23154 14196 23156
rect 13860 23102 14030 23154
rect 14082 23102 14196 23154
rect 13860 23100 14196 23102
rect 13804 23090 13860 23100
rect 14028 23090 14084 23100
rect 13188 22484 13244 23046
rect 13748 22932 13804 22942
rect 13748 22930 14084 22932
rect 13748 22878 13750 22930
rect 13802 22878 14084 22930
rect 13748 22876 14084 22878
rect 13748 22866 13804 22876
rect 13686 22764 13950 22774
rect 13742 22708 13790 22764
rect 13846 22708 13894 22764
rect 13686 22698 13950 22708
rect 14028 22596 14084 22876
rect 13804 22540 14084 22596
rect 13188 22428 13300 22484
rect 13132 21588 13188 21598
rect 13132 21494 13188 21532
rect 13244 21374 13300 22428
rect 13804 22370 13860 22540
rect 13804 22318 13806 22370
rect 13858 22318 13860 22370
rect 13804 22306 13860 22318
rect 14028 22372 14084 22382
rect 14028 22278 14084 22316
rect 13524 22260 13580 22270
rect 13524 22166 13580 22204
rect 14028 21588 14084 21598
rect 13244 21364 13356 21374
rect 13244 21362 13412 21364
rect 13244 21310 13302 21362
rect 13354 21310 13412 21362
rect 13244 21308 13412 21310
rect 13300 21298 13412 21308
rect 12684 20066 12740 20076
rect 12796 20188 12964 20244
rect 13020 20804 13076 20814
rect 12516 20010 12572 20022
rect 12012 19906 12404 19908
rect 12012 19854 12126 19906
rect 12178 19854 12404 19906
rect 12012 19852 12404 19854
rect 12684 19908 12740 19918
rect 12124 19842 12180 19852
rect 11900 19292 12180 19348
rect 11788 19236 11844 19246
rect 11676 19234 11844 19236
rect 11676 19182 11790 19234
rect 11842 19182 11844 19234
rect 11676 19180 11844 19182
rect 11788 19170 11844 19180
rect 9528 18844 9792 18854
rect 9584 18788 9632 18844
rect 9688 18788 9736 18844
rect 9528 18778 9792 18788
rect 9100 18610 9156 18620
rect 8988 18274 9044 18284
rect 11228 18340 11284 18350
rect 10892 17666 10948 17678
rect 10892 17614 10894 17666
rect 10946 17614 10948 17666
rect 10892 17556 10948 17614
rect 11228 17666 11284 18284
rect 12012 18228 12068 19292
rect 12124 19290 12180 19292
rect 12124 19238 12126 19290
rect 12178 19238 12180 19290
rect 12124 19226 12180 19238
rect 12236 19196 12292 19852
rect 12684 19814 12740 19852
rect 12796 19348 12852 20188
rect 12908 20020 12964 20030
rect 13020 20020 13076 20748
rect 13356 20356 13412 21298
rect 13686 21196 13950 21206
rect 13742 21140 13790 21196
rect 13846 21140 13894 21196
rect 13686 21130 13950 21140
rect 14028 20802 14084 21532
rect 14028 20750 14030 20802
rect 14082 20750 14084 20802
rect 14028 20738 14084 20750
rect 13356 20290 13412 20300
rect 13468 20132 13524 20142
rect 12908 20018 13076 20020
rect 12908 19966 12910 20018
rect 12962 19966 13076 20018
rect 12908 19964 13076 19966
rect 12908 19954 12964 19964
rect 13020 19796 13076 19964
rect 13020 19730 13076 19740
rect 13132 20046 13188 20058
rect 13132 19994 13134 20046
rect 13186 19994 13188 20046
rect 12236 19144 12238 19196
rect 12290 19144 12292 19196
rect 12236 19132 12292 19144
rect 12684 19292 12852 19348
rect 12012 17780 12068 18172
rect 12124 18900 12180 18910
rect 12124 17902 12180 18844
rect 12236 18450 12292 18462
rect 12236 18398 12238 18450
rect 12290 18398 12292 18450
rect 12236 18340 12292 18398
rect 12236 18274 12292 18284
rect 12348 18452 12404 18462
rect 12124 17890 12198 17902
rect 12124 17838 12144 17890
rect 12196 17838 12198 17890
rect 12124 17836 12198 17838
rect 12142 17826 12198 17836
rect 11228 17614 11230 17666
rect 11282 17614 11284 17666
rect 11900 17668 11956 17678
rect 11228 17602 11284 17614
rect 11396 17610 11452 17622
rect 10892 17490 10948 17500
rect 11396 17558 11398 17610
rect 11450 17558 11452 17610
rect 11900 17574 11956 17612
rect 10556 17444 10612 17454
rect 8764 17378 8820 17388
rect 10220 17442 10612 17444
rect 10220 17390 10558 17442
rect 10610 17390 10612 17442
rect 10220 17388 10612 17390
rect 9528 17276 9792 17286
rect 9584 17220 9632 17276
rect 9688 17220 9736 17276
rect 9528 17210 9792 17220
rect 8708 17108 8764 17118
rect 8092 16942 8094 16994
rect 8146 16942 8148 16994
rect 8092 16930 8148 16942
rect 8540 17106 8764 17108
rect 8540 17054 8710 17106
rect 8762 17054 8764 17106
rect 8540 17052 8764 17054
rect 4508 16210 4788 16212
rect 4508 16158 4510 16210
rect 4562 16158 4788 16210
rect 4508 16156 4788 16158
rect 5180 16604 5460 16660
rect 6188 16770 6244 16782
rect 6188 16718 6190 16770
rect 6242 16718 6244 16770
rect 4508 16146 4564 16156
rect 5180 16110 5236 16604
rect 5370 16492 5634 16502
rect 5426 16436 5474 16492
rect 5530 16436 5578 16492
rect 5370 16426 5634 16436
rect 4900 16100 4956 16110
rect 4900 15538 4956 16044
rect 5124 16100 5236 16110
rect 5180 16044 5236 16100
rect 5852 16100 5908 16110
rect 5124 16006 5180 16044
rect 4900 15486 4902 15538
rect 4954 15486 4956 15538
rect 4900 15474 4956 15486
rect 4284 15374 4286 15426
rect 4338 15374 4340 15426
rect 4284 15362 4340 15374
rect 2380 15204 2436 15214
rect 2380 15202 2660 15204
rect 2380 15150 2382 15202
rect 2434 15150 2660 15202
rect 2380 15148 2660 15150
rect 2380 15138 2436 15148
rect 2604 14868 2660 15148
rect 5370 14924 5634 14934
rect 5426 14868 5474 14924
rect 5530 14868 5578 14924
rect 2604 14812 3108 14868
rect 5370 14858 5634 14868
rect 3052 14754 3108 14812
rect 3052 14702 3054 14754
rect 3106 14702 3108 14754
rect 3052 14690 3108 14702
rect 3388 14532 3444 14542
rect 3388 14438 3444 14476
rect 2940 13860 2996 13870
rect 2940 13746 2996 13804
rect 3612 13860 3668 13870
rect 3612 13802 3668 13804
rect 2940 13694 2942 13746
rect 2994 13694 2996 13746
rect 2940 13682 2996 13694
rect 3052 13748 3108 13758
rect 3612 13750 3614 13802
rect 3666 13750 3668 13802
rect 4956 13860 5012 13870
rect 3612 13738 3668 13750
rect 3836 13748 3892 13758
rect 2828 13636 2884 13646
rect 2660 13524 2716 13534
rect 2268 13458 2324 13468
rect 2380 13522 2716 13524
rect 2380 13470 2662 13522
rect 2714 13470 2716 13522
rect 2380 13468 2716 13470
rect 2380 12962 2436 13468
rect 2660 13458 2716 13468
rect 2828 13300 2884 13580
rect 2380 12910 2382 12962
rect 2434 12910 2436 12962
rect 2380 12898 2436 12910
rect 2604 13244 2884 13300
rect 2604 12962 2660 13244
rect 3052 13188 3108 13692
rect 4844 13746 4900 13758
rect 3836 13654 3892 13692
rect 4228 13690 4284 13702
rect 4060 13636 4116 13646
rect 4060 13542 4116 13580
rect 4228 13638 4230 13690
rect 4282 13638 4284 13690
rect 2604 12910 2606 12962
rect 2658 12910 2660 12962
rect 2604 12898 2660 12910
rect 2716 13130 2772 13142
rect 2716 13078 2718 13130
rect 2770 13078 2772 13130
rect 2716 12964 2772 13078
rect 2716 12898 2772 12908
rect 2828 13132 3108 13188
rect 3612 13524 3668 13534
rect 2828 12290 2884 13132
rect 3612 13074 3668 13468
rect 4228 13412 4284 13638
rect 4452 13690 4508 13702
rect 4452 13638 4454 13690
rect 4506 13638 4508 13690
rect 4844 13694 4846 13746
rect 4898 13694 4900 13746
rect 4452 13636 4508 13638
rect 4452 13570 4508 13580
rect 4620 13634 4676 13646
rect 4620 13582 4622 13634
rect 4674 13582 4676 13634
rect 3612 13022 3614 13074
rect 3666 13022 3668 13074
rect 3612 13010 3668 13022
rect 4060 13356 4284 13412
rect 3052 12964 3108 12974
rect 2828 12238 2830 12290
rect 2882 12238 2884 12290
rect 2828 12226 2884 12238
rect 2940 12962 3108 12964
rect 2940 12910 3054 12962
rect 3106 12910 3108 12962
rect 2940 12908 3108 12910
rect 2660 12180 2716 12190
rect 2660 12086 2716 12124
rect 2716 11172 2772 11182
rect 2716 10386 2772 11116
rect 2716 10334 2718 10386
rect 2770 10334 2772 10386
rect 2716 9828 2772 10334
rect 2940 10388 2996 12908
rect 3052 12898 3108 12908
rect 3388 12964 3444 12974
rect 3836 12964 3892 12974
rect 3388 12870 3444 12908
rect 3724 12962 3892 12964
rect 3724 12910 3838 12962
rect 3890 12910 3892 12962
rect 3724 12908 3892 12910
rect 3276 12206 3332 12218
rect 3052 12178 3108 12190
rect 3052 12126 3054 12178
rect 3106 12126 3108 12178
rect 3052 11956 3108 12126
rect 3276 12154 3278 12206
rect 3330 12154 3332 12206
rect 3276 12068 3332 12154
rect 3276 12002 3332 12012
rect 3052 11890 3108 11900
rect 3556 11620 3612 11630
rect 3724 11620 3780 12908
rect 3836 12898 3892 12908
rect 4060 12964 4116 13356
rect 4620 13300 4676 13582
rect 4060 12898 4116 12908
rect 4284 13244 4676 13300
rect 4284 12962 4340 13244
rect 4284 12910 4286 12962
rect 4338 12910 4340 12962
rect 4284 12898 4340 12910
rect 4620 13130 4676 13142
rect 4620 13078 4622 13130
rect 4674 13078 4676 13130
rect 4620 12404 4676 13078
rect 4004 12348 4676 12404
rect 4732 12962 4788 12974
rect 4732 12910 4734 12962
rect 4786 12910 4788 12962
rect 4732 12404 4788 12910
rect 4004 12234 4116 12348
rect 4732 12338 4788 12348
rect 3836 12180 3892 12190
rect 4004 12182 4006 12234
rect 4058 12182 4116 12234
rect 4004 12170 4116 12182
rect 3836 12086 3892 12124
rect 4060 11956 4116 12170
rect 4284 12180 4340 12190
rect 4508 12180 4564 12190
rect 4844 12180 4900 13694
rect 4340 12124 4452 12180
rect 4284 12114 4340 12124
rect 4060 11900 4172 11956
rect 3556 11618 3780 11620
rect 3556 11566 3558 11618
rect 3610 11566 3780 11618
rect 3556 11564 3780 11566
rect 3836 11844 3892 11854
rect 3556 11554 3612 11564
rect 3836 11394 3892 11788
rect 3836 11342 3838 11394
rect 3890 11342 3892 11394
rect 4116 11450 4172 11900
rect 4116 11398 4118 11450
rect 4170 11398 4172 11450
rect 4116 11386 4172 11398
rect 4284 11394 4340 11406
rect 3836 11330 3892 11342
rect 4284 11342 4286 11394
rect 4338 11342 4340 11394
rect 3948 11282 4004 11294
rect 3948 11230 3950 11282
rect 4002 11230 4004 11282
rect 3220 11172 3276 11182
rect 3220 11078 3276 11116
rect 3724 11060 3780 11070
rect 3052 10612 3108 10622
rect 3052 10518 3108 10556
rect 3612 10610 3668 10622
rect 3612 10558 3614 10610
rect 3666 10558 3668 10610
rect 2940 10332 3164 10388
rect 3108 10050 3164 10332
rect 3108 9998 3110 10050
rect 3162 9998 3164 10050
rect 3108 9986 3164 9998
rect 3332 10386 3388 10398
rect 3332 10334 3334 10386
rect 3386 10334 3388 10386
rect 3332 9940 3388 10334
rect 3612 10164 3668 10558
rect 3612 10098 3668 10108
rect 3332 9884 3556 9940
rect 3500 9828 3556 9884
rect 3500 9791 3612 9828
rect 2716 9614 2772 9772
rect 3388 9770 3444 9782
rect 3500 9772 3558 9791
rect 3276 9716 3332 9726
rect 2716 9602 2828 9614
rect 2716 9550 2774 9602
rect 2826 9550 2828 9602
rect 2716 9538 2828 9550
rect 3052 9604 3108 9614
rect 2492 8148 2548 8158
rect 2492 5684 2548 8092
rect 2492 5590 2548 5628
rect 2604 7476 2660 7486
rect 2604 5684 2660 7420
rect 2716 6814 2772 9538
rect 3052 9070 3108 9548
rect 3052 9018 3054 9070
rect 3106 9018 3108 9070
rect 3052 8484 3108 9018
rect 3276 9042 3332 9660
rect 3388 9718 3390 9770
rect 3442 9718 3444 9770
rect 3556 9739 3558 9772
rect 3610 9739 3612 9791
rect 3556 9727 3612 9739
rect 3388 9380 3444 9718
rect 3724 9604 3780 11004
rect 3836 10610 3892 10622
rect 3836 10558 3838 10610
rect 3890 10558 3892 10610
rect 3836 10388 3892 10558
rect 3836 10322 3892 10332
rect 3948 10052 4004 11230
rect 4284 11172 4340 11342
rect 4284 11106 4340 11116
rect 4172 10388 4228 10398
rect 4396 10388 4452 12124
rect 4508 12086 4564 12124
rect 4750 12124 4900 12180
rect 4956 12180 5012 13804
rect 5180 13784 5236 13796
rect 5180 13732 5182 13784
rect 5234 13732 5236 13784
rect 5180 13076 5236 13732
rect 5370 13356 5634 13366
rect 5426 13300 5474 13356
rect 5530 13300 5578 13356
rect 5370 13290 5634 13300
rect 5628 13076 5684 13086
rect 5180 13074 5684 13076
rect 5180 13022 5630 13074
rect 5682 13022 5684 13074
rect 5180 13020 5684 13022
rect 5628 13010 5684 13020
rect 5740 13076 5796 13086
rect 5068 12962 5124 12974
rect 5068 12910 5070 12962
rect 5122 12910 5124 12962
rect 5068 12852 5124 12910
rect 5740 12947 5796 13020
rect 5740 12895 5742 12947
rect 5794 12895 5796 12947
rect 5740 12883 5796 12895
rect 5068 12786 5124 12796
rect 5852 12740 5908 16044
rect 6188 14756 6244 16718
rect 6300 15426 6356 16828
rect 8540 16772 8596 17052
rect 8708 17042 8764 17052
rect 7868 16100 7924 16110
rect 8540 16100 8596 16716
rect 9436 16882 9492 16894
rect 9436 16830 9438 16882
rect 9490 16830 9492 16882
rect 9436 16772 9492 16830
rect 10220 16882 10276 17388
rect 10556 17378 10612 17388
rect 11396 17108 11452 17558
rect 11340 17052 11452 17108
rect 10220 16830 10222 16882
rect 10274 16830 10276 16882
rect 10220 16818 10276 16830
rect 10444 16884 10500 16894
rect 9436 16706 9492 16716
rect 10444 16212 10500 16828
rect 11340 16884 11396 17052
rect 12012 16996 12068 17724
rect 12124 16996 12180 17006
rect 12012 16994 12180 16996
rect 12012 16942 12126 16994
rect 12178 16942 12180 16994
rect 12012 16940 12180 16942
rect 12124 16930 12180 16940
rect 11340 16818 11396 16828
rect 10556 16212 10612 16222
rect 10444 16210 10612 16212
rect 10444 16158 10558 16210
rect 10610 16158 10612 16210
rect 10444 16156 10612 16158
rect 10556 16146 10612 16156
rect 7924 16044 8036 16100
rect 7868 16006 7924 16044
rect 6300 15374 6302 15426
rect 6354 15374 6356 15426
rect 6300 15362 6356 15374
rect 7980 15316 8036 16044
rect 8540 16034 8596 16044
rect 8652 16098 8708 16110
rect 8652 16046 8654 16098
rect 8706 16046 8708 16098
rect 6188 14690 6244 14700
rect 6748 14756 6804 14766
rect 6748 14662 6804 14700
rect 7308 14756 7364 14766
rect 7308 14662 7364 14700
rect 6412 14530 6468 14542
rect 7644 14532 7700 14542
rect 6412 14478 6414 14530
rect 6466 14478 6468 14530
rect 6412 13198 6468 14478
rect 7532 14530 7700 14532
rect 7532 14478 7646 14530
rect 7698 14478 7700 14530
rect 7532 14476 7700 14478
rect 7084 13636 7140 13646
rect 6412 13186 6524 13198
rect 6412 13134 6470 13186
rect 6522 13134 6524 13186
rect 6412 13132 6524 13134
rect 6468 13122 6524 13132
rect 5964 12964 6020 12974
rect 5964 12870 6020 12908
rect 6300 12964 6356 12974
rect 6972 12964 7028 12974
rect 5852 12684 6020 12740
rect 5516 12516 5572 12526
rect 5292 12180 5348 12190
rect 4956 12178 5348 12180
rect 4956 12126 5294 12178
rect 5346 12126 5348 12178
rect 4956 12124 5348 12126
rect 4750 12066 4806 12124
rect 4750 12014 4752 12066
rect 4804 12014 4806 12066
rect 4750 12002 4806 12014
rect 4172 10386 4452 10388
rect 4172 10334 4174 10386
rect 4226 10334 4452 10386
rect 4172 10332 4452 10334
rect 4172 10322 4228 10332
rect 3948 9986 4004 9996
rect 3836 9828 3892 9838
rect 4284 9828 4340 9838
rect 3836 9746 3838 9772
rect 3890 9746 3892 9772
rect 4004 9826 4340 9828
rect 4004 9810 4286 9826
rect 4004 9758 4006 9810
rect 4058 9774 4286 9810
rect 4338 9774 4340 9826
rect 4058 9772 4340 9774
rect 4058 9758 4060 9772
rect 4004 9746 4060 9758
rect 3836 9734 3892 9746
rect 3724 9538 3780 9548
rect 3388 9324 4116 9380
rect 3276 8990 3278 9042
rect 3330 8990 3332 9042
rect 3276 8978 3332 8990
rect 3668 9156 3724 9166
rect 3668 9098 3724 9100
rect 3668 9046 3670 9098
rect 3722 9046 3724 9098
rect 3500 8932 3556 8942
rect 3388 8930 3556 8932
rect 3388 8878 3502 8930
rect 3554 8878 3556 8930
rect 3388 8876 3556 8878
rect 3388 8708 3444 8876
rect 3500 8866 3556 8876
rect 3052 8418 3108 8428
rect 3276 8652 3444 8708
rect 3276 8230 3332 8652
rect 3668 8428 3724 9046
rect 4060 8930 4116 9324
rect 4060 8878 4062 8930
rect 4114 8878 4116 8930
rect 4060 8866 4116 8878
rect 4172 9057 4228 9069
rect 4172 9005 4174 9057
rect 4226 9005 4228 9057
rect 4172 8708 4228 9005
rect 3052 8202 3108 8214
rect 3052 8150 3054 8202
rect 3106 8150 3108 8202
rect 3276 8178 3278 8230
rect 3330 8178 3332 8230
rect 3276 8166 3332 8178
rect 3388 8372 3724 8428
rect 4060 8652 4228 8708
rect 3892 8372 3948 8382
rect 3052 8148 3108 8150
rect 3052 8082 3108 8092
rect 3164 7476 3220 7486
rect 3388 7476 3444 8372
rect 3892 8314 3948 8316
rect 3892 8262 3894 8314
rect 3946 8262 3948 8314
rect 3892 8250 3948 8262
rect 3724 8148 3780 8158
rect 3164 7474 3444 7476
rect 3164 7422 3166 7474
rect 3218 7422 3444 7474
rect 3164 7420 3444 7422
rect 3612 8146 3780 8148
rect 3612 8094 3726 8146
rect 3778 8094 3780 8146
rect 3612 8092 3780 8094
rect 3164 7410 3220 7420
rect 3612 7364 3668 8092
rect 3724 8082 3780 8092
rect 4060 8148 4116 8652
rect 4172 8484 4228 8494
rect 4172 8426 4228 8428
rect 4172 8374 4174 8426
rect 4226 8374 4228 8426
rect 4172 8362 4228 8374
rect 4284 8428 4340 9772
rect 4396 9716 4452 10332
rect 4508 11396 4564 11406
rect 4508 10610 4564 11340
rect 4732 11284 4788 11294
rect 4732 10722 4788 11228
rect 4956 11060 5012 12124
rect 5292 12114 5348 12124
rect 5516 12178 5572 12460
rect 5516 12126 5518 12178
rect 5570 12126 5572 12178
rect 5516 12114 5572 12126
rect 5180 12010 5236 12022
rect 4956 10994 5012 11004
rect 5068 11956 5124 11966
rect 5068 10836 5124 11900
rect 5180 11958 5182 12010
rect 5234 11958 5236 12010
rect 5180 11844 5236 11958
rect 5180 11778 5236 11788
rect 5370 11788 5634 11798
rect 5426 11732 5474 11788
rect 5530 11732 5578 11788
rect 5370 11722 5634 11732
rect 5180 10836 5236 10846
rect 5068 10780 5180 10836
rect 4732 10670 4734 10722
rect 4786 10670 4788 10722
rect 4732 10658 4788 10670
rect 5180 10666 5236 10780
rect 4870 10643 4926 10655
rect 4508 10558 4510 10610
rect 4562 10558 4564 10610
rect 4508 10164 4564 10558
rect 4508 10098 4564 10108
rect 4620 10612 4676 10622
rect 4620 9828 4676 10556
rect 4870 10591 4872 10643
rect 4924 10591 4926 10643
rect 5180 10614 5182 10666
rect 5234 10614 5236 10666
rect 5852 10724 5908 10734
rect 5852 10666 5908 10668
rect 5180 10602 5236 10614
rect 5628 10643 5684 10655
rect 4870 10276 4926 10591
rect 5628 10591 5630 10643
rect 5682 10591 5684 10643
rect 5852 10614 5854 10666
rect 5906 10614 5908 10666
rect 5852 10602 5908 10614
rect 4732 10220 4926 10276
rect 5068 10388 5124 10398
rect 4732 9994 4788 10220
rect 5068 10164 5124 10332
rect 5628 10388 5684 10591
rect 5964 10500 6020 12684
rect 6300 12234 6356 12908
rect 6748 12906 6804 12918
rect 6748 12854 6750 12906
rect 6802 12854 6804 12906
rect 6972 12882 6974 12908
rect 7026 12882 7028 12908
rect 6972 12870 7028 12882
rect 6300 12182 6302 12234
rect 6354 12182 6356 12234
rect 5628 10322 5684 10332
rect 5852 10444 6020 10500
rect 6188 11732 6244 11742
rect 4732 9942 4734 9994
rect 4786 9942 4788 9994
rect 4732 9930 4788 9942
rect 4956 10108 5124 10164
rect 5370 10220 5634 10230
rect 5426 10164 5474 10220
rect 5530 10164 5578 10220
rect 5370 10154 5634 10164
rect 4844 9828 4900 9838
rect 4620 9826 4788 9828
rect 4620 9774 4622 9826
rect 4674 9774 4788 9826
rect 4620 9772 4788 9774
rect 4620 9762 4676 9772
rect 4396 9650 4452 9660
rect 4620 9604 4676 9614
rect 4508 9042 4564 9054
rect 4508 8990 4510 9042
rect 4562 8990 4564 9042
rect 4508 8820 4564 8990
rect 4508 8754 4564 8764
rect 4284 8372 4452 8428
rect 4284 8260 4340 8270
rect 4284 8166 4340 8204
rect 4060 8082 4116 8092
rect 3724 7476 3780 7486
rect 4284 7476 4340 7486
rect 3724 7474 4340 7476
rect 3724 7422 3726 7474
rect 3778 7422 4286 7474
rect 4338 7422 4340 7474
rect 3724 7420 4340 7422
rect 3724 7410 3780 7420
rect 4284 7410 4340 7420
rect 2940 7306 2996 7318
rect 2940 7254 2942 7306
rect 2994 7254 2996 7306
rect 2716 6804 2828 6814
rect 2716 6748 2772 6804
rect 2772 6690 2828 6748
rect 2772 6638 2774 6690
rect 2826 6638 2828 6690
rect 2772 6626 2828 6638
rect 2940 6020 2996 7254
rect 3388 7308 3668 7364
rect 3108 6692 3164 6702
rect 3108 6598 3164 6636
rect 3388 6662 3444 7308
rect 3388 6610 3390 6662
rect 3442 6610 3444 6662
rect 3948 6804 4004 6814
rect 4396 6804 4452 8372
rect 4508 8258 4564 8270
rect 4508 8206 4510 8258
rect 4562 8206 4564 8258
rect 4508 7698 4564 8206
rect 4508 7646 4510 7698
rect 4562 7646 4564 7698
rect 4508 7634 4564 7646
rect 4620 7474 4676 9548
rect 4732 8372 4788 9772
rect 4732 8306 4788 8316
rect 4620 7422 4622 7474
rect 4674 7422 4676 7474
rect 4620 7410 4676 7422
rect 4732 7698 4788 7710
rect 4732 7646 4734 7698
rect 4786 7646 4788 7698
rect 4396 6748 4564 6804
rect 3388 6598 3444 6610
rect 3612 6634 3668 6646
rect 3500 6580 3556 6590
rect 2940 5954 2996 5964
rect 3108 6468 3164 6478
rect 3108 6018 3164 6412
rect 3500 6020 3556 6524
rect 3612 6582 3614 6634
rect 3666 6582 3668 6634
rect 3612 6244 3668 6582
rect 3836 6634 3892 6646
rect 3836 6582 3838 6634
rect 3890 6582 3892 6634
rect 3836 6468 3892 6582
rect 3948 6634 4004 6748
rect 3948 6582 3950 6634
rect 4002 6582 4004 6634
rect 4228 6692 4284 6702
rect 4228 6598 4284 6636
rect 3948 6468 4004 6582
rect 4396 6578 4452 6590
rect 4396 6526 4398 6578
rect 4450 6526 4452 6578
rect 4060 6468 4116 6478
rect 3948 6412 4060 6468
rect 3836 6402 3892 6412
rect 4060 6402 4116 6412
rect 3612 6178 3668 6188
rect 3724 6356 3780 6366
rect 3108 5966 3110 6018
rect 3162 5966 3164 6018
rect 3108 5954 3164 5966
rect 3388 5964 3556 6020
rect 3612 6020 3668 6030
rect 3388 5962 3444 5964
rect 2828 5908 2884 5918
rect 3388 5910 3390 5962
rect 3442 5910 3444 5962
rect 3388 5908 3444 5910
rect 2828 5814 2884 5852
rect 3276 5852 3388 5908
rect 3612 5962 3668 5964
rect 3612 5910 3614 5962
rect 3666 5910 3668 5962
rect 3612 5898 3668 5910
rect 2604 5628 2828 5684
rect 1596 4340 1652 4350
rect 1596 4246 1652 4284
rect 2380 4340 2436 4350
rect 2604 4340 2660 5628
rect 2772 5346 2828 5628
rect 2772 5294 2774 5346
rect 2826 5294 2828 5346
rect 2772 5282 2828 5294
rect 3276 5346 3332 5852
rect 3388 5832 3444 5852
rect 3276 5294 3278 5346
rect 3330 5294 3332 5346
rect 3276 5282 3332 5294
rect 2940 5124 2996 5134
rect 2940 5030 2996 5068
rect 3612 5124 3668 5134
rect 3724 5124 3780 6300
rect 4396 6244 4452 6526
rect 3836 6188 4452 6244
rect 4508 6244 4564 6748
rect 4732 6356 4788 7646
rect 4732 6290 4788 6300
rect 4508 6188 4620 6244
rect 3836 5962 3892 6188
rect 3836 5910 3838 5962
rect 3890 5910 3892 5962
rect 4172 6020 4228 6030
rect 4564 6020 4620 6188
rect 4844 6132 4900 9772
rect 4956 9604 5012 10108
rect 5740 10052 5796 10062
rect 5740 9994 5796 9996
rect 5740 9942 5742 9994
rect 5794 9942 5796 9994
rect 5740 9930 5796 9942
rect 4956 9538 5012 9548
rect 5740 9826 5796 9838
rect 5740 9774 5742 9826
rect 5794 9774 5796 9826
rect 5068 9268 5124 9278
rect 4956 8036 5012 8046
rect 4956 6652 5012 7980
rect 5068 6746 5124 9212
rect 5740 9268 5796 9774
rect 5740 9202 5796 9212
rect 5370 8652 5634 8662
rect 5426 8596 5474 8652
rect 5530 8596 5578 8652
rect 5370 8586 5634 8596
rect 5852 8428 5908 10444
rect 6076 10052 6132 10062
rect 5964 9828 6020 9838
rect 5964 9734 6020 9772
rect 6076 9098 6132 9996
rect 6076 9046 6078 9098
rect 6130 9046 6132 9098
rect 6188 9156 6244 11676
rect 6300 9380 6356 12182
rect 6524 12516 6580 12526
rect 6748 12516 6804 12854
rect 6748 12460 7028 12516
rect 6524 12234 6580 12460
rect 6524 12182 6526 12234
rect 6578 12182 6580 12234
rect 6524 12170 6580 12182
rect 6860 12292 6916 12302
rect 6748 11844 6804 11854
rect 6748 9604 6804 11788
rect 6748 9538 6804 9548
rect 6300 9324 6748 9380
rect 6188 9090 6244 9100
rect 6692 9098 6748 9324
rect 6076 9034 6132 9046
rect 6300 9042 6356 9054
rect 5740 8372 5908 8428
rect 6300 8990 6302 9042
rect 6354 8990 6356 9042
rect 6300 8484 6356 8990
rect 6524 9044 6580 9054
rect 6692 9046 6694 9098
rect 6746 9046 6748 9098
rect 6692 9044 6748 9046
rect 6692 8988 6804 9044
rect 6524 8950 6580 8988
rect 6300 8418 6356 8428
rect 6636 8820 6692 8830
rect 5370 7084 5634 7094
rect 5426 7028 5474 7084
rect 5530 7028 5578 7084
rect 5370 7018 5634 7028
rect 5068 6694 5070 6746
rect 5122 6694 5124 6746
rect 5068 6682 5124 6694
rect 5516 6692 5572 6702
rect 4956 6600 4958 6652
rect 5010 6600 5012 6652
rect 4956 6588 5012 6600
rect 5516 6598 5572 6636
rect 4844 6066 4900 6076
rect 5236 6020 5292 6030
rect 4564 5964 4676 6020
rect 3836 5898 3892 5910
rect 3948 5941 4004 5953
rect 3948 5889 3950 5941
rect 4002 5889 4004 5941
rect 3948 5796 4004 5889
rect 3948 5730 4004 5740
rect 3836 5124 3892 5134
rect 3724 5122 3892 5124
rect 3724 5070 3838 5122
rect 3890 5070 3892 5122
rect 3724 5068 3892 5070
rect 3612 4676 3668 5068
rect 3836 5058 3892 5068
rect 4172 5122 4228 5964
rect 4172 5070 4174 5122
rect 4226 5070 4228 5122
rect 4172 5058 4228 5070
rect 4284 5290 4340 5302
rect 4284 5238 4286 5290
rect 4338 5238 4340 5290
rect 4284 5124 4340 5238
rect 4284 5058 4340 5068
rect 3612 4620 4452 4676
rect 4284 4452 4340 4462
rect 4284 4358 4340 4396
rect 2380 4338 2660 4340
rect 2380 4286 2382 4338
rect 2434 4286 2660 4338
rect 2380 4284 2660 4286
rect 2380 4274 2436 4284
rect 3612 4228 3668 4238
rect 3612 800 3668 4172
rect 4396 3722 4452 4620
rect 4620 4452 4676 5964
rect 5236 5926 5292 5964
rect 4732 5908 4788 5918
rect 4956 5908 5012 5918
rect 4732 5814 4788 5852
rect 4844 5906 5012 5908
rect 4844 5854 4958 5906
rect 5010 5854 5012 5906
rect 4844 5852 5012 5854
rect 4732 5124 4788 5134
rect 4844 5124 4900 5852
rect 4956 5842 5012 5852
rect 5370 5516 5634 5526
rect 5426 5460 5474 5516
rect 5530 5460 5578 5516
rect 5370 5450 5634 5460
rect 4956 5348 5012 5358
rect 4956 5290 5012 5292
rect 4956 5238 4958 5290
rect 5010 5238 5012 5290
rect 4956 5226 5012 5238
rect 4788 5068 4900 5124
rect 4956 5124 5012 5134
rect 4732 5030 4788 5068
rect 4956 5030 5012 5068
rect 4620 4340 4676 4396
rect 5608 4564 5664 4574
rect 5608 4394 5664 4508
rect 4732 4340 4788 4350
rect 4620 4338 4788 4340
rect 4620 4286 4734 4338
rect 4786 4286 4788 4338
rect 5608 4342 5610 4394
rect 5662 4342 5664 4394
rect 5608 4330 5664 4342
rect 5740 4340 5796 8372
rect 5852 7924 5908 7934
rect 5852 6914 5908 7868
rect 5852 6862 5854 6914
rect 5906 6862 5908 6914
rect 5852 6850 5908 6862
rect 6636 6692 6692 8764
rect 6748 8596 6804 8988
rect 6748 8530 6804 8540
rect 6748 8260 6804 8270
rect 6748 6916 6804 8204
rect 6748 6850 6804 6860
rect 6636 6636 6804 6692
rect 5852 6244 5908 6254
rect 5852 5794 5908 6188
rect 5852 5742 5854 5794
rect 5906 5742 5908 5794
rect 5852 5730 5908 5742
rect 6246 5906 6302 5918
rect 6246 5854 6248 5906
rect 6300 5854 6302 5906
rect 6246 5684 6302 5854
rect 6412 5908 6468 5918
rect 6412 5814 6468 5852
rect 6524 5906 6580 5918
rect 6524 5854 6526 5906
rect 6578 5854 6580 5906
rect 6246 5618 6302 5628
rect 6412 5236 6468 5246
rect 6524 5236 6580 5854
rect 6748 5460 6804 6636
rect 6860 5572 6916 12236
rect 6972 12290 7028 12460
rect 6972 12238 6974 12290
rect 7026 12238 7028 12290
rect 6972 12226 7028 12238
rect 7084 12292 7140 13580
rect 7364 12927 7420 12939
rect 7196 12906 7252 12918
rect 7196 12854 7198 12906
rect 7250 12854 7252 12906
rect 7364 12875 7366 12927
rect 7418 12926 7420 12927
rect 7418 12875 7476 12926
rect 7364 12863 7476 12875
rect 7196 12404 7252 12854
rect 7196 12348 7364 12404
rect 7084 12236 7196 12292
rect 7140 12122 7196 12236
rect 7140 12070 7142 12122
rect 7194 12070 7196 12122
rect 6972 11956 7028 11966
rect 6972 11359 7028 11900
rect 7140 11844 7196 12070
rect 7140 11778 7196 11788
rect 7308 11508 7364 12348
rect 7420 11956 7476 12863
rect 7532 12628 7588 14476
rect 7644 14466 7700 14476
rect 7868 14532 7924 14542
rect 7980 14532 8036 15260
rect 8204 15202 8260 15214
rect 8204 15150 8206 15202
rect 8258 15150 8260 15202
rect 8204 14756 8260 15150
rect 8204 14690 8260 14700
rect 7868 14530 8036 14532
rect 7868 14478 7870 14530
rect 7922 14478 8036 14530
rect 7868 14476 8036 14478
rect 7868 14466 7924 14476
rect 7756 13188 7812 13198
rect 7644 13130 7700 13142
rect 7644 13078 7646 13130
rect 7698 13078 7700 13130
rect 7644 12964 7700 13078
rect 7644 12898 7700 12908
rect 7756 12962 7812 13132
rect 7756 12910 7758 12962
rect 7810 12910 7812 12962
rect 7756 12898 7812 12910
rect 8432 12924 8488 12936
rect 8432 12872 8434 12924
rect 8486 12872 8488 12924
rect 8432 12628 8488 12872
rect 7532 12572 7700 12628
rect 7532 12292 7588 12302
rect 7532 12211 7588 12236
rect 7532 12159 7534 12211
rect 7586 12159 7588 12211
rect 7532 12147 7588 12159
rect 7420 11900 7588 11956
rect 6972 11307 6974 11359
rect 7026 11307 7028 11359
rect 7196 11452 7364 11508
rect 7420 11508 7476 11518
rect 6972 11295 7028 11307
rect 7084 11338 7140 11350
rect 7084 11286 7086 11338
rect 7138 11286 7140 11338
rect 7084 11284 7140 11286
rect 7084 11218 7140 11228
rect 7084 9828 7140 9838
rect 7084 9156 7140 9772
rect 7084 9090 7140 9100
rect 7084 8596 7140 8606
rect 7084 8370 7140 8540
rect 7084 8318 7086 8370
rect 7138 8318 7140 8370
rect 7084 8306 7140 8318
rect 7196 6804 7252 11452
rect 7420 11396 7476 11452
rect 7308 11366 7476 11396
rect 7308 11314 7310 11366
rect 7362 11340 7476 11366
rect 7362 11314 7364 11340
rect 7308 11302 7364 11314
rect 7532 11338 7588 11900
rect 7532 11286 7534 11338
rect 7586 11286 7588 11338
rect 7532 10948 7588 11286
rect 7420 10892 7588 10948
rect 7308 9826 7364 9838
rect 7308 9774 7310 9826
rect 7362 9774 7364 9826
rect 7308 9492 7364 9774
rect 7308 9426 7364 9436
rect 7308 9080 7364 9092
rect 7308 9044 7310 9080
rect 7362 9044 7364 9080
rect 7308 8978 7364 8988
rect 7420 8428 7476 10892
rect 7644 10734 7700 12572
rect 8432 12562 8488 12572
rect 8652 12404 8708 16046
rect 11172 15876 11228 15886
rect 9528 15708 9792 15718
rect 9584 15652 9632 15708
rect 9688 15652 9736 15708
rect 9528 15642 9792 15652
rect 8988 15316 9044 15326
rect 8988 13982 9044 15260
rect 9772 15316 9828 15326
rect 9772 15222 9828 15260
rect 11172 15316 11228 15820
rect 12348 15540 12404 18396
rect 12460 18450 12516 18462
rect 12460 18398 12462 18450
rect 12514 18398 12516 18450
rect 12460 17444 12516 18398
rect 12684 18452 12740 19292
rect 12964 19236 13020 19246
rect 12964 19142 13020 19180
rect 12796 19122 12852 19134
rect 12796 19070 12798 19122
rect 12850 19070 12852 19122
rect 12796 18676 12852 19070
rect 13132 18900 13188 19994
rect 13468 19460 13524 20076
rect 13860 20020 13916 20030
rect 13860 19926 13916 19964
rect 14028 20020 14084 20030
rect 14140 20020 14196 23100
rect 14364 23380 14420 23390
rect 14364 22594 14420 23324
rect 14812 23156 14868 23166
rect 14924 23156 14980 25230
rect 15708 24500 15764 25452
rect 15820 24836 15876 26124
rect 15988 26114 16044 26124
rect 16156 25620 16212 25630
rect 16044 25508 16100 25518
rect 16044 25450 16100 25452
rect 15932 25396 15988 25406
rect 16044 25398 16046 25450
rect 16098 25398 16100 25450
rect 16156 25478 16212 25564
rect 16156 25426 16158 25478
rect 16210 25426 16212 25478
rect 16156 25414 16212 25426
rect 16044 25386 16100 25398
rect 15932 24836 15988 25340
rect 16100 24836 16156 24846
rect 15932 24834 16156 24836
rect 15932 24782 16102 24834
rect 16154 24782 16156 24834
rect 15932 24780 16156 24782
rect 15820 24770 15876 24780
rect 16100 24770 16156 24780
rect 16268 24724 16324 26908
rect 16436 26898 16492 26908
rect 17612 26852 17668 27134
rect 17612 26786 17668 26796
rect 18172 26852 18228 26862
rect 17844 26684 18108 26694
rect 17900 26628 17948 26684
rect 18004 26628 18052 26684
rect 17844 26618 18108 26628
rect 17276 26292 17332 26302
rect 17276 26198 17332 26236
rect 16436 26180 16492 26190
rect 18060 26180 18116 26190
rect 16436 26178 16548 26180
rect 16436 26126 16438 26178
rect 16490 26126 16548 26178
rect 16436 26114 16548 26126
rect 16380 25450 16436 25462
rect 16380 25398 16382 25450
rect 16434 25398 16436 25450
rect 16380 25284 16436 25398
rect 16380 25218 16436 25228
rect 16380 24724 16436 24734
rect 16268 24668 16380 24724
rect 16380 24630 16436 24668
rect 16492 24722 16548 26114
rect 17500 26178 18116 26180
rect 17500 26126 18062 26178
rect 18114 26126 18116 26178
rect 17500 26124 18116 26126
rect 17500 25730 17556 26124
rect 18060 26114 18116 26124
rect 17500 25678 17502 25730
rect 17554 25678 17556 25730
rect 17500 25666 17556 25678
rect 18172 25620 18228 26796
rect 19180 25674 19236 28364
rect 20188 27074 20244 27086
rect 20188 27022 20190 27074
rect 20242 27022 20244 27074
rect 19180 25622 19182 25674
rect 19234 25622 19236 25674
rect 19180 25610 19236 25622
rect 19852 26292 19908 26302
rect 16884 25508 16940 25518
rect 17164 25508 17220 25518
rect 16884 25506 17220 25508
rect 16604 25450 16660 25462
rect 16604 25398 16606 25450
rect 16658 25398 16660 25450
rect 16884 25454 16886 25506
rect 16938 25454 17166 25506
rect 17218 25454 17220 25506
rect 16884 25452 17220 25454
rect 16884 25442 16940 25452
rect 17164 25442 17220 25452
rect 16604 24836 16660 25398
rect 17844 25116 18108 25126
rect 17900 25060 17948 25116
rect 18004 25060 18052 25116
rect 17844 25050 18108 25060
rect 16604 24770 16660 24780
rect 17612 24948 17668 24958
rect 17276 24724 17332 24734
rect 16492 24670 16494 24722
rect 16546 24670 16548 24722
rect 15708 24444 16380 24500
rect 16324 24162 16380 24444
rect 16324 24110 16326 24162
rect 16378 24110 16380 24162
rect 16324 24098 16380 24110
rect 16492 24164 16548 24670
rect 17164 24668 17276 24724
rect 16492 24108 16772 24164
rect 16604 23938 16660 23950
rect 16604 23886 16606 23938
rect 16658 23886 16660 23938
rect 16604 23828 16660 23886
rect 16604 23762 16660 23772
rect 16716 23938 16772 24108
rect 16716 23886 16718 23938
rect 16770 23886 16772 23938
rect 16716 23380 16772 23886
rect 16940 23938 16996 23950
rect 16940 23886 16942 23938
rect 16994 23886 16996 23938
rect 16940 23828 16996 23886
rect 16940 23762 16996 23772
rect 14812 23154 14980 23156
rect 14812 23102 14814 23154
rect 14866 23102 14980 23154
rect 14812 23100 14980 23102
rect 16604 23324 16716 23380
rect 14812 23090 14868 23100
rect 14364 22542 14366 22594
rect 14418 22542 14420 22594
rect 14364 22530 14420 22542
rect 14700 22484 14756 22494
rect 14700 22370 14756 22428
rect 14700 22318 14702 22370
rect 14754 22318 14756 22370
rect 14420 20774 14476 20784
rect 14420 20772 14644 20774
rect 14420 20720 14422 20772
rect 14474 20720 14644 20772
rect 14420 20718 14644 20720
rect 14420 20708 14476 20718
rect 14364 20636 14420 20646
rect 14364 20634 14532 20636
rect 14364 20582 14366 20634
rect 14418 20582 14532 20634
rect 14364 20580 14532 20582
rect 14364 20570 14420 20580
rect 14084 19964 14196 20020
rect 14028 19926 14084 19964
rect 14364 19684 14420 19694
rect 13686 19628 13950 19638
rect 13742 19572 13790 19628
rect 13846 19572 13894 19628
rect 13686 19562 13950 19572
rect 13916 19460 13972 19470
rect 13468 19404 13860 19460
rect 13804 19348 13860 19404
rect 13524 19236 13580 19246
rect 13524 19142 13580 19180
rect 13804 19234 13860 19292
rect 13804 19182 13806 19234
rect 13858 19182 13860 19234
rect 13804 19170 13860 19182
rect 13916 19234 13972 19404
rect 13916 19182 13918 19234
rect 13970 19182 13972 19234
rect 13916 19170 13972 19182
rect 14364 19234 14420 19628
rect 14476 19302 14532 20580
rect 14588 19460 14644 20718
rect 14588 19394 14644 19404
rect 14476 19290 14588 19302
rect 14476 19238 14534 19290
rect 14586 19238 14588 19290
rect 14476 19236 14588 19238
rect 14364 19182 14366 19234
rect 14418 19182 14420 19234
rect 14532 19226 14588 19236
rect 14364 19170 14420 19182
rect 14700 19124 14756 22318
rect 15988 22146 16044 22158
rect 15988 22094 15990 22146
rect 16042 22094 16044 22146
rect 15988 21924 16044 22094
rect 15988 21858 16044 21868
rect 16604 21924 16660 23324
rect 16716 23286 16772 23324
rect 16604 21858 16660 21868
rect 16716 23042 16772 23054
rect 16716 22990 16718 23042
rect 16770 22990 16772 23042
rect 16716 21588 16772 22990
rect 17164 22370 17220 24668
rect 17276 24630 17332 24668
rect 17612 23940 17668 24892
rect 17612 23874 17668 23884
rect 18172 23940 18228 25564
rect 18732 25508 18788 25518
rect 18396 24836 18452 24846
rect 18396 24722 18452 24780
rect 18396 24670 18398 24722
rect 18450 24670 18452 24722
rect 18396 24658 18452 24670
rect 18564 24500 18620 24510
rect 18732 24500 18788 25452
rect 18956 25506 19012 25518
rect 18956 25454 18958 25506
rect 19010 25454 19012 25506
rect 18956 24948 19012 25454
rect 19292 25506 19348 25518
rect 19292 25454 19294 25506
rect 19346 25454 19348 25506
rect 19852 25468 19908 26236
rect 19292 25396 19348 25454
rect 19292 25330 19348 25340
rect 19740 25450 19796 25462
rect 19740 25398 19742 25450
rect 19794 25398 19796 25450
rect 19852 25416 19854 25468
rect 19906 25416 19908 25468
rect 19964 26178 20020 26190
rect 19964 26126 19966 26178
rect 20018 26126 20020 26178
rect 19964 25508 20020 26126
rect 19964 25442 20020 25452
rect 19852 25404 19908 25416
rect 18956 24882 19012 24892
rect 19068 24836 19124 24846
rect 19068 24742 19124 24780
rect 19740 24612 19796 25398
rect 20188 25396 20244 27022
rect 20412 27076 20468 27086
rect 20860 27076 20916 28590
rect 21196 27860 21252 27870
rect 21196 27858 21364 27860
rect 21196 27806 21198 27858
rect 21250 27806 21364 27858
rect 21196 27804 21364 27806
rect 21196 27794 21252 27804
rect 21196 27076 21252 27086
rect 20860 27074 21252 27076
rect 20860 27022 21198 27074
rect 21250 27022 21252 27074
rect 20860 27020 21252 27022
rect 20412 26982 20468 27020
rect 20692 26964 20748 26974
rect 20692 26962 20916 26964
rect 20692 26910 20694 26962
rect 20746 26910 20916 26962
rect 20692 26908 20916 26910
rect 20692 26898 20748 26908
rect 20860 26290 20916 26908
rect 20860 26238 20862 26290
rect 20914 26238 20916 26290
rect 20860 26226 20916 26238
rect 20972 26292 21028 26302
rect 20972 26198 21028 26236
rect 20412 25620 20468 25630
rect 20412 25618 21028 25620
rect 20412 25566 20414 25618
rect 20466 25566 21028 25618
rect 20412 25564 21028 25566
rect 20412 25554 20468 25564
rect 20188 25330 20244 25340
rect 20580 25450 20636 25462
rect 20580 25398 20582 25450
rect 20634 25398 20636 25450
rect 20580 24948 20636 25398
rect 20860 25396 20916 25406
rect 20580 24892 20804 24948
rect 19628 24556 19796 24612
rect 19852 24836 19908 24846
rect 19628 24500 19684 24556
rect 18732 24444 18844 24500
rect 18564 24406 18620 24444
rect 18788 23994 18844 24444
rect 18788 23942 18790 23994
rect 18842 23942 18844 23994
rect 18172 23938 18340 23940
rect 18172 23886 18174 23938
rect 18226 23886 18340 23938
rect 18788 23930 18844 23942
rect 19292 24164 19348 24174
rect 18172 23884 18340 23886
rect 18172 23874 18228 23884
rect 17836 23828 17892 23838
rect 17836 23734 17892 23772
rect 17276 23716 17332 23726
rect 17276 23622 17332 23660
rect 17844 23548 18108 23558
rect 17900 23492 17948 23548
rect 18004 23492 18052 23548
rect 17844 23482 18108 23492
rect 18172 23156 18228 23166
rect 17780 23098 17836 23110
rect 17780 23046 17782 23098
rect 17834 23046 17836 23098
rect 17780 22932 17836 23046
rect 17780 22866 17836 22876
rect 17948 23042 18004 23054
rect 17948 22990 17950 23042
rect 18002 22990 18004 23042
rect 17948 22708 18004 22990
rect 17164 22318 17166 22370
rect 17218 22318 17220 22370
rect 17164 22306 17220 22318
rect 17612 22652 18004 22708
rect 18060 22932 18116 22942
rect 17612 22331 17668 22652
rect 17836 22372 17892 22382
rect 17612 22279 17614 22331
rect 17666 22279 17668 22331
rect 17612 22267 17668 22279
rect 17724 22370 17892 22372
rect 17724 22318 17838 22370
rect 17890 22318 17892 22370
rect 17724 22316 17892 22318
rect 16716 21522 16772 21532
rect 17276 22202 17332 22214
rect 17276 22150 17278 22202
rect 17330 22150 17332 22202
rect 15036 20916 15092 20926
rect 14812 20914 15092 20916
rect 14812 20862 15038 20914
rect 15090 20862 15092 20914
rect 14812 20860 15092 20862
rect 14812 20018 14868 20860
rect 15036 20850 15092 20860
rect 15484 20802 15540 20814
rect 15148 20758 15204 20770
rect 15148 20706 15150 20758
rect 15202 20706 15204 20758
rect 15148 20188 15204 20706
rect 14812 19966 14814 20018
rect 14866 19966 14868 20018
rect 14812 19954 14868 19966
rect 15036 20132 15204 20188
rect 15484 20750 15486 20802
rect 15538 20750 15540 20802
rect 15484 20188 15540 20750
rect 16156 20804 16212 20814
rect 16156 20802 16660 20804
rect 16156 20750 16158 20802
rect 16210 20750 16660 20802
rect 16156 20748 16660 20750
rect 16156 20738 16212 20748
rect 15988 20580 16044 20590
rect 15988 20578 16548 20580
rect 15988 20526 15990 20578
rect 16042 20526 16548 20578
rect 15988 20524 16548 20526
rect 15988 20514 16044 20524
rect 16044 20356 16100 20366
rect 15484 20132 15988 20188
rect 13132 18834 13188 18844
rect 14476 19068 14756 19124
rect 14812 19684 14868 19694
rect 15036 19684 15092 20132
rect 15932 19684 15988 20132
rect 15036 19628 15204 19684
rect 12796 18620 13300 18676
rect 13244 18564 13300 18620
rect 14046 18564 14102 18574
rect 13244 18508 13524 18564
rect 12684 18386 12740 18396
rect 13132 18450 13188 18462
rect 13132 18398 13134 18450
rect 13186 18398 13188 18450
rect 12740 18226 12796 18238
rect 12740 18174 12742 18226
rect 12794 18174 12796 18226
rect 12740 18116 12796 18174
rect 12740 18050 12796 18060
rect 12628 17834 12684 17846
rect 12628 17782 12630 17834
rect 12682 17782 12684 17834
rect 12628 17668 12684 17782
rect 12628 17602 12684 17612
rect 12796 17780 12852 17790
rect 12796 17666 12852 17724
rect 12796 17614 12798 17666
rect 12850 17614 12852 17666
rect 12796 17602 12852 17614
rect 13132 17668 13188 18398
rect 13300 18394 13356 18406
rect 13300 18342 13302 18394
rect 13354 18342 13356 18394
rect 13300 18116 13356 18342
rect 13300 18050 13356 18060
rect 13468 17892 13524 18508
rect 14046 18470 14102 18508
rect 13804 18450 13860 18462
rect 13804 18398 13806 18450
rect 13858 18398 13860 18450
rect 13804 18228 13860 18398
rect 13804 18162 13860 18172
rect 14476 18450 14532 19068
rect 14476 18398 14478 18450
rect 14530 18398 14532 18450
rect 14812 18562 14868 19628
rect 15036 19236 15092 19246
rect 15036 19142 15092 19180
rect 14812 18510 14814 18562
rect 14866 18510 14868 18562
rect 14476 18116 14532 18398
rect 13686 18060 13950 18070
rect 13742 18004 13790 18060
rect 13846 18004 13894 18060
rect 14476 18050 14532 18060
rect 14644 18394 14700 18406
rect 14644 18342 14646 18394
rect 14698 18342 14700 18394
rect 13686 17994 13950 18004
rect 14252 18004 14308 18014
rect 13468 17836 13804 17892
rect 13748 17722 13804 17836
rect 13132 17602 13188 17612
rect 13580 17668 13636 17678
rect 13748 17670 13750 17722
rect 13802 17670 13804 17722
rect 13748 17658 13804 17670
rect 14252 17666 14308 17948
rect 14644 17780 14700 18342
rect 14812 18004 14868 18510
rect 15148 18462 15204 19628
rect 15278 19628 15988 19684
rect 15278 19458 15334 19628
rect 15278 19406 15280 19458
rect 15332 19406 15334 19458
rect 15278 19394 15334 19406
rect 16044 19124 16100 20300
rect 16156 20244 16212 20254
rect 16156 19234 16212 20188
rect 16156 19182 16158 19234
rect 16210 19182 16212 19234
rect 16324 19460 16380 19470
rect 16324 19290 16380 19404
rect 16324 19238 16326 19290
rect 16378 19238 16380 19290
rect 16324 19226 16380 19238
rect 16492 19236 16548 20524
rect 16604 20188 16660 20748
rect 17276 20188 17332 22150
rect 17724 21812 17780 22316
rect 17836 22306 17892 22316
rect 18060 22148 18116 22876
rect 18172 22372 18228 23100
rect 18172 22306 18228 22316
rect 18060 22092 18228 22148
rect 17844 21980 18108 21990
rect 17900 21924 17948 21980
rect 18004 21924 18052 21980
rect 17844 21914 18108 21924
rect 17724 21746 17780 21756
rect 18060 21812 18116 21822
rect 18172 21812 18228 22092
rect 18060 21810 18228 21812
rect 18060 21758 18062 21810
rect 18114 21758 18228 21810
rect 18060 21756 18228 21758
rect 18060 21746 18116 21756
rect 16604 20132 16772 20188
rect 16716 19906 16772 20132
rect 16716 19854 16718 19906
rect 16770 19854 16772 19906
rect 16156 19170 16212 19182
rect 16492 19142 16548 19180
rect 16604 19348 16660 19358
rect 16604 19234 16660 19292
rect 16604 19182 16606 19234
rect 16658 19182 16660 19234
rect 16604 19170 16660 19182
rect 15764 19068 16100 19124
rect 15596 18564 15652 18574
rect 14924 18450 14980 18462
rect 14924 18398 14926 18450
rect 14978 18398 14980 18450
rect 14924 18340 14980 18398
rect 15148 18450 15260 18462
rect 15148 18398 15206 18450
rect 15258 18398 15260 18450
rect 15148 18396 15260 18398
rect 15204 18386 15260 18396
rect 15596 18450 15652 18508
rect 15596 18398 15598 18450
rect 15650 18398 15652 18450
rect 15596 18386 15652 18398
rect 15764 18394 15820 19068
rect 16716 19012 16772 19854
rect 17164 20132 17332 20188
rect 17724 21588 17780 21598
rect 17724 20244 17780 21532
rect 18172 21364 18228 21374
rect 17844 20412 18108 20422
rect 17900 20356 17948 20412
rect 18004 20356 18052 20412
rect 17844 20346 18108 20356
rect 17724 20178 17780 20188
rect 16884 19236 16940 19246
rect 16884 19142 16940 19180
rect 15932 18956 16772 19012
rect 15932 18562 15988 18956
rect 15932 18510 15934 18562
rect 15986 18510 15988 18562
rect 15932 18498 15988 18510
rect 16604 18788 16660 18798
rect 14924 18274 14980 18284
rect 15764 18342 15766 18394
rect 15818 18342 15820 18394
rect 16044 18452 16100 18462
rect 16044 18450 16212 18452
rect 16044 18398 16046 18450
rect 16098 18398 16212 18450
rect 16044 18396 16212 18398
rect 16044 18386 16100 18396
rect 15260 18228 15316 18238
rect 14812 17948 14980 18004
rect 14924 17892 14980 17948
rect 14924 17826 14980 17836
rect 13580 17574 13636 17612
rect 14252 17614 14254 17666
rect 14306 17614 14308 17666
rect 12460 17388 12740 17444
rect 12684 16994 12740 17388
rect 12684 16942 12686 16994
rect 12738 16942 12740 16994
rect 12684 16930 12740 16942
rect 12927 16884 12983 16894
rect 12927 16790 12983 16828
rect 13804 16884 13860 16894
rect 13804 16882 14084 16884
rect 13804 16830 13806 16882
rect 13858 16830 14084 16882
rect 13804 16828 14084 16830
rect 13804 16818 13860 16828
rect 14028 16772 14084 16828
rect 13686 16492 13950 16502
rect 13742 16436 13790 16492
rect 13846 16436 13894 16492
rect 13686 16426 13950 16436
rect 12516 15876 12572 15886
rect 12516 15782 12572 15820
rect 12516 15540 12572 15550
rect 12012 15538 12572 15540
rect 12012 15486 12518 15538
rect 12570 15486 12572 15538
rect 12012 15484 12572 15486
rect 12012 15341 12068 15484
rect 12012 15289 12014 15341
rect 12066 15289 12068 15341
rect 12012 15277 12068 15289
rect 12460 15474 12572 15484
rect 11172 15250 11228 15260
rect 11452 14530 11508 14542
rect 11452 14478 11454 14530
rect 11506 14478 11508 14530
rect 9548 14420 9604 14430
rect 9548 14418 9940 14420
rect 9548 14366 9550 14418
rect 9602 14366 9940 14418
rect 9548 14364 9940 14366
rect 9548 14354 9604 14364
rect 9528 14140 9792 14150
rect 9584 14084 9632 14140
rect 9688 14084 9736 14140
rect 9528 14074 9792 14084
rect 8988 13972 9100 13982
rect 9716 13972 9772 13982
rect 8988 13970 9772 13972
rect 8988 13918 9046 13970
rect 9098 13918 9718 13970
rect 9770 13918 9772 13970
rect 8988 13916 9772 13918
rect 9044 13906 9100 13916
rect 9716 13906 9772 13916
rect 9884 13300 9940 14364
rect 9884 13234 9940 13244
rect 11340 13300 11396 13310
rect 10332 13132 11060 13188
rect 9324 13076 9380 13086
rect 8428 12348 8708 12404
rect 8876 12516 8932 12526
rect 7756 12292 7812 12302
rect 7756 11508 7812 12236
rect 7980 12214 8036 12226
rect 7980 12180 7982 12214
rect 8034 12180 8036 12214
rect 7980 12114 8036 12124
rect 8316 12211 8372 12223
rect 8316 12159 8318 12211
rect 8370 12159 8372 12211
rect 8316 12068 8372 12159
rect 8428 12068 8484 12348
rect 8764 12292 8820 12302
rect 8626 12213 8682 12223
rect 8626 12211 8708 12213
rect 8626 12159 8628 12211
rect 8680 12159 8708 12211
rect 8764 12198 8820 12236
rect 8626 12147 8708 12159
rect 8428 12012 8596 12068
rect 8316 12002 8372 12012
rect 7756 11442 7812 11452
rect 7812 11284 7868 11294
rect 7812 11282 8372 11284
rect 7812 11230 7814 11282
rect 7866 11230 8372 11282
rect 7812 11228 8372 11230
rect 7812 11218 7868 11228
rect 7588 10722 7700 10734
rect 7588 10670 7590 10722
rect 7642 10670 7700 10722
rect 7588 10668 7700 10670
rect 7756 10780 8204 10836
rect 7588 10658 7644 10668
rect 7588 9716 7644 9726
rect 7588 9622 7644 9660
rect 7644 9492 7700 9502
rect 7532 9380 7588 9390
rect 7532 8820 7588 9324
rect 7644 9042 7700 9436
rect 7756 9380 7812 10780
rect 8148 10666 8204 10780
rect 7868 10610 7924 10622
rect 7868 10558 7870 10610
rect 7922 10558 7924 10610
rect 7868 10164 7924 10558
rect 7980 10610 8036 10622
rect 7980 10558 7982 10610
rect 8034 10558 8036 10610
rect 8148 10614 8150 10666
rect 8202 10614 8204 10666
rect 8148 10602 8204 10614
rect 8316 10610 8372 11228
rect 7980 10276 8036 10558
rect 8316 10558 8318 10610
rect 8370 10558 8372 10610
rect 8316 10546 8372 10558
rect 7980 10220 8260 10276
rect 7868 10108 8092 10164
rect 8036 10050 8092 10108
rect 8036 9998 8038 10050
rect 8090 9998 8092 10050
rect 8036 9986 8092 9998
rect 7756 9324 8092 9380
rect 7644 8990 7646 9042
rect 7698 8990 7700 9042
rect 7644 8978 7700 8990
rect 8036 9098 8092 9324
rect 8036 9046 8038 9098
rect 8090 9046 8092 9098
rect 7868 8932 7924 8942
rect 7756 8930 7924 8932
rect 7756 8878 7870 8930
rect 7922 8878 7924 8930
rect 7756 8876 7924 8878
rect 7532 8764 7700 8820
rect 7308 8372 7476 8428
rect 7532 8484 7588 8494
rect 7308 7598 7364 8372
rect 7420 8258 7476 8270
rect 7420 8206 7422 8258
rect 7474 8206 7476 8258
rect 7420 8148 7476 8206
rect 7420 8082 7476 8092
rect 7308 7586 7420 7598
rect 7308 7534 7366 7586
rect 7418 7534 7420 7586
rect 7308 7532 7420 7534
rect 7364 7522 7420 7532
rect 6860 5506 6916 5516
rect 6972 6748 7252 6804
rect 7532 6804 7588 8428
rect 7644 7476 7700 8764
rect 7756 8260 7812 8876
rect 7868 8866 7924 8876
rect 8036 8428 8092 9046
rect 8204 8820 8260 10220
rect 8316 9826 8372 9838
rect 8316 9774 8318 9826
rect 8370 9774 8372 9826
rect 8316 9044 8372 9774
rect 8428 9828 8484 9838
rect 8428 9734 8484 9772
rect 8316 8978 8372 8988
rect 8428 9042 8484 9054
rect 8428 8990 8430 9042
rect 8482 8990 8484 9042
rect 8316 8874 8372 8886
rect 8316 8822 8318 8874
rect 8370 8822 8372 8874
rect 8316 8820 8372 8822
rect 8204 8764 8372 8820
rect 8428 8484 8484 8990
rect 7756 8194 7812 8204
rect 7868 8372 8092 8428
rect 8316 8428 8484 8484
rect 7868 8258 7924 8372
rect 8204 8260 8260 8270
rect 7868 8206 7870 8258
rect 7922 8206 7924 8258
rect 7868 7924 7924 8206
rect 7644 7382 7700 7420
rect 7756 7868 7868 7924
rect 7756 7252 7812 7868
rect 7868 7858 7924 7868
rect 7980 8258 8260 8260
rect 7980 8206 8206 8258
rect 8258 8206 8260 8258
rect 7980 8204 8260 8206
rect 7756 7186 7812 7196
rect 7868 7474 7924 7486
rect 7868 7422 7870 7474
rect 7922 7422 7924 7474
rect 7868 7140 7924 7422
rect 7868 7074 7924 7084
rect 7532 6748 7700 6804
rect 6412 5234 6580 5236
rect 6412 5182 6414 5234
rect 6466 5182 6580 5234
rect 6412 5180 6580 5182
rect 6636 5404 6748 5460
rect 6412 5124 6468 5180
rect 6412 5058 6468 5068
rect 6636 4900 6692 5404
rect 6748 5394 6804 5404
rect 6972 5348 7028 6748
rect 7644 6692 7700 6748
rect 7868 6692 7924 6702
rect 7644 6690 7924 6692
rect 7532 6634 7588 6646
rect 7644 6638 7870 6690
rect 7922 6638 7924 6690
rect 7644 6636 7924 6638
rect 7084 6580 7140 6590
rect 7084 6018 7140 6524
rect 7532 6582 7534 6634
rect 7586 6582 7588 6634
rect 7084 5966 7086 6018
rect 7138 5966 7140 6018
rect 7084 5954 7140 5966
rect 7252 6020 7308 6030
rect 7252 5962 7308 5964
rect 7252 5910 7254 5962
rect 7306 5910 7308 5962
rect 7252 5898 7308 5910
rect 7532 5460 7588 6582
rect 7868 6244 7924 6636
rect 7868 6178 7924 6188
rect 7980 6030 8036 8204
rect 8204 8194 8260 8204
rect 8316 7476 8372 8428
rect 8428 8260 8484 8270
rect 8540 8260 8596 12012
rect 8652 11732 8708 12147
rect 8876 11844 8932 12460
rect 8876 11778 8932 11788
rect 8652 11666 8708 11676
rect 9212 11732 9268 11742
rect 9100 11394 9156 11406
rect 9100 11342 9102 11394
rect 9154 11342 9156 11394
rect 9100 9828 9156 11342
rect 9212 11226 9268 11676
rect 9324 11355 9380 13020
rect 9772 13076 9828 13086
rect 10164 13076 10220 13086
rect 9772 13074 9940 13076
rect 9772 13022 9774 13074
rect 9826 13022 9940 13074
rect 9772 13020 9940 13022
rect 9772 13010 9828 13020
rect 9528 12572 9792 12582
rect 9584 12516 9632 12572
rect 9688 12516 9736 12572
rect 9528 12506 9792 12516
rect 9884 11956 9940 13020
rect 10164 12962 10220 13020
rect 10164 12910 10166 12962
rect 10218 12910 10220 12962
rect 10164 12898 10220 12910
rect 10332 12962 10388 13132
rect 10332 12910 10334 12962
rect 10386 12910 10388 12962
rect 10332 12898 10388 12910
rect 10444 12962 10500 12974
rect 10444 12910 10446 12962
rect 10498 12910 10500 12962
rect 9884 11890 9940 11900
rect 10332 12206 10388 12218
rect 10332 12154 10334 12206
rect 10386 12154 10388 12206
rect 10332 11620 10388 12154
rect 10332 11554 10388 11564
rect 9324 11303 9326 11355
rect 9378 11303 9380 11355
rect 9324 11291 9380 11303
rect 9660 11396 9716 11406
rect 10444 11396 10500 12910
rect 10556 12852 10612 12862
rect 10556 12292 10612 12796
rect 10556 12178 10612 12236
rect 10556 12126 10558 12178
rect 10610 12126 10612 12178
rect 10556 12114 10612 12126
rect 9660 11302 9716 11340
rect 10108 11340 10500 11396
rect 9212 11174 9214 11226
rect 9266 11174 9268 11226
rect 9212 10276 9268 11174
rect 9528 11004 9792 11014
rect 9584 10948 9632 11004
rect 9688 10948 9736 11004
rect 9528 10938 9792 10948
rect 10108 10610 10164 11340
rect 10220 11172 10276 11182
rect 10220 10836 10276 11116
rect 10220 10770 10276 10780
rect 10108 10558 10110 10610
rect 10162 10558 10164 10610
rect 10108 10546 10164 10558
rect 10444 10612 10500 11340
rect 10556 11396 10612 11406
rect 10668 11396 10724 13132
rect 11004 13130 11060 13132
rect 11004 13078 11006 13130
rect 11058 13078 11060 13130
rect 11004 13066 11060 13078
rect 11340 13076 11396 13244
rect 10780 12964 10836 12974
rect 10780 12290 10836 12908
rect 10780 12238 10782 12290
rect 10834 12238 10836 12290
rect 10780 12226 10836 12238
rect 11116 12962 11172 12974
rect 11116 12910 11118 12962
rect 11170 12910 11172 12962
rect 10948 12180 11004 12190
rect 10948 12086 11004 12124
rect 11116 11620 11172 12910
rect 11340 12962 11396 13020
rect 11340 12910 11342 12962
rect 11394 12910 11396 12962
rect 11340 12898 11396 12910
rect 11116 11554 11172 11564
rect 11228 12180 11284 12190
rect 10556 11394 10724 11396
rect 10556 11342 10558 11394
rect 10610 11342 10724 11394
rect 10556 11340 10724 11342
rect 11228 11394 11284 12124
rect 11340 12068 11396 12078
rect 11340 11974 11396 12012
rect 11452 11844 11508 14478
rect 12236 14530 12292 14542
rect 12236 14478 12238 14530
rect 12290 14478 12292 14530
rect 11788 13746 11844 13758
rect 11788 13694 11790 13746
rect 11842 13694 11844 13746
rect 11788 12964 11844 13694
rect 12012 12964 12068 12974
rect 11788 12908 12012 12964
rect 12012 12870 12068 12908
rect 12236 12964 12292 14478
rect 12236 12898 12292 12908
rect 12012 12404 12068 12414
rect 11754 12215 11810 12227
rect 11754 12163 11756 12215
rect 11808 12163 11810 12215
rect 11228 11342 11230 11394
rect 11282 11342 11284 11394
rect 10556 11330 10612 11340
rect 11228 11330 11284 11342
rect 11340 11788 11508 11844
rect 11564 11844 11620 11854
rect 10948 11284 11004 11294
rect 10948 11282 11060 11284
rect 10948 11230 10950 11282
rect 11002 11230 11060 11282
rect 10948 11218 11060 11230
rect 10444 10556 10612 10612
rect 9772 10388 9828 10398
rect 9772 10294 9828 10332
rect 10444 10388 10500 10398
rect 9212 10210 9268 10220
rect 9100 9762 9156 9772
rect 8652 9716 8708 9726
rect 8652 9042 8708 9660
rect 9528 9436 9792 9446
rect 9584 9380 9632 9436
rect 9688 9380 9736 9436
rect 9528 9370 9792 9380
rect 10220 9380 10276 9390
rect 10220 9156 10276 9324
rect 8652 8990 8654 9042
rect 8706 8990 8708 9042
rect 8652 8978 8708 8990
rect 9548 9044 9604 9054
rect 9548 8370 9604 8988
rect 9548 8318 9550 8370
rect 9602 8318 9604 8370
rect 9548 8306 9604 8318
rect 8428 8258 8596 8260
rect 8428 8206 8430 8258
rect 8482 8206 8596 8258
rect 8428 8204 8596 8206
rect 8652 8260 8708 8270
rect 8428 8194 8484 8204
rect 8652 8166 8708 8204
rect 9100 8258 9156 8270
rect 9436 8260 9492 8270
rect 9100 8206 9102 8258
rect 9154 8206 9156 8258
rect 8092 7420 8372 7476
rect 8540 8036 8596 8046
rect 8092 6690 8148 7420
rect 8540 6916 8596 7980
rect 9100 7364 9156 8206
rect 9100 7298 9156 7308
rect 9324 8258 9492 8260
rect 9324 8206 9438 8258
rect 9490 8206 9492 8258
rect 10108 8260 10164 8270
rect 9324 8204 9492 8206
rect 8988 7140 9044 7150
rect 8652 6916 8708 6926
rect 8092 6638 8094 6690
rect 8146 6638 8148 6690
rect 8092 6626 8148 6638
rect 8260 6914 8708 6916
rect 8260 6862 8654 6914
rect 8706 6862 8708 6914
rect 8260 6860 8708 6862
rect 8260 6634 8316 6860
rect 8652 6850 8708 6860
rect 8260 6582 8262 6634
rect 8314 6582 8316 6634
rect 8988 6690 9044 7084
rect 8988 6638 8990 6690
rect 9042 6638 9044 6690
rect 8988 6626 9044 6638
rect 8260 6580 8316 6582
rect 8260 6514 8316 6524
rect 8204 6356 8260 6366
rect 7980 6018 8054 6030
rect 7980 5966 8000 6018
rect 8052 5966 8054 6018
rect 7980 5964 8054 5966
rect 7998 5954 8054 5964
rect 6972 5282 7028 5292
rect 7308 5404 7588 5460
rect 7756 5906 7812 5918
rect 7756 5854 7758 5906
rect 7810 5854 7812 5906
rect 6806 5236 6862 5246
rect 6806 5122 6862 5180
rect 6806 5070 6808 5122
rect 6860 5070 6862 5122
rect 6806 5058 6862 5070
rect 6972 5122 7028 5134
rect 6972 5070 6974 5122
rect 7026 5070 7028 5122
rect 6972 4900 7028 5070
rect 7084 5124 7140 5134
rect 7084 5030 7140 5068
rect 6636 4844 7252 4900
rect 4620 4284 4788 4286
rect 4732 4274 4788 4284
rect 5370 3948 5634 3958
rect 5426 3892 5474 3948
rect 5530 3892 5578 3948
rect 5370 3882 5634 3892
rect 4396 3670 4398 3722
rect 4450 3670 4452 3722
rect 5740 3678 5796 4284
rect 7196 4228 7252 4844
rect 7308 4450 7364 5404
rect 7532 5236 7588 5246
rect 7756 5236 7812 5854
rect 8092 5796 8148 5806
rect 7532 5234 7812 5236
rect 7532 5182 7534 5234
rect 7586 5182 7812 5234
rect 7532 5180 7812 5182
rect 7980 5740 8092 5796
rect 7532 5170 7588 5180
rect 7980 5134 8036 5740
rect 8092 5730 8148 5740
rect 7924 5122 8036 5134
rect 7924 5070 7926 5122
rect 7978 5070 8036 5122
rect 7924 5068 8036 5070
rect 8092 5572 8148 5582
rect 8092 5122 8148 5516
rect 8092 5070 8094 5122
rect 8146 5070 8148 5122
rect 7924 5058 7980 5068
rect 8092 5058 8148 5070
rect 8204 5122 8260 6300
rect 8204 5070 8206 5122
rect 8258 5070 8260 5122
rect 8204 5012 8260 5070
rect 8204 4946 8260 4956
rect 8316 6244 8372 6254
rect 7308 4398 7310 4450
rect 7362 4398 7364 4450
rect 7308 4386 7364 4398
rect 8316 4452 8372 6188
rect 9324 6132 9380 8204
rect 9436 8194 9492 8204
rect 9772 8202 9828 8214
rect 9772 8150 9774 8202
rect 9826 8150 9828 8202
rect 10108 8166 10164 8204
rect 9772 8148 9828 8150
rect 9772 8082 9828 8092
rect 9528 7868 9792 7878
rect 9584 7812 9632 7868
rect 9688 7812 9736 7868
rect 9528 7802 9792 7812
rect 9996 7364 10052 7374
rect 9996 7270 10052 7308
rect 9528 6300 9792 6310
rect 9584 6244 9632 6300
rect 9688 6244 9736 6300
rect 9528 6234 9792 6244
rect 9324 6066 9380 6076
rect 9996 6132 10052 6142
rect 8316 4386 8372 4396
rect 8428 5348 8484 5358
rect 8428 5124 8484 5292
rect 7551 4338 7607 4350
rect 7551 4286 7553 4338
rect 7605 4286 7607 4338
rect 7551 4228 7607 4286
rect 8428 4338 8484 5068
rect 9996 5236 10052 6076
rect 10108 5908 10164 5918
rect 10108 5290 10164 5852
rect 10220 5684 10276 9100
rect 10444 8428 10500 10332
rect 10556 9994 10612 10556
rect 10556 9942 10558 9994
rect 10610 9942 10612 9994
rect 10556 9930 10612 9942
rect 10668 9828 10724 9838
rect 10668 9826 10836 9828
rect 10668 9774 10670 9826
rect 10722 9774 10836 9826
rect 10668 9772 10836 9774
rect 10668 9762 10724 9772
rect 10444 8372 10724 8428
rect 10390 7474 10446 7486
rect 10390 7422 10392 7474
rect 10444 7422 10446 7474
rect 10390 6916 10446 7422
rect 10390 6850 10446 6860
rect 10556 7476 10612 7486
rect 10556 6804 10612 7420
rect 10668 7474 10724 8372
rect 10668 7422 10670 7474
rect 10722 7422 10724 7474
rect 10668 7410 10724 7422
rect 10556 6738 10612 6748
rect 10780 6580 10836 9772
rect 10780 6514 10836 6524
rect 10892 9826 10948 9838
rect 10892 9774 10894 9826
rect 10946 9774 10948 9826
rect 10892 9716 10948 9774
rect 10220 5618 10276 5628
rect 10444 6244 10500 6254
rect 10892 6244 10948 9660
rect 11004 7476 11060 11218
rect 11116 11172 11172 11182
rect 11116 9042 11172 11116
rect 11340 10052 11396 11788
rect 11452 11620 11508 11630
rect 11452 11394 11508 11564
rect 11452 11342 11454 11394
rect 11506 11342 11508 11394
rect 11452 11330 11508 11342
rect 11228 9996 11396 10052
rect 11228 9492 11284 9996
rect 11396 9828 11452 9838
rect 11396 9734 11452 9772
rect 11228 9268 11284 9436
rect 11228 9202 11284 9212
rect 11116 8990 11118 9042
rect 11170 8990 11172 9042
rect 11116 8978 11172 8990
rect 11284 8818 11340 8830
rect 11284 8766 11286 8818
rect 11338 8766 11340 8818
rect 11284 8428 11340 8766
rect 11284 8372 11508 8428
rect 11340 8260 11396 8270
rect 11116 8202 11172 8214
rect 11116 8150 11118 8202
rect 11170 8150 11172 8202
rect 11116 8036 11172 8150
rect 11116 7970 11172 7980
rect 11004 7410 11060 7420
rect 11172 6916 11228 6926
rect 11172 6822 11228 6860
rect 11340 6692 11396 8204
rect 11452 7474 11508 8372
rect 11564 8258 11620 11788
rect 11754 11732 11810 12163
rect 11900 12180 11956 12190
rect 11754 11676 11844 11732
rect 11788 10052 11844 11676
rect 11900 11618 11956 12124
rect 12012 12178 12068 12348
rect 12012 12126 12014 12178
rect 12066 12126 12068 12178
rect 12460 12404 12516 15474
rect 14028 15428 14084 16716
rect 14252 16210 14308 17614
rect 14364 17724 14700 17780
rect 14812 17780 14868 17790
rect 14364 16772 14420 17724
rect 14494 17556 14550 17566
rect 14364 16706 14420 16716
rect 14476 17554 14550 17556
rect 14476 17502 14496 17554
rect 14548 17502 14550 17554
rect 14476 17490 14550 17502
rect 14252 16158 14254 16210
rect 14306 16158 14308 16210
rect 14252 16146 14308 16158
rect 14028 15362 14084 15372
rect 14476 15314 14532 17490
rect 14812 17332 14868 17724
rect 15260 17666 15316 18172
rect 15764 18004 15820 18342
rect 15764 17938 15820 17948
rect 15932 17892 15988 17902
rect 15260 17614 15262 17666
rect 15314 17614 15316 17666
rect 15260 17602 15316 17614
rect 15484 17780 15540 17790
rect 15484 17666 15540 17724
rect 15820 17780 15876 17790
rect 15932 17780 15988 17836
rect 15820 17778 15988 17780
rect 15820 17726 15822 17778
rect 15874 17726 15988 17778
rect 15820 17724 15988 17726
rect 15820 17714 15876 17724
rect 15484 17614 15486 17666
rect 15538 17614 15540 17666
rect 15484 17602 15540 17614
rect 16156 17668 16212 18396
rect 16324 18228 16380 18238
rect 16324 18134 16380 18172
rect 16156 17574 16212 17612
rect 14980 17556 15036 17566
rect 14980 17462 15036 17500
rect 14588 17276 14868 17332
rect 14588 16882 14644 17276
rect 14588 16830 14590 16882
rect 14642 16830 14644 16882
rect 14588 16818 14644 16830
rect 14700 16884 14756 16894
rect 14700 15764 14756 16828
rect 14812 16882 14868 16894
rect 14812 16830 14814 16882
rect 14866 16830 14868 16882
rect 14812 15876 14868 16830
rect 15092 16884 15148 16894
rect 15372 16884 15428 16894
rect 15092 16882 15428 16884
rect 15092 16830 15094 16882
rect 15146 16830 15374 16882
rect 15426 16830 15428 16882
rect 15092 16828 15428 16830
rect 15092 16818 15148 16828
rect 15372 16818 15428 16828
rect 15708 16660 15764 16670
rect 15708 16658 16212 16660
rect 15708 16606 15710 16658
rect 15762 16606 16212 16658
rect 15708 16604 16212 16606
rect 15708 16594 15764 16604
rect 16156 16210 16212 16604
rect 16156 16158 16158 16210
rect 16210 16158 16212 16210
rect 16156 16146 16212 16158
rect 14812 15820 15260 15876
rect 14700 15708 14868 15764
rect 14476 15262 14478 15314
rect 14530 15262 14532 15314
rect 14644 15428 14700 15438
rect 14644 15370 14700 15372
rect 14644 15318 14646 15370
rect 14698 15318 14700 15370
rect 14812 15426 14868 15708
rect 14812 15374 14814 15426
rect 14866 15374 14868 15426
rect 14812 15362 14868 15374
rect 15204 15426 15260 15820
rect 15204 15374 15206 15426
rect 15258 15374 15260 15426
rect 15204 15362 15260 15374
rect 15932 15540 15988 15550
rect 14644 15306 14700 15318
rect 14924 15314 14980 15326
rect 14476 15250 14532 15262
rect 14924 15262 14926 15314
rect 14978 15262 14980 15314
rect 14924 15204 14980 15262
rect 14924 15138 14980 15148
rect 13686 14924 13950 14934
rect 13742 14868 13790 14924
rect 13846 14868 13894 14924
rect 13686 14858 13950 14868
rect 14644 14306 14700 14318
rect 14644 14254 14646 14306
rect 14698 14254 14700 14306
rect 14644 13748 14700 14254
rect 15148 13972 15204 13982
rect 15148 13878 15204 13916
rect 14812 13748 14868 13758
rect 14644 13746 14868 13748
rect 14644 13694 14814 13746
rect 14866 13694 14868 13746
rect 14644 13692 14868 13694
rect 12572 13634 12628 13646
rect 12572 13582 12574 13634
rect 12626 13582 12628 13634
rect 12572 12516 12628 13582
rect 14476 13636 14532 13646
rect 14476 13542 14532 13580
rect 13686 13356 13950 13366
rect 13742 13300 13790 13356
rect 13846 13300 13894 13356
rect 13686 13290 13950 13300
rect 14028 13188 14084 13198
rect 12572 12450 12628 12460
rect 13356 12962 13412 12974
rect 13356 12910 13358 12962
rect 13410 12910 13412 12962
rect 12460 12205 12516 12348
rect 12460 12153 12462 12205
rect 12514 12153 12516 12205
rect 12460 12141 12516 12153
rect 12012 12114 12068 12126
rect 11900 11566 11902 11618
rect 11954 11566 11956 11618
rect 11900 10612 11956 11566
rect 12572 11620 12628 11630
rect 12572 11526 12628 11564
rect 13356 11620 13412 12910
rect 13692 12738 13748 12750
rect 13692 12686 13694 12738
rect 13746 12686 13748 12738
rect 13692 12516 13748 12686
rect 13692 12450 13748 12460
rect 14028 11844 14084 13132
rect 14364 13076 14420 13086
rect 14364 12962 14420 13020
rect 14364 12910 14366 12962
rect 14418 12910 14420 12962
rect 14364 12898 14420 12910
rect 14588 12964 14644 12974
rect 14812 12964 14868 13692
rect 15820 13074 15876 13086
rect 15820 13022 15822 13074
rect 15874 13022 15876 13074
rect 15036 12964 15092 12974
rect 14812 12962 15092 12964
rect 14812 12910 15038 12962
rect 15090 12910 15092 12962
rect 14812 12908 15092 12910
rect 14196 12738 14252 12750
rect 14196 12686 14198 12738
rect 14250 12686 14252 12738
rect 14196 12180 14252 12686
rect 14196 12114 14252 12124
rect 14588 12178 14644 12908
rect 14868 12740 14924 12908
rect 15036 12898 15092 12908
rect 15596 12964 15652 12974
rect 15596 12870 15652 12908
rect 14588 12126 14590 12178
rect 14642 12126 14644 12178
rect 13686 11788 13950 11798
rect 13742 11732 13790 11788
rect 13846 11732 13894 11788
rect 14028 11778 14084 11788
rect 13686 11722 13950 11732
rect 14588 11732 14644 12126
rect 14588 11666 14644 11676
rect 14700 12738 14924 12740
rect 14700 12686 14870 12738
rect 14922 12686 14924 12738
rect 15204 12852 15260 12862
rect 15204 12794 15260 12796
rect 15204 12742 15206 12794
rect 15258 12742 15260 12794
rect 15204 12730 15260 12742
rect 14700 12684 14924 12686
rect 13356 11554 13412 11564
rect 14700 11508 14756 12684
rect 14868 12674 14924 12684
rect 15316 12404 15372 12414
rect 15316 12310 15372 12348
rect 14980 11844 15036 11854
rect 14588 11452 14756 11508
rect 14812 11620 14868 11630
rect 12236 11394 12292 11406
rect 12236 11342 12238 11394
rect 12290 11342 12292 11394
rect 12236 10724 12292 11342
rect 12908 11394 12964 11406
rect 12908 11342 12910 11394
rect 12962 11342 12964 11394
rect 12908 11172 12964 11342
rect 13692 11396 13748 11406
rect 13692 11394 13972 11396
rect 13692 11342 13694 11394
rect 13746 11342 13972 11394
rect 13692 11340 13972 11342
rect 13692 11330 13748 11340
rect 12236 10658 12292 10668
rect 12460 10724 12516 10734
rect 12012 10612 12068 10622
rect 11900 10610 12068 10612
rect 11900 10558 12014 10610
rect 12066 10558 12068 10610
rect 11900 10556 12068 10558
rect 12012 10546 12068 10556
rect 12180 10500 12236 10510
rect 12180 10442 12236 10444
rect 12180 10390 12182 10442
rect 12234 10390 12236 10442
rect 12180 10378 12236 10390
rect 11788 9986 11844 9996
rect 12012 10276 12068 10286
rect 11676 9826 11732 9838
rect 11676 9774 11678 9826
rect 11730 9774 11732 9826
rect 11676 9268 11732 9774
rect 11676 9202 11732 9212
rect 11788 9826 11844 9838
rect 11788 9774 11790 9826
rect 11842 9774 11844 9826
rect 11788 9716 11844 9774
rect 11788 8932 11844 9660
rect 11788 8866 11844 8876
rect 11900 9156 11956 9166
rect 11564 8206 11566 8258
rect 11618 8206 11620 8258
rect 11564 8194 11620 8206
rect 11788 8708 11844 8718
rect 11788 8148 11844 8652
rect 11788 8082 11844 8092
rect 11564 8036 11620 8046
rect 11564 7642 11620 7980
rect 11564 7590 11566 7642
rect 11618 7590 11620 7642
rect 11564 7578 11620 7590
rect 11452 7422 11454 7474
rect 11506 7422 11508 7474
rect 11452 7410 11508 7422
rect 11676 7513 11732 7525
rect 11676 7461 11678 7513
rect 11730 7461 11732 7513
rect 11676 6916 11732 7461
rect 11900 7252 11956 9100
rect 12012 8484 12068 10220
rect 12348 10052 12404 10062
rect 12180 9714 12236 9726
rect 12180 9662 12182 9714
rect 12234 9662 12236 9714
rect 12180 9156 12236 9662
rect 12180 9090 12236 9100
rect 12348 9044 12404 9996
rect 12012 8418 12068 8428
rect 12180 8818 12236 8830
rect 12180 8766 12182 8818
rect 12234 8766 12236 8818
rect 12180 8428 12236 8766
rect 12348 8708 12404 8988
rect 12460 9826 12516 10668
rect 12796 10724 12852 10734
rect 12796 10654 12852 10668
rect 12796 10602 12798 10654
rect 12850 10602 12852 10654
rect 12796 10590 12852 10602
rect 12684 10500 12740 10510
rect 12460 9774 12462 9826
rect 12514 9774 12516 9826
rect 12460 9042 12516 9774
rect 12572 10498 12740 10500
rect 12572 10446 12686 10498
rect 12738 10446 12740 10498
rect 12572 10444 12740 10446
rect 12572 9380 12628 10444
rect 12684 10434 12740 10444
rect 12684 9828 12740 9838
rect 12908 9828 12964 11116
rect 13524 11172 13580 11182
rect 13524 11078 13580 11116
rect 13132 10612 13188 10622
rect 13132 10518 13188 10556
rect 13916 10612 13972 11340
rect 14476 11394 14532 11406
rect 14476 11342 14478 11394
rect 14530 11342 14532 11394
rect 14476 11284 14532 11342
rect 14476 11218 14532 11228
rect 14140 11170 14196 11182
rect 14140 11118 14142 11170
rect 14194 11118 14196 11170
rect 14140 10724 14196 11118
rect 14140 10658 14196 10668
rect 13916 10518 13972 10556
rect 12684 9826 12964 9828
rect 12684 9774 12686 9826
rect 12738 9774 12964 9826
rect 12684 9772 12964 9774
rect 13132 10388 13188 10398
rect 13580 10388 13636 10398
rect 13132 9940 13188 10332
rect 12684 9762 12740 9772
rect 13020 9604 13076 9614
rect 12572 9314 12628 9324
rect 12908 9492 12964 9502
rect 12460 8990 12462 9042
rect 12514 8990 12516 9042
rect 12460 8978 12516 8990
rect 12684 9268 12740 9278
rect 12684 9042 12740 9212
rect 12684 8990 12686 9042
rect 12738 8990 12740 9042
rect 12348 8642 12404 8652
rect 12348 8484 12404 8494
rect 12180 8372 12292 8428
rect 12236 8260 12292 8372
rect 12124 8202 12180 8214
rect 12124 8150 12126 8202
rect 12178 8150 12180 8202
rect 12236 8194 12292 8204
rect 12124 8148 12180 8150
rect 12012 7924 12068 7934
rect 12012 7474 12068 7868
rect 12012 7422 12014 7474
rect 12066 7422 12068 7474
rect 12012 7410 12068 7422
rect 11900 7196 12068 7252
rect 11676 6850 11732 6860
rect 11452 6692 11508 6702
rect 11340 6690 11508 6692
rect 11340 6638 11454 6690
rect 11506 6638 11508 6690
rect 11900 6690 11956 6702
rect 11340 6636 11508 6638
rect 11452 6626 11508 6636
rect 11732 6634 11788 6646
rect 11564 6580 11620 6590
rect 10108 5238 10110 5290
rect 10162 5238 10164 5290
rect 10108 5226 10164 5238
rect 10332 5572 10388 5582
rect 10332 5236 10388 5516
rect 9528 4732 9792 4742
rect 9584 4676 9632 4732
rect 9688 4676 9736 4732
rect 9528 4666 9792 4676
rect 8428 4286 8430 4338
rect 8482 4286 8484 4338
rect 8428 4274 8484 4286
rect 9660 4340 9716 4350
rect 9660 4246 9716 4284
rect 9996 4338 10052 5180
rect 10332 5170 10388 5180
rect 10220 5122 10276 5134
rect 10220 5070 10222 5122
rect 10274 5070 10276 5122
rect 10220 4900 10276 5070
rect 10220 4834 10276 4844
rect 10444 5124 10500 6188
rect 10780 6188 11284 6244
rect 10668 6132 10724 6142
rect 10444 4562 10500 5068
rect 10556 5124 10612 5134
rect 10668 5124 10724 6076
rect 10556 5122 10724 5124
rect 10556 5070 10558 5122
rect 10610 5070 10724 5122
rect 10556 5068 10724 5070
rect 10556 5058 10612 5068
rect 10444 4510 10446 4562
rect 10498 4510 10500 4562
rect 10444 4498 10500 4510
rect 9996 4286 9998 4338
rect 10050 4286 10052 4338
rect 9996 4274 10052 4286
rect 10780 4338 10836 6188
rect 11004 6020 11060 6030
rect 11004 5906 11060 5964
rect 11004 5854 11006 5906
rect 11058 5854 11060 5906
rect 11004 5842 11060 5854
rect 11116 5908 11172 5918
rect 10986 5122 11042 5134
rect 10986 5070 10988 5122
rect 11040 5070 11042 5122
rect 10986 4900 11042 5070
rect 10986 4834 11042 4844
rect 11116 4562 11172 5852
rect 11228 5906 11284 6188
rect 11564 6020 11620 6524
rect 11732 6582 11734 6634
rect 11786 6582 11788 6634
rect 11732 6244 11788 6582
rect 11732 6178 11788 6188
rect 11900 6638 11902 6690
rect 11954 6638 11956 6690
rect 11900 6580 11956 6638
rect 11564 5954 11620 5964
rect 11228 5854 11230 5906
rect 11282 5854 11284 5906
rect 11228 5842 11284 5854
rect 11676 5908 11732 5918
rect 11676 5814 11732 5852
rect 11228 5684 11284 5694
rect 11228 5122 11284 5628
rect 11396 5684 11452 5694
rect 11396 5682 11620 5684
rect 11396 5630 11398 5682
rect 11450 5630 11620 5682
rect 11396 5628 11620 5630
rect 11396 5618 11452 5628
rect 11228 5070 11230 5122
rect 11282 5070 11284 5122
rect 11228 5058 11284 5070
rect 11116 4510 11118 4562
rect 11170 4510 11172 4562
rect 11116 4498 11172 4510
rect 11564 4954 11620 5628
rect 11732 5460 11788 5470
rect 11732 5178 11788 5404
rect 11732 5126 11734 5178
rect 11786 5126 11788 5178
rect 11732 5114 11788 5126
rect 11564 4902 11566 4954
rect 11618 4902 11620 4954
rect 10780 4286 10782 4338
rect 10834 4286 10836 4338
rect 10780 4274 10836 4286
rect 11452 4340 11508 4350
rect 11564 4340 11620 4902
rect 11452 4338 11620 4340
rect 11452 4286 11454 4338
rect 11506 4286 11620 4338
rect 11452 4284 11620 4286
rect 11676 5012 11732 5022
rect 11676 4338 11732 4956
rect 11676 4286 11678 4338
rect 11730 4286 11732 4338
rect 11452 4274 11508 4284
rect 11676 4274 11732 4286
rect 11788 4900 11844 4910
rect 11900 4900 11956 6524
rect 12012 6356 12068 7196
rect 12012 6290 12068 6300
rect 12012 6132 12068 6142
rect 12012 5348 12068 6076
rect 12124 5908 12180 8092
rect 12348 7812 12404 8428
rect 12684 8428 12740 8990
rect 12684 8372 12852 8428
rect 12572 8260 12628 8270
rect 12572 8202 12628 8204
rect 12572 8150 12574 8202
rect 12626 8150 12628 8202
rect 12572 8138 12628 8150
rect 12348 7746 12404 7756
rect 12348 7588 12404 7598
rect 12348 6466 12404 7532
rect 12460 7476 12516 7486
rect 12628 7476 12684 7486
rect 12460 7028 12516 7420
rect 12460 6962 12516 6972
rect 12572 7474 12684 7476
rect 12572 7422 12630 7474
rect 12682 7422 12684 7474
rect 12572 7410 12684 7422
rect 12796 7474 12852 8372
rect 12908 7700 12964 9436
rect 13020 8930 13076 9548
rect 13020 8878 13022 8930
rect 13074 8878 13076 8930
rect 13020 8866 13076 8878
rect 13132 8428 13188 9884
rect 13468 10386 13636 10388
rect 13468 10334 13582 10386
rect 13634 10334 13636 10386
rect 13468 10332 13636 10334
rect 13468 9268 13524 10332
rect 13580 10322 13636 10332
rect 14420 10386 14476 10398
rect 14420 10334 14422 10386
rect 14474 10334 14476 10386
rect 13686 10220 13950 10230
rect 13742 10164 13790 10220
rect 13846 10164 13894 10220
rect 13686 10154 13950 10164
rect 13468 9202 13524 9212
rect 13580 9938 13636 9950
rect 14420 9940 14476 10334
rect 13580 9886 13582 9938
rect 13634 9886 13636 9938
rect 13434 9079 13490 9091
rect 13434 9027 13436 9079
rect 13488 9027 13490 9079
rect 13434 8596 13490 9027
rect 13580 9042 13636 9886
rect 14364 9938 14476 9940
rect 14364 9886 14422 9938
rect 14474 9886 14476 9938
rect 14364 9874 14476 9886
rect 13580 8990 13582 9042
rect 13634 8990 13636 9042
rect 13580 8978 13636 8990
rect 13692 9044 13748 9054
rect 13692 8950 13748 8988
rect 14196 9044 14252 9054
rect 14196 8950 14252 8988
rect 14364 9042 14420 9874
rect 14364 8990 14366 9042
rect 14418 8990 14420 9042
rect 14364 8978 14420 8990
rect 14588 9044 14644 11452
rect 14700 11284 14756 11294
rect 14700 10610 14756 11228
rect 14700 10558 14702 10610
rect 14754 10558 14756 10610
rect 14700 10546 14756 10558
rect 14812 10612 14868 11564
rect 14980 11618 15036 11788
rect 14980 11566 14982 11618
rect 15034 11566 15036 11618
rect 14980 11554 15036 11566
rect 15820 11508 15876 13022
rect 15932 12935 15988 15484
rect 16380 15314 16436 15326
rect 16380 15262 16382 15314
rect 16434 15262 16436 15314
rect 16268 15204 16324 15214
rect 16100 13524 16156 13534
rect 16100 13522 16212 13524
rect 16100 13470 16102 13522
rect 16154 13470 16212 13522
rect 16100 13458 16212 13470
rect 15932 12883 15934 12935
rect 15986 12883 15988 12935
rect 15932 12292 15988 12883
rect 15932 12226 15988 12236
rect 16156 12180 16212 13458
rect 16268 13076 16324 15148
rect 16380 15148 16436 15262
rect 16380 15092 16548 15148
rect 16380 13746 16436 13758
rect 16380 13694 16382 13746
rect 16434 13694 16436 13746
rect 16380 13636 16436 13694
rect 16492 13748 16548 15036
rect 16604 13972 16660 18732
rect 17052 17668 17108 17678
rect 17052 17574 17108 17612
rect 16716 16772 16772 16782
rect 16716 15204 16772 16716
rect 16940 16100 16996 16110
rect 16940 16098 17108 16100
rect 16940 16046 16942 16098
rect 16994 16046 17108 16098
rect 16940 16044 17108 16046
rect 16940 16034 16996 16044
rect 16716 15110 16772 15148
rect 16604 13906 16660 13916
rect 16492 13654 16548 13692
rect 16660 13748 16716 13758
rect 16660 13654 16716 13692
rect 16828 13746 16884 13758
rect 16828 13694 16830 13746
rect 16882 13694 16884 13746
rect 16380 13524 16436 13580
rect 16716 13524 16772 13534
rect 16380 13468 16660 13524
rect 16268 12962 16324 13020
rect 16268 12910 16270 12962
rect 16322 12910 16324 12962
rect 16268 12898 16324 12910
rect 16604 12962 16660 13468
rect 16604 12910 16606 12962
rect 16658 12910 16660 12962
rect 16604 12898 16660 12910
rect 16380 12740 16436 12750
rect 16716 12740 16772 13468
rect 16828 12964 16884 13694
rect 16828 12898 16884 12908
rect 16940 13524 16996 13534
rect 16716 12684 16884 12740
rect 16156 12124 16324 12180
rect 16100 11956 16156 11966
rect 16100 11954 16212 11956
rect 16100 11902 16102 11954
rect 16154 11902 16212 11954
rect 16100 11890 16212 11902
rect 16044 11620 16100 11630
rect 16044 11562 16100 11564
rect 16044 11510 16046 11562
rect 16098 11510 16100 11562
rect 16044 11498 16100 11510
rect 15820 11442 15876 11452
rect 16156 11406 16212 11890
rect 15148 11396 15204 11406
rect 15148 10836 15204 11340
rect 15148 10770 15204 10780
rect 15260 11394 15316 11406
rect 15260 11342 15262 11394
rect 15314 11342 15316 11394
rect 14812 10518 14868 10556
rect 15260 9156 15316 11342
rect 15540 11396 15596 11406
rect 15540 11302 15596 11340
rect 15708 11394 15764 11406
rect 16100 11396 16212 11406
rect 15708 11342 15710 11394
rect 15762 11342 15764 11394
rect 15372 11282 15428 11294
rect 15372 11230 15374 11282
rect 15426 11230 15428 11282
rect 15372 10834 15428 11230
rect 15708 11060 15764 11342
rect 15372 10782 15374 10834
rect 15426 10782 15428 10834
rect 15372 10770 15428 10782
rect 15484 11004 15764 11060
rect 16044 11394 16212 11396
rect 16044 11342 16102 11394
rect 16154 11342 16212 11394
rect 16044 11340 16212 11342
rect 16044 11330 16156 11340
rect 15260 9100 15428 9156
rect 14588 8978 14644 8988
rect 15036 9044 15092 9054
rect 15148 9044 15204 9054
rect 15092 9042 15204 9044
rect 15092 8990 15150 9042
rect 15202 8990 15204 9042
rect 15092 8988 15204 8990
rect 14700 8818 14756 8830
rect 14700 8766 14702 8818
rect 14754 8766 14756 8818
rect 13686 8652 13950 8662
rect 13742 8596 13790 8652
rect 13846 8596 13894 8652
rect 13434 8540 13524 8596
rect 13686 8586 13950 8596
rect 12908 7634 12964 7644
rect 13020 8372 13188 8428
rect 13468 8428 13524 8540
rect 13468 8372 13748 8428
rect 12796 7422 12798 7474
rect 12850 7422 12852 7474
rect 12348 6414 12350 6466
rect 12402 6414 12404 6466
rect 12348 6402 12404 6414
rect 12124 5842 12180 5852
rect 12236 6356 12292 6366
rect 12236 5460 12292 6300
rect 12572 6244 12628 7410
rect 12796 7252 12852 7422
rect 12908 7476 12964 7486
rect 13020 7476 13076 8372
rect 13580 8258 13636 8270
rect 13580 8206 13582 8258
rect 13634 8206 13636 8258
rect 12908 7474 13076 7476
rect 12908 7422 12910 7474
rect 12962 7422 13076 7474
rect 12908 7420 13076 7422
rect 13356 7812 13412 7822
rect 12908 7410 12964 7420
rect 12796 7196 12964 7252
rect 12460 6188 12628 6244
rect 12740 6466 12796 6478
rect 12740 6414 12742 6466
rect 12794 6414 12796 6466
rect 12460 6132 12516 6188
rect 12460 6066 12516 6076
rect 12572 5908 12628 5918
rect 12740 5908 12796 6414
rect 12908 6018 12964 7196
rect 13188 7250 13244 7262
rect 13188 7198 13190 7250
rect 13242 7198 13244 7250
rect 13188 6692 13244 7198
rect 13188 6626 13244 6636
rect 13356 6690 13412 7756
rect 13580 7364 13636 8206
rect 13692 7812 13748 8372
rect 13916 8370 13972 8382
rect 13916 8318 13918 8370
rect 13970 8318 13972 8370
rect 13804 8214 13860 8226
rect 13804 8162 13806 8214
rect 13858 8162 13860 8214
rect 13804 8036 13860 8162
rect 13804 7970 13860 7980
rect 13916 7924 13972 8318
rect 14700 7924 14756 8766
rect 13916 7868 14644 7924
rect 13692 7756 14532 7812
rect 13580 7298 13636 7308
rect 14028 7509 14084 7521
rect 14028 7457 14030 7509
rect 14082 7457 14084 7509
rect 13356 6638 13358 6690
rect 13410 6638 13412 6690
rect 13356 6626 13412 6638
rect 13468 7252 13524 7262
rect 13468 6468 13524 7196
rect 14028 7252 14084 7457
rect 14196 7509 14252 7521
rect 14196 7457 14198 7509
rect 14250 7476 14252 7509
rect 14364 7502 14420 7514
rect 14250 7457 14308 7476
rect 14196 7420 14308 7457
rect 14028 7186 14084 7196
rect 13686 7084 13950 7094
rect 13742 7028 13790 7084
rect 13846 7028 13894 7084
rect 13686 7018 13950 7028
rect 13860 6916 13916 6926
rect 13860 6822 13916 6860
rect 14028 6804 14084 6814
rect 13580 6692 13636 6702
rect 13580 6598 13636 6636
rect 13804 6692 13860 6702
rect 12908 5966 12910 6018
rect 12962 5966 12964 6018
rect 12908 5954 12964 5966
rect 13300 6412 13524 6468
rect 13300 6018 13356 6412
rect 13300 5966 13302 6018
rect 13354 5966 13356 6018
rect 13300 5954 13356 5966
rect 13468 6244 13524 6254
rect 12236 5394 12292 5404
rect 12348 5906 12628 5908
rect 12348 5854 12574 5906
rect 12626 5854 12628 5906
rect 12348 5852 12628 5854
rect 12012 5124 12068 5292
rect 12124 5124 12180 5134
rect 12012 5122 12180 5124
rect 12012 5070 12126 5122
rect 12178 5070 12180 5122
rect 12012 5068 12180 5070
rect 12124 5058 12180 5068
rect 11900 4844 11990 4900
rect 11788 4338 11844 4844
rect 11788 4286 11790 4338
rect 11842 4286 11844 4338
rect 11934 4376 11990 4844
rect 11934 4324 11936 4376
rect 11988 4324 11990 4376
rect 11934 4312 11990 4324
rect 11788 4274 11844 4286
rect 7196 4172 7607 4228
rect 12348 4226 12404 5852
rect 12572 5842 12628 5852
rect 12684 5906 12796 5908
rect 12684 5854 12742 5906
rect 12794 5854 12796 5906
rect 12684 5842 12796 5854
rect 13020 5906 13076 5918
rect 13020 5854 13022 5906
rect 13074 5854 13076 5906
rect 12684 5684 12740 5842
rect 12460 5628 12740 5684
rect 12460 5346 12516 5628
rect 12460 5294 12462 5346
rect 12514 5294 12516 5346
rect 12460 5282 12516 5294
rect 13020 4340 13076 5854
rect 13468 5348 13524 6188
rect 13804 5796 13860 6636
rect 13804 5730 13860 5740
rect 13686 5516 13950 5526
rect 13742 5460 13790 5516
rect 13846 5460 13894 5516
rect 13686 5450 13950 5460
rect 14028 5348 14084 6748
rect 14252 6468 14308 7420
rect 14364 7450 14366 7502
rect 14418 7450 14420 7502
rect 14364 6916 14420 7450
rect 14364 6850 14420 6860
rect 14364 6692 14420 6702
rect 14364 6598 14420 6636
rect 14364 6468 14420 6478
rect 14252 6412 14364 6468
rect 14364 6402 14420 6412
rect 14476 6020 14532 7756
rect 14588 7530 14644 7868
rect 14700 7858 14756 7868
rect 14868 7924 14924 7934
rect 14588 7478 14590 7530
rect 14642 7478 14644 7530
rect 14868 7586 14924 7868
rect 14868 7534 14870 7586
rect 14922 7534 14924 7586
rect 14868 7522 14924 7534
rect 14588 7466 14644 7478
rect 14588 7252 14644 7262
rect 14588 6690 14644 7196
rect 15036 6916 15092 8988
rect 15148 8978 15204 8988
rect 15260 8932 15316 8942
rect 15260 8838 15316 8876
rect 15372 8708 15428 9100
rect 15148 8652 15428 8708
rect 15148 8372 15204 8652
rect 15484 8484 15540 11004
rect 16044 10948 16100 11330
rect 15820 10892 16100 10948
rect 15708 10836 15764 10846
rect 15596 9828 15652 9838
rect 15596 9098 15652 9772
rect 15596 9046 15598 9098
rect 15650 9046 15652 9098
rect 15596 9034 15652 9046
rect 15708 9826 15764 10780
rect 15820 10834 15876 10892
rect 15820 10782 15822 10834
rect 15874 10782 15876 10834
rect 15820 10770 15876 10782
rect 16268 10780 16324 12124
rect 16380 12178 16436 12684
rect 16492 12292 16548 12302
rect 16492 12198 16548 12236
rect 16660 12292 16716 12302
rect 16660 12234 16716 12236
rect 16380 12126 16382 12178
rect 16434 12126 16436 12178
rect 16660 12182 16662 12234
rect 16714 12182 16716 12234
rect 16660 12170 16716 12182
rect 16828 12178 16884 12684
rect 16380 12114 16436 12126
rect 16828 12126 16830 12178
rect 16882 12126 16884 12178
rect 16828 12068 16884 12126
rect 16828 12002 16884 12012
rect 16940 11844 16996 13468
rect 16896 11788 16996 11844
rect 15708 9774 15710 9826
rect 15762 9774 15764 9826
rect 15148 8278 15204 8316
rect 15260 8428 15540 8484
rect 14588 6638 14590 6690
rect 14642 6638 14644 6690
rect 14588 6626 14644 6638
rect 14700 6860 15092 6916
rect 14476 5954 14532 5964
rect 13468 5292 13692 5348
rect 13636 5236 13692 5292
rect 13636 5142 13692 5180
rect 13804 5292 14084 5348
rect 13804 5122 13860 5292
rect 13804 5070 13806 5122
rect 13858 5070 13860 5122
rect 13804 5058 13860 5070
rect 13020 4274 13076 4284
rect 14028 4338 14084 5292
rect 14588 5236 14644 5246
rect 14588 5142 14644 5180
rect 14028 4286 14030 4338
rect 14082 4286 14084 4338
rect 14028 4274 14084 4286
rect 12348 4174 12350 4226
rect 12402 4174 12404 4226
rect 12348 4162 12404 4174
rect 4396 3658 4452 3670
rect 5684 3666 5796 3678
rect 5684 3614 5686 3666
rect 5738 3614 5796 3666
rect 5684 3612 5796 3614
rect 5852 4114 5908 4126
rect 5852 4062 5854 4114
rect 5906 4062 5908 4114
rect 5684 3602 5740 3612
rect 4508 3556 4564 3566
rect 4508 3462 4564 3500
rect 4844 3554 4900 3566
rect 4844 3502 4846 3554
rect 4898 3502 4900 3554
rect 4844 3444 4900 3502
rect 5852 3556 5908 4062
rect 13686 3948 13950 3958
rect 13742 3892 13790 3948
rect 13846 3892 13894 3948
rect 13686 3882 13950 3892
rect 11228 3780 11284 3790
rect 10892 3556 10948 3566
rect 5852 3490 5908 3500
rect 10780 3554 10948 3556
rect 10780 3502 10894 3554
rect 10946 3502 10948 3554
rect 10780 3500 10948 3502
rect 10780 3454 10836 3500
rect 10892 3490 10948 3500
rect 4844 3378 4900 3388
rect 6132 3444 6188 3454
rect 6132 3350 6188 3388
rect 10724 3442 10836 3454
rect 10724 3390 10726 3442
rect 10778 3390 10836 3442
rect 10724 3378 10836 3390
rect 11228 3444 11284 3724
rect 14700 3780 14756 6860
rect 15036 6692 15092 6702
rect 14868 6578 14924 6590
rect 14868 6526 14870 6578
rect 14922 6526 14924 6578
rect 14868 6468 14924 6526
rect 14868 6402 14924 6412
rect 14868 6074 14924 6086
rect 14868 6022 14870 6074
rect 14922 6022 14924 6074
rect 14868 6020 14924 6022
rect 14868 5954 14924 5964
rect 15036 5906 15092 6636
rect 15036 5854 15038 5906
rect 15090 5854 15092 5906
rect 15036 5842 15092 5854
rect 15260 6244 15316 8428
rect 15596 8258 15652 8270
rect 15484 8202 15540 8214
rect 15484 8150 15486 8202
rect 15538 8150 15540 8202
rect 15372 7252 15428 7262
rect 15372 7158 15428 7196
rect 15372 6692 15428 6702
rect 15372 6598 15428 6636
rect 15484 6468 15540 8150
rect 15596 8206 15598 8258
rect 15650 8206 15652 8258
rect 15596 7924 15652 8206
rect 15596 7858 15652 7868
rect 15708 7700 15764 9774
rect 15932 10724 16324 10780
rect 16380 11508 16436 11518
rect 15932 9787 15988 10724
rect 15932 9735 15934 9787
rect 15986 9735 15988 9787
rect 15820 9044 15876 9054
rect 15932 9044 15988 9735
rect 15820 9042 15988 9044
rect 15820 8990 15822 9042
rect 15874 8990 15988 9042
rect 15820 8988 15988 8990
rect 16044 9938 16100 9950
rect 16044 9886 16046 9938
rect 16098 9886 16100 9938
rect 15820 8978 15876 8988
rect 15932 8260 15988 8270
rect 15932 8166 15988 8204
rect 15596 7644 15764 7700
rect 15932 7812 15988 7822
rect 15596 6916 15652 7644
rect 15764 7476 15820 7486
rect 15764 7382 15820 7420
rect 15932 7474 15988 7756
rect 15932 7422 15934 7474
rect 15986 7422 15988 7474
rect 15932 7410 15988 7422
rect 16044 7474 16100 9886
rect 16380 9828 16436 11452
rect 16896 11356 16952 11788
rect 16896 11304 16898 11356
rect 16950 11304 16952 11356
rect 16896 11292 16952 11304
rect 17052 11732 17108 16044
rect 17164 15092 17220 20132
rect 18172 20018 18228 21308
rect 18284 20188 18340 23884
rect 18956 23826 19012 23838
rect 18956 23774 18958 23826
rect 19010 23774 19012 23826
rect 18508 23192 18564 23204
rect 18508 23140 18510 23192
rect 18562 23140 18564 23192
rect 18508 23044 18564 23140
rect 18956 23156 19012 23774
rect 18956 23090 19012 23100
rect 19292 23154 19348 24108
rect 19516 24052 19572 24062
rect 19516 23900 19572 23996
rect 19628 23994 19684 24444
rect 19628 23942 19630 23994
rect 19682 23942 19684 23994
rect 19628 23930 19684 23942
rect 19852 24388 19908 24780
rect 20412 24388 20468 24398
rect 19852 24332 20188 24388
rect 19516 23848 19518 23900
rect 19570 23848 19572 23900
rect 19516 23836 19572 23848
rect 19292 23102 19294 23154
rect 19346 23102 19348 23154
rect 19292 23090 19348 23102
rect 19628 23156 19684 23166
rect 19852 23156 19908 24332
rect 20132 23994 20188 24332
rect 19628 23154 19908 23156
rect 19628 23102 19630 23154
rect 19682 23102 19908 23154
rect 19628 23100 19908 23102
rect 19964 23938 20020 23950
rect 19964 23886 19966 23938
rect 20018 23886 20020 23938
rect 20132 23942 20134 23994
rect 20186 23942 20188 23994
rect 20132 23930 20188 23942
rect 20412 23938 20468 24332
rect 20748 24174 20804 24892
rect 20692 24162 20804 24174
rect 20692 24110 20694 24162
rect 20746 24110 20804 24162
rect 20692 24108 20804 24110
rect 20692 24098 20748 24108
rect 19628 23090 19684 23100
rect 18508 22978 18564 22988
rect 19180 23044 19236 23054
rect 19180 22986 19236 22988
rect 19180 22934 19182 22986
rect 19234 22934 19236 22986
rect 19180 22820 19236 22934
rect 19068 22764 19236 22820
rect 18508 22482 18564 22494
rect 18508 22430 18510 22482
rect 18562 22430 18564 22482
rect 18508 22036 18564 22430
rect 19068 22370 19124 22764
rect 19964 22484 20020 23886
rect 20412 23886 20414 23938
rect 20466 23886 20468 23938
rect 20412 23874 20468 23886
rect 20300 23828 20356 23838
rect 20300 23734 20356 23772
rect 20860 23548 20916 25340
rect 20972 24722 21028 25564
rect 20972 24670 20974 24722
rect 21026 24670 21028 24722
rect 20972 24658 21028 24670
rect 21084 24724 21140 27020
rect 21196 27010 21252 27020
rect 21308 26414 21364 27804
rect 21532 27634 21588 27646
rect 21532 27582 21534 27634
rect 21586 27582 21588 27634
rect 21532 27188 21588 27582
rect 22002 27468 22266 27478
rect 22058 27412 22106 27468
rect 22162 27412 22210 27468
rect 22002 27402 22266 27412
rect 21532 27122 21588 27132
rect 21980 27188 22036 27198
rect 21980 27094 22036 27132
rect 23212 26514 23268 29372
rect 23324 29362 23380 29372
rect 23436 29542 23438 29594
rect 23490 29542 23492 29594
rect 23324 28644 23380 28654
rect 23436 28644 23492 29542
rect 23660 29453 23716 29465
rect 23660 29401 23662 29453
rect 23714 29401 23716 29453
rect 23996 29428 24052 30044
rect 24332 30098 24388 30156
rect 24332 30046 24334 30098
rect 24386 30046 24388 30098
rect 23660 29316 23716 29401
rect 23660 29250 23716 29260
rect 23884 29426 24052 29428
rect 23884 29374 23998 29426
rect 24050 29374 24052 29426
rect 23884 29372 24052 29374
rect 23884 28868 23940 29372
rect 23996 29362 24052 29372
rect 24108 29428 24164 29438
rect 24332 29428 24388 30046
rect 24164 29372 24388 29428
rect 23324 28642 23492 28644
rect 23324 28590 23326 28642
rect 23378 28590 23492 28642
rect 23324 28588 23492 28590
rect 23660 28812 23940 28868
rect 23324 28578 23380 28588
rect 23660 27860 23716 28812
rect 23996 28754 24052 28766
rect 23996 28702 23998 28754
rect 24050 28702 24052 28754
rect 23772 28642 23828 28654
rect 23772 28590 23774 28642
rect 23826 28590 23828 28642
rect 23772 28084 23828 28590
rect 23772 28028 23940 28084
rect 23772 27860 23828 27870
rect 23660 27858 23828 27860
rect 23660 27806 23774 27858
rect 23826 27806 23828 27858
rect 23660 27804 23828 27806
rect 23772 27794 23828 27804
rect 23884 27858 23940 28028
rect 23884 27806 23886 27858
rect 23938 27806 23940 27858
rect 23492 27634 23548 27646
rect 23492 27582 23494 27634
rect 23546 27582 23548 27634
rect 23492 27076 23548 27582
rect 23884 27186 23940 27806
rect 23884 27134 23886 27186
rect 23938 27134 23940 27186
rect 23884 27122 23940 27134
rect 23492 27010 23548 27020
rect 23212 26462 23214 26514
rect 23266 26462 23268 26514
rect 23212 26450 23268 26462
rect 21252 26402 21364 26414
rect 21252 26350 21254 26402
rect 21306 26350 21364 26402
rect 21252 26348 21364 26350
rect 21252 26338 21308 26348
rect 23884 26305 23940 26317
rect 21868 26292 21924 26302
rect 22876 26292 22932 26302
rect 21868 25732 21924 26236
rect 22764 26290 22932 26292
rect 22764 26238 22878 26290
rect 22930 26238 22932 26290
rect 22764 26236 22932 26238
rect 22002 25900 22266 25910
rect 22058 25844 22106 25900
rect 22162 25844 22210 25900
rect 22002 25834 22266 25844
rect 21868 25676 22036 25732
rect 21084 24658 21140 24668
rect 21756 24724 21812 24734
rect 21756 24630 21812 24668
rect 21980 24554 22036 25676
rect 21980 24502 21982 24554
rect 22034 24502 22036 24554
rect 21980 24490 22036 24502
rect 22092 25060 22148 25070
rect 22092 24722 22148 25004
rect 22092 24670 22094 24722
rect 22146 24670 22148 24722
rect 22092 24500 22148 24670
rect 22092 24434 22148 24444
rect 22428 24836 22484 24846
rect 22428 24722 22484 24780
rect 22428 24670 22430 24722
rect 22482 24670 22484 24722
rect 22002 24332 22266 24342
rect 22058 24276 22106 24332
rect 22162 24276 22210 24332
rect 22002 24266 22266 24276
rect 22428 23828 22484 24670
rect 22652 23940 22708 23950
rect 22764 23940 22820 26236
rect 22876 26226 22932 26236
rect 23884 26253 23886 26305
rect 23938 26253 23940 26305
rect 23772 26180 23828 26190
rect 23548 26178 23828 26180
rect 23548 26126 23774 26178
rect 23826 26126 23828 26178
rect 23548 26124 23828 26126
rect 23380 25282 23436 25294
rect 23380 25230 23382 25282
rect 23434 25230 23436 25282
rect 23380 25172 23436 25230
rect 23212 25116 23436 25172
rect 22988 24836 23044 24846
rect 22988 24766 23044 24780
rect 22988 24714 22990 24766
rect 23042 24714 23044 24766
rect 22988 24702 23044 24714
rect 22876 24612 22932 24622
rect 22876 24518 22932 24556
rect 22652 23938 22820 23940
rect 22652 23886 22654 23938
rect 22706 23886 22820 23938
rect 22652 23884 22820 23886
rect 22652 23874 22708 23884
rect 22428 23762 22484 23772
rect 20636 23492 21588 23548
rect 20132 23380 20188 23390
rect 20636 23380 20692 23492
rect 20188 23324 20356 23380
rect 20132 23314 20188 23324
rect 20300 23154 20356 23324
rect 20300 23102 20302 23154
rect 20354 23102 20356 23154
rect 20300 23090 20356 23102
rect 20412 23378 20692 23380
rect 20412 23326 20638 23378
rect 20690 23326 20692 23378
rect 20412 23324 20692 23326
rect 19964 22418 20020 22428
rect 18396 21980 18564 22036
rect 18902 22314 18958 22326
rect 18902 22262 18904 22314
rect 18956 22262 18958 22314
rect 19068 22318 19070 22370
rect 19122 22318 19124 22370
rect 19068 22306 19124 22318
rect 19180 22372 19236 22382
rect 19180 22278 19236 22316
rect 18396 21364 18452 21980
rect 18564 21812 18620 21822
rect 18564 21718 18620 21756
rect 18902 21812 18958 22262
rect 18902 21746 18958 21756
rect 19852 21812 19908 21822
rect 18396 21298 18452 21308
rect 18732 21586 18788 21598
rect 18732 21534 18734 21586
rect 18786 21534 18788 21586
rect 18284 20132 18452 20188
rect 18172 19966 18174 20018
rect 18226 19966 18228 20018
rect 17892 19796 17948 19806
rect 17500 19794 17948 19796
rect 17500 19742 17894 19794
rect 17946 19742 17948 19794
rect 17500 19740 17948 19742
rect 17276 19234 17332 19246
rect 17276 19182 17278 19234
rect 17330 19182 17332 19234
rect 17276 17892 17332 19182
rect 17500 18452 17556 19740
rect 17892 19730 17948 19740
rect 17276 17826 17332 17836
rect 17388 18450 17556 18452
rect 17388 18398 17502 18450
rect 17554 18398 17556 18450
rect 17388 18396 17556 18398
rect 17388 17666 17444 18396
rect 17500 18386 17556 18396
rect 17612 19346 17668 19358
rect 17612 19294 17614 19346
rect 17666 19294 17668 19346
rect 17388 17614 17390 17666
rect 17442 17614 17444 17666
rect 17388 17602 17444 17614
rect 17500 17892 17556 17902
rect 17164 15026 17220 15036
rect 17500 15314 17556 17836
rect 17500 15262 17502 15314
rect 17554 15262 17556 15314
rect 17052 9828 17108 11676
rect 16380 9734 16436 9772
rect 16828 9826 17108 9828
rect 16828 9774 17054 9826
rect 17106 9774 17108 9826
rect 16828 9772 17108 9774
rect 16828 8428 16884 9772
rect 17052 9762 17108 9772
rect 17276 14308 17332 14318
rect 17276 9268 17332 14252
rect 17500 13748 17556 15262
rect 17500 13682 17556 13692
rect 17444 13524 17500 13534
rect 17444 13430 17500 13468
rect 17612 13188 17668 19294
rect 17948 19236 18004 19246
rect 18172 19236 18228 19966
rect 18396 20018 18452 20132
rect 18396 19966 18398 20018
rect 18450 19966 18452 20018
rect 17948 19234 18228 19236
rect 17724 19178 17780 19190
rect 17724 19126 17726 19178
rect 17778 19126 17780 19178
rect 17948 19182 17950 19234
rect 18002 19182 18228 19234
rect 17948 19180 18228 19182
rect 18284 19236 18340 19246
rect 17948 19170 18004 19180
rect 18284 19142 18340 19180
rect 17724 19012 17780 19126
rect 18396 19012 18452 19966
rect 18732 19236 18788 21534
rect 19740 20578 19796 20590
rect 19740 20526 19742 20578
rect 19794 20526 19796 20578
rect 19740 20188 19796 20526
rect 19628 20132 19796 20188
rect 18844 20020 18900 20030
rect 18844 19926 18900 19964
rect 19628 20018 19684 20132
rect 19628 19966 19630 20018
rect 19682 19966 19684 20018
rect 19628 19954 19684 19966
rect 18732 19170 18788 19180
rect 19404 19908 19460 19918
rect 19404 19219 19460 19852
rect 17724 18956 18452 19012
rect 19404 19167 19406 19219
rect 19458 19167 19460 19219
rect 17844 18844 18108 18854
rect 17900 18788 17948 18844
rect 18004 18788 18052 18844
rect 17844 18778 18108 18788
rect 17724 18676 17780 18686
rect 17724 18450 17780 18620
rect 18844 18564 18900 18574
rect 17724 18398 17726 18450
rect 17778 18398 17780 18450
rect 17724 18340 17780 18398
rect 18172 18477 18228 18489
rect 18172 18425 18174 18477
rect 18226 18425 18228 18477
rect 17724 18274 17780 18284
rect 17836 18282 17892 18294
rect 17836 18230 17838 18282
rect 17890 18230 17892 18282
rect 17724 18116 17780 18126
rect 17724 17108 17780 18060
rect 17836 17668 17892 18230
rect 17836 17602 17892 17612
rect 17892 17444 17948 17454
rect 18172 17444 18228 18425
rect 18508 18004 18564 18014
rect 18508 17666 18564 17948
rect 18508 17614 18510 17666
rect 18562 17614 18564 17666
rect 18508 17602 18564 17614
rect 18620 17834 18676 17846
rect 18620 17782 18622 17834
rect 18674 17782 18676 17834
rect 17892 17442 18228 17444
rect 17892 17390 17894 17442
rect 17946 17390 18228 17442
rect 17892 17388 18228 17390
rect 17892 17378 17948 17388
rect 18172 17332 18228 17388
rect 18620 17332 18676 17782
rect 18844 17666 18900 18508
rect 19404 18564 19460 19167
rect 19740 19236 19796 19246
rect 19740 19142 19796 19180
rect 19404 18498 19460 18508
rect 19628 19066 19684 19078
rect 19628 19014 19630 19066
rect 19682 19014 19684 19066
rect 19516 18452 19572 18462
rect 19516 18226 19572 18396
rect 19516 18174 19518 18226
rect 19570 18174 19572 18226
rect 19348 17892 19404 17902
rect 19348 17798 19404 17836
rect 18844 17614 18846 17666
rect 18898 17614 18900 17666
rect 18844 17602 18900 17614
rect 18956 17668 19012 17678
rect 17844 17276 18108 17286
rect 18172 17276 18340 17332
rect 17900 17220 17948 17276
rect 18004 17220 18052 17276
rect 17844 17210 18108 17220
rect 17836 17108 17892 17118
rect 17724 17052 17836 17108
rect 17836 17014 17892 17052
rect 18172 16884 18228 16894
rect 17724 16882 18228 16884
rect 17724 16830 18174 16882
rect 18226 16830 18228 16882
rect 17724 16828 18228 16830
rect 17724 16100 17780 16828
rect 18172 16818 18228 16828
rect 18284 16660 18340 17276
rect 18508 17276 18676 17332
rect 18732 17332 18788 17342
rect 18396 16882 18452 16894
rect 18396 16830 18398 16882
rect 18450 16830 18452 16882
rect 18396 16772 18452 16830
rect 18508 16882 18564 17276
rect 18732 16940 18788 17276
rect 18508 16830 18510 16882
rect 18562 16830 18564 16882
rect 18694 16920 18788 16940
rect 18694 16868 18696 16920
rect 18748 16884 18788 16920
rect 18748 16868 18750 16884
rect 18694 16856 18750 16868
rect 18508 16818 18564 16830
rect 18396 16706 18452 16716
rect 17724 14308 17780 16044
rect 18172 16604 18340 16660
rect 17844 15708 18108 15718
rect 17900 15652 17948 15708
rect 18004 15652 18052 15708
rect 17844 15642 18108 15652
rect 17836 15540 17892 15550
rect 17836 15446 17892 15484
rect 18172 15204 18228 16604
rect 18844 16098 18900 16110
rect 18844 16046 18846 16098
rect 18898 16046 18900 16098
rect 18844 15540 18900 16046
rect 18956 16100 19012 17612
rect 19516 17668 19572 18174
rect 19516 17602 19572 17612
rect 19628 17666 19684 19014
rect 19852 18900 19908 21756
rect 20412 21364 20468 23324
rect 20636 23314 20692 23324
rect 21420 21812 21476 21822
rect 21420 21586 21476 21756
rect 21420 21534 21422 21586
rect 21474 21534 21476 21586
rect 21420 21522 21476 21534
rect 21532 21586 21588 23492
rect 22204 23181 22260 23193
rect 22204 23129 22206 23181
rect 22258 23129 22260 23181
rect 21924 23044 21980 23054
rect 22204 23044 22260 23129
rect 21868 23042 22260 23044
rect 21868 22990 21926 23042
rect 21978 22990 22260 23042
rect 21868 22988 22260 22990
rect 21868 22978 21980 22988
rect 21868 22596 21924 22978
rect 22002 22764 22266 22774
rect 22058 22708 22106 22764
rect 22162 22708 22210 22764
rect 22002 22698 22266 22708
rect 22764 22596 22820 23884
rect 21868 22540 22036 22596
rect 21868 21812 21924 21822
rect 21532 21534 21534 21586
rect 21586 21534 21588 21586
rect 21532 21522 21588 21534
rect 21756 21756 21868 21812
rect 20300 21308 20468 21364
rect 21084 21362 21140 21374
rect 21084 21310 21086 21362
rect 21138 21310 21140 21362
rect 20076 20804 20132 20814
rect 20076 20710 20132 20748
rect 20300 20802 20356 21308
rect 20300 20750 20302 20802
rect 20354 20750 20356 20802
rect 20300 20738 20356 20750
rect 20412 20802 20468 20814
rect 20412 20750 20414 20802
rect 20466 20750 20468 20802
rect 20412 20188 20468 20750
rect 20692 20690 20748 20702
rect 20692 20638 20694 20690
rect 20746 20638 20748 20690
rect 20692 20580 20748 20638
rect 20692 20514 20748 20524
rect 20412 20132 20804 20188
rect 19964 19234 20020 19246
rect 19964 19182 19966 19234
rect 20018 19182 20020 19234
rect 19964 19124 20020 19182
rect 19964 19058 20020 19068
rect 20300 19010 20356 19022
rect 20300 18958 20302 19010
rect 20354 18958 20356 19010
rect 19852 18844 20132 18900
rect 19628 17614 19630 17666
rect 19682 17614 19684 17666
rect 20076 17666 20132 18844
rect 20300 18564 20356 18958
rect 20300 18498 20356 18508
rect 20748 18452 20804 20132
rect 21084 19460 21140 21310
rect 21644 21028 21700 21038
rect 21364 20804 21420 20814
rect 21364 20710 21420 20748
rect 21644 20802 21700 20972
rect 21644 20750 21646 20802
rect 21698 20750 21700 20802
rect 21644 20738 21700 20750
rect 21756 20802 21812 21756
rect 21868 21718 21924 21756
rect 21980 21364 22036 22540
rect 22540 22540 22820 22596
rect 22988 24500 23044 24510
rect 22988 23714 23044 24444
rect 23212 24500 23268 25116
rect 23548 25060 23604 26124
rect 23772 26114 23828 26124
rect 23884 25508 23940 26253
rect 23996 26292 24052 28702
rect 24108 28615 24164 29372
rect 24108 28563 24110 28615
rect 24162 28563 24164 28615
rect 24444 28644 24500 28654
rect 24556 28644 24612 30830
rect 25340 30884 25396 30894
rect 25340 30790 25396 30828
rect 24668 30212 24724 30222
rect 24668 30118 24724 30156
rect 24892 30210 24948 30222
rect 24892 30158 24894 30210
rect 24946 30158 24948 30210
rect 24892 29988 24948 30158
rect 25172 30100 25228 30110
rect 25172 30006 25228 30044
rect 24892 29922 24948 29932
rect 25788 29594 25844 30940
rect 27244 30994 27300 31006
rect 27244 30942 27246 30994
rect 27298 30942 27300 30994
rect 27244 30548 27300 30942
rect 27580 30772 27636 30782
rect 27580 30770 27972 30772
rect 27580 30718 27582 30770
rect 27634 30718 27972 30770
rect 27580 30716 27972 30718
rect 27580 30706 27636 30716
rect 27244 30492 27748 30548
rect 26012 30098 26068 30110
rect 26012 30046 26014 30098
rect 26066 30046 26068 30098
rect 25228 29540 25284 29550
rect 25788 29542 25790 29594
rect 25842 29542 25844 29594
rect 25788 29530 25844 29542
rect 25900 29988 25956 29998
rect 25228 29426 25284 29484
rect 25564 29453 25620 29465
rect 25228 29374 25230 29426
rect 25282 29374 25284 29426
rect 25228 29362 25284 29374
rect 25452 29428 25508 29438
rect 24444 28642 24556 28644
rect 24444 28590 24446 28642
rect 24498 28590 24556 28642
rect 24444 28588 24556 28590
rect 24444 28578 24500 28588
rect 24108 28551 24164 28563
rect 24556 28550 24612 28588
rect 24780 28756 24836 28766
rect 24780 28642 24836 28700
rect 24780 28590 24782 28642
rect 24834 28590 24836 28642
rect 24780 28578 24836 28590
rect 25228 28644 25284 28654
rect 25228 27858 25284 28588
rect 25452 28642 25508 29372
rect 25452 28590 25454 28642
rect 25506 28590 25508 28642
rect 25452 27972 25508 28590
rect 25564 29401 25566 29453
rect 25618 29401 25620 29453
rect 25564 28308 25620 29401
rect 25900 29426 25956 29932
rect 25900 29374 25902 29426
rect 25954 29374 25956 29426
rect 25732 28868 25788 28878
rect 25900 28868 25956 29374
rect 25732 28866 25956 28868
rect 25732 28814 25734 28866
rect 25786 28814 25956 28866
rect 25732 28812 25956 28814
rect 25732 28802 25788 28812
rect 26012 28756 26068 30046
rect 26160 29820 26424 29830
rect 26216 29764 26264 29820
rect 26320 29764 26368 29820
rect 26160 29754 26424 29764
rect 27692 29594 27748 30492
rect 27916 30322 27972 30716
rect 30318 30604 30582 30614
rect 30374 30548 30422 30604
rect 30478 30548 30526 30604
rect 30318 30538 30582 30548
rect 27916 30270 27918 30322
rect 27970 30270 27972 30322
rect 27916 30258 27972 30270
rect 28700 30212 28756 30222
rect 29316 30212 29372 30222
rect 28700 30210 29540 30212
rect 28700 30158 28702 30210
rect 28754 30158 29318 30210
rect 29370 30158 29540 30210
rect 28700 30156 29540 30158
rect 28700 30146 28756 30156
rect 29316 30146 29372 30156
rect 26796 29540 26852 29550
rect 27692 29542 27694 29594
rect 27746 29542 27748 29594
rect 27692 29530 27748 29542
rect 26796 29428 26852 29484
rect 27244 29453 27300 29465
rect 26908 29428 26964 29438
rect 26796 29426 26964 29428
rect 26796 29374 26910 29426
rect 26962 29374 26964 29426
rect 26796 29372 26964 29374
rect 26012 28690 26068 28700
rect 26684 28756 26740 28766
rect 26684 28642 26740 28700
rect 26684 28590 26686 28642
rect 26738 28590 26740 28642
rect 26684 28578 26740 28590
rect 25564 28252 25732 28308
rect 25452 27916 25564 27972
rect 25228 27806 25230 27858
rect 25282 27806 25284 27858
rect 25508 27914 25564 27916
rect 25508 27862 25510 27914
rect 25562 27862 25564 27914
rect 25508 27850 25564 27862
rect 25228 27794 25284 27806
rect 25676 27746 25732 28252
rect 26160 28252 26424 28262
rect 26216 28196 26264 28252
rect 26320 28196 26368 28252
rect 26160 28186 26424 28196
rect 26796 27858 26852 29372
rect 26908 29362 26964 29372
rect 27244 29401 27246 29453
rect 27298 29401 27300 29453
rect 27132 28756 27188 28766
rect 27244 28756 27300 29401
rect 27580 29428 27636 29438
rect 27580 29334 27636 29372
rect 29036 29428 29092 29438
rect 27132 28754 27300 28756
rect 27132 28702 27134 28754
rect 27186 28702 27300 28754
rect 27132 28700 27300 28702
rect 27356 28756 27412 28766
rect 27132 28690 27188 28700
rect 27356 28642 27412 28700
rect 27020 28598 27076 28610
rect 27020 28546 27022 28598
rect 27074 28546 27076 28598
rect 27356 28590 27358 28642
rect 27410 28590 27412 28642
rect 27356 28578 27412 28590
rect 27580 28642 27636 28654
rect 27580 28590 27582 28642
rect 27634 28590 27636 28642
rect 27020 28196 27076 28546
rect 27580 28196 27636 28590
rect 27860 28532 27916 28542
rect 27860 28438 27916 28476
rect 28700 28532 28756 28542
rect 27020 28140 27524 28196
rect 26796 27806 26798 27858
rect 26850 27806 26852 27858
rect 26796 27794 26852 27806
rect 27020 28026 27076 28038
rect 27020 27974 27022 28026
rect 27074 27974 27076 28026
rect 25676 27694 25678 27746
rect 25730 27694 25732 27746
rect 25676 27682 25732 27694
rect 25116 27076 25172 27086
rect 25004 27074 25172 27076
rect 25004 27022 25118 27074
rect 25170 27022 25172 27074
rect 25004 27020 25172 27022
rect 24108 26292 24164 26302
rect 23996 26290 24164 26292
rect 23996 26238 24110 26290
rect 24162 26238 24164 26290
rect 23996 26236 24164 26238
rect 23996 25508 24052 25518
rect 23884 25452 23996 25508
rect 23996 25414 24052 25452
rect 24108 25506 24164 26236
rect 24556 25620 24612 25630
rect 24108 25454 24110 25506
rect 24162 25454 24164 25506
rect 24108 25442 24164 25454
rect 24444 25506 24500 25518
rect 24444 25454 24446 25506
rect 24498 25454 24500 25506
rect 23716 25396 23772 25406
rect 23716 25394 23828 25396
rect 23716 25342 23718 25394
rect 23770 25342 23828 25394
rect 23716 25330 23828 25342
rect 23548 24994 23604 25004
rect 23324 24948 23380 24958
rect 23324 24722 23380 24892
rect 23324 24670 23326 24722
rect 23378 24670 23380 24722
rect 23324 24658 23380 24670
rect 23436 24724 23492 24734
rect 23212 24434 23268 24444
rect 22988 23662 22990 23714
rect 23042 23662 23044 23714
rect 22428 22370 22484 22382
rect 22428 22318 22430 22370
rect 22482 22318 22484 22370
rect 22428 21812 22484 22318
rect 22428 21746 22484 21756
rect 21980 21298 22036 21308
rect 22002 21196 22266 21206
rect 22058 21140 22106 21196
rect 22162 21140 22210 21196
rect 22540 21140 22596 22540
rect 22876 22538 22932 22550
rect 22876 22486 22878 22538
rect 22930 22486 22932 22538
rect 22764 22372 22820 22382
rect 22764 22278 22820 22316
rect 22876 22036 22932 22486
rect 22876 21970 22932 21980
rect 22988 21700 23044 23662
rect 23436 23940 23492 24668
rect 23660 24722 23716 24734
rect 23660 24670 23662 24722
rect 23714 24670 23716 24722
rect 23660 24500 23716 24670
rect 23660 24434 23716 24444
rect 23660 24052 23716 24062
rect 23772 24052 23828 25330
rect 24444 25060 24500 25454
rect 24556 25506 24612 25564
rect 24556 25454 24558 25506
rect 24610 25454 24612 25506
rect 24556 25442 24612 25454
rect 24444 24994 24500 25004
rect 24836 25394 24892 25406
rect 24836 25342 24838 25394
rect 24890 25342 24892 25394
rect 24444 24890 24500 24902
rect 24332 24836 24388 24846
rect 23996 24749 24052 24761
rect 23996 24697 23998 24749
rect 24050 24697 24052 24749
rect 23996 24612 24052 24697
rect 24332 24722 24388 24780
rect 24332 24670 24334 24722
rect 24386 24670 24388 24722
rect 24332 24658 24388 24670
rect 24444 24838 24446 24890
rect 24498 24838 24500 24890
rect 23996 24546 24052 24556
rect 24444 24500 24500 24838
rect 24836 24836 24892 25342
rect 24836 24770 24892 24780
rect 25004 24724 25060 27020
rect 25116 27010 25172 27020
rect 25900 27074 25956 27086
rect 25900 27022 25902 27074
rect 25954 27022 25956 27074
rect 25900 26516 25956 27022
rect 26160 26684 26424 26694
rect 26216 26628 26264 26684
rect 26320 26628 26368 26684
rect 26160 26618 26424 26628
rect 26572 26516 26628 26526
rect 25900 26514 26628 26516
rect 25900 26462 26574 26514
rect 26626 26462 26628 26514
rect 25900 26460 26628 26462
rect 26572 26450 26628 26460
rect 26908 26292 26964 26302
rect 27020 26292 27076 27974
rect 27468 27972 27524 28140
rect 27580 28130 27636 28140
rect 28476 28196 28532 28206
rect 28084 27972 28140 27982
rect 27468 27970 28140 27972
rect 27468 27918 28086 27970
rect 28138 27918 28140 27970
rect 27468 27916 28140 27918
rect 26908 26290 27076 26292
rect 26908 26238 26910 26290
rect 26962 26238 27076 26290
rect 26908 26236 27076 26238
rect 27244 27897 27300 27909
rect 27244 27845 27246 27897
rect 27298 27845 27300 27897
rect 26908 26226 26964 26236
rect 27244 26180 27300 27845
rect 27468 27858 27524 27916
rect 28084 27906 28140 27916
rect 27468 27806 27470 27858
rect 27522 27806 27524 27858
rect 27468 27794 27524 27806
rect 28364 27860 28420 27870
rect 28364 27300 28420 27804
rect 28140 27244 28420 27300
rect 28476 27858 28532 28140
rect 28476 27806 28478 27858
rect 28530 27806 28532 27858
rect 27804 27188 27860 27198
rect 27580 26305 27636 26317
rect 27580 26253 27582 26305
rect 27634 26253 27636 26305
rect 27468 26180 27524 26190
rect 27244 26178 27524 26180
rect 27244 26126 27470 26178
rect 27522 26126 27524 26178
rect 27244 26124 27524 26126
rect 27468 26114 27524 26124
rect 27580 26068 27636 26253
rect 27804 26290 27860 27132
rect 27804 26238 27806 26290
rect 27858 26238 27860 26290
rect 27804 26226 27860 26238
rect 27580 26002 27636 26012
rect 28140 26068 28196 27244
rect 28476 27188 28532 27806
rect 28700 27858 28756 28476
rect 29036 27972 29092 29372
rect 29204 27972 29260 27982
rect 29036 27970 29260 27972
rect 29036 27918 29206 27970
rect 29258 27918 29260 27970
rect 29036 27916 29260 27918
rect 29204 27906 29260 27916
rect 28700 27806 28702 27858
rect 28754 27806 28756 27858
rect 28700 27794 28756 27806
rect 28924 27860 28980 27870
rect 28924 27766 28980 27804
rect 28364 27132 28476 27188
rect 28140 26002 28196 26012
rect 28252 26404 28308 26414
rect 28140 25618 28196 25630
rect 28140 25566 28142 25618
rect 28194 25566 28196 25618
rect 27356 25506 27412 25518
rect 27692 25508 27748 25518
rect 27356 25454 27358 25506
rect 27410 25454 27412 25506
rect 26160 25116 26424 25126
rect 26216 25060 26264 25116
rect 26320 25060 26368 25116
rect 26160 25050 26424 25060
rect 26236 24948 26292 24958
rect 25004 24658 25060 24668
rect 25116 24722 25172 24734
rect 25116 24670 25118 24722
rect 25170 24670 25172 24722
rect 25116 24500 25172 24670
rect 24444 24444 25172 24500
rect 25452 24498 25508 24510
rect 25452 24446 25454 24498
rect 25506 24446 25508 24498
rect 23716 23996 23828 24052
rect 24332 24052 24388 24062
rect 23660 23986 23716 23996
rect 24332 23958 24388 23996
rect 25452 24052 25508 24446
rect 25452 23986 25508 23996
rect 26236 24050 26292 24892
rect 27356 24948 27412 25454
rect 27356 24882 27412 24892
rect 27468 25506 27748 25508
rect 27468 25454 27694 25506
rect 27746 25454 27748 25506
rect 28140 25508 28196 25566
rect 27468 25452 27748 25454
rect 27020 24836 27076 24846
rect 26740 24610 26796 24622
rect 26740 24558 26742 24610
rect 26794 24558 26796 24610
rect 26740 24500 26796 24558
rect 26740 24434 26796 24444
rect 26236 23998 26238 24050
rect 26290 23998 26292 24050
rect 26236 23986 26292 23998
rect 23548 23940 23604 23950
rect 23436 23938 23604 23940
rect 23436 23886 23550 23938
rect 23602 23886 23604 23938
rect 23436 23884 23604 23886
rect 23212 22930 23268 22942
rect 23212 22878 23214 22930
rect 23266 22878 23268 22930
rect 23100 22370 23156 22382
rect 23100 22318 23102 22370
rect 23154 22318 23156 22370
rect 23100 22260 23156 22318
rect 23212 22260 23268 22878
rect 23436 22260 23492 23884
rect 23548 23874 23604 23884
rect 26796 23940 26852 23950
rect 26160 23548 26424 23558
rect 26216 23492 26264 23548
rect 26320 23492 26368 23548
rect 26160 23482 26424 23492
rect 26180 23380 26236 23390
rect 25564 23378 26236 23380
rect 25564 23326 26182 23378
rect 26234 23326 26236 23378
rect 25564 23324 26236 23326
rect 25564 23154 25620 23324
rect 26180 23314 26236 23324
rect 26796 23266 26852 23884
rect 27020 23923 27076 24780
rect 27356 24724 27412 24734
rect 27468 24724 27524 25452
rect 27692 25442 27748 25452
rect 28028 25450 28084 25462
rect 28028 25398 28030 25450
rect 28082 25398 28084 25450
rect 28140 25442 28196 25452
rect 28028 25396 28084 25398
rect 28028 25330 28084 25340
rect 28252 24948 28308 26348
rect 28364 25506 28420 27132
rect 28476 27122 28532 27132
rect 28588 26404 28644 26414
rect 28588 26334 28644 26348
rect 28588 26282 28590 26334
rect 28642 26282 28644 26334
rect 29372 26404 29428 26414
rect 28588 26270 28644 26282
rect 28924 26292 28980 26302
rect 29260 26292 29316 26302
rect 28924 26290 29316 26292
rect 28924 26238 28926 26290
rect 28978 26238 29262 26290
rect 29314 26238 29316 26290
rect 28924 26236 29316 26238
rect 28924 26226 28980 26236
rect 28476 26180 28532 26190
rect 28476 26178 28644 26180
rect 28476 26126 28478 26178
rect 28530 26126 28644 26178
rect 28476 26124 28644 26126
rect 28476 26114 28532 26124
rect 28364 25454 28366 25506
rect 28418 25454 28420 25506
rect 28364 25442 28420 25454
rect 27860 24892 28420 24948
rect 27356 24722 27524 24724
rect 27356 24670 27358 24722
rect 27410 24670 27524 24722
rect 27356 24668 27524 24670
rect 27580 24836 27636 24846
rect 27580 24722 27636 24780
rect 27860 24834 27916 24892
rect 27860 24782 27862 24834
rect 27914 24782 27916 24834
rect 27860 24770 27916 24782
rect 27580 24670 27582 24722
rect 27634 24670 27636 24722
rect 27188 24610 27244 24622
rect 27188 24558 27190 24610
rect 27242 24558 27244 24610
rect 27188 24500 27244 24558
rect 27188 24434 27244 24444
rect 27020 23871 27022 23923
rect 27074 23871 27076 23923
rect 27244 23940 27300 23978
rect 27356 23940 27412 24668
rect 27580 24658 27636 24670
rect 28252 24722 28308 24734
rect 28252 24670 28254 24722
rect 28306 24670 28308 24722
rect 27300 23884 27412 23940
rect 27692 24500 27748 24510
rect 27692 23938 27748 24444
rect 28252 24500 28308 24670
rect 28252 24434 28308 24444
rect 27692 23886 27694 23938
rect 27746 23886 27748 23938
rect 28364 23938 28420 24892
rect 28588 24778 28644 26124
rect 28588 24726 28590 24778
rect 28642 24726 28644 24778
rect 28588 24714 28644 24726
rect 28924 26068 28980 26078
rect 28924 24722 28980 26012
rect 29260 25396 29316 26236
rect 29372 26290 29428 26348
rect 29372 26238 29374 26290
rect 29426 26238 29428 26290
rect 29372 26226 29428 26238
rect 29260 25302 29316 25340
rect 28924 24670 28926 24722
rect 28978 24670 28980 24722
rect 28924 24658 28980 24670
rect 29036 24890 29092 24902
rect 29036 24838 29038 24890
rect 29090 24838 29092 24890
rect 29036 24724 29092 24838
rect 29372 24724 29428 24734
rect 29036 24722 29428 24724
rect 29036 24670 29374 24722
rect 29426 24670 29428 24722
rect 29036 24668 29428 24670
rect 29372 24658 29428 24668
rect 27244 23874 27300 23884
rect 27692 23874 27748 23886
rect 27972 23882 28028 23894
rect 27020 23859 27076 23871
rect 27972 23830 27974 23882
rect 28026 23830 28028 23882
rect 28364 23886 28366 23938
rect 28418 23886 28420 23938
rect 28364 23874 28420 23886
rect 28476 23940 28532 23950
rect 27972 23828 28028 23830
rect 27244 23770 27300 23782
rect 27244 23718 27246 23770
rect 27298 23718 27300 23770
rect 27244 23716 27300 23718
rect 27804 23772 28028 23828
rect 27804 23716 27860 23772
rect 27244 23660 27860 23716
rect 28476 23770 28532 23884
rect 29036 23940 29092 23950
rect 29036 23846 29092 23884
rect 28476 23718 28478 23770
rect 28530 23718 28532 23770
rect 28476 23706 28532 23718
rect 29372 23716 29428 23726
rect 28700 23714 29428 23716
rect 28700 23662 29374 23714
rect 29426 23662 29428 23714
rect 28700 23660 29428 23662
rect 26796 23214 26798 23266
rect 26850 23214 26852 23266
rect 26796 23202 26852 23214
rect 25564 23102 25566 23154
rect 25618 23102 25620 23154
rect 25284 22930 25340 22942
rect 25284 22878 25286 22930
rect 25338 22878 25340 22930
rect 23100 22204 23492 22260
rect 23156 22036 23212 22046
rect 22988 21644 23100 21700
rect 22932 21476 22988 21486
rect 23044 21476 23100 21644
rect 23156 21642 23212 21980
rect 23156 21590 23158 21642
rect 23210 21590 23212 21642
rect 23324 21924 23380 21934
rect 23324 21698 23380 21868
rect 23324 21646 23326 21698
rect 23378 21646 23380 21698
rect 23324 21634 23380 21646
rect 23156 21578 23212 21590
rect 23044 21420 23380 21476
rect 22932 21382 22988 21420
rect 22002 21130 22266 21140
rect 22372 21084 22596 21140
rect 22988 21252 23044 21262
rect 22372 21028 22428 21084
rect 22204 20972 22428 21028
rect 22876 21028 22932 21038
rect 21756 20750 21758 20802
rect 21810 20750 21812 20802
rect 22092 20804 22148 20842
rect 21756 20692 21812 20750
rect 21756 20626 21812 20636
rect 21924 20746 21980 20758
rect 21924 20694 21926 20746
rect 21978 20694 21980 20746
rect 22092 20738 22148 20748
rect 21924 20188 21980 20694
rect 22092 20580 22148 20590
rect 21924 20132 22036 20188
rect 21868 20018 21924 20030
rect 21868 19966 21870 20018
rect 21922 19966 21924 20018
rect 21532 19908 21588 19918
rect 21532 19814 21588 19852
rect 19628 17602 19684 17614
rect 19908 17610 19964 17622
rect 19740 17556 19796 17566
rect 19740 17462 19796 17500
rect 19908 17558 19910 17610
rect 19962 17558 19964 17610
rect 20076 17614 20078 17666
rect 20130 17614 20132 17666
rect 20076 17602 20132 17614
rect 20188 17892 20244 17902
rect 19908 17220 19964 17558
rect 19852 17164 19908 17220
rect 19852 17154 19964 17164
rect 20076 17332 20132 17342
rect 19460 16884 19516 16894
rect 19068 16882 19516 16884
rect 19068 16830 19462 16882
rect 19514 16830 19516 16882
rect 19068 16828 19516 16830
rect 19068 16770 19124 16828
rect 19460 16818 19516 16828
rect 19852 16882 19908 17154
rect 19852 16830 19854 16882
rect 19906 16830 19908 16882
rect 19852 16818 19908 16830
rect 19068 16718 19070 16770
rect 19122 16718 19124 16770
rect 19068 16706 19124 16718
rect 19628 16772 19684 16782
rect 19628 16770 19796 16772
rect 19628 16718 19630 16770
rect 19682 16718 19796 16770
rect 19628 16716 19796 16718
rect 19628 16706 19684 16716
rect 19292 16660 19348 16670
rect 19292 16210 19348 16604
rect 19292 16158 19294 16210
rect 19346 16158 19348 16210
rect 19292 16146 19348 16158
rect 19516 16100 19572 16110
rect 18956 16068 19180 16100
rect 18956 16044 19126 16068
rect 19124 16016 19126 16044
rect 19178 16016 19180 16068
rect 19124 16004 19180 16016
rect 19516 16006 19572 16044
rect 18340 15482 18396 15494
rect 18340 15430 18342 15482
rect 18394 15430 18396 15482
rect 18340 15428 18396 15430
rect 18340 15362 18396 15372
rect 18732 15484 18844 15540
rect 18508 15314 18564 15326
rect 18508 15262 18510 15314
rect 18562 15262 18564 15314
rect 18172 15148 18452 15204
rect 17836 14532 17892 14542
rect 17836 14530 18340 14532
rect 17836 14478 17838 14530
rect 17890 14478 18340 14530
rect 17836 14476 18340 14478
rect 17836 14466 17892 14476
rect 17724 14242 17780 14252
rect 18172 14308 18228 14318
rect 18172 14214 18228 14252
rect 17844 14140 18108 14150
rect 17900 14084 17948 14140
rect 18004 14084 18052 14140
rect 17844 14074 18108 14084
rect 17836 13860 17892 13870
rect 17836 13766 17892 13804
rect 17724 13746 17780 13758
rect 17724 13694 17726 13746
rect 17778 13694 17780 13746
rect 17724 13524 17780 13694
rect 18004 13748 18060 13758
rect 18004 13654 18060 13692
rect 18172 13748 18228 13758
rect 18284 13748 18340 14476
rect 18172 13746 18340 13748
rect 18172 13694 18174 13746
rect 18226 13694 18340 13746
rect 18172 13692 18340 13694
rect 18172 13682 18228 13692
rect 17724 13458 17780 13468
rect 17612 13132 18116 13188
rect 17500 13074 17556 13086
rect 17500 13022 17502 13074
rect 17554 13022 17556 13074
rect 17500 12964 17556 13022
rect 17500 12898 17556 12908
rect 17500 12346 17556 12358
rect 17500 12294 17502 12346
rect 17554 12294 17556 12346
rect 17388 12180 17444 12190
rect 17388 12086 17444 12124
rect 17276 9202 17332 9212
rect 17500 8596 17556 12294
rect 17724 12234 17780 13132
rect 18060 12962 18116 13132
rect 17892 12906 17948 12918
rect 17892 12854 17894 12906
rect 17946 12854 17948 12906
rect 18060 12910 18062 12962
rect 18114 12910 18116 12962
rect 18060 12898 18116 12910
rect 18172 12962 18228 12974
rect 18172 12910 18174 12962
rect 18226 12910 18228 12962
rect 17892 12852 17948 12854
rect 17892 12786 17948 12796
rect 18172 12852 18228 12910
rect 18172 12786 18228 12796
rect 18284 12740 18340 13692
rect 18284 12674 18340 12684
rect 17844 12572 18108 12582
rect 17900 12516 17948 12572
rect 18004 12516 18052 12572
rect 17844 12506 18108 12516
rect 17724 12182 17726 12234
rect 17778 12182 17780 12234
rect 17724 11620 17780 12182
rect 18060 12180 18116 12190
rect 17948 12124 18060 12180
rect 17724 11564 17892 11620
rect 17668 11396 17724 11406
rect 17668 11302 17724 11340
rect 17836 11172 17892 11564
rect 17948 11394 18004 12124
rect 18060 12086 18116 12124
rect 17948 11342 17950 11394
rect 18002 11342 18004 11394
rect 17948 11330 18004 11342
rect 18060 11394 18116 11406
rect 18060 11342 18062 11394
rect 18114 11342 18116 11394
rect 18060 11172 18116 11342
rect 17836 11116 18116 11172
rect 17844 11004 18108 11014
rect 17900 10948 17948 11004
rect 18004 10948 18052 11004
rect 17844 10938 18108 10948
rect 18396 10164 18452 15148
rect 18508 13748 18564 15262
rect 18508 13682 18564 13692
rect 18564 13524 18620 13534
rect 18732 13524 18788 15484
rect 18844 15474 18900 15484
rect 19068 15314 19124 15326
rect 19068 15262 19070 15314
rect 19122 15262 19124 15314
rect 19068 15204 19124 15262
rect 19740 15316 19796 16716
rect 19852 16324 19908 16334
rect 20076 16324 20132 17276
rect 20188 16938 20244 17836
rect 20636 17892 20692 17902
rect 20636 17798 20692 17836
rect 20300 17780 20356 17790
rect 20300 17666 20356 17724
rect 20300 17614 20302 17666
rect 20354 17614 20356 17666
rect 20300 17602 20356 17614
rect 20188 16886 20190 16938
rect 20242 16886 20244 16938
rect 20188 16874 20244 16886
rect 20748 16884 20804 18396
rect 20860 19404 21140 19460
rect 20860 18004 20916 19404
rect 21868 19348 21924 19966
rect 21980 19908 22036 20132
rect 22092 20018 22148 20524
rect 22092 19966 22094 20018
rect 22146 19966 22148 20018
rect 22092 19954 22148 19966
rect 21980 19842 22036 19852
rect 22204 19796 22260 20972
rect 22316 20804 22372 20814
rect 22316 20142 22372 20748
rect 22428 20802 22484 20814
rect 22428 20750 22430 20802
rect 22482 20750 22484 20802
rect 22428 20580 22484 20750
rect 22596 20804 22652 20814
rect 22596 20710 22652 20748
rect 22876 20802 22932 20972
rect 22876 20750 22878 20802
rect 22930 20750 22932 20802
rect 22764 20692 22820 20702
rect 22764 20598 22820 20636
rect 22428 20514 22484 20524
rect 22540 20468 22596 20478
rect 22316 20130 22428 20142
rect 22316 20078 22374 20130
rect 22426 20078 22428 20130
rect 22316 20076 22428 20078
rect 22372 20066 22428 20076
rect 22540 20020 22596 20412
rect 22876 20188 22932 20750
rect 22540 19954 22596 19964
rect 22652 20132 22932 20188
rect 22988 20244 23044 21196
rect 22988 20178 23044 20188
rect 23156 20690 23212 20702
rect 23156 20638 23158 20690
rect 23210 20638 23212 20690
rect 23156 20188 23212 20638
rect 23324 20468 23380 21420
rect 23436 20802 23492 22204
rect 23884 22370 23940 22382
rect 23884 22318 23886 22370
rect 23938 22318 23940 22370
rect 23884 21924 23940 22318
rect 25284 22372 25340 22878
rect 25284 22306 25340 22316
rect 23884 21858 23940 21868
rect 23548 21812 23604 21822
rect 23548 21586 23604 21756
rect 23548 21534 23550 21586
rect 23602 21534 23604 21586
rect 23548 21522 23604 21534
rect 23772 21614 23828 21626
rect 23772 21562 23774 21614
rect 23826 21562 23828 21614
rect 23772 21476 23828 21562
rect 23772 21410 23828 21420
rect 25564 21476 25620 23102
rect 25788 23154 25844 23166
rect 25788 23102 25790 23154
rect 25842 23102 25844 23154
rect 25788 22258 25844 23102
rect 28700 23154 28756 23660
rect 29372 23650 29428 23660
rect 28700 23102 28702 23154
rect 28754 23102 28756 23154
rect 28700 23090 28756 23102
rect 29484 23380 29540 30156
rect 34476 29820 34740 29830
rect 34532 29764 34580 29820
rect 34636 29764 34684 29820
rect 34476 29754 34740 29764
rect 30318 29036 30582 29046
rect 30374 28980 30422 29036
rect 30478 28980 30526 29036
rect 30318 28970 30582 28980
rect 34476 28252 34740 28262
rect 34532 28196 34580 28252
rect 34636 28196 34684 28252
rect 34476 28186 34740 28196
rect 30318 27468 30582 27478
rect 30374 27412 30422 27468
rect 30478 27412 30526 27468
rect 30318 27402 30582 27412
rect 34476 26684 34740 26694
rect 34532 26628 34580 26684
rect 34636 26628 34684 26684
rect 34476 26618 34740 26628
rect 29652 26068 29708 26078
rect 29652 25974 29708 26012
rect 30318 25900 30582 25910
rect 30374 25844 30422 25900
rect 30478 25844 30526 25900
rect 30318 25834 30582 25844
rect 29708 25508 29764 25518
rect 29708 24946 29764 25452
rect 31164 25508 31220 25518
rect 31164 25414 31220 25452
rect 31948 25508 32004 25518
rect 32340 25508 32396 25518
rect 31948 25506 32396 25508
rect 31948 25454 31950 25506
rect 32002 25454 32342 25506
rect 32394 25454 32396 25506
rect 31948 25452 32396 25454
rect 31948 25442 32004 25452
rect 29708 24894 29710 24946
rect 29762 24894 29764 24946
rect 29708 24882 29764 24894
rect 30318 24332 30582 24342
rect 30374 24276 30422 24332
rect 30478 24276 30526 24332
rect 30318 24266 30582 24276
rect 29876 23380 29932 23390
rect 29484 23378 29932 23380
rect 29484 23326 29878 23378
rect 29930 23326 29932 23378
rect 29484 23324 29932 23326
rect 29484 23154 29540 23324
rect 29876 23314 29932 23324
rect 29484 23102 29486 23154
rect 29538 23102 29540 23154
rect 25788 22206 25790 22258
rect 25842 22206 25844 22258
rect 25788 21812 25844 22206
rect 29484 22342 29540 23102
rect 30940 23154 30996 23166
rect 30940 23102 30942 23154
rect 30994 23102 30996 23154
rect 30604 22932 30660 22942
rect 30604 22930 30772 22932
rect 30604 22878 30606 22930
rect 30658 22878 30772 22930
rect 30604 22876 30772 22878
rect 30604 22866 30660 22876
rect 30318 22764 30582 22774
rect 30374 22708 30422 22764
rect 30478 22708 30526 22764
rect 30318 22698 30582 22708
rect 29484 22290 29486 22342
rect 29538 22290 29540 22342
rect 29484 22260 29540 22290
rect 29484 22204 29764 22260
rect 26160 21980 26424 21990
rect 26216 21924 26264 21980
rect 26320 21924 26368 21980
rect 26160 21914 26424 21924
rect 25788 21746 25844 21756
rect 26460 21812 26516 21822
rect 25564 21410 25620 21420
rect 23436 20750 23438 20802
rect 23490 20750 23492 20802
rect 23436 20692 23492 20750
rect 24220 20802 24276 20814
rect 24220 20750 24222 20802
rect 24274 20750 24276 20802
rect 23436 20636 24052 20692
rect 23324 20402 23380 20412
rect 23884 20356 23940 20366
rect 23884 20242 23940 20300
rect 23884 20190 23886 20242
rect 23938 20190 23940 20242
rect 23156 20132 23604 20188
rect 23884 20178 23940 20190
rect 23996 20188 24052 20636
rect 24220 20356 24276 20750
rect 26124 20804 26180 20814
rect 26124 20710 26180 20748
rect 26460 20802 26516 21756
rect 29372 21586 29428 21598
rect 29372 21534 29374 21586
rect 29426 21534 29428 21586
rect 29092 21362 29148 21374
rect 29092 21310 29094 21362
rect 29146 21310 29148 21362
rect 29092 21028 29148 21310
rect 29092 20962 29148 20972
rect 26460 20750 26462 20802
rect 26514 20750 26516 20802
rect 26460 20738 26516 20750
rect 26684 20804 26740 20814
rect 26684 20710 26740 20748
rect 27748 20804 27804 20814
rect 26964 20692 27020 20702
rect 26964 20690 27300 20692
rect 26964 20638 26966 20690
rect 27018 20638 27300 20690
rect 26964 20636 27300 20638
rect 26964 20626 27020 20636
rect 26160 20412 26424 20422
rect 26216 20356 26264 20412
rect 26320 20356 26368 20412
rect 26160 20346 26424 20356
rect 24220 20290 24276 20300
rect 23996 20132 24724 20188
rect 22204 19740 22596 19796
rect 22002 19628 22266 19638
rect 22058 19572 22106 19628
rect 22162 19572 22210 19628
rect 22002 19562 22266 19572
rect 21980 19348 22036 19358
rect 21532 19346 22036 19348
rect 21532 19294 21982 19346
rect 22034 19294 22036 19346
rect 21532 19292 22036 19294
rect 20972 19236 21028 19246
rect 20972 18450 21028 19180
rect 21364 19236 21420 19246
rect 21364 19066 21420 19180
rect 21532 19234 21588 19292
rect 21980 19282 22036 19292
rect 21532 19182 21534 19234
rect 21586 19182 21588 19234
rect 21532 19170 21588 19182
rect 22204 19236 22260 19246
rect 21364 19014 21366 19066
rect 21418 19014 21420 19066
rect 21364 19002 21420 19014
rect 21230 18487 21286 18499
rect 20972 18398 20974 18450
rect 21026 18398 21028 18450
rect 20972 18386 21028 18398
rect 21084 18450 21140 18462
rect 21084 18398 21086 18450
rect 21138 18398 21140 18450
rect 20860 17612 20916 17948
rect 21084 17780 21140 18398
rect 21230 18435 21232 18487
rect 21284 18435 21286 18487
rect 21230 18004 21286 18435
rect 22036 18450 22092 18462
rect 22036 18398 22038 18450
rect 22090 18398 22092 18450
rect 21644 18340 21700 18350
rect 22036 18340 22092 18398
rect 22204 18450 22260 19180
rect 22204 18398 22206 18450
rect 22258 18398 22260 18450
rect 22204 18386 22260 18398
rect 22428 18452 22484 18462
rect 22428 18358 22484 18396
rect 21644 18338 22092 18340
rect 21644 18286 21646 18338
rect 21698 18286 22092 18338
rect 21644 18284 22092 18286
rect 21644 18274 21700 18284
rect 21084 17714 21140 17724
rect 21196 17948 21286 18004
rect 22002 18060 22266 18070
rect 22058 18004 22106 18060
rect 22162 18004 22210 18060
rect 22002 17994 22266 18004
rect 20860 17556 21140 17612
rect 20972 16920 21028 16932
rect 20972 16884 20974 16920
rect 20804 16868 20974 16884
rect 21026 16868 21028 16920
rect 20804 16828 21028 16868
rect 20748 16818 20804 16828
rect 19852 16322 20132 16324
rect 19852 16270 19854 16322
rect 19906 16270 20132 16322
rect 19852 16268 20132 16270
rect 19852 16258 19908 16268
rect 19852 15316 19908 15326
rect 19740 15314 19908 15316
rect 19740 15262 19854 15314
rect 19906 15262 19908 15314
rect 19740 15260 19908 15262
rect 19852 15250 19908 15260
rect 19068 15138 19124 15148
rect 18844 13916 19124 13972
rect 18844 13746 18900 13916
rect 18844 13694 18846 13746
rect 18898 13694 18900 13746
rect 18844 13682 18900 13694
rect 18956 13746 19012 13758
rect 18956 13694 18958 13746
rect 19010 13694 19012 13746
rect 18956 13636 19012 13694
rect 18956 13570 19012 13580
rect 18732 13468 18900 13524
rect 18564 13430 18620 13468
rect 18508 12964 18564 12974
rect 18844 12962 18900 13468
rect 18508 12870 18564 12908
rect 18676 12906 18732 12918
rect 18676 12854 18678 12906
rect 18730 12854 18732 12906
rect 18844 12910 18846 12962
rect 18898 12910 18900 12962
rect 18844 12898 18900 12910
rect 18956 13076 19012 13086
rect 18956 12962 19012 13020
rect 18956 12910 18958 12962
rect 19010 12910 19012 12962
rect 18956 12898 19012 12910
rect 18676 12404 18732 12854
rect 18676 12338 18732 12348
rect 18844 12740 18900 12750
rect 18620 12178 18676 12190
rect 18620 12126 18622 12178
rect 18674 12126 18676 12178
rect 18620 12068 18676 12126
rect 18620 12002 18676 12012
rect 18732 12180 18788 12190
rect 18732 12010 18788 12124
rect 18732 11958 18734 12010
rect 18786 11958 18788 12010
rect 18732 11946 18788 11958
rect 18732 11844 18788 11854
rect 18732 11618 18788 11788
rect 18732 11566 18734 11618
rect 18786 11566 18788 11618
rect 18732 11554 18788 11566
rect 18844 11620 18900 12684
rect 18956 12292 19012 12302
rect 18956 12178 19012 12236
rect 18956 12126 18958 12178
rect 19010 12126 19012 12178
rect 18956 11844 19012 12126
rect 18956 11778 19012 11788
rect 18844 11564 19012 11620
rect 18060 10108 18452 10164
rect 17836 9940 17892 9950
rect 17836 9846 17892 9884
rect 18060 9604 18116 10108
rect 18060 9548 18340 9604
rect 17844 9436 18108 9446
rect 17900 9380 17948 9436
rect 18004 9380 18052 9436
rect 17844 9370 18108 9380
rect 16268 8372 16884 8428
rect 17164 8540 17556 8596
rect 18172 9268 18228 9278
rect 16268 8258 16324 8372
rect 16268 8206 16270 8258
rect 16322 8206 16324 8258
rect 16044 7422 16046 7474
rect 16098 7422 16100 7474
rect 16044 7410 16100 7422
rect 16156 7476 16212 7486
rect 15708 6916 15764 6926
rect 15596 6914 15764 6916
rect 15596 6862 15710 6914
rect 15762 6862 15764 6914
rect 15596 6860 15764 6862
rect 15708 6850 15764 6860
rect 15484 6402 15540 6412
rect 15932 6692 15988 6702
rect 15260 6188 15652 6244
rect 15260 5460 15316 6188
rect 15596 6130 15652 6188
rect 15596 6078 15598 6130
rect 15650 6078 15652 6130
rect 15596 6066 15652 6078
rect 15932 5906 15988 6636
rect 16156 6580 16212 7420
rect 16268 6804 16324 8206
rect 17052 8260 17108 8270
rect 17052 8166 17108 8204
rect 16268 6738 16324 6748
rect 16604 6692 16660 6702
rect 17052 6692 17108 6702
rect 16604 6690 17108 6692
rect 16604 6638 16606 6690
rect 16658 6638 17054 6690
rect 17106 6638 17108 6690
rect 16604 6636 17108 6638
rect 16604 6626 16660 6636
rect 16268 6580 16324 6590
rect 16156 6578 16324 6580
rect 16156 6526 16270 6578
rect 16322 6526 16324 6578
rect 16156 6524 16324 6526
rect 16268 6514 16324 6524
rect 16884 6468 16940 6478
rect 16884 6374 16940 6412
rect 16436 6132 16492 6142
rect 16436 6018 16492 6076
rect 16436 5966 16438 6018
rect 16490 5966 16492 6018
rect 16436 5954 16492 5966
rect 17052 6020 17108 6636
rect 17052 5954 17108 5964
rect 15932 5854 15934 5906
rect 15986 5854 15988 5906
rect 15932 5842 15988 5854
rect 16716 5908 16772 5918
rect 16716 5814 16772 5852
rect 16828 5906 16884 5918
rect 16828 5854 16830 5906
rect 16882 5854 16884 5906
rect 15260 5394 15316 5404
rect 16492 5124 16548 5134
rect 16492 5030 16548 5068
rect 16716 4452 16772 4462
rect 16828 4452 16884 5854
rect 17164 5908 17220 8540
rect 17844 7868 18108 7878
rect 17900 7812 17948 7868
rect 18004 7812 18052 7868
rect 17844 7802 18108 7812
rect 18172 7700 18228 9212
rect 18060 7644 18228 7700
rect 17388 6858 17444 6870
rect 17388 6806 17390 6858
rect 17442 6806 17444 6858
rect 17276 6690 17332 6702
rect 17276 6638 17278 6690
rect 17330 6638 17332 6690
rect 17276 6132 17332 6638
rect 17388 6692 17444 6806
rect 18060 6702 18116 7644
rect 17388 6626 17444 6636
rect 17612 6690 17668 6702
rect 17612 6638 17614 6690
rect 17666 6638 17668 6690
rect 17612 6468 17668 6638
rect 18004 6692 18116 6702
rect 18060 6636 18116 6692
rect 18004 6598 18060 6636
rect 18172 6578 18228 6590
rect 18172 6526 18174 6578
rect 18226 6526 18228 6578
rect 18172 6468 18228 6526
rect 17612 6412 18228 6468
rect 17844 6300 18108 6310
rect 17900 6244 17948 6300
rect 18004 6244 18052 6300
rect 17844 6234 18108 6244
rect 17276 6066 17332 6076
rect 18060 6020 18116 6030
rect 17276 5908 17332 5918
rect 17220 5906 17332 5908
rect 17220 5854 17278 5906
rect 17330 5854 17332 5906
rect 17220 5852 17332 5854
rect 17164 5814 17220 5852
rect 17276 5842 17332 5852
rect 17836 5908 17892 5918
rect 17612 5684 17668 5694
rect 17836 5684 17892 5852
rect 17612 5682 17892 5684
rect 17612 5630 17614 5682
rect 17666 5630 17892 5682
rect 18060 5738 18116 5964
rect 18060 5686 18062 5738
rect 18114 5686 18116 5738
rect 18172 5906 18228 5918
rect 18172 5854 18174 5906
rect 18226 5854 18228 5906
rect 18172 5796 18228 5854
rect 18172 5730 18228 5740
rect 18060 5674 18116 5686
rect 17612 5628 17892 5630
rect 17612 5618 17668 5628
rect 17836 5122 17892 5628
rect 17836 5070 17838 5122
rect 17890 5070 17892 5122
rect 17836 5058 17892 5070
rect 18060 5236 18116 5246
rect 18060 5066 18116 5180
rect 18060 5014 18062 5066
rect 18114 5014 18116 5066
rect 18060 4900 18116 5014
rect 17724 4844 18116 4900
rect 18172 5234 18228 5246
rect 18172 5182 18174 5234
rect 18226 5182 18228 5234
rect 17724 4564 17780 4844
rect 17844 4732 18108 4742
rect 17900 4676 17948 4732
rect 18004 4676 18052 4732
rect 17844 4666 18108 4676
rect 18172 4564 18228 5182
rect 17724 4508 18116 4564
rect 16716 4450 16884 4452
rect 16716 4398 16718 4450
rect 16770 4398 16884 4450
rect 16716 4396 16884 4398
rect 16716 4386 16772 4396
rect 14812 4340 14868 4350
rect 14812 4246 14868 4284
rect 16828 4340 16884 4396
rect 16828 4274 16884 4284
rect 17836 4340 17892 4350
rect 18060 4340 18116 4508
rect 18172 4498 18228 4508
rect 18172 4340 18228 4350
rect 18060 4338 18228 4340
rect 18060 4286 18174 4338
rect 18226 4286 18228 4338
rect 18060 4284 18228 4286
rect 17836 4246 17892 4284
rect 18172 4274 18228 4284
rect 18284 4228 18340 9548
rect 18956 8370 19012 11564
rect 19068 11396 19124 13916
rect 21084 13746 21140 17556
rect 21196 17108 21252 17948
rect 22092 17780 22148 17790
rect 21756 17778 22148 17780
rect 21756 17726 22094 17778
rect 22146 17726 22148 17778
rect 21756 17724 22148 17726
rect 21196 17042 21252 17052
rect 21308 17220 21364 17230
rect 21308 16996 21364 17164
rect 21756 17052 21812 17724
rect 22092 17714 22148 17724
rect 22540 17622 22596 19740
rect 22484 17610 22596 17622
rect 22484 17558 22486 17610
rect 22538 17558 22596 17610
rect 22652 17892 22708 20132
rect 22764 20020 22820 20030
rect 22764 18676 22820 19964
rect 23548 20018 23604 20132
rect 23548 19966 23550 20018
rect 23602 19966 23604 20018
rect 23548 19954 23604 19966
rect 23884 19236 23940 19246
rect 23884 19142 23940 19180
rect 24668 19236 24724 20132
rect 26908 20018 26964 20030
rect 26908 19966 26910 20018
rect 26962 19966 26964 20018
rect 26572 19796 26628 19806
rect 25900 19794 26628 19796
rect 25900 19742 26574 19794
rect 26626 19742 26628 19794
rect 25900 19740 26628 19742
rect 25900 19346 25956 19740
rect 26572 19730 26628 19740
rect 26908 19684 26964 19966
rect 27020 20020 27076 20030
rect 27020 19926 27076 19964
rect 26908 19628 27188 19684
rect 25900 19294 25902 19346
rect 25954 19294 25956 19346
rect 25900 19282 25956 19294
rect 25116 19236 25172 19246
rect 24668 19234 25172 19236
rect 24668 19182 24670 19234
rect 24722 19182 25118 19234
rect 25170 19182 25172 19234
rect 24668 19180 25172 19182
rect 24668 19170 24724 19180
rect 25116 19170 25172 19180
rect 26160 18844 26424 18854
rect 26216 18788 26264 18844
rect 26320 18788 26368 18844
rect 26160 18778 26424 18788
rect 22764 18620 22932 18676
rect 22764 18488 22820 18500
rect 22764 18436 22766 18488
rect 22818 18436 22820 18488
rect 22764 18004 22820 18436
rect 22764 17938 22820 17948
rect 22652 17666 22708 17836
rect 22652 17614 22654 17666
rect 22706 17614 22708 17666
rect 22652 17602 22708 17614
rect 22764 17666 22820 17678
rect 22764 17614 22766 17666
rect 22818 17614 22820 17666
rect 22484 17556 22596 17558
rect 22764 17556 22820 17614
rect 22484 17332 22540 17556
rect 22764 17490 22820 17500
rect 22484 17266 22540 17276
rect 22876 17052 22932 18620
rect 27132 18618 27188 19628
rect 27132 18566 27134 18618
rect 27186 18566 27188 18618
rect 27132 18554 27188 18566
rect 27132 18450 27188 18462
rect 27132 18398 27134 18450
rect 27186 18398 27188 18450
rect 27132 18340 27188 18398
rect 27132 18274 27188 18284
rect 21308 16882 21364 16940
rect 21308 16830 21310 16882
rect 21362 16830 21364 16882
rect 21700 16996 21812 17052
rect 22652 16996 22932 17052
rect 22988 18004 23044 18014
rect 22988 16996 23044 17948
rect 23324 17666 23380 17678
rect 23324 17614 23326 17666
rect 23378 17614 23380 17666
rect 23156 17556 23212 17566
rect 23156 17498 23212 17500
rect 23156 17446 23158 17498
rect 23210 17446 23212 17498
rect 23156 17434 23212 17446
rect 23100 16996 23156 17006
rect 21700 16938 21756 16996
rect 21700 16886 21702 16938
rect 21754 16886 21756 16938
rect 21700 16874 21756 16886
rect 21980 16884 22036 16922
rect 21308 16818 21364 16830
rect 21812 16828 21980 16884
rect 21532 16770 21588 16782
rect 21812 16772 21868 16828
rect 21980 16818 22036 16828
rect 21532 16718 21534 16770
rect 21586 16718 21588 16770
rect 21532 16324 21588 16718
rect 21532 16258 21588 16268
rect 21756 16716 21868 16772
rect 21532 16098 21588 16110
rect 21532 16046 21534 16098
rect 21586 16046 21588 16098
rect 21532 15204 21588 16046
rect 21756 15426 21812 16716
rect 22002 16492 22266 16502
rect 22058 16436 22106 16492
rect 22162 16436 22210 16492
rect 22652 16436 22708 16996
rect 22988 16994 23156 16996
rect 22988 16942 23102 16994
rect 23154 16942 23156 16994
rect 22988 16940 23156 16942
rect 23100 16930 23156 16940
rect 22856 16882 22912 16894
rect 22856 16830 22858 16882
rect 22910 16830 22912 16882
rect 22856 16772 22912 16830
rect 22856 16706 22912 16716
rect 23324 16772 23380 17614
rect 25452 17668 25508 17678
rect 23604 17050 23660 17062
rect 23604 16998 23606 17050
rect 23658 16998 23660 17050
rect 23604 16996 23660 16998
rect 23604 16930 23660 16940
rect 23436 16884 23492 16894
rect 23436 16790 23492 16828
rect 23324 16706 23380 16716
rect 24220 16772 24276 16782
rect 22002 16426 22266 16436
rect 22540 16380 22708 16436
rect 22316 16324 22372 16334
rect 22316 16210 22372 16268
rect 22316 16158 22318 16210
rect 22370 16158 22372 16210
rect 22316 16146 22372 16158
rect 21756 15374 21758 15426
rect 21810 15374 21812 15426
rect 21756 15362 21812 15374
rect 21532 15138 21588 15148
rect 22372 15204 22428 15214
rect 22372 15110 22428 15148
rect 22002 14924 22266 14934
rect 22058 14868 22106 14924
rect 22162 14868 22210 14924
rect 22002 14858 22266 14868
rect 21084 13694 21086 13746
rect 21138 13694 21140 13746
rect 21084 13682 21140 13694
rect 21308 13746 21364 13758
rect 21308 13694 21310 13746
rect 21362 13694 21364 13746
rect 21308 13188 21364 13694
rect 21588 13748 21644 13758
rect 21868 13748 21924 13758
rect 21588 13746 21924 13748
rect 21588 13694 21590 13746
rect 21642 13694 21870 13746
rect 21922 13694 21924 13746
rect 21588 13692 21924 13694
rect 21588 13682 21644 13692
rect 21868 13682 21924 13692
rect 22204 13524 22260 13534
rect 22204 13522 22484 13524
rect 22204 13470 22206 13522
rect 22258 13470 22484 13522
rect 22204 13468 22484 13470
rect 22204 13458 22260 13468
rect 22002 13356 22266 13366
rect 22058 13300 22106 13356
rect 22162 13300 22210 13356
rect 22002 13290 22266 13300
rect 22428 13188 22484 13468
rect 21308 13122 21364 13132
rect 22204 13132 22484 13188
rect 19516 12962 19572 12974
rect 19516 12910 19518 12962
rect 19570 12910 19572 12962
rect 19236 12852 19292 12862
rect 19236 12850 19460 12852
rect 19236 12798 19238 12850
rect 19290 12798 19460 12850
rect 19236 12796 19460 12798
rect 19236 12786 19292 12796
rect 19404 11620 19460 12796
rect 19516 12292 19572 12910
rect 20188 12964 20244 12974
rect 19684 12852 19740 12862
rect 19684 12794 19740 12796
rect 19684 12742 19686 12794
rect 19738 12742 19740 12794
rect 19684 12730 19740 12742
rect 19516 12226 19572 12236
rect 19964 12066 20020 12078
rect 19964 12014 19966 12066
rect 20018 12014 20020 12066
rect 19964 11956 20020 12014
rect 20188 11956 20244 12908
rect 21532 12964 21588 12974
rect 21532 12870 21588 12908
rect 22204 12628 22260 13132
rect 22408 12964 22464 12974
rect 22408 12870 22464 12908
rect 21868 12572 22260 12628
rect 21868 12178 21924 12572
rect 21868 12126 21870 12178
rect 21922 12126 21924 12178
rect 21868 12114 21924 12126
rect 19964 11900 20244 11956
rect 19404 11554 19460 11564
rect 19068 11394 19796 11396
rect 19068 11342 19070 11394
rect 19122 11342 19796 11394
rect 19068 11340 19796 11342
rect 19068 11330 19124 11340
rect 19740 9938 19796 11340
rect 19740 9886 19742 9938
rect 19794 9886 19796 9938
rect 19740 9874 19796 9886
rect 18956 8318 18958 8370
rect 19010 8318 19012 8370
rect 18956 8306 19012 8318
rect 19516 9042 19572 9054
rect 19516 8990 19518 9042
rect 19570 8990 19572 9042
rect 19516 8484 19572 8990
rect 19404 7474 19460 7486
rect 19404 7422 19406 7474
rect 19458 7422 19460 7474
rect 19404 7364 19460 7422
rect 19516 7364 19572 8428
rect 20188 7700 20244 11900
rect 22002 11788 22266 11798
rect 22058 11732 22106 11788
rect 22162 11732 22210 11788
rect 22002 11722 22266 11732
rect 22428 11396 22484 11406
rect 21868 11394 22484 11396
rect 21868 11342 22430 11394
rect 22482 11342 22484 11394
rect 21868 11340 22484 11342
rect 21308 10610 21364 10622
rect 21308 10558 21310 10610
rect 21362 10558 21364 10610
rect 20972 10388 21028 10398
rect 20300 10386 21028 10388
rect 20300 10334 20974 10386
rect 21026 10334 21028 10386
rect 20300 10332 21028 10334
rect 20300 9042 20356 10332
rect 20972 10322 21028 10332
rect 21308 10052 21364 10558
rect 21308 9986 21364 9996
rect 21868 9940 21924 11340
rect 22428 11330 22484 11340
rect 22036 11170 22092 11182
rect 22036 11118 22038 11170
rect 22090 11118 22092 11170
rect 22036 10780 22092 11118
rect 22540 10948 22596 16380
rect 24220 16210 24276 16716
rect 24220 16158 24222 16210
rect 24274 16158 24276 16210
rect 24220 16146 24276 16158
rect 25340 16770 25396 16782
rect 25340 16718 25342 16770
rect 25394 16718 25396 16770
rect 25340 16100 25396 16718
rect 25340 16034 25396 16044
rect 24836 15876 24892 15886
rect 24780 15874 24892 15876
rect 24780 15822 24838 15874
rect 24890 15822 24892 15874
rect 24780 15810 24892 15822
rect 23436 15204 23492 15214
rect 22932 13972 22988 13982
rect 22932 13878 22988 13916
rect 23212 13972 23268 13982
rect 23212 13746 23268 13916
rect 23212 13694 23214 13746
rect 23266 13694 23268 13746
rect 23212 13682 23268 13694
rect 23324 13748 23380 13758
rect 23100 13636 23156 13646
rect 22652 13188 22708 13198
rect 22652 13094 22708 13132
rect 23100 12962 23156 13580
rect 23324 13578 23380 13692
rect 23324 13526 23326 13578
rect 23378 13526 23380 13578
rect 23436 13636 23492 15148
rect 24780 15204 24836 15810
rect 24780 15138 24836 15148
rect 25340 14420 25396 14430
rect 25340 13790 25396 14364
rect 23436 13570 23492 13580
rect 23548 13746 23604 13758
rect 23548 13694 23550 13746
rect 23602 13694 23604 13746
rect 25340 13738 25342 13790
rect 25394 13738 25396 13790
rect 25340 13726 25396 13738
rect 23324 13514 23380 13526
rect 23100 12910 23102 12962
rect 23154 12910 23156 12962
rect 22540 10882 22596 10892
rect 22652 12180 22708 12190
rect 22876 12180 22932 12190
rect 23100 12180 23156 12910
rect 23548 12964 23604 13694
rect 24164 13636 24220 13646
rect 24164 13542 24220 13580
rect 25228 13634 25284 13646
rect 25228 13582 25230 13634
rect 25282 13582 25284 13634
rect 25228 13524 25284 13582
rect 25228 13458 25284 13468
rect 23884 13300 23940 13310
rect 23884 13074 23940 13244
rect 23884 13022 23886 13074
rect 23938 13022 23940 13074
rect 23884 13010 23940 13022
rect 23548 12852 23604 12908
rect 23548 12796 23940 12852
rect 22652 12178 23156 12180
rect 22652 12126 22654 12178
rect 22706 12126 22878 12178
rect 22930 12126 23156 12178
rect 22652 12124 23156 12126
rect 23772 12178 23828 12190
rect 23772 12126 23774 12178
rect 23826 12126 23828 12178
rect 22652 10780 22708 12124
rect 22876 12114 22932 12124
rect 23772 11732 23828 12126
rect 23884 12066 23940 12796
rect 24220 12292 24276 12302
rect 24220 12234 24276 12236
rect 24220 12182 24222 12234
rect 24274 12182 24276 12234
rect 25452 12205 25508 17612
rect 26684 17610 26740 17622
rect 26684 17558 26686 17610
rect 26738 17558 26740 17610
rect 26160 17276 26424 17286
rect 26216 17220 26264 17276
rect 26320 17220 26368 17276
rect 26160 17210 26424 17220
rect 26684 17052 26740 17558
rect 27132 17610 27188 17622
rect 27132 17558 27134 17610
rect 27186 17558 27188 17610
rect 27132 17332 27188 17558
rect 27132 17266 27188 17276
rect 26124 16996 26740 17052
rect 27244 16996 27300 20636
rect 27748 20244 27804 20748
rect 28476 20802 28532 20814
rect 28476 20750 28478 20802
rect 28530 20750 28532 20802
rect 28140 20578 28196 20590
rect 28140 20526 28142 20578
rect 28194 20526 28196 20578
rect 28140 20188 28196 20526
rect 27748 20178 27804 20188
rect 27916 20132 28196 20188
rect 28476 20244 28532 20750
rect 29148 20804 29204 20814
rect 29148 20722 29150 20748
rect 29202 20722 29204 20748
rect 29148 20710 29204 20722
rect 28476 20178 28532 20188
rect 28924 20132 28980 20142
rect 27804 20020 27860 20030
rect 27916 20020 27972 20132
rect 27804 20018 27972 20020
rect 27804 19966 27806 20018
rect 27858 19966 27972 20018
rect 27804 19964 27972 19966
rect 28028 20020 28084 20030
rect 27804 19954 27860 19964
rect 27804 19124 27860 19134
rect 27804 19122 27972 19124
rect 27804 19070 27806 19122
rect 27858 19070 27972 19122
rect 27804 19068 27972 19070
rect 27804 19058 27860 19068
rect 27468 18489 27524 18501
rect 27468 18437 27470 18489
rect 27522 18437 27524 18489
rect 27468 18004 27524 18437
rect 27692 18452 27748 18462
rect 27692 18358 27748 18396
rect 27468 17948 27860 18004
rect 27804 17778 27860 17948
rect 27804 17726 27806 17778
rect 27858 17726 27860 17778
rect 27804 17714 27860 17726
rect 27580 17668 27636 17678
rect 27580 17577 27582 17612
rect 27634 17577 27636 17612
rect 27580 17565 27636 17577
rect 27778 17626 27834 17638
rect 27778 17574 27780 17626
rect 27832 17612 27834 17626
rect 27916 17612 27972 19068
rect 27832 17574 27972 17612
rect 27778 17556 27972 17574
rect 27778 17490 27834 17500
rect 26124 16100 26180 16996
rect 27020 16940 27300 16996
rect 27692 17332 27748 17342
rect 26908 16548 26964 16558
rect 26292 16324 26348 16334
rect 26292 16230 26348 16268
rect 26124 16006 26180 16044
rect 26908 16070 26964 16492
rect 26908 16018 26910 16070
rect 26962 16018 26964 16070
rect 26160 15708 26424 15718
rect 26216 15652 26264 15708
rect 26320 15652 26368 15708
rect 26160 15642 26424 15652
rect 26908 15204 26964 16018
rect 26908 15138 26964 15148
rect 27020 14980 27076 16940
rect 27244 16770 27300 16782
rect 27244 16718 27246 16770
rect 27298 16718 27300 16770
rect 27132 16660 27188 16670
rect 27132 16324 27188 16604
rect 27132 16098 27188 16268
rect 27244 16212 27300 16718
rect 27356 16212 27412 16222
rect 27244 16210 27412 16212
rect 27244 16158 27358 16210
rect 27410 16158 27412 16210
rect 27244 16156 27412 16158
rect 27356 16146 27412 16156
rect 27132 16046 27134 16098
rect 27186 16046 27188 16098
rect 27132 16034 27188 16046
rect 27524 16042 27580 16054
rect 27524 15990 27526 16042
rect 27578 15990 27580 16042
rect 27524 15988 27580 15990
rect 27524 15922 27580 15932
rect 27244 15314 27300 15326
rect 27244 15262 27246 15314
rect 27298 15262 27300 15314
rect 27244 14980 27300 15262
rect 27580 15316 27636 15326
rect 27580 15222 27636 15260
rect 27356 15204 27412 15214
rect 27356 15146 27412 15148
rect 27356 15094 27358 15146
rect 27410 15094 27412 15146
rect 27356 15082 27412 15094
rect 27692 14980 27748 17276
rect 28028 16882 28084 19964
rect 28812 19348 28868 19358
rect 28812 18477 28868 19292
rect 28924 18618 28980 20076
rect 29372 19908 29428 21534
rect 29484 21588 29540 21598
rect 29484 21494 29540 21532
rect 29708 20188 29764 22204
rect 29596 20132 29764 20188
rect 29932 21588 29988 21598
rect 29932 21474 29988 21532
rect 29932 21422 29934 21474
rect 29986 21422 29988 21474
rect 29932 20132 29988 21422
rect 30716 21476 30772 22876
rect 30940 21812 30996 23102
rect 30940 21746 30996 21756
rect 32060 22494 32116 25452
rect 32340 25442 32396 25452
rect 34476 25116 34740 25126
rect 34532 25060 34580 25116
rect 34636 25060 34684 25116
rect 34476 25050 34740 25060
rect 34476 23548 34740 23558
rect 34532 23492 34580 23548
rect 34636 23492 34684 23548
rect 34476 23482 34740 23492
rect 32060 22482 32172 22494
rect 32060 22430 32118 22482
rect 32170 22430 32172 22482
rect 32060 22418 32172 22430
rect 32060 21700 32116 22418
rect 34476 21980 34740 21990
rect 34532 21924 34580 21980
rect 34636 21924 34684 21980
rect 34476 21914 34740 21924
rect 33236 21700 33292 21710
rect 30716 21410 30772 21420
rect 31612 21698 33292 21700
rect 31612 21646 33238 21698
rect 33290 21646 33292 21698
rect 31612 21644 33292 21646
rect 30318 21196 30582 21206
rect 30374 21140 30422 21196
rect 30478 21140 30526 21196
rect 30318 21130 30582 21140
rect 30828 20804 30884 20814
rect 29596 20020 29652 20132
rect 29596 19954 29652 19964
rect 29428 19852 29540 19908
rect 29372 19842 29428 19852
rect 29148 19348 29204 19358
rect 29148 19254 29204 19292
rect 29316 19178 29372 19190
rect 29316 19126 29318 19178
rect 29370 19126 29372 19178
rect 29316 19124 29372 19126
rect 29316 19068 29428 19124
rect 28924 18566 28926 18618
rect 28978 18566 28980 18618
rect 28924 18554 28980 18566
rect 28476 18452 28532 18462
rect 28364 18450 28532 18452
rect 28364 18398 28478 18450
rect 28530 18398 28532 18450
rect 28364 18396 28532 18398
rect 28028 16830 28030 16882
rect 28082 16830 28084 16882
rect 28028 16772 28084 16830
rect 28028 16706 28084 16716
rect 28140 17668 28196 17678
rect 28140 16436 28196 17612
rect 28364 17668 28420 18396
rect 28476 18386 28532 18396
rect 28700 18452 28756 18462
rect 28812 18425 28814 18477
rect 28866 18425 28868 18477
rect 28812 18413 28868 18425
rect 29036 18452 29092 18462
rect 29036 18450 29316 18452
rect 28364 17602 28420 17612
rect 28476 17666 28532 17678
rect 28476 17614 28478 17666
rect 28530 17614 28532 17666
rect 28476 17556 28532 17614
rect 28308 17444 28364 17454
rect 28252 17442 28364 17444
rect 28252 17390 28310 17442
rect 28362 17390 28364 17442
rect 28252 17378 28364 17390
rect 28252 16884 28308 17378
rect 28364 16884 28420 16894
rect 28252 16882 28420 16884
rect 28252 16830 28366 16882
rect 28418 16830 28420 16882
rect 28252 16828 28420 16830
rect 28364 16818 28420 16828
rect 28476 16884 28532 17500
rect 28476 16818 28532 16828
rect 28588 17668 28644 17678
rect 28588 16938 28644 17612
rect 28700 17052 28756 18396
rect 29036 18398 29038 18450
rect 29090 18398 29316 18450
rect 29036 18396 29316 18398
rect 29036 18386 29092 18396
rect 29260 18228 29316 18396
rect 29260 17780 29316 18172
rect 29036 17724 29316 17780
rect 28812 17052 28868 17062
rect 28700 17050 28868 17052
rect 28700 16998 28814 17050
rect 28866 16998 28868 17050
rect 28700 16996 28868 16998
rect 28812 16986 28868 16996
rect 28924 16996 28980 17006
rect 28588 16886 28590 16938
rect 28642 16886 28644 16938
rect 28476 16660 28532 16670
rect 28588 16660 28644 16886
rect 28924 16882 28980 16940
rect 28924 16830 28926 16882
rect 28978 16830 28980 16882
rect 28924 16818 28980 16830
rect 28532 16604 28644 16660
rect 28476 16594 28532 16604
rect 28140 16380 28308 16436
rect 27804 16098 27860 16110
rect 27804 16046 27806 16098
rect 27858 16046 27860 16098
rect 27804 15764 27860 16046
rect 27972 16100 28028 16110
rect 27972 16006 28028 16044
rect 28252 16098 28308 16380
rect 28252 16046 28254 16098
rect 28306 16046 28308 16098
rect 27804 15698 27860 15708
rect 28140 15986 28196 15998
rect 28140 15934 28142 15986
rect 28194 15934 28196 15986
rect 28140 15540 28196 15934
rect 27916 15484 28196 15540
rect 28252 15540 28308 16046
rect 28532 15988 28588 15998
rect 28532 15894 28588 15932
rect 27916 14980 27972 15484
rect 28252 15428 28308 15484
rect 28196 15372 28308 15428
rect 28700 15764 28756 15774
rect 28196 15370 28252 15372
rect 28196 15318 28198 15370
rect 28250 15318 28252 15370
rect 28196 15306 28252 15318
rect 28476 15314 28532 15326
rect 28476 15262 28478 15314
rect 28530 15262 28532 15314
rect 27020 14924 27132 14980
rect 27244 14924 27972 14980
rect 28028 15202 28084 15214
rect 28028 15150 28030 15202
rect 28082 15150 28084 15202
rect 27076 14868 27132 14924
rect 27076 14812 27300 14868
rect 27132 14644 27188 14654
rect 26031 14532 26087 14542
rect 26031 14438 26087 14476
rect 26908 14530 26964 14542
rect 26908 14478 26910 14530
rect 26962 14478 26964 14530
rect 25788 14420 25844 14430
rect 25788 14326 25844 14364
rect 26160 14140 26424 14150
rect 26216 14084 26264 14140
rect 26320 14084 26368 14140
rect 26160 14074 26424 14084
rect 26460 13860 26516 13870
rect 24220 12170 24276 12182
rect 24444 12178 24500 12190
rect 23884 12014 23886 12066
rect 23938 12014 23940 12066
rect 23884 12002 23940 12014
rect 24444 12126 24446 12178
rect 24498 12126 24500 12178
rect 23772 11676 24164 11732
rect 22036 10724 22708 10780
rect 23324 10948 23380 10958
rect 22002 10220 22266 10230
rect 22058 10164 22106 10220
rect 22162 10164 22210 10220
rect 22002 10154 22266 10164
rect 21868 9874 21924 9884
rect 21980 9828 22036 9838
rect 20300 8990 20302 9042
rect 20354 8990 20356 9042
rect 20300 8978 20356 8990
rect 21868 9782 21924 9794
rect 21868 9730 21870 9782
rect 21922 9730 21924 9782
rect 21868 9044 21924 9730
rect 21980 9658 22036 9772
rect 21980 9606 21982 9658
rect 22034 9606 22036 9658
rect 21980 9594 22036 9606
rect 22204 9826 22260 9838
rect 22204 9774 22206 9826
rect 22258 9774 22260 9826
rect 21308 8370 21364 8382
rect 21308 8318 21310 8370
rect 21362 8318 21364 8370
rect 21308 7812 21364 8318
rect 21756 8260 21812 8270
rect 21868 8260 21924 8988
rect 22204 8932 22260 9774
rect 22204 8838 22260 8876
rect 22002 8652 22266 8662
rect 22058 8596 22106 8652
rect 22162 8596 22210 8652
rect 22002 8586 22266 8596
rect 22428 8484 22484 10724
rect 23119 10612 23175 10622
rect 22764 10610 23175 10612
rect 22764 10558 23121 10610
rect 23173 10558 23175 10610
rect 22764 10556 23175 10558
rect 22652 10052 22708 10062
rect 22652 9658 22708 9996
rect 22764 9828 22820 10556
rect 23119 10546 23175 10556
rect 22876 10388 22932 10398
rect 22876 10294 22932 10332
rect 23212 10052 23268 10062
rect 23100 9828 23156 9838
rect 22764 9826 22932 9828
rect 22764 9774 22766 9826
rect 22818 9774 22932 9826
rect 22764 9772 22932 9774
rect 22764 9762 22820 9772
rect 22652 9606 22654 9658
rect 22706 9606 22708 9658
rect 22652 9594 22708 9606
rect 22876 9156 22932 9772
rect 23100 9747 23102 9772
rect 23154 9747 23156 9772
rect 23100 9734 23156 9747
rect 23212 9492 23268 9996
rect 23324 9940 23380 10892
rect 24108 10724 24164 11676
rect 24332 11508 24388 11518
rect 24332 11414 24388 11452
rect 24108 10668 24388 10724
rect 23996 10612 24052 10622
rect 23996 10610 24276 10612
rect 23996 10558 23998 10610
rect 24050 10558 24276 10610
rect 23996 10556 24276 10558
rect 23996 10546 24052 10556
rect 23324 9826 23380 9884
rect 23940 9940 23996 9950
rect 23940 9846 23996 9884
rect 23324 9774 23326 9826
rect 23378 9774 23380 9826
rect 23324 9762 23380 9774
rect 24220 9604 24276 10556
rect 24220 9538 24276 9548
rect 23212 9436 23380 9492
rect 23044 9156 23100 9166
rect 22876 9154 23100 9156
rect 22876 9102 23046 9154
rect 23098 9102 23100 9154
rect 22876 9100 23100 9102
rect 23044 9090 23100 9100
rect 22652 9042 22708 9054
rect 22652 8990 22654 9042
rect 22706 8990 22708 9042
rect 22652 8932 22708 8990
rect 22652 8708 22708 8876
rect 22764 9044 22820 9054
rect 22764 8820 22820 8988
rect 22764 8764 23268 8820
rect 22652 8652 22932 8708
rect 22428 8418 22484 8428
rect 22652 8484 22708 8494
rect 21756 8258 21924 8260
rect 20076 7644 20244 7700
rect 20412 7756 21364 7812
rect 21420 8214 21476 8226
rect 21420 8162 21422 8214
rect 21474 8162 21476 8214
rect 21756 8206 21758 8258
rect 21810 8206 21924 8258
rect 21756 8204 21924 8206
rect 21756 8194 21812 8204
rect 19404 7308 19796 7364
rect 18396 6690 18452 6702
rect 18396 6638 18398 6690
rect 18450 6638 18452 6690
rect 19180 6692 19236 6702
rect 18396 6132 18452 6638
rect 18396 6066 18452 6076
rect 18732 6634 18788 6646
rect 18732 6582 18734 6634
rect 18786 6582 18788 6634
rect 18732 5908 18788 6582
rect 19068 6132 19124 6142
rect 18912 6020 18968 6030
rect 18912 5944 18968 5964
rect 18912 5892 18914 5944
rect 18966 5892 18968 5944
rect 18912 5880 18968 5892
rect 18732 5842 18788 5852
rect 18956 5796 19012 5806
rect 18956 5346 19012 5740
rect 18956 5294 18958 5346
rect 19010 5294 19012 5346
rect 18956 5282 19012 5294
rect 19068 5236 19124 6076
rect 19180 5906 19236 6636
rect 19516 6132 19572 6142
rect 19516 6018 19572 6076
rect 19516 5966 19518 6018
rect 19570 5966 19572 6018
rect 19516 5954 19572 5966
rect 19180 5854 19182 5906
rect 19234 5854 19236 5906
rect 19628 5908 19684 5918
rect 19180 5842 19236 5854
rect 19348 5850 19404 5862
rect 19068 5170 19124 5180
rect 19348 5798 19350 5850
rect 19402 5798 19404 5850
rect 18508 5124 18564 5134
rect 18508 5030 18564 5068
rect 19348 5124 19404 5798
rect 19628 5684 19684 5852
rect 19348 5030 19404 5068
rect 19516 5628 19684 5684
rect 19516 5122 19572 5628
rect 19516 5070 19518 5122
rect 19570 5070 19572 5122
rect 19516 5058 19572 5070
rect 19628 5236 19684 5246
rect 19628 5122 19684 5180
rect 19628 5070 19630 5122
rect 19682 5070 19684 5122
rect 19628 5058 19684 5070
rect 19628 4340 19684 4350
rect 19740 4340 19796 7308
rect 20076 7252 20132 7644
rect 20188 7476 20244 7486
rect 20412 7476 20468 7756
rect 20188 7474 20468 7476
rect 20188 7422 20190 7474
rect 20242 7422 20468 7474
rect 20188 7420 20468 7422
rect 20188 7410 20244 7420
rect 20076 7196 20244 7252
rect 19908 6020 19964 6030
rect 19908 5926 19964 5964
rect 20188 5124 20244 7196
rect 21420 6804 21476 8162
rect 21868 6916 21924 8204
rect 22428 8258 22484 8270
rect 22428 8206 22430 8258
rect 22482 8206 22484 8258
rect 22428 8036 22484 8206
rect 22428 7970 22484 7980
rect 22092 7588 22148 7598
rect 22092 7494 22148 7532
rect 22540 7588 22596 7598
rect 22002 7084 22266 7094
rect 22058 7028 22106 7084
rect 22162 7028 22210 7084
rect 22002 7018 22266 7028
rect 22204 6916 22260 6926
rect 21868 6914 22260 6916
rect 21868 6862 22206 6914
rect 22258 6862 22260 6914
rect 21868 6860 22260 6862
rect 22204 6850 22260 6860
rect 21420 6738 21476 6748
rect 21756 6804 21812 6814
rect 21364 5796 21420 5806
rect 21364 5346 21420 5740
rect 21364 5294 21366 5346
rect 21418 5294 21420 5346
rect 21364 5282 21420 5294
rect 21532 5348 21588 5358
rect 20412 5124 20468 5134
rect 20188 5122 20468 5124
rect 20188 5070 20414 5122
rect 20466 5070 20468 5122
rect 20188 5068 20468 5070
rect 20412 5058 20468 5068
rect 21532 5122 21588 5292
rect 21532 5070 21534 5122
rect 21586 5070 21588 5122
rect 21532 5058 21588 5070
rect 21756 5122 21812 6748
rect 22540 6690 22596 7532
rect 22652 7252 22708 8428
rect 22764 8372 22820 8410
rect 22764 8306 22820 8316
rect 22764 8202 22820 8214
rect 22764 8150 22766 8202
rect 22818 8150 22820 8202
rect 22764 7588 22820 8150
rect 22876 8036 22932 8652
rect 23100 8260 23156 8298
rect 23100 8194 23156 8204
rect 22876 7970 22932 7980
rect 23044 8036 23100 8046
rect 22764 7522 22820 7532
rect 22876 7812 22932 7822
rect 22876 7474 22932 7756
rect 22876 7422 22878 7474
rect 22930 7422 22932 7474
rect 23044 7530 23100 7980
rect 23044 7478 23046 7530
rect 23098 7478 23100 7530
rect 23212 7586 23268 8764
rect 23212 7534 23214 7586
rect 23266 7534 23268 7586
rect 23212 7522 23268 7534
rect 23044 7466 23100 7478
rect 23324 7474 23380 9436
rect 23604 8930 23660 8942
rect 23604 8878 23606 8930
rect 23658 8878 23660 8930
rect 23604 8484 23660 8878
rect 24332 8428 24388 10668
rect 24444 10500 24500 12126
rect 25452 12153 25454 12205
rect 25506 12153 25508 12205
rect 25452 11844 25508 12153
rect 25452 11778 25508 11788
rect 25676 13748 25732 13758
rect 26124 13748 26180 13758
rect 25676 13746 26180 13748
rect 25676 13694 25678 13746
rect 25730 13694 26126 13746
rect 26178 13694 26180 13746
rect 25676 13692 26180 13694
rect 25340 11508 25396 11518
rect 25340 11414 25396 11452
rect 24724 11396 24780 11406
rect 24724 10834 24780 11340
rect 25116 11396 25172 11406
rect 25676 11396 25732 13692
rect 26124 13682 26180 13692
rect 26460 13746 26516 13804
rect 26460 13694 26462 13746
rect 26514 13694 26516 13746
rect 26460 13682 26516 13694
rect 26572 13746 26628 13758
rect 26572 13694 26574 13746
rect 26626 13694 26628 13746
rect 25788 13524 25844 13534
rect 25788 13074 25844 13468
rect 25788 13022 25790 13074
rect 25842 13022 25844 13074
rect 25788 13010 25844 13022
rect 26460 13524 26516 13534
rect 26460 12962 26516 13468
rect 26460 12910 26462 12962
rect 26514 12910 26516 12962
rect 26460 12898 26516 12910
rect 26160 12572 26424 12582
rect 26216 12516 26264 12572
rect 26320 12516 26368 12572
rect 26160 12506 26424 12516
rect 26236 11954 26292 11966
rect 26236 11902 26238 11954
rect 26290 11902 26292 11954
rect 26124 11844 26180 11854
rect 26012 11620 26068 11630
rect 25788 11396 25844 11406
rect 25676 11394 25844 11396
rect 25116 11302 25172 11340
rect 25452 11350 25508 11362
rect 24724 10782 24726 10834
rect 24778 10782 24780 10834
rect 24724 10770 24780 10782
rect 25452 11298 25454 11350
rect 25506 11298 25508 11350
rect 25676 11342 25790 11394
rect 25842 11342 25844 11394
rect 25676 11340 25844 11342
rect 25340 10625 25396 10637
rect 25340 10612 25342 10625
rect 25394 10612 25396 10625
rect 25340 10533 25396 10556
rect 24444 10434 24500 10444
rect 25228 10500 25284 10510
rect 25228 10406 25284 10444
rect 25452 10388 25508 11298
rect 25452 10322 25508 10332
rect 25676 10610 25732 10622
rect 25676 10558 25678 10610
rect 25730 10558 25732 10610
rect 24780 10052 24836 10062
rect 24780 9826 24836 9996
rect 25676 9938 25732 10558
rect 25676 9886 25678 9938
rect 25730 9886 25732 9938
rect 25676 9874 25732 9886
rect 24780 9774 24782 9826
rect 24834 9774 24836 9826
rect 24780 9762 24836 9774
rect 25564 9826 25620 9838
rect 25564 9774 25566 9826
rect 25618 9774 25620 9826
rect 23604 8418 23660 8428
rect 23772 8372 24388 8428
rect 25116 9604 25172 9614
rect 25116 9044 25172 9548
rect 25564 9380 25620 9774
rect 25564 9324 25732 9380
rect 25564 9057 25620 9082
rect 24444 8372 24500 8382
rect 23436 8258 23492 8270
rect 23436 8206 23438 8258
rect 23490 8206 23492 8258
rect 23436 8148 23492 8206
rect 23436 8082 23492 8092
rect 22876 7410 22932 7422
rect 23324 7422 23326 7474
rect 23378 7422 23380 7474
rect 23324 7410 23380 7422
rect 23604 7476 23660 7486
rect 23604 7382 23660 7420
rect 22652 7196 22988 7252
rect 22540 6638 22542 6690
rect 22594 6638 22596 6690
rect 22540 6626 22596 6638
rect 22932 6692 22988 7196
rect 23212 7140 23268 7150
rect 23212 6804 23268 7084
rect 23100 6692 23156 6702
rect 22932 6690 23156 6692
rect 22932 6638 22934 6690
rect 22986 6638 23102 6690
rect 23154 6638 23156 6690
rect 22932 6636 23156 6638
rect 22932 6626 23044 6636
rect 23100 6626 23156 6636
rect 22652 6020 22708 6030
rect 22652 5950 22708 5964
rect 22316 5906 22372 5918
rect 22316 5854 22318 5906
rect 22370 5854 22372 5906
rect 22652 5898 22654 5950
rect 22706 5898 22708 5950
rect 22652 5886 22708 5898
rect 22316 5684 22372 5854
rect 22764 5796 22820 5806
rect 22316 5618 22372 5628
rect 22428 5794 22820 5796
rect 22428 5742 22766 5794
rect 22818 5742 22820 5794
rect 22428 5740 22820 5742
rect 22002 5516 22266 5526
rect 22058 5460 22106 5516
rect 22162 5460 22210 5516
rect 22002 5450 22266 5460
rect 22316 5348 22372 5358
rect 21756 5070 21758 5122
rect 21810 5070 21812 5122
rect 21756 5058 21812 5070
rect 22204 5124 22260 5134
rect 22204 5031 22206 5068
rect 22258 5031 22260 5068
rect 22204 5019 22260 5031
rect 21868 4954 21924 4966
rect 19628 4338 19796 4340
rect 19628 4286 19630 4338
rect 19682 4286 19796 4338
rect 19628 4284 19796 4286
rect 20076 4898 20132 4910
rect 20076 4846 20078 4898
rect 20130 4846 20132 4898
rect 19628 4274 19684 4284
rect 18284 4162 18340 4172
rect 14700 3714 14756 3724
rect 11228 3378 11284 3388
rect 18172 3554 18228 3566
rect 18172 3502 18174 3554
rect 18226 3502 18228 3554
rect 9528 3164 9792 3174
rect 9584 3108 9632 3164
rect 9688 3108 9736 3164
rect 9528 3098 9792 3108
rect 10780 800 10836 3378
rect 17844 3164 18108 3174
rect 17900 3108 17948 3164
rect 18004 3108 18052 3164
rect 17844 3098 18108 3108
rect 18172 1652 18228 3502
rect 20076 3526 20132 4846
rect 21868 4902 21870 4954
rect 21922 4902 21924 4954
rect 20412 4228 20468 4238
rect 20412 4226 20692 4228
rect 20412 4174 20414 4226
rect 20466 4174 20692 4226
rect 20412 4172 20692 4174
rect 20412 4162 20468 4172
rect 20636 3892 20692 4172
rect 20636 3836 21140 3892
rect 21084 3778 21140 3836
rect 21084 3726 21086 3778
rect 21138 3726 21140 3778
rect 21084 3714 21140 3726
rect 20076 3474 20078 3526
rect 20130 3474 20132 3526
rect 20076 3462 20132 3474
rect 21420 3556 21476 3566
rect 21420 3462 21476 3500
rect 21868 3556 21924 4902
rect 22316 4450 22372 5292
rect 22428 5122 22484 5740
rect 22764 5730 22820 5740
rect 22988 5124 23044 6626
rect 23212 6468 23268 6748
rect 22428 5070 22430 5122
rect 22482 5070 22484 5122
rect 22428 5058 22484 5070
rect 22764 5122 23044 5124
rect 22764 5070 22990 5122
rect 23042 5070 23044 5122
rect 22764 5068 23044 5070
rect 22316 4398 22318 4450
rect 22370 4398 22372 4450
rect 22316 4386 22372 4398
rect 22002 3948 22266 3958
rect 22058 3892 22106 3948
rect 22162 3892 22210 3948
rect 22002 3882 22266 3892
rect 22764 3678 22820 5068
rect 22988 5058 23044 5068
rect 23100 6412 23268 6468
rect 22988 4340 23044 4350
rect 23100 4340 23156 6412
rect 23212 6244 23268 6254
rect 23212 5906 23268 6188
rect 23772 6244 23828 8372
rect 24332 8258 24388 8270
rect 24108 8214 24164 8226
rect 24108 8162 24110 8214
rect 24162 8162 24164 8214
rect 24108 7812 24164 8162
rect 24332 8206 24334 8258
rect 24386 8206 24388 8258
rect 23996 7756 24164 7812
rect 24220 8090 24276 8102
rect 24220 8038 24222 8090
rect 24274 8038 24276 8090
rect 23996 7306 24052 7756
rect 24108 7476 24164 7486
rect 24108 7382 24164 7420
rect 23996 7254 23998 7306
rect 24050 7254 24052 7306
rect 23996 7242 24052 7254
rect 24220 7028 24276 8038
rect 24332 7476 24388 8206
rect 24332 7410 24388 7420
rect 24444 7474 24500 8316
rect 24444 7422 24446 7474
rect 24498 7422 24500 7474
rect 23884 6972 24276 7028
rect 24444 7028 24500 7422
rect 23884 6802 23940 6972
rect 24444 6962 24500 6972
rect 25116 8148 25172 8988
rect 23884 6750 23886 6802
rect 23938 6750 23940 6802
rect 23884 6738 23940 6750
rect 23996 6804 24052 6814
rect 23772 6178 23828 6188
rect 23884 6580 23940 6590
rect 23436 6132 23492 6142
rect 23884 6076 23940 6524
rect 23212 5854 23214 5906
rect 23266 5854 23268 5906
rect 23212 5796 23268 5854
rect 23212 5730 23268 5740
rect 23324 6020 23380 6030
rect 22988 4338 23156 4340
rect 22988 4286 22990 4338
rect 23042 4286 23156 4338
rect 22988 4284 23156 4286
rect 23324 4394 23380 5964
rect 23436 5962 23492 6076
rect 23436 5910 23438 5962
rect 23490 5910 23492 5962
rect 23436 5898 23492 5910
rect 23660 6074 23940 6076
rect 23660 6022 23886 6074
rect 23938 6022 23940 6074
rect 23660 6020 23940 6022
rect 23436 5796 23492 5806
rect 23436 4506 23492 5740
rect 23660 5124 23716 6020
rect 23884 6010 23940 6020
rect 23772 5908 23828 5918
rect 23996 5908 24052 6748
rect 24892 6132 24948 6142
rect 23772 5906 24052 5908
rect 23772 5854 23774 5906
rect 23826 5854 24052 5906
rect 23772 5852 24052 5854
rect 23772 5842 23828 5852
rect 23772 5684 23828 5694
rect 23772 5234 23828 5628
rect 23772 5182 23774 5234
rect 23826 5182 23828 5234
rect 23772 5170 23828 5182
rect 23660 5058 23716 5068
rect 23996 4900 24052 5852
rect 24220 5908 24276 5918
rect 24220 5814 24276 5852
rect 24556 5684 24612 5694
rect 24556 5590 24612 5628
rect 24892 4900 24948 6076
rect 23436 4454 23438 4506
rect 23490 4454 23492 4506
rect 23436 4442 23492 4454
rect 23772 4844 24276 4900
rect 23324 4342 23326 4394
rect 23378 4342 23380 4394
rect 22988 4274 23044 4284
rect 23324 4228 23380 4342
rect 23548 4340 23604 4350
rect 23324 4162 23380 4172
rect 23492 4338 23604 4340
rect 23492 4286 23550 4338
rect 23602 4286 23604 4338
rect 23492 4274 23604 4286
rect 23492 3778 23548 4274
rect 23492 3726 23494 3778
rect 23546 3726 23548 3778
rect 23492 3714 23548 3726
rect 22708 3666 22820 3678
rect 22708 3614 22710 3666
rect 22762 3614 22820 3666
rect 22708 3612 22820 3614
rect 22708 3602 22764 3612
rect 21868 3490 21924 3500
rect 23772 3554 23828 4844
rect 24220 4382 24276 4844
rect 24220 4330 24222 4382
rect 24274 4330 24276 4382
rect 24556 4844 24948 4900
rect 24556 4340 24612 4844
rect 24220 4318 24276 4330
rect 24332 4338 24612 4340
rect 24332 4286 24558 4338
rect 24610 4286 24612 4338
rect 24332 4284 24612 4286
rect 24108 4228 24164 4238
rect 24108 4134 24164 4172
rect 24332 4004 24388 4284
rect 24556 4274 24612 4284
rect 25116 4338 25172 8092
rect 25340 9042 25396 9054
rect 25340 8990 25342 9042
rect 25394 8990 25396 9042
rect 25340 8260 25396 8990
rect 25564 9044 25566 9057
rect 25618 9044 25620 9057
rect 25564 8978 25620 8988
rect 25676 8930 25732 9324
rect 25676 8878 25678 8930
rect 25730 8878 25732 8930
rect 25676 8866 25732 8878
rect 25340 6804 25396 8204
rect 25788 7476 25844 11340
rect 25900 11396 25956 11406
rect 25900 10610 25956 11340
rect 25900 10558 25902 10610
rect 25954 10558 25956 10610
rect 25900 10546 25956 10558
rect 26012 9787 26068 11564
rect 26124 11172 26180 11788
rect 26236 11396 26292 11902
rect 26572 11956 26628 13694
rect 26684 13636 26740 13646
rect 26684 12962 26740 13580
rect 26908 13524 26964 14478
rect 26908 13458 26964 13468
rect 26964 13188 27020 13198
rect 27132 13188 27188 14588
rect 26964 13186 27188 13188
rect 26964 13134 26966 13186
rect 27018 13134 27188 13186
rect 26964 13132 27188 13134
rect 26964 13122 27020 13132
rect 26684 12910 26686 12962
rect 26738 12910 26740 12962
rect 26684 12898 26740 12910
rect 26572 11900 26964 11956
rect 26740 11396 26796 11406
rect 26236 11394 26796 11396
rect 26236 11342 26742 11394
rect 26794 11342 26796 11394
rect 26236 11340 26796 11342
rect 26292 11172 26348 11182
rect 26124 11170 26348 11172
rect 26124 11118 26294 11170
rect 26346 11118 26348 11170
rect 26124 11116 26348 11118
rect 26292 11106 26348 11116
rect 26160 11004 26424 11014
rect 26216 10948 26264 11004
rect 26320 10948 26368 11004
rect 26160 10938 26424 10948
rect 26572 10052 26628 11340
rect 26740 11330 26796 11340
rect 26908 11396 26964 11900
rect 27132 11620 27188 13132
rect 27132 11554 27188 11564
rect 26908 11330 26964 11340
rect 27132 11172 27188 11182
rect 26684 11170 27188 11172
rect 26684 11118 27134 11170
rect 27186 11118 27188 11170
rect 26684 11116 27188 11118
rect 26684 10610 26740 11116
rect 27132 11106 27188 11116
rect 27244 10780 27300 14812
rect 27356 14644 27412 14924
rect 27356 14578 27412 14588
rect 27692 14532 27748 14542
rect 27692 14438 27748 14476
rect 28028 14503 28084 15150
rect 28476 15092 28532 15262
rect 28476 15026 28532 15036
rect 28028 14451 28030 14503
rect 28082 14451 28084 14503
rect 28364 14644 28420 14654
rect 28364 14530 28420 14588
rect 28364 14478 28366 14530
rect 28418 14478 28420 14530
rect 28364 14466 28420 14478
rect 28028 14439 28084 14451
rect 28252 14362 28308 14374
rect 28252 14310 28254 14362
rect 28306 14310 28308 14362
rect 28252 13972 28308 14310
rect 28252 13916 28532 13972
rect 27356 13636 27412 13646
rect 27356 13634 27636 13636
rect 27356 13582 27358 13634
rect 27410 13582 27636 13634
rect 27356 13580 27636 13582
rect 27356 13570 27412 13580
rect 27580 13188 27636 13580
rect 28476 13412 28532 13916
rect 28028 13356 28532 13412
rect 28700 13748 28756 15708
rect 28924 15540 28980 15550
rect 28924 15446 28980 15484
rect 29036 14644 29092 17724
rect 29372 17668 29428 19068
rect 29484 18452 29540 19852
rect 29708 19906 29764 19918
rect 29708 19854 29710 19906
rect 29762 19854 29764 19906
rect 29484 18386 29540 18396
rect 29596 19236 29652 19246
rect 29708 19236 29764 19854
rect 29932 19348 29988 20076
rect 30604 20132 30660 20142
rect 30268 20056 30324 20068
rect 30268 20004 30270 20056
rect 30322 20004 30324 20056
rect 30268 19908 30324 20004
rect 30604 20018 30660 20076
rect 30828 20130 30884 20748
rect 30828 20078 30830 20130
rect 30882 20078 30884 20130
rect 30828 20066 30884 20078
rect 31388 20804 31444 20814
rect 31612 20804 31668 21644
rect 32620 21586 32676 21644
rect 33236 21634 33292 21644
rect 32620 21534 32622 21586
rect 32674 21534 32676 21586
rect 32620 21522 32676 21534
rect 31836 21476 31892 21486
rect 31836 21382 31892 21420
rect 32340 21476 32396 21486
rect 31388 20802 31668 20804
rect 31388 20750 31390 20802
rect 31442 20750 31668 20802
rect 31388 20748 31668 20750
rect 31836 21028 31892 21038
rect 31836 20802 31892 20972
rect 32340 21026 32396 21420
rect 32340 20974 32342 21026
rect 32394 20974 32396 21026
rect 32340 20962 32396 20974
rect 31836 20750 31838 20802
rect 31890 20750 31892 20802
rect 31388 20020 31444 20748
rect 31836 20738 31892 20750
rect 32060 20804 32116 20814
rect 32060 20710 32116 20748
rect 34476 20412 34740 20422
rect 34532 20356 34580 20412
rect 34636 20356 34684 20412
rect 34476 20346 34740 20356
rect 30604 19966 30606 20018
rect 30658 19966 30660 20018
rect 30604 19954 30660 19966
rect 30996 19962 31052 19974
rect 30268 19842 30324 19852
rect 30996 19910 30998 19962
rect 31050 19910 31052 19962
rect 30318 19628 30582 19638
rect 30374 19572 30422 19628
rect 30478 19572 30526 19628
rect 30318 19562 30582 19572
rect 30996 19460 31052 19910
rect 30604 19404 31052 19460
rect 31276 19964 31388 20020
rect 29932 19292 30324 19348
rect 29596 19234 29988 19236
rect 29596 19182 29598 19234
rect 29650 19182 29988 19234
rect 29596 19180 29988 19182
rect 29484 17668 29540 17678
rect 29372 17666 29540 17668
rect 29372 17614 29486 17666
rect 29538 17614 29540 17666
rect 29372 17612 29540 17614
rect 29204 17556 29260 17566
rect 29148 17554 29260 17556
rect 29148 17502 29206 17554
rect 29258 17502 29260 17554
rect 29148 17490 29260 17502
rect 29484 17556 29540 17612
rect 29596 17666 29652 19180
rect 29932 18452 29988 19180
rect 30100 19012 30156 19022
rect 30100 18918 30156 18956
rect 30044 18452 30100 18462
rect 29932 18450 30100 18452
rect 29932 18398 30046 18450
rect 30098 18398 30100 18450
rect 29932 18396 30100 18398
rect 30044 18386 30100 18396
rect 30156 18452 30212 18462
rect 30156 18358 30212 18396
rect 29764 18228 29820 18238
rect 30268 18228 30324 19292
rect 29596 17614 29598 17666
rect 29650 17614 29652 17666
rect 29596 17602 29652 17614
rect 29708 18226 29820 18228
rect 29708 18174 29766 18226
rect 29818 18174 29820 18226
rect 29708 18162 29820 18174
rect 30156 18172 30324 18228
rect 30604 18340 30660 19404
rect 31276 19358 31332 19964
rect 31388 19954 31444 19964
rect 31948 20033 32004 20045
rect 31948 19981 31950 20033
rect 32002 19981 32004 20033
rect 31220 19346 31332 19358
rect 31220 19294 31222 19346
rect 31274 19294 31332 19346
rect 31220 19282 31332 19294
rect 31276 19012 31332 19282
rect 31836 19906 31892 19918
rect 31836 19854 31838 19906
rect 31890 19854 31892 19906
rect 31612 19124 31668 19134
rect 31612 19030 31668 19068
rect 31276 18946 31332 18956
rect 31052 18564 31108 18574
rect 30940 18465 30996 18477
rect 30716 18452 30772 18462
rect 30716 18450 30884 18452
rect 30716 18398 30718 18450
rect 30770 18398 30884 18450
rect 30716 18396 30884 18398
rect 30716 18386 30772 18396
rect 30604 18228 30660 18284
rect 30604 18172 30772 18228
rect 29484 17490 29540 17500
rect 29148 15316 29204 17490
rect 29596 17050 29652 17062
rect 29596 16998 29598 17050
rect 29650 16998 29652 17050
rect 29484 16884 29540 16894
rect 29484 16790 29540 16828
rect 29316 16772 29372 16782
rect 29316 16212 29372 16716
rect 29316 16118 29372 16156
rect 29260 15316 29316 15326
rect 29204 15314 29316 15316
rect 29204 15262 29262 15314
rect 29314 15262 29316 15314
rect 29204 15260 29316 15262
rect 29148 15222 29204 15260
rect 29036 14578 29092 14588
rect 29148 15092 29204 15102
rect 27692 13188 27748 13198
rect 27580 13186 27748 13188
rect 27580 13134 27694 13186
rect 27746 13134 27748 13186
rect 27580 13132 27748 13134
rect 27692 13122 27748 13132
rect 28028 12962 28084 13356
rect 28028 12910 28030 12962
rect 28082 12910 28084 12962
rect 28028 12898 28084 12910
rect 28364 12964 28420 12974
rect 28364 12740 28420 12908
rect 28700 12962 28756 13692
rect 29148 14530 29204 15036
rect 29148 14478 29150 14530
rect 29202 14478 29204 14530
rect 29148 13636 29204 14478
rect 29260 14530 29316 15260
rect 29596 14756 29652 16998
rect 29708 16996 29764 18162
rect 30156 17666 30212 18172
rect 30318 18060 30582 18070
rect 30374 18004 30422 18060
rect 30478 18004 30526 18060
rect 30318 17994 30582 18004
rect 30716 17892 30772 18172
rect 30828 18004 30884 18396
rect 30940 18413 30942 18465
rect 30994 18413 30996 18465
rect 30940 18340 30996 18413
rect 30940 18274 30996 18284
rect 31052 18338 31108 18508
rect 31836 18506 31892 19854
rect 31052 18286 31054 18338
rect 31106 18286 31108 18338
rect 31052 18274 31108 18286
rect 31388 18450 31444 18462
rect 31388 18398 31390 18450
rect 31442 18398 31444 18450
rect 31388 18228 31444 18398
rect 31388 18162 31444 18172
rect 31612 18452 31668 18462
rect 31836 18454 31838 18506
rect 31890 18454 31892 18506
rect 31948 18564 32004 19981
rect 32284 20018 32340 20030
rect 32284 19966 32286 20018
rect 32338 19966 32340 20018
rect 32172 19572 32228 19582
rect 32172 18618 32228 19516
rect 32284 19124 32340 19966
rect 32956 20018 33012 20030
rect 32956 19966 32958 20018
rect 33010 19966 33012 20018
rect 32956 19572 33012 19966
rect 33292 19796 33348 19806
rect 33292 19794 33572 19796
rect 33292 19742 33294 19794
rect 33346 19742 33572 19794
rect 33292 19740 33572 19742
rect 33292 19730 33348 19740
rect 32956 19506 33012 19516
rect 33516 19346 33572 19740
rect 33516 19294 33518 19346
rect 33570 19294 33572 19346
rect 33516 19282 33572 19294
rect 34300 19234 34356 19246
rect 34300 19182 34302 19234
rect 34354 19182 34356 19234
rect 32284 19058 32340 19068
rect 33292 19124 33348 19134
rect 32172 18566 32174 18618
rect 32226 18566 32228 18618
rect 32172 18554 32228 18566
rect 31948 18498 32004 18508
rect 31836 18442 31892 18454
rect 32060 18450 32116 18462
rect 30828 17948 30996 18004
rect 30604 17836 30772 17892
rect 30940 17892 30996 17948
rect 30940 17836 31332 17892
rect 30156 17614 30158 17666
rect 30210 17614 30212 17666
rect 30156 17602 30212 17614
rect 30492 17668 30548 17678
rect 30492 17574 30548 17612
rect 29708 16940 29820 16996
rect 29764 16938 29820 16940
rect 29764 16886 29766 16938
rect 29818 16886 29820 16938
rect 29764 16874 29820 16886
rect 30156 16884 30212 16894
rect 30156 16790 30212 16828
rect 30604 16660 30660 17836
rect 30828 17778 30884 17790
rect 30828 17726 30830 17778
rect 30882 17726 30884 17778
rect 30716 17668 30772 17678
rect 30716 17575 30718 17612
rect 30770 17575 30772 17612
rect 30716 17563 30772 17575
rect 30828 16884 30884 17726
rect 30828 16818 30884 16828
rect 30940 16670 30996 17836
rect 31164 17666 31220 17678
rect 31164 17614 31166 17666
rect 31218 17614 31220 17666
rect 31052 16884 31108 16894
rect 31052 16790 31108 16828
rect 30604 16604 30772 16660
rect 30318 16492 30582 16502
rect 30374 16436 30422 16492
rect 30478 16436 30526 16492
rect 30318 16426 30582 16436
rect 30716 16324 30772 16604
rect 30884 16658 30996 16670
rect 30884 16606 30886 16658
rect 30938 16606 30996 16658
rect 30884 16604 30996 16606
rect 30884 16594 30940 16604
rect 31164 16436 31220 17614
rect 31276 16884 31332 17836
rect 31612 17778 31668 18396
rect 32060 18398 32062 18450
rect 32114 18398 32116 18450
rect 31948 18340 32004 18350
rect 31612 17726 31614 17778
rect 31666 17726 31668 17778
rect 31612 17108 31668 17726
rect 31612 17042 31668 17052
rect 31724 18228 31780 18238
rect 31724 17668 31780 18172
rect 31724 16938 31780 17612
rect 31724 16886 31726 16938
rect 31778 16886 31780 16938
rect 31276 16882 31668 16884
rect 31276 16830 31278 16882
rect 31330 16830 31668 16882
rect 31724 16874 31780 16886
rect 31836 16884 31892 16894
rect 31276 16828 31668 16830
rect 31276 16818 31332 16828
rect 30492 16268 30772 16324
rect 30940 16380 31220 16436
rect 30156 15764 30212 15774
rect 30156 15428 30212 15708
rect 30492 15540 30548 16268
rect 30492 15538 30772 15540
rect 30492 15486 30494 15538
rect 30546 15486 30772 15538
rect 30492 15484 30772 15486
rect 30492 15474 30548 15484
rect 30156 15314 30212 15372
rect 30156 15262 30158 15314
rect 30210 15262 30212 15314
rect 30156 15250 30212 15262
rect 30318 14924 30582 14934
rect 30374 14868 30422 14924
rect 30478 14868 30526 14924
rect 30318 14858 30582 14868
rect 29596 14700 29764 14756
rect 29260 14478 29262 14530
rect 29314 14478 29316 14530
rect 29260 14466 29316 14478
rect 29372 14644 29428 14654
rect 29260 13636 29316 13646
rect 29148 13580 29260 13636
rect 29260 13542 29316 13580
rect 29372 13186 29428 14588
rect 29540 14532 29596 14542
rect 29540 14438 29596 14476
rect 29372 13134 29374 13186
rect 29426 13134 29428 13186
rect 28700 12910 28702 12962
rect 28754 12910 28756 12962
rect 28700 12898 28756 12910
rect 29036 12964 29092 12974
rect 29036 12870 29092 12908
rect 28140 12738 28420 12740
rect 28140 12686 28366 12738
rect 28418 12686 28420 12738
rect 28140 12684 28420 12686
rect 28028 12205 28084 12217
rect 28028 12153 28030 12205
rect 28082 12153 28084 12205
rect 28028 11844 28084 12153
rect 28028 11778 28084 11788
rect 26684 10558 26686 10610
rect 26738 10558 26740 10610
rect 26684 10546 26740 10558
rect 26908 10724 27300 10780
rect 27468 11394 27524 11406
rect 27468 11342 27470 11394
rect 27522 11342 27524 11394
rect 27468 10780 27524 11342
rect 27580 11396 27636 11406
rect 27580 11302 27636 11340
rect 27468 10724 28084 10780
rect 26572 9996 26740 10052
rect 26012 9735 26014 9787
rect 26066 9735 26068 9787
rect 26012 9723 26068 9735
rect 26236 9828 26292 9838
rect 26236 9734 26292 9772
rect 26572 9826 26628 9838
rect 26572 9774 26574 9826
rect 26626 9774 26628 9826
rect 26160 9436 26424 9446
rect 26216 9380 26264 9436
rect 26320 9380 26368 9436
rect 26160 9370 26424 9380
rect 26572 8820 26628 9774
rect 26460 8764 26628 8820
rect 26460 8036 26516 8764
rect 26460 7970 26516 7980
rect 26572 8484 26628 8494
rect 26684 8484 26740 9996
rect 26628 8428 26740 8484
rect 26908 8428 26964 10724
rect 27300 10052 27356 10062
rect 28028 10052 28084 10724
rect 27300 10050 27972 10052
rect 27300 9998 27302 10050
rect 27354 9998 27972 10050
rect 27300 9996 27972 9998
rect 27300 9986 27356 9996
rect 27468 9828 27524 9838
rect 27468 9734 27524 9772
rect 27804 9826 27860 9838
rect 27804 9774 27806 9826
rect 27858 9774 27860 9826
rect 27804 9044 27860 9774
rect 27916 9828 27972 9996
rect 28028 9986 28084 9996
rect 27916 9772 28028 9828
rect 27972 9770 28028 9772
rect 27972 9718 27974 9770
rect 28026 9718 28028 9770
rect 27972 9706 28028 9718
rect 28028 9044 28084 9054
rect 27804 8988 28028 9044
rect 28028 8950 28084 8988
rect 26160 7868 26424 7878
rect 26216 7812 26264 7868
rect 26320 7812 26368 7868
rect 26160 7802 26424 7812
rect 25788 7410 25844 7420
rect 25788 6804 25844 6814
rect 25340 6802 25844 6804
rect 25340 6750 25790 6802
rect 25842 6750 25844 6802
rect 25340 6748 25844 6750
rect 25788 6738 25844 6748
rect 26404 6692 26460 6702
rect 26572 6692 26628 8428
rect 26908 8372 27076 8428
rect 27020 7700 27076 8372
rect 27916 8260 27972 8270
rect 27916 8166 27972 8204
rect 28140 8260 28196 12684
rect 28364 12674 28420 12684
rect 29372 12180 29428 13134
rect 29708 12292 29764 14700
rect 30436 14532 30492 14542
rect 30324 14476 30436 14532
rect 29876 13972 29932 13982
rect 30324 13972 30380 14476
rect 30436 14438 30492 14476
rect 30716 14530 30772 15484
rect 30716 14478 30718 14530
rect 30770 14478 30772 14530
rect 29876 13970 30380 13972
rect 29876 13918 29878 13970
rect 29930 13918 30326 13970
rect 30378 13918 30380 13970
rect 29876 13916 30380 13918
rect 29876 13906 29932 13916
rect 30156 13188 30212 13916
rect 30324 13906 30380 13916
rect 30716 13860 30772 14478
rect 30716 13794 30772 13804
rect 30940 14420 30996 16380
rect 31220 16212 31276 16222
rect 31220 16118 31276 16156
rect 31612 16154 31668 16828
rect 31612 16102 31614 16154
rect 31666 16102 31668 16154
rect 31612 16090 31668 16102
rect 31836 16070 31892 16828
rect 31948 16884 32004 18284
rect 32060 17556 32116 18398
rect 33292 18450 33348 19068
rect 34300 19012 34356 19182
rect 33292 18398 33294 18450
rect 33346 18398 33348 18450
rect 33292 18386 33348 18398
rect 33404 18564 33460 18574
rect 33124 18228 33180 18238
rect 33124 18134 33180 18172
rect 32060 17050 32116 17500
rect 32060 16998 32062 17050
rect 32114 16998 32116 17050
rect 32060 16986 32116 16998
rect 32284 17668 32340 17678
rect 31948 16790 32004 16828
rect 32284 16210 32340 17612
rect 32956 16882 33012 16894
rect 32956 16830 32958 16882
rect 33010 16830 33012 16882
rect 32844 16324 32900 16334
rect 32284 16158 32286 16210
rect 32338 16158 32340 16210
rect 32284 16146 32340 16158
rect 32452 16322 32900 16324
rect 32452 16270 32846 16322
rect 32898 16270 32900 16322
rect 32452 16268 32900 16270
rect 32452 16154 32508 16268
rect 32844 16258 32900 16268
rect 32452 16102 32454 16154
rect 32506 16102 32508 16154
rect 32452 16090 32508 16102
rect 31836 16018 31838 16070
rect 31890 16018 31892 16070
rect 31836 15764 31892 16018
rect 31612 15708 31892 15764
rect 31612 15314 31668 15708
rect 31612 15262 31614 15314
rect 31666 15262 31668 15314
rect 31612 15250 31668 15262
rect 31724 15314 31780 15326
rect 31724 15262 31726 15314
rect 31778 15262 31780 15314
rect 31164 14644 31220 14654
rect 31724 14644 31780 15262
rect 31836 14868 31892 15708
rect 32956 15428 33012 16830
rect 33180 16884 33236 16894
rect 33404 16884 33460 18508
rect 33516 17668 33572 17678
rect 33516 17574 33572 17612
rect 34300 17666 34356 18956
rect 34476 18844 34740 18854
rect 34532 18788 34580 18844
rect 34636 18788 34684 18844
rect 34476 18778 34740 18788
rect 34300 17614 34302 17666
rect 34354 17614 34356 17666
rect 34300 17602 34356 17614
rect 34476 17276 34740 17286
rect 34532 17220 34580 17276
rect 34636 17220 34684 17276
rect 34476 17210 34740 17220
rect 33180 16882 33460 16884
rect 33180 16830 33182 16882
rect 33234 16830 33460 16882
rect 33180 16828 33460 16830
rect 33180 16818 33236 16828
rect 33460 16658 33516 16670
rect 33460 16606 33462 16658
rect 33514 16606 33516 16658
rect 33460 16322 33516 16606
rect 33460 16270 33462 16322
rect 33514 16270 33516 16322
rect 33460 16258 33516 16270
rect 34476 15708 34740 15718
rect 34532 15652 34580 15708
rect 34636 15652 34684 15708
rect 34476 15642 34740 15652
rect 32956 15362 33012 15372
rect 32004 15092 32060 15102
rect 32004 15090 32452 15092
rect 32004 15038 32006 15090
rect 32058 15038 32452 15090
rect 32004 15036 32452 15038
rect 32004 15026 32060 15036
rect 31836 14802 31892 14812
rect 31164 14642 31780 14644
rect 31164 14590 31166 14642
rect 31218 14590 31780 14642
rect 31164 14588 31780 14590
rect 32060 14756 32116 14766
rect 31164 14578 31220 14588
rect 30940 13746 30996 14364
rect 31052 14486 31108 14498
rect 31052 14434 31054 14486
rect 31106 14434 31108 14486
rect 31052 13914 31108 14434
rect 31612 14420 31668 14430
rect 31668 14364 32004 14420
rect 31612 14326 31668 14364
rect 31052 13862 31054 13914
rect 31106 13862 31108 13914
rect 31052 13850 31108 13862
rect 31948 13802 32004 14364
rect 30940 13694 30942 13746
rect 30994 13694 30996 13746
rect 30940 13682 30996 13694
rect 31220 13775 31276 13787
rect 31220 13723 31222 13775
rect 31274 13748 31276 13775
rect 31274 13723 31444 13748
rect 31220 13692 31444 13723
rect 30318 13356 30582 13366
rect 30374 13300 30422 13356
rect 30478 13300 30526 13356
rect 30318 13290 30582 13300
rect 30156 13132 30436 13188
rect 29932 12964 29988 12974
rect 29932 12870 29988 12908
rect 30268 12962 30324 12974
rect 30268 12910 30270 12962
rect 30322 12910 30324 12962
rect 30268 12852 30324 12910
rect 30268 12786 30324 12796
rect 30380 12962 30436 13132
rect 30380 12910 30382 12962
rect 30434 12910 30436 12962
rect 29708 12226 29764 12236
rect 30268 12180 30324 12190
rect 30380 12180 30436 12910
rect 31164 12964 31220 12974
rect 31164 12870 31220 12908
rect 31276 12852 31332 12862
rect 31276 12346 31332 12796
rect 31276 12294 31278 12346
rect 31330 12294 31332 12346
rect 31276 12282 31332 12294
rect 29372 12114 29428 12124
rect 30156 12178 30436 12180
rect 30156 12126 30270 12178
rect 30322 12126 30436 12178
rect 30156 12124 30436 12126
rect 31164 12180 31220 12190
rect 29316 11844 29372 11854
rect 29316 11506 29372 11788
rect 30156 11518 30212 12124
rect 30268 12114 30324 12124
rect 31164 12086 31220 12124
rect 31388 12180 31444 13692
rect 31724 13746 31780 13758
rect 31724 13694 31726 13746
rect 31778 13694 31780 13746
rect 31948 13750 31950 13802
rect 32002 13750 32004 13802
rect 31948 13738 32004 13750
rect 31724 13412 31780 13694
rect 31948 13636 32004 13646
rect 32060 13636 32116 14700
rect 32396 14308 32452 15036
rect 33516 14532 33572 14542
rect 33292 14530 33572 14532
rect 33292 14478 33518 14530
rect 33570 14478 33572 14530
rect 33292 14476 33572 14478
rect 32396 14252 33012 14308
rect 32284 13748 32340 13758
rect 32284 13746 32452 13748
rect 32284 13694 32286 13746
rect 32338 13694 32452 13746
rect 32284 13692 32452 13694
rect 32284 13682 32340 13692
rect 31948 13634 32116 13636
rect 31948 13582 31950 13634
rect 32002 13582 32116 13634
rect 31948 13580 32116 13582
rect 31948 13570 32004 13580
rect 31724 13346 31780 13356
rect 32284 13412 32340 13422
rect 31612 12740 31668 12750
rect 31612 12234 31668 12684
rect 31612 12182 31614 12234
rect 31666 12182 31668 12234
rect 31612 12170 31668 12182
rect 31836 12180 31892 12190
rect 31388 12114 31444 12124
rect 31276 11844 31332 11854
rect 30318 11788 30582 11798
rect 30374 11732 30422 11788
rect 30478 11732 30526 11788
rect 30318 11722 30582 11732
rect 29316 11454 29318 11506
rect 29370 11454 29372 11506
rect 29316 11442 29372 11454
rect 29764 11508 29820 11518
rect 30156 11508 30268 11518
rect 29764 11506 30268 11508
rect 29764 11454 29766 11506
rect 29818 11454 30214 11506
rect 30266 11454 30268 11506
rect 29764 11452 30268 11454
rect 29764 11396 29820 11452
rect 30212 11442 30268 11452
rect 29708 11340 29764 11396
rect 29708 11330 29820 11340
rect 29260 10612 29316 10622
rect 29036 10610 29316 10612
rect 29036 10558 29262 10610
rect 29314 10558 29316 10610
rect 29036 10556 29316 10558
rect 28588 10498 28644 10510
rect 28588 10446 28590 10498
rect 28642 10446 28644 10498
rect 28364 9828 28420 9838
rect 28252 9826 28420 9828
rect 28252 9774 28366 9826
rect 28418 9774 28420 9826
rect 28252 9772 28420 9774
rect 28252 9057 28308 9772
rect 28364 9762 28420 9772
rect 28588 9828 28644 10446
rect 28588 9762 28644 9772
rect 28476 9716 28532 9726
rect 28476 9658 28532 9660
rect 28476 9606 28478 9658
rect 28530 9606 28532 9658
rect 28476 9594 28532 9606
rect 28588 9604 28644 9614
rect 28252 9005 28254 9057
rect 28306 9005 28308 9057
rect 28252 8820 28308 9005
rect 28364 9268 28420 9278
rect 28364 8930 28420 9212
rect 28364 8878 28366 8930
rect 28418 8878 28420 8930
rect 28364 8866 28420 8878
rect 28252 8754 28308 8764
rect 28476 8372 28532 8382
rect 28588 8372 28644 9548
rect 28924 9070 28980 9082
rect 28924 9018 28926 9070
rect 28978 9018 28980 9070
rect 28924 8820 28980 9018
rect 28924 8754 28980 8764
rect 29036 8428 29092 10556
rect 29260 10546 29316 10556
rect 29596 10610 29652 10622
rect 29596 10558 29598 10610
rect 29650 10558 29652 10610
rect 29596 10500 29652 10558
rect 29596 10434 29652 10444
rect 29260 10052 29316 10062
rect 29260 9658 29316 9996
rect 29596 9940 29652 9950
rect 29260 9606 29262 9658
rect 29314 9606 29316 9658
rect 29372 9826 29428 9838
rect 29372 9774 29374 9826
rect 29426 9774 29428 9826
rect 29372 9716 29428 9774
rect 29596 9787 29652 9884
rect 29596 9735 29598 9787
rect 29650 9735 29652 9787
rect 29596 9723 29652 9735
rect 29372 9650 29428 9660
rect 29260 9594 29316 9606
rect 29260 9268 29316 9278
rect 29148 9044 29204 9054
rect 29148 8950 29204 8988
rect 29036 8372 29204 8428
rect 28476 8370 28644 8372
rect 28476 8318 28478 8370
rect 28530 8318 28644 8370
rect 28476 8316 28644 8318
rect 28476 8306 28532 8316
rect 28140 8166 28196 8204
rect 29036 8260 29092 8270
rect 29036 8166 29092 8204
rect 27580 8036 27636 8046
rect 27580 7942 27636 7980
rect 28252 8036 28308 8046
rect 25956 6690 26628 6692
rect 25956 6638 26406 6690
rect 26458 6638 26628 6690
rect 25956 6636 26628 6638
rect 26796 7644 27076 7700
rect 25284 6132 25340 6142
rect 25284 6038 25340 6076
rect 25956 6130 26012 6636
rect 26404 6626 26460 6636
rect 26160 6300 26424 6310
rect 26216 6244 26264 6300
rect 26320 6244 26368 6300
rect 26160 6234 26424 6244
rect 25956 6078 25958 6130
rect 26010 6078 26012 6130
rect 25956 6066 26012 6078
rect 25452 5906 25508 5918
rect 25452 5854 25454 5906
rect 25506 5854 25508 5906
rect 25452 5124 25508 5854
rect 26124 5908 26180 5918
rect 26124 5906 26628 5908
rect 26124 5854 26126 5906
rect 26178 5854 26628 5906
rect 26124 5852 26628 5854
rect 26124 5842 26180 5852
rect 26348 5348 26404 5358
rect 26348 5254 26404 5292
rect 25676 5124 25732 5134
rect 25452 5068 25676 5124
rect 25676 5030 25732 5068
rect 26160 4732 26424 4742
rect 26216 4676 26264 4732
rect 26320 4676 26368 4732
rect 26160 4666 26424 4676
rect 26572 4564 26628 5852
rect 26684 5124 26740 5134
rect 26796 5124 26852 7644
rect 27300 7503 27356 7515
rect 26908 7476 26964 7486
rect 27300 7451 27302 7503
rect 27354 7491 27356 7503
rect 27354 7451 27524 7491
rect 27300 7435 27524 7451
rect 26908 7382 26964 7420
rect 27356 7364 27412 7374
rect 27020 7362 27412 7364
rect 27020 7310 27358 7362
rect 27410 7310 27412 7362
rect 27020 7308 27412 7310
rect 26908 5908 26964 5918
rect 27020 5908 27076 7308
rect 27356 7298 27412 7308
rect 27468 6244 27524 7435
rect 27468 6178 27524 6188
rect 28028 6802 28084 6814
rect 28028 6750 28030 6802
rect 28082 6750 28084 6802
rect 26908 5906 27076 5908
rect 26908 5854 26910 5906
rect 26962 5854 27076 5906
rect 26908 5852 27076 5854
rect 26908 5842 26964 5852
rect 27244 5572 27300 5582
rect 26684 5122 26852 5124
rect 26684 5070 26686 5122
rect 26738 5070 26852 5122
rect 26684 5068 26852 5070
rect 26908 5124 26964 5134
rect 26684 5058 26740 5068
rect 26908 5030 26964 5068
rect 27244 5107 27300 5516
rect 27244 5055 27246 5107
rect 27298 5055 27300 5107
rect 27356 5234 27412 5246
rect 27356 5182 27358 5234
rect 27410 5182 27412 5234
rect 27356 5124 27412 5182
rect 27356 5058 27412 5068
rect 27804 5236 27860 5246
rect 27804 5122 27860 5180
rect 27804 5070 27806 5122
rect 27858 5070 27860 5122
rect 27804 5058 27860 5070
rect 28028 5095 28084 6750
rect 28252 6804 28308 7980
rect 28140 6646 28196 6658
rect 28140 6594 28142 6646
rect 28194 6594 28196 6646
rect 28140 6580 28196 6594
rect 28140 5908 28196 6524
rect 28140 5842 28196 5852
rect 28252 5236 28308 6748
rect 28476 6690 28532 6702
rect 28476 6638 28478 6690
rect 28530 6638 28532 6690
rect 28476 6020 28532 6638
rect 29036 6578 29092 6590
rect 29036 6526 29038 6578
rect 29090 6526 29092 6578
rect 28476 5954 28532 5964
rect 28812 6020 28868 6030
rect 29036 6020 29092 6526
rect 28812 6018 29092 6020
rect 28812 5966 28814 6018
rect 28866 5966 29092 6018
rect 28812 5964 29092 5966
rect 28812 5954 28868 5964
rect 28700 5908 28756 5918
rect 28700 5460 28756 5852
rect 28700 5404 28980 5460
rect 28252 5170 28308 5180
rect 27244 5043 27300 5055
rect 28028 5043 28030 5095
rect 28082 5043 28084 5095
rect 28364 5124 28420 5134
rect 28364 5122 28532 5124
rect 28364 5070 28366 5122
rect 28418 5070 28532 5122
rect 28364 5068 28532 5070
rect 28364 5058 28420 5068
rect 28028 5031 28084 5043
rect 25116 4286 25118 4338
rect 25170 4286 25172 4338
rect 25116 4274 25172 4286
rect 26348 4340 26404 4350
rect 26348 4246 26404 4284
rect 26460 4340 26516 4350
rect 26572 4340 26628 4508
rect 26460 4338 26628 4340
rect 26460 4286 26462 4338
rect 26514 4286 26628 4338
rect 26460 4284 26628 4286
rect 28364 4954 28420 4966
rect 28364 4902 28366 4954
rect 28418 4902 28420 4954
rect 28364 4340 28420 4902
rect 26460 4274 26516 4284
rect 28364 4274 28420 4284
rect 26012 4228 26068 4238
rect 26012 4134 26068 4172
rect 27244 4228 27300 4238
rect 27244 4134 27300 4172
rect 23772 3502 23774 3554
rect 23826 3502 23828 3554
rect 23772 3490 23828 3502
rect 23996 3948 24388 4004
rect 25452 4114 25508 4126
rect 25452 4062 25454 4114
rect 25506 4062 25508 4114
rect 23996 3554 24052 3948
rect 23996 3502 23998 3554
rect 24050 3502 24052 3554
rect 23996 3490 24052 3502
rect 25116 3668 25172 3678
rect 17948 1596 18228 1652
rect 17948 800 18004 1596
rect 25116 800 25172 3612
rect 25452 3526 25508 4062
rect 28476 3892 28532 5068
rect 28476 3836 28700 3892
rect 28644 3778 28700 3836
rect 28644 3726 28646 3778
rect 28698 3726 28700 3778
rect 26348 3668 26404 3678
rect 26348 3574 26404 3612
rect 25452 3474 25454 3526
rect 25506 3474 25508 3526
rect 28644 3556 28700 3726
rect 28644 3490 28700 3500
rect 28924 3554 28980 5404
rect 29148 5358 29204 8372
rect 29260 8258 29316 9212
rect 29708 9044 29764 11330
rect 29820 10649 29876 10661
rect 29820 10597 29822 10649
rect 29874 10597 29876 10649
rect 30940 10625 30996 10637
rect 29820 9828 29876 10597
rect 29932 10612 29988 10622
rect 29932 10498 29988 10556
rect 29932 10446 29934 10498
rect 29986 10446 29988 10498
rect 29932 10434 29988 10446
rect 30268 10610 30324 10622
rect 30268 10558 30270 10610
rect 30322 10558 30324 10610
rect 30268 10388 30324 10558
rect 30940 10612 30942 10625
rect 30994 10612 30996 10625
rect 30940 10533 30996 10556
rect 31276 10610 31332 11788
rect 31836 11788 31892 12124
rect 32284 11844 32340 13356
rect 32396 12964 32452 13692
rect 32956 13746 33012 14252
rect 33292 13970 33348 14476
rect 33516 14466 33572 14476
rect 34300 14532 34356 14542
rect 34300 14438 34356 14476
rect 34476 14140 34740 14150
rect 34532 14084 34580 14140
rect 34636 14084 34684 14140
rect 34476 14074 34740 14084
rect 33292 13918 33294 13970
rect 33346 13918 33348 13970
rect 33292 13906 33348 13918
rect 32956 13694 32958 13746
rect 33010 13694 33012 13746
rect 32956 13682 33012 13694
rect 33068 13412 33124 13422
rect 33068 13074 33124 13356
rect 33068 13022 33070 13074
rect 33122 13022 33124 13074
rect 33068 13010 33124 13022
rect 33852 13412 33908 13422
rect 33628 12964 33684 12987
rect 32452 12908 32564 12964
rect 32396 12898 32452 12908
rect 32340 11788 32452 11844
rect 31836 11732 32060 11788
rect 32284 11778 32340 11788
rect 32004 11618 32060 11732
rect 32004 11566 32006 11618
rect 32058 11566 32060 11618
rect 32004 11554 32060 11566
rect 32284 11394 32340 11406
rect 32284 11342 32286 11394
rect 32338 11342 32340 11394
rect 32284 11172 32340 11342
rect 32396 11394 32452 11788
rect 32396 11342 32398 11394
rect 32450 11342 32452 11394
rect 32396 11330 32452 11342
rect 32508 11172 32564 12908
rect 33516 12908 33628 12964
rect 32284 11116 32564 11172
rect 32732 11506 32788 11518
rect 32732 11454 32734 11506
rect 32786 11454 32788 11506
rect 31948 10778 32004 10790
rect 31948 10726 31950 10778
rect 32002 10726 32004 10778
rect 31276 10558 31278 10610
rect 31330 10558 31332 10610
rect 31276 10546 31332 10558
rect 31724 10610 31780 10622
rect 31724 10558 31726 10610
rect 31778 10558 31780 10610
rect 30828 10500 30884 10510
rect 30828 10406 30884 10444
rect 30156 10332 30324 10388
rect 29820 9762 29876 9772
rect 29932 9826 29988 9838
rect 29932 9774 29934 9826
rect 29986 9774 29988 9826
rect 29932 9604 29988 9774
rect 29932 9538 29988 9548
rect 30156 9044 30212 10332
rect 30318 10220 30582 10230
rect 30374 10164 30422 10220
rect 30478 10164 30526 10220
rect 30318 10154 30582 10164
rect 30380 9940 30436 9950
rect 30380 9846 30436 9884
rect 30716 9828 30772 9838
rect 30492 9782 30548 9794
rect 30492 9730 30494 9782
rect 30546 9730 30548 9782
rect 30716 9734 30772 9772
rect 31388 9826 31444 9838
rect 31388 9774 31390 9826
rect 31442 9774 31444 9826
rect 30492 9268 30548 9730
rect 31388 9268 31444 9774
rect 31724 9604 31780 10558
rect 31388 9212 31668 9268
rect 30492 9202 30548 9212
rect 29708 9042 30100 9044
rect 29540 8986 29596 8998
rect 29372 8932 29428 8942
rect 29372 8838 29428 8876
rect 29540 8934 29542 8986
rect 29594 8934 29596 8986
rect 29708 8990 29710 9042
rect 29762 8990 30100 9042
rect 29708 8988 30100 8990
rect 29708 8978 29764 8988
rect 29540 8482 29596 8934
rect 29540 8430 29542 8482
rect 29594 8430 29596 8482
rect 29540 8418 29596 8430
rect 29932 8820 29988 8830
rect 29260 8206 29262 8258
rect 29314 8206 29316 8258
rect 29260 8194 29316 8206
rect 29764 7588 29820 7598
rect 29260 7474 29316 7486
rect 29260 7422 29262 7474
rect 29314 7422 29316 7474
rect 29260 6580 29316 7422
rect 29484 7476 29540 7486
rect 29484 7382 29540 7420
rect 29764 7140 29820 7532
rect 29764 7074 29820 7084
rect 29932 7140 29988 8764
rect 30044 8428 30100 8988
rect 30156 8978 30212 8988
rect 30492 8932 30548 8942
rect 30492 8838 30548 8876
rect 30318 8652 30582 8662
rect 30374 8596 30422 8652
rect 30478 8596 30526 8652
rect 30318 8586 30582 8596
rect 30044 8372 30212 8428
rect 30100 8370 30212 8372
rect 30100 8318 30102 8370
rect 30154 8318 30212 8370
rect 30100 8296 30212 8318
rect 29932 7074 29988 7084
rect 29484 6690 29540 6702
rect 29484 6638 29486 6690
rect 29538 6638 29540 6690
rect 29484 6580 29540 6638
rect 29260 6578 29540 6580
rect 29260 6526 29262 6578
rect 29314 6526 29540 6578
rect 29260 6524 29540 6526
rect 29596 6692 29652 6702
rect 29260 6514 29316 6524
rect 29596 6356 29652 6636
rect 30156 6580 30212 8296
rect 31220 8036 31276 8046
rect 31612 8036 31668 9212
rect 31220 8034 31668 8036
rect 31220 7982 31222 8034
rect 31274 7982 31668 8034
rect 31220 7980 31668 7982
rect 30318 7084 30582 7094
rect 30374 7028 30422 7084
rect 30478 7028 30526 7084
rect 30318 7018 30582 7028
rect 30360 6692 30416 6702
rect 30360 6690 30436 6692
rect 30360 6638 30362 6690
rect 30414 6638 30436 6690
rect 30360 6626 30436 6638
rect 30156 6524 30324 6580
rect 30156 6356 30212 6366
rect 29596 6300 29876 6356
rect 29596 6020 29652 6030
rect 29484 5908 29540 5918
rect 29484 5814 29540 5852
rect 29148 5346 29260 5358
rect 29148 5294 29206 5346
rect 29258 5294 29260 5346
rect 29148 5292 29260 5294
rect 29204 5282 29260 5292
rect 29484 5124 29540 5134
rect 29484 5030 29540 5068
rect 29596 5122 29652 5964
rect 29820 5906 29876 6300
rect 29820 5854 29822 5906
rect 29874 5854 29876 5906
rect 30044 6020 30100 6030
rect 30044 5962 30100 5964
rect 30044 5910 30046 5962
rect 30098 5910 30100 5962
rect 30044 5898 30100 5910
rect 29820 5842 29876 5854
rect 30156 5794 30212 6300
rect 30156 5742 30158 5794
rect 30210 5742 30212 5794
rect 30156 5730 30212 5742
rect 29596 5070 29598 5122
rect 29650 5070 29652 5122
rect 29596 4676 29652 5070
rect 28924 3502 28926 3554
rect 28978 3502 28980 3554
rect 28924 3490 28980 3502
rect 29148 4620 29652 4676
rect 29820 5684 29876 5694
rect 29148 4450 29204 4620
rect 29820 4574 29876 5628
rect 30268 5684 30324 6524
rect 30380 6132 30436 6626
rect 30604 6578 30660 6590
rect 30604 6526 30606 6578
rect 30658 6526 30660 6578
rect 30604 6244 30660 6526
rect 31220 6468 31276 7980
rect 31612 7476 31668 7486
rect 31612 7382 31668 7420
rect 31388 6690 31444 6702
rect 31388 6638 31390 6690
rect 31442 6638 31444 6690
rect 31388 6468 31444 6638
rect 31220 6466 31444 6468
rect 31220 6414 31222 6466
rect 31274 6414 31444 6466
rect 31220 6412 31444 6414
rect 31220 6402 31276 6412
rect 30604 6178 30660 6188
rect 30380 6066 30436 6076
rect 30380 5906 30436 5918
rect 30380 5854 30382 5906
rect 30434 5854 30436 5906
rect 30380 5796 30436 5854
rect 30380 5730 30436 5740
rect 30996 5794 31052 5806
rect 30996 5742 30998 5794
rect 31050 5742 31052 5794
rect 30268 5618 30324 5628
rect 30716 5684 30772 5694
rect 30318 5516 30582 5526
rect 30374 5460 30422 5516
rect 30478 5460 30526 5516
rect 30318 5450 30582 5460
rect 30380 5124 30436 5134
rect 30380 5030 30436 5068
rect 30604 5066 30660 5078
rect 30604 5014 30606 5066
rect 30658 5014 30660 5066
rect 30604 4900 30660 5014
rect 30604 4834 30660 4844
rect 29764 4564 29876 4574
rect 29820 4508 29876 4564
rect 29764 4470 29820 4508
rect 29148 4398 29150 4450
rect 29202 4398 29204 4450
rect 29148 3554 29204 4398
rect 30318 3948 30582 3958
rect 30374 3892 30422 3948
rect 30478 3892 30526 3948
rect 30318 3882 30582 3892
rect 30716 3678 30772 5628
rect 30996 5684 31052 5742
rect 30996 5618 31052 5628
rect 31276 5796 31332 5806
rect 30940 5236 30996 5246
rect 30940 5122 30996 5180
rect 30940 5070 30942 5122
rect 30994 5070 30996 5122
rect 30940 5058 30996 5070
rect 31052 4954 31108 4966
rect 30660 3666 30772 3678
rect 30660 3614 30662 3666
rect 30714 3614 30772 3666
rect 30660 3612 30772 3614
rect 30940 4900 30996 4910
rect 30940 3666 30996 4844
rect 31052 4902 31054 4954
rect 31106 4902 31108 4954
rect 31052 3892 31108 4902
rect 31052 3826 31108 3836
rect 30940 3614 30942 3666
rect 30994 3614 30996 3666
rect 30660 3602 30716 3612
rect 30940 3602 30996 3614
rect 29148 3502 29150 3554
rect 29202 3502 29204 3554
rect 29148 3490 29204 3502
rect 31052 3556 31108 3566
rect 25452 3462 25508 3474
rect 31052 3487 31054 3500
rect 31106 3487 31108 3500
rect 31276 3556 31332 5740
rect 31388 5684 31444 6412
rect 31388 5122 31444 5628
rect 31388 5070 31390 5122
rect 31442 5070 31444 5122
rect 31388 5058 31444 5070
rect 31612 5908 31668 5918
rect 31724 5908 31780 9548
rect 31948 9268 32004 10726
rect 32060 10666 32116 10678
rect 32060 10614 32062 10666
rect 32114 10614 32116 10666
rect 32060 10388 32116 10614
rect 32284 10610 32340 11116
rect 32284 10558 32286 10610
rect 32338 10558 32340 10610
rect 32284 10546 32340 10558
rect 32732 10388 32788 11454
rect 33180 11394 33236 11406
rect 32900 11338 32956 11350
rect 32900 11286 32902 11338
rect 32954 11286 32956 11338
rect 32900 11284 32956 11286
rect 33180 11342 33182 11394
rect 33234 11342 33236 11394
rect 32900 11228 33012 11284
rect 32956 11172 33012 11228
rect 32956 11116 33124 11172
rect 32956 10612 33012 10622
rect 33068 10612 33124 11116
rect 33180 10836 33236 11342
rect 33180 10770 33236 10780
rect 33516 10734 33572 12908
rect 33628 12895 33630 12908
rect 33682 12895 33684 12908
rect 33852 12962 33908 13356
rect 33852 12910 33854 12962
rect 33906 12910 33908 12962
rect 33852 12898 33908 12910
rect 33628 12883 33684 12895
rect 33628 12794 33684 12806
rect 33628 12742 33630 12794
rect 33682 12742 33684 12794
rect 33628 12740 33684 12742
rect 33628 12674 33684 12684
rect 34476 12572 34740 12582
rect 34532 12516 34580 12572
rect 34636 12516 34684 12572
rect 34476 12506 34740 12516
rect 34476 11004 34740 11014
rect 34532 10948 34580 11004
rect 34636 10948 34684 11004
rect 34476 10938 34740 10948
rect 33460 10722 33572 10734
rect 33460 10670 33462 10722
rect 33514 10670 33572 10722
rect 33460 10668 33572 10670
rect 33460 10658 33516 10668
rect 33180 10612 33236 10622
rect 34076 10612 34132 10622
rect 33068 10610 33348 10612
rect 33068 10558 33182 10610
rect 33234 10558 33348 10610
rect 33068 10556 33348 10558
rect 32956 10518 33012 10556
rect 33180 10546 33236 10556
rect 32060 10332 32788 10388
rect 32172 9828 32228 9838
rect 32172 9826 32452 9828
rect 32172 9774 32174 9826
rect 32226 9774 32452 9826
rect 32172 9772 32452 9774
rect 32172 9762 32228 9772
rect 32396 9380 32452 9772
rect 33292 9716 33348 10556
rect 34076 9938 34132 10556
rect 34076 9886 34078 9938
rect 34130 9886 34132 9938
rect 34076 9874 34132 9886
rect 33292 9650 33348 9660
rect 34476 9436 34740 9446
rect 34532 9380 34580 9436
rect 34636 9380 34684 9436
rect 32396 9324 33348 9380
rect 34476 9370 34740 9380
rect 31948 9212 33012 9268
rect 31892 9044 31948 9054
rect 31892 8482 31948 8988
rect 32956 9042 33012 9212
rect 33292 9266 33348 9324
rect 33292 9214 33294 9266
rect 33346 9214 33348 9266
rect 33292 9202 33348 9214
rect 32956 8990 32958 9042
rect 33010 8990 33012 9042
rect 32956 8978 33012 8990
rect 31892 8430 31894 8482
rect 31946 8430 31948 8482
rect 31892 8418 31948 8430
rect 32396 8930 32452 8942
rect 32396 8878 32398 8930
rect 32450 8878 32452 8930
rect 32396 8428 32452 8878
rect 32060 8372 32452 8428
rect 32060 8258 32116 8372
rect 32060 8206 32062 8258
rect 32114 8206 32116 8258
rect 32060 8194 32116 8206
rect 34476 7868 34740 7878
rect 34532 7812 34580 7868
rect 34636 7812 34684 7868
rect 34476 7802 34740 7812
rect 31948 7489 32004 7501
rect 31948 7437 31950 7489
rect 32002 7437 32004 7489
rect 31612 5906 31780 5908
rect 31612 5854 31614 5906
rect 31666 5854 31780 5906
rect 31836 7364 31892 7374
rect 31836 5962 31892 7308
rect 31836 5910 31838 5962
rect 31890 5910 31892 5962
rect 31836 5898 31892 5910
rect 31948 5908 32004 7437
rect 32956 7474 33012 7486
rect 32956 7422 32958 7474
rect 33010 7422 33012 7474
rect 32060 7364 32116 7374
rect 32060 7270 32116 7308
rect 32956 7028 33012 7422
rect 33628 7476 33684 7486
rect 32284 6972 33012 7028
rect 33292 7250 33348 7262
rect 33292 7198 33294 7250
rect 33346 7198 33348 7250
rect 32172 6804 32228 6814
rect 32172 6710 32228 6748
rect 31612 5852 31780 5854
rect 31612 5124 31668 5852
rect 31612 5058 31668 5068
rect 31948 5236 32004 5852
rect 32172 6132 32228 6142
rect 32172 5906 32228 6076
rect 32284 6074 32340 6972
rect 33292 6804 33348 7198
rect 33292 6738 33348 6748
rect 32284 6022 32286 6074
rect 32338 6022 32340 6074
rect 32284 6010 32340 6022
rect 33124 6132 33180 6142
rect 33124 6018 33180 6076
rect 33124 5966 33126 6018
rect 33178 5966 33180 6018
rect 33124 5954 33180 5966
rect 32172 5854 32174 5906
rect 32226 5854 32228 5906
rect 32172 5842 32228 5854
rect 33404 5908 33460 5918
rect 33404 5814 33460 5852
rect 33628 5906 33684 7420
rect 34076 7476 34132 7486
rect 34076 6690 34132 7420
rect 34076 6638 34078 6690
rect 34130 6638 34132 6690
rect 34076 6626 34132 6638
rect 34476 6300 34740 6310
rect 34532 6244 34580 6300
rect 34636 6244 34684 6300
rect 34476 6234 34740 6244
rect 33628 5854 33630 5906
rect 33682 5854 33684 5906
rect 33628 5842 33684 5854
rect 34076 5796 34132 5806
rect 31500 4116 31556 4126
rect 31500 4022 31556 4060
rect 31948 3780 32004 5180
rect 32396 5348 32452 5358
rect 32172 5124 32228 5134
rect 32172 5122 32340 5124
rect 32172 5070 32174 5122
rect 32226 5070 32340 5122
rect 32172 5068 32340 5070
rect 32172 5058 32228 5068
rect 31948 3714 32004 3724
rect 32172 4116 32228 4126
rect 32284 4116 32340 5068
rect 32396 4228 32452 5292
rect 34076 5234 34132 5740
rect 34076 5182 34078 5234
rect 34130 5182 34132 5234
rect 34076 5170 34132 5182
rect 34476 4732 34740 4742
rect 34532 4676 34580 4732
rect 34636 4676 34684 4732
rect 34476 4666 34740 4676
rect 33292 4564 33348 4574
rect 32508 4562 33348 4564
rect 32508 4510 33294 4562
rect 33346 4510 33348 4562
rect 32508 4508 33348 4510
rect 32508 4365 32564 4508
rect 33292 4498 33348 4508
rect 32508 4313 32510 4365
rect 32562 4313 32564 4365
rect 32508 4301 32564 4313
rect 32956 4338 33012 4350
rect 32956 4286 32958 4338
rect 33010 4286 33012 4338
rect 32956 4228 33012 4286
rect 32396 4172 33012 4228
rect 32284 4060 33236 4116
rect 32060 3556 32116 3566
rect 31276 3554 32116 3556
rect 31276 3502 31278 3554
rect 31330 3502 32062 3554
rect 32114 3502 32116 3554
rect 31276 3500 32116 3502
rect 31276 3490 31332 3500
rect 32060 3490 32116 3500
rect 31052 3462 31108 3487
rect 26160 3164 26424 3174
rect 26216 3108 26264 3164
rect 26320 3108 26368 3164
rect 26160 3098 26424 3108
rect 32172 2100 32228 4060
rect 32844 3892 32900 3902
rect 32564 3780 32620 3790
rect 32564 3686 32620 3724
rect 32284 3556 32340 3566
rect 32284 3462 32340 3500
rect 32844 3554 32900 3836
rect 33180 3778 33236 4060
rect 33180 3726 33182 3778
rect 33234 3726 33236 3778
rect 33180 3714 33236 3726
rect 32844 3502 32846 3554
rect 32898 3502 32900 3554
rect 32844 3490 32900 3502
rect 34476 3164 34740 3174
rect 34532 3108 34580 3164
rect 34636 3108 34684 3164
rect 34476 3098 34740 3108
rect 32172 2044 32340 2100
rect 32284 800 32340 2044
rect 3584 0 3696 800
rect 10752 0 10864 800
rect 17920 0 18032 800
rect 25088 0 25200 800
rect 32256 0 32368 800
<< via2 >>
rect 5370 32170 5426 32172
rect 5370 32118 5372 32170
rect 5372 32118 5424 32170
rect 5424 32118 5426 32170
rect 5370 32116 5426 32118
rect 5474 32170 5530 32172
rect 5474 32118 5476 32170
rect 5476 32118 5528 32170
rect 5528 32118 5530 32170
rect 5474 32116 5530 32118
rect 5578 32170 5634 32172
rect 5578 32118 5580 32170
rect 5580 32118 5632 32170
rect 5632 32118 5634 32170
rect 5578 32116 5634 32118
rect 13686 32170 13742 32172
rect 13686 32118 13688 32170
rect 13688 32118 13740 32170
rect 13740 32118 13742 32170
rect 13686 32116 13742 32118
rect 13790 32170 13846 32172
rect 13790 32118 13792 32170
rect 13792 32118 13844 32170
rect 13844 32118 13846 32170
rect 13790 32116 13846 32118
rect 13894 32170 13950 32172
rect 13894 32118 13896 32170
rect 13896 32118 13948 32170
rect 13948 32118 13950 32170
rect 13894 32116 13950 32118
rect 22002 32170 22058 32172
rect 22002 32118 22004 32170
rect 22004 32118 22056 32170
rect 22056 32118 22058 32170
rect 22002 32116 22058 32118
rect 22106 32170 22162 32172
rect 22106 32118 22108 32170
rect 22108 32118 22160 32170
rect 22160 32118 22162 32170
rect 22106 32116 22162 32118
rect 22210 32170 22266 32172
rect 22210 32118 22212 32170
rect 22212 32118 22264 32170
rect 22264 32118 22266 32170
rect 22210 32116 22266 32118
rect 30318 32170 30374 32172
rect 30318 32118 30320 32170
rect 30320 32118 30372 32170
rect 30372 32118 30374 32170
rect 30318 32116 30374 32118
rect 30422 32170 30478 32172
rect 30422 32118 30424 32170
rect 30424 32118 30476 32170
rect 30476 32118 30478 32170
rect 30422 32116 30478 32118
rect 30526 32170 30582 32172
rect 30526 32118 30528 32170
rect 30528 32118 30580 32170
rect 30580 32118 30582 32170
rect 30526 32116 30582 32118
rect 9528 31386 9584 31388
rect 9528 31334 9530 31386
rect 9530 31334 9582 31386
rect 9582 31334 9584 31386
rect 9528 31332 9584 31334
rect 9632 31386 9688 31388
rect 9632 31334 9634 31386
rect 9634 31334 9686 31386
rect 9686 31334 9688 31386
rect 9632 31332 9688 31334
rect 9736 31386 9792 31388
rect 9736 31334 9738 31386
rect 9738 31334 9790 31386
rect 9790 31334 9792 31386
rect 9736 31332 9792 31334
rect 19628 31890 19684 31892
rect 19628 31838 19630 31890
rect 19630 31838 19682 31890
rect 19682 31838 19684 31890
rect 19628 31836 19684 31838
rect 20524 31836 20580 31892
rect 5370 30602 5426 30604
rect 5370 30550 5372 30602
rect 5372 30550 5424 30602
rect 5424 30550 5426 30602
rect 5370 30548 5426 30550
rect 5474 30602 5530 30604
rect 5474 30550 5476 30602
rect 5476 30550 5528 30602
rect 5528 30550 5530 30602
rect 5474 30548 5530 30550
rect 5578 30602 5634 30604
rect 5578 30550 5580 30602
rect 5580 30550 5632 30602
rect 5632 30550 5634 30602
rect 5578 30548 5634 30550
rect 10444 30210 10500 30212
rect 10444 30158 10446 30210
rect 10446 30158 10498 30210
rect 10498 30158 10500 30210
rect 10444 30156 10500 30158
rect 11564 30044 11620 30100
rect 11676 30156 11732 30212
rect 14812 31500 14868 31556
rect 13686 30602 13742 30604
rect 13686 30550 13688 30602
rect 13688 30550 13740 30602
rect 13740 30550 13742 30602
rect 13686 30548 13742 30550
rect 13790 30602 13846 30604
rect 13790 30550 13792 30602
rect 13792 30550 13844 30602
rect 13844 30550 13846 30602
rect 13790 30548 13846 30550
rect 13894 30602 13950 30604
rect 13894 30550 13896 30602
rect 13896 30550 13948 30602
rect 13948 30550 13950 30602
rect 13894 30548 13950 30550
rect 9528 29818 9584 29820
rect 9528 29766 9530 29818
rect 9530 29766 9582 29818
rect 9582 29766 9584 29818
rect 9528 29764 9584 29766
rect 9632 29818 9688 29820
rect 9632 29766 9634 29818
rect 9634 29766 9686 29818
rect 9686 29766 9688 29818
rect 9632 29764 9688 29766
rect 9736 29818 9792 29820
rect 9736 29766 9738 29818
rect 9738 29766 9790 29818
rect 9790 29766 9792 29818
rect 9736 29764 9792 29766
rect 5370 29034 5426 29036
rect 5370 28982 5372 29034
rect 5372 28982 5424 29034
rect 5424 28982 5426 29034
rect 5370 28980 5426 28982
rect 5474 29034 5530 29036
rect 5474 28982 5476 29034
rect 5476 28982 5528 29034
rect 5528 28982 5530 29034
rect 5474 28980 5530 28982
rect 5578 29034 5634 29036
rect 5578 28982 5580 29034
rect 5580 28982 5632 29034
rect 5632 28982 5634 29034
rect 5578 28980 5634 28982
rect 11788 29932 11844 29988
rect 12124 29260 12180 29316
rect 13692 29932 13748 29988
rect 12348 29260 12404 29316
rect 12684 29389 12686 29428
rect 12686 29389 12738 29428
rect 12738 29389 12740 29428
rect 12684 29372 12740 29389
rect 9528 28250 9584 28252
rect 9528 28198 9530 28250
rect 9530 28198 9582 28250
rect 9582 28198 9584 28250
rect 9528 28196 9584 28198
rect 9632 28250 9688 28252
rect 9632 28198 9634 28250
rect 9634 28198 9686 28250
rect 9686 28198 9688 28250
rect 9632 28196 9688 28198
rect 9736 28250 9792 28252
rect 9736 28198 9738 28250
rect 9738 28198 9790 28250
rect 9790 28198 9792 28250
rect 9736 28196 9792 28198
rect 5370 27466 5426 27468
rect 5370 27414 5372 27466
rect 5372 27414 5424 27466
rect 5424 27414 5426 27466
rect 5370 27412 5426 27414
rect 5474 27466 5530 27468
rect 5474 27414 5476 27466
rect 5476 27414 5528 27466
rect 5528 27414 5530 27466
rect 5474 27412 5530 27414
rect 5578 27466 5634 27468
rect 5578 27414 5580 27466
rect 5580 27414 5632 27466
rect 5632 27414 5634 27466
rect 5578 27412 5634 27414
rect 6076 26908 6132 26964
rect 5796 26850 5852 26852
rect 5796 26798 5798 26850
rect 5798 26798 5850 26850
rect 5850 26798 5852 26850
rect 5796 26796 5852 26798
rect 1596 25228 1652 25284
rect 4620 26236 4676 26292
rect 3052 26178 3108 26180
rect 3052 26126 3054 26178
rect 3054 26126 3106 26178
rect 3106 26126 3108 26178
rect 3052 26124 3108 26126
rect 2268 25228 2324 25284
rect 5292 26290 5348 26292
rect 5292 26238 5294 26290
rect 5294 26238 5346 26290
rect 5346 26238 5348 26290
rect 5292 26236 5348 26238
rect 5796 26236 5852 26292
rect 4844 26124 4900 26180
rect 4620 25228 4676 25284
rect 3052 24108 3108 24164
rect 4396 24780 4452 24836
rect 3388 22428 3444 22484
rect 3612 23436 3668 23492
rect 3052 22370 3108 22372
rect 3052 22318 3054 22370
rect 3054 22318 3106 22370
rect 3106 22318 3108 22370
rect 3052 22316 3108 22318
rect 3948 23548 4004 23604
rect 3836 23436 3892 23492
rect 5370 25898 5426 25900
rect 5370 25846 5372 25898
rect 5372 25846 5424 25898
rect 5424 25846 5426 25898
rect 5370 25844 5426 25846
rect 5474 25898 5530 25900
rect 5474 25846 5476 25898
rect 5476 25846 5528 25898
rect 5528 25846 5530 25898
rect 5474 25844 5530 25846
rect 5578 25898 5634 25900
rect 5578 25846 5580 25898
rect 5580 25846 5632 25898
rect 5632 25846 5634 25898
rect 5578 25844 5634 25846
rect 6972 26962 7028 26964
rect 6972 26910 6974 26962
rect 6974 26910 7026 26962
rect 7026 26910 7028 26962
rect 6972 26908 7028 26910
rect 6748 25788 6804 25844
rect 6524 25564 6580 25620
rect 4956 24668 5012 24724
rect 5068 25004 5124 25060
rect 7420 25676 7476 25732
rect 7532 26796 7588 26852
rect 6860 25564 6916 25620
rect 5180 24892 5236 24948
rect 5068 24780 5124 24836
rect 6748 25116 6804 25172
rect 6244 24780 6300 24836
rect 6524 24892 6580 24948
rect 4340 24162 4396 24164
rect 4340 24110 4342 24162
rect 4342 24110 4394 24162
rect 4394 24110 4396 24162
rect 4340 24108 4396 24110
rect 4396 23772 4452 23828
rect 4284 23266 4340 23268
rect 4284 23214 4286 23266
rect 4286 23214 4338 23266
rect 4338 23214 4340 23266
rect 4284 23212 4340 23214
rect 4172 22988 4228 23044
rect 4060 22428 4116 22484
rect 4900 23996 4956 24052
rect 4620 23938 4676 23940
rect 4620 23886 4622 23938
rect 4622 23886 4674 23938
rect 4674 23886 4676 23938
rect 4620 23884 4676 23886
rect 4732 23826 4788 23828
rect 4732 23774 4734 23826
rect 4734 23774 4786 23826
rect 4786 23774 4788 23826
rect 4732 23772 4788 23774
rect 4732 23548 4788 23604
rect 6300 24556 6356 24612
rect 5370 24330 5426 24332
rect 5370 24278 5372 24330
rect 5372 24278 5424 24330
rect 5424 24278 5426 24330
rect 5370 24276 5426 24278
rect 5474 24330 5530 24332
rect 5474 24278 5476 24330
rect 5476 24278 5528 24330
rect 5528 24278 5530 24330
rect 5474 24276 5530 24278
rect 5578 24330 5634 24332
rect 5578 24278 5580 24330
rect 5580 24278 5632 24330
rect 5632 24278 5634 24330
rect 5578 24276 5634 24278
rect 5796 23938 5852 23940
rect 5796 23886 5798 23938
rect 5798 23886 5850 23938
rect 5850 23886 5852 23938
rect 5796 23884 5852 23886
rect 6636 24722 6692 24724
rect 6636 24670 6638 24722
rect 6638 24670 6690 24722
rect 6690 24670 6692 24722
rect 6636 24668 6692 24670
rect 6300 23772 6356 23828
rect 6076 23660 6132 23716
rect 7308 25228 7364 25284
rect 7980 26236 8036 26292
rect 7532 25452 7588 25508
rect 9528 26682 9584 26684
rect 9528 26630 9530 26682
rect 9530 26630 9582 26682
rect 9582 26630 9584 26682
rect 9528 26628 9584 26630
rect 9632 26682 9688 26684
rect 9632 26630 9634 26682
rect 9634 26630 9686 26682
rect 9686 26630 9688 26682
rect 9632 26628 9688 26630
rect 9736 26682 9792 26684
rect 9736 26630 9738 26682
rect 9738 26630 9790 26682
rect 9790 26630 9792 26682
rect 9736 26628 9792 26630
rect 12908 29260 12964 29316
rect 13356 29260 13412 29316
rect 13244 29148 13300 29204
rect 11452 27858 11508 27860
rect 11452 27806 11454 27858
rect 11454 27806 11506 27858
rect 11506 27806 11508 27858
rect 11452 27804 11508 27806
rect 7812 25730 7868 25732
rect 7812 25678 7814 25730
rect 7814 25678 7866 25730
rect 7866 25678 7868 25730
rect 7812 25676 7868 25678
rect 8204 26012 8260 26068
rect 8652 25788 8708 25844
rect 7980 25228 8036 25284
rect 8372 25228 8428 25284
rect 7532 24780 7588 24836
rect 7700 24780 7756 24836
rect 7140 24220 7196 24276
rect 7140 23996 7196 24052
rect 6860 23938 6916 23940
rect 6860 23886 6862 23938
rect 6862 23886 6914 23938
rect 6914 23886 6916 23938
rect 6860 23884 6916 23886
rect 6860 23660 6916 23716
rect 5180 23548 5236 23604
rect 6300 23548 6356 23604
rect 4844 23100 4900 23156
rect 5608 23212 5664 23268
rect 6636 23212 6692 23268
rect 6412 23100 6468 23156
rect 5852 22930 5908 22932
rect 5852 22878 5854 22930
rect 5854 22878 5906 22930
rect 5906 22878 5908 22930
rect 5852 22876 5908 22878
rect 5370 22762 5426 22764
rect 5370 22710 5372 22762
rect 5372 22710 5424 22762
rect 5424 22710 5426 22762
rect 5370 22708 5426 22710
rect 5474 22762 5530 22764
rect 5474 22710 5476 22762
rect 5476 22710 5528 22762
rect 5528 22710 5530 22762
rect 5474 22708 5530 22710
rect 5578 22762 5634 22764
rect 5578 22710 5580 22762
rect 5580 22710 5632 22762
rect 5632 22710 5634 22762
rect 5578 22708 5634 22710
rect 4452 22370 4508 22372
rect 4452 22318 4454 22370
rect 4454 22318 4506 22370
rect 4506 22318 4508 22370
rect 4452 22316 4508 22318
rect 3612 21532 3668 21588
rect 3668 20914 3724 20916
rect 3668 20862 3670 20914
rect 3670 20862 3722 20914
rect 3722 20862 3724 20914
rect 3668 20860 3724 20862
rect 2828 20076 2884 20132
rect 3612 20076 3668 20132
rect 2604 18396 2660 18452
rect 3276 18844 3332 18900
rect 3388 18284 3444 18340
rect 3724 19852 3780 19908
rect 4060 21532 4116 21588
rect 4172 20860 4228 20916
rect 3948 20636 4004 20692
rect 3966 20018 4022 20020
rect 3966 19966 3968 20018
rect 3968 19966 4020 20018
rect 4020 19966 4022 20018
rect 3966 19964 4022 19966
rect 4844 21586 4900 21588
rect 4844 21534 4846 21586
rect 4846 21534 4898 21586
rect 4898 21534 4900 21586
rect 4844 21532 4900 21534
rect 5370 21194 5426 21196
rect 5370 21142 5372 21194
rect 5372 21142 5424 21194
rect 5424 21142 5426 21194
rect 5370 21140 5426 21142
rect 5474 21194 5530 21196
rect 5474 21142 5476 21194
rect 5476 21142 5528 21194
rect 5528 21142 5530 21194
rect 5474 21140 5530 21142
rect 5578 21194 5634 21196
rect 5578 21142 5580 21194
rect 5580 21142 5632 21194
rect 5632 21142 5634 21194
rect 5578 21140 5634 21142
rect 6748 23042 6804 23044
rect 6748 22990 6750 23042
rect 6750 22990 6802 23042
rect 6802 22990 6804 23042
rect 6748 22988 6804 22990
rect 5012 20972 5068 21028
rect 5628 20972 5684 21028
rect 6860 22540 6916 22596
rect 5964 20802 6020 20804
rect 5964 20750 5966 20802
rect 5966 20750 6018 20802
rect 6018 20750 6020 20802
rect 5964 20748 6020 20750
rect 4508 20300 4564 20356
rect 5796 20300 5852 20356
rect 5516 20076 5572 20132
rect 4284 19964 4340 20020
rect 4732 20018 4788 20020
rect 4732 19966 4734 20018
rect 4734 19966 4786 20018
rect 4786 19966 4788 20018
rect 4732 19964 4788 19966
rect 4508 19852 4564 19908
rect 5852 20018 5908 20020
rect 5852 19966 5854 20018
rect 5854 19966 5906 20018
rect 5906 19966 5908 20018
rect 5852 19964 5908 19966
rect 5370 19626 5426 19628
rect 5370 19574 5372 19626
rect 5372 19574 5424 19626
rect 5424 19574 5426 19626
rect 5370 19572 5426 19574
rect 5474 19626 5530 19628
rect 5474 19574 5476 19626
rect 5476 19574 5528 19626
rect 5528 19574 5530 19626
rect 5474 19572 5530 19574
rect 5578 19626 5634 19628
rect 5578 19574 5580 19626
rect 5580 19574 5632 19626
rect 5632 19574 5634 19626
rect 5578 19572 5634 19574
rect 3612 17836 3668 17892
rect 3836 18732 3892 18788
rect 3948 18844 4004 18900
rect 4060 18450 4116 18452
rect 4060 18398 4062 18450
rect 4062 18398 4114 18450
rect 4114 18398 4116 18450
rect 4060 18396 4116 18398
rect 4060 18172 4116 18228
rect 4060 17836 4116 17892
rect 4508 18284 4564 18340
rect 4396 17836 4452 17892
rect 4284 17666 4340 17668
rect 4284 17614 4286 17666
rect 4286 17614 4338 17666
rect 4338 17614 4340 17666
rect 4284 17612 4340 17614
rect 7868 23772 7924 23828
rect 8428 24780 8484 24836
rect 8260 24722 8316 24724
rect 8260 24670 8262 24722
rect 8262 24670 8314 24722
rect 8314 24670 8316 24722
rect 8260 24668 8316 24670
rect 8316 24108 8372 24164
rect 8204 23996 8260 24052
rect 7532 23100 7588 23156
rect 8876 26290 8932 26292
rect 8876 26238 8878 26290
rect 8878 26238 8930 26290
rect 8930 26238 8932 26290
rect 8876 26236 8932 26238
rect 9660 26253 9662 26292
rect 9662 26253 9714 26292
rect 9714 26253 9716 26292
rect 9660 26236 9716 26253
rect 8764 25676 8820 25732
rect 8764 25506 8820 25508
rect 8764 25454 8766 25506
rect 8766 25454 8818 25506
rect 8818 25454 8820 25506
rect 8764 25452 8820 25454
rect 9212 24220 9268 24276
rect 8540 23660 8596 23716
rect 8876 23772 8932 23828
rect 7532 22876 7588 22932
rect 8484 22988 8540 23044
rect 7924 22930 7980 22932
rect 7924 22878 7926 22930
rect 7926 22878 7978 22930
rect 7978 22878 7980 22930
rect 7924 22876 7980 22878
rect 8428 22764 8484 22820
rect 7868 22428 7924 22484
rect 8092 22370 8148 22372
rect 8092 22318 8094 22370
rect 8094 22318 8146 22370
rect 8146 22318 8148 22370
rect 8092 22316 8148 22318
rect 8652 22652 8708 22708
rect 8988 22764 9044 22820
rect 8876 22428 8932 22484
rect 9828 25452 9884 25508
rect 10220 25788 10276 25844
rect 10500 26178 10556 26180
rect 10500 26126 10502 26178
rect 10502 26126 10554 26178
rect 10554 26126 10556 26178
rect 10500 26124 10556 26126
rect 10892 26124 10948 26180
rect 9996 25452 10052 25508
rect 12124 26236 12180 26292
rect 12348 27804 12404 27860
rect 12908 27858 12964 27860
rect 12908 27806 12910 27858
rect 12910 27806 12962 27858
rect 12962 27806 12964 27858
rect 12908 27804 12964 27806
rect 12684 27020 12740 27076
rect 9528 25114 9584 25116
rect 9528 25062 9530 25114
rect 9530 25062 9582 25114
rect 9582 25062 9584 25114
rect 9528 25060 9584 25062
rect 9632 25114 9688 25116
rect 9632 25062 9634 25114
rect 9634 25062 9686 25114
rect 9686 25062 9688 25114
rect 9632 25060 9688 25062
rect 9736 25114 9792 25116
rect 9736 25062 9738 25114
rect 9738 25062 9790 25114
rect 9790 25062 9792 25114
rect 9736 25060 9792 25062
rect 11004 25340 11060 25396
rect 9324 24108 9380 24164
rect 10220 23996 10276 24052
rect 9828 23938 9884 23940
rect 9828 23886 9830 23938
rect 9830 23886 9882 23938
rect 9882 23886 9884 23938
rect 9828 23884 9884 23886
rect 9548 23772 9604 23828
rect 9528 23546 9584 23548
rect 9528 23494 9530 23546
rect 9530 23494 9582 23546
rect 9582 23494 9584 23546
rect 9528 23492 9584 23494
rect 9632 23546 9688 23548
rect 9632 23494 9634 23546
rect 9634 23494 9686 23546
rect 9686 23494 9688 23546
rect 9632 23492 9688 23494
rect 9736 23546 9792 23548
rect 9736 23494 9738 23546
rect 9738 23494 9790 23546
rect 9790 23494 9792 23546
rect 9736 23492 9792 23494
rect 9324 22876 9380 22932
rect 8540 22370 8596 22372
rect 8540 22318 8542 22370
rect 8542 22318 8594 22370
rect 8594 22318 8596 22370
rect 8540 22316 8596 22318
rect 8316 21586 8372 21588
rect 8316 21534 8318 21586
rect 8318 21534 8370 21586
rect 8370 21534 8372 21586
rect 8316 21532 8372 21534
rect 8652 22092 8708 22148
rect 8764 21532 8820 21588
rect 8876 22258 8932 22260
rect 8876 22206 8878 22258
rect 8878 22206 8930 22258
rect 8930 22206 8932 22258
rect 8876 22204 8932 22206
rect 8428 21420 8484 21476
rect 7196 20860 7252 20916
rect 9884 22594 9940 22596
rect 9884 22542 9886 22594
rect 9886 22542 9938 22594
rect 9938 22542 9940 22594
rect 9884 22540 9940 22542
rect 9548 22092 9604 22148
rect 9528 21978 9584 21980
rect 9528 21926 9530 21978
rect 9530 21926 9582 21978
rect 9582 21926 9584 21978
rect 9528 21924 9584 21926
rect 9632 21978 9688 21980
rect 9632 21926 9634 21978
rect 9634 21926 9686 21978
rect 9686 21926 9688 21978
rect 9632 21924 9688 21926
rect 9736 21978 9792 21980
rect 9736 21926 9738 21978
rect 9738 21926 9790 21978
rect 9790 21926 9792 21978
rect 9736 21924 9792 21926
rect 9044 21474 9100 21476
rect 9044 21422 9046 21474
rect 9046 21422 9098 21474
rect 9098 21422 9100 21474
rect 9044 21420 9100 21422
rect 7084 20076 7140 20132
rect 4956 19180 5012 19236
rect 4900 18732 4956 18788
rect 5292 18284 5348 18340
rect 6416 18844 6472 18900
rect 6412 18620 6468 18676
rect 6300 18508 6356 18564
rect 5740 18284 5796 18340
rect 5370 18058 5426 18060
rect 5370 18006 5372 18058
rect 5372 18006 5424 18058
rect 5424 18006 5426 18058
rect 5370 18004 5426 18006
rect 5474 18058 5530 18060
rect 5474 18006 5476 18058
rect 5476 18006 5528 18058
rect 5528 18006 5530 18058
rect 5474 18004 5530 18006
rect 5578 18058 5634 18060
rect 5578 18006 5580 18058
rect 5580 18006 5632 18058
rect 5632 18006 5634 18058
rect 5578 18004 5634 18006
rect 5964 17836 6020 17892
rect 4172 17500 4228 17556
rect 3948 17276 4004 17332
rect 4172 16882 4228 16884
rect 4172 16830 4174 16882
rect 4174 16830 4226 16882
rect 4226 16830 4228 16882
rect 4172 16828 4228 16830
rect 1820 16098 1876 16100
rect 1820 16046 1822 16098
rect 1822 16046 1874 16098
rect 1874 16046 1876 16098
rect 1820 16044 1876 16046
rect 4508 16882 4564 16884
rect 4508 16830 4510 16882
rect 4510 16830 4562 16882
rect 4562 16830 4564 16882
rect 4508 16828 4564 16830
rect 5740 17666 5796 17668
rect 5740 17614 5742 17666
rect 5742 17614 5794 17666
rect 5794 17614 5796 17666
rect 5740 17612 5796 17614
rect 7196 19292 7252 19348
rect 7532 20018 7588 20020
rect 7532 19966 7534 20018
rect 7534 19966 7586 20018
rect 7586 19966 7588 20018
rect 7532 19964 7588 19966
rect 7308 19234 7364 19236
rect 7308 19182 7310 19234
rect 7310 19182 7362 19234
rect 7362 19182 7364 19234
rect 7308 19180 7364 19182
rect 7196 18732 7252 18788
rect 7084 18562 7140 18564
rect 7084 18510 7086 18562
rect 7086 18510 7138 18562
rect 7138 18510 7140 18562
rect 7084 18508 7140 18510
rect 6300 17612 6356 17668
rect 4956 17500 5012 17556
rect 7756 18450 7812 18452
rect 7756 18398 7758 18450
rect 7758 18398 7810 18450
rect 7810 18398 7812 18450
rect 7756 18396 7812 18398
rect 7644 18172 7700 18228
rect 7644 17724 7700 17780
rect 6972 17500 7028 17556
rect 7998 18338 8054 18340
rect 7998 18286 8000 18338
rect 8000 18286 8052 18338
rect 8052 18286 8054 18338
rect 7998 18284 8054 18286
rect 7756 17612 7812 17668
rect 8092 17724 8148 17780
rect 7308 17388 7364 17444
rect 7812 17442 7868 17444
rect 7812 17390 7814 17442
rect 7814 17390 7866 17442
rect 7866 17390 7868 17442
rect 7812 17388 7868 17390
rect 8820 20018 8876 20020
rect 8820 19966 8822 20018
rect 8822 19966 8874 20018
rect 8874 19966 8876 20018
rect 8820 19964 8876 19966
rect 8540 19292 8596 19348
rect 8428 18844 8484 18900
rect 8540 18620 8596 18676
rect 8428 18450 8484 18452
rect 8428 18398 8430 18450
rect 8430 18398 8482 18450
rect 8482 18398 8484 18450
rect 8428 18396 8484 18398
rect 8316 17724 8372 17780
rect 9212 20748 9268 20804
rect 9528 20410 9584 20412
rect 9528 20358 9530 20410
rect 9530 20358 9582 20410
rect 9582 20358 9584 20410
rect 9528 20356 9584 20358
rect 9632 20410 9688 20412
rect 9632 20358 9634 20410
rect 9634 20358 9686 20410
rect 9686 20358 9688 20410
rect 9632 20356 9688 20358
rect 9736 20410 9792 20412
rect 9736 20358 9738 20410
rect 9738 20358 9790 20410
rect 9790 20358 9792 20410
rect 9736 20356 9792 20358
rect 9436 20018 9492 20020
rect 9436 19966 9438 20018
rect 9438 19966 9490 20018
rect 9490 19966 9492 20018
rect 9436 19964 9492 19966
rect 10892 23996 10948 24052
rect 11116 24892 11172 24948
rect 12012 24780 12068 24836
rect 11676 24668 11732 24724
rect 11844 23996 11900 24052
rect 11228 23910 11284 23940
rect 11228 23884 11230 23910
rect 11230 23884 11282 23910
rect 11282 23884 11284 23910
rect 11564 23884 11620 23940
rect 12292 26066 12348 26068
rect 12292 26014 12294 26066
rect 12294 26014 12346 26066
rect 12346 26014 12348 26066
rect 12292 26012 12348 26014
rect 12684 26290 12740 26292
rect 12684 26238 12686 26290
rect 12686 26238 12738 26290
rect 12738 26238 12740 26290
rect 12684 26236 12740 26238
rect 13468 29426 13524 29428
rect 13468 29374 13470 29426
rect 13470 29374 13522 29426
rect 13522 29374 13524 29426
rect 13468 29372 13524 29374
rect 13748 29202 13804 29204
rect 13748 29150 13750 29202
rect 13750 29150 13802 29202
rect 13802 29150 13804 29202
rect 13748 29148 13804 29150
rect 13686 29034 13742 29036
rect 13686 28982 13688 29034
rect 13688 28982 13740 29034
rect 13740 28982 13742 29034
rect 13686 28980 13742 28982
rect 13790 29034 13846 29036
rect 13790 28982 13792 29034
rect 13792 28982 13844 29034
rect 13844 28982 13846 29034
rect 13790 28980 13846 28982
rect 13894 29034 13950 29036
rect 13894 28982 13896 29034
rect 13896 28982 13948 29034
rect 13948 28982 13950 29034
rect 13894 28980 13950 28982
rect 13356 28588 13412 28644
rect 13636 28642 13692 28644
rect 13636 28590 13638 28642
rect 13638 28590 13690 28642
rect 13690 28590 13692 28642
rect 13636 28588 13692 28590
rect 13916 28812 13972 28868
rect 13468 28476 13524 28532
rect 13244 27804 13300 27860
rect 15820 31554 15876 31556
rect 15820 31502 15822 31554
rect 15822 31502 15874 31554
rect 15874 31502 15876 31554
rect 15820 31500 15876 31502
rect 14700 30044 14756 30100
rect 14644 29538 14700 29540
rect 14644 29486 14646 29538
rect 14646 29486 14698 29538
rect 14698 29486 14700 29538
rect 14644 29484 14700 29486
rect 14252 29426 14308 29428
rect 14252 29374 14254 29426
rect 14254 29374 14306 29426
rect 14306 29374 14308 29426
rect 14252 29372 14308 29374
rect 14364 29148 14420 29204
rect 15708 29932 15764 29988
rect 17844 31386 17900 31388
rect 17844 31334 17846 31386
rect 17846 31334 17898 31386
rect 17898 31334 17900 31386
rect 17844 31332 17900 31334
rect 17948 31386 18004 31388
rect 17948 31334 17950 31386
rect 17950 31334 18002 31386
rect 18002 31334 18004 31386
rect 17948 31332 18004 31334
rect 18052 31386 18108 31388
rect 18052 31334 18054 31386
rect 18054 31334 18106 31386
rect 18106 31334 18108 31386
rect 18052 31332 18108 31334
rect 15932 29484 15988 29540
rect 16828 30210 16884 30212
rect 16828 30158 16830 30210
rect 16830 30158 16882 30210
rect 16882 30158 16884 30210
rect 16828 30156 16884 30158
rect 16380 29596 16436 29652
rect 14812 29148 14868 29204
rect 15428 29372 15484 29428
rect 14364 28700 14420 28756
rect 13686 27466 13742 27468
rect 13686 27414 13688 27466
rect 13688 27414 13740 27466
rect 13740 27414 13742 27466
rect 13686 27412 13742 27414
rect 13790 27466 13846 27468
rect 13790 27414 13792 27466
rect 13792 27414 13844 27466
rect 13844 27414 13846 27466
rect 13790 27412 13846 27414
rect 13894 27466 13950 27468
rect 13894 27414 13896 27466
rect 13896 27414 13948 27466
rect 13948 27414 13950 27466
rect 13894 27412 13950 27414
rect 14028 27074 14084 27076
rect 14028 27022 14030 27074
rect 14030 27022 14082 27074
rect 14082 27022 14084 27074
rect 14028 27020 14084 27022
rect 14476 27020 14532 27076
rect 14252 26236 14308 26292
rect 13188 26178 13244 26180
rect 13188 26126 13190 26178
rect 13190 26126 13242 26178
rect 13242 26126 13244 26178
rect 13188 26124 13244 26126
rect 13686 25898 13742 25900
rect 13686 25846 13688 25898
rect 13688 25846 13740 25898
rect 13740 25846 13742 25898
rect 13686 25844 13742 25846
rect 13790 25898 13846 25900
rect 13790 25846 13792 25898
rect 13792 25846 13844 25898
rect 13844 25846 13846 25898
rect 13790 25844 13846 25846
rect 13894 25898 13950 25900
rect 13894 25846 13896 25898
rect 13896 25846 13948 25898
rect 13948 25846 13950 25898
rect 13894 25844 13950 25846
rect 13692 25564 13748 25620
rect 13524 25452 13580 25508
rect 12572 25340 12628 25396
rect 12236 24220 12292 24276
rect 12460 24722 12516 24724
rect 12460 24670 12462 24722
rect 12462 24670 12514 24722
rect 12514 24670 12516 24722
rect 12460 24668 12516 24670
rect 13468 25116 13524 25172
rect 12740 24892 12796 24948
rect 12908 24780 12964 24836
rect 12348 23996 12404 24052
rect 10948 22146 11004 22148
rect 10948 22094 10950 22146
rect 10950 22094 11002 22146
rect 11002 22094 11004 22146
rect 10948 22092 11004 22094
rect 11788 22204 11844 22260
rect 11564 22092 11620 22148
rect 12236 23938 12292 23940
rect 12236 23886 12238 23938
rect 12238 23886 12290 23938
rect 12290 23886 12292 23938
rect 12236 23884 12292 23886
rect 12402 23324 12458 23380
rect 12684 23324 12740 23380
rect 12068 22594 12124 22596
rect 12068 22542 12070 22594
rect 12070 22542 12122 22594
rect 12122 22542 12124 22594
rect 12068 22540 12124 22542
rect 12236 22428 12292 22484
rect 12460 22652 12516 22708
rect 12124 22204 12180 22260
rect 11564 21420 11620 21476
rect 12796 23154 12852 23156
rect 12796 23102 12798 23154
rect 12798 23102 12850 23154
rect 12850 23102 12852 23154
rect 12796 23100 12852 23102
rect 12796 22482 12852 22484
rect 12796 22430 12798 22482
rect 12798 22430 12850 22482
rect 12850 22430 12852 22482
rect 12796 22428 12852 22430
rect 12796 21532 12852 21588
rect 11788 20802 11844 20804
rect 11788 20750 11790 20802
rect 11790 20750 11842 20802
rect 11842 20750 11844 20802
rect 11788 20748 11844 20750
rect 10332 19964 10388 20020
rect 11564 19852 11620 19908
rect 12516 20412 12572 20468
rect 12796 20412 12852 20468
rect 13244 24780 13300 24836
rect 14140 25116 14196 25172
rect 13692 25004 13748 25060
rect 15428 28700 15484 28756
rect 15708 28812 15764 28868
rect 15820 28642 15876 28644
rect 15820 28590 15822 28642
rect 15822 28590 15874 28642
rect 15874 28590 15876 28642
rect 15820 28588 15876 28590
rect 16268 29426 16324 29428
rect 16268 29374 16270 29426
rect 16270 29374 16322 29426
rect 16322 29374 16324 29426
rect 16268 29372 16324 29374
rect 17724 30210 17780 30212
rect 17724 30158 17726 30210
rect 17726 30158 17778 30210
rect 17778 30158 17780 30210
rect 17724 30156 17780 30158
rect 18060 30210 18116 30212
rect 18060 30158 18062 30210
rect 18062 30158 18114 30210
rect 18114 30158 18116 30210
rect 18060 30156 18116 30158
rect 17332 29596 17388 29652
rect 26160 31386 26216 31388
rect 26160 31334 26162 31386
rect 26162 31334 26214 31386
rect 26214 31334 26216 31386
rect 26160 31332 26216 31334
rect 26264 31386 26320 31388
rect 26264 31334 26266 31386
rect 26266 31334 26318 31386
rect 26318 31334 26320 31386
rect 26264 31332 26320 31334
rect 26368 31386 26424 31388
rect 26368 31334 26370 31386
rect 26370 31334 26422 31386
rect 26422 31334 26424 31386
rect 26368 31332 26424 31334
rect 34476 31386 34532 31388
rect 34476 31334 34478 31386
rect 34478 31334 34530 31386
rect 34530 31334 34532 31386
rect 34476 31332 34532 31334
rect 34580 31386 34636 31388
rect 34580 31334 34582 31386
rect 34582 31334 34634 31386
rect 34634 31334 34636 31386
rect 34580 31332 34636 31334
rect 34684 31386 34740 31388
rect 34684 31334 34686 31386
rect 34686 31334 34738 31386
rect 34738 31334 34740 31386
rect 34684 31332 34740 31334
rect 20860 30268 20916 30324
rect 18620 30156 18676 30212
rect 18956 30156 19012 30212
rect 20300 30210 20356 30212
rect 18508 29932 18564 29988
rect 17052 29484 17108 29540
rect 16828 29372 16884 29428
rect 16716 28588 16772 28644
rect 17844 29818 17900 29820
rect 17844 29766 17846 29818
rect 17846 29766 17898 29818
rect 17898 29766 17900 29818
rect 17844 29764 17900 29766
rect 17948 29818 18004 29820
rect 17948 29766 17950 29818
rect 17950 29766 18002 29818
rect 18002 29766 18004 29818
rect 17948 29764 18004 29766
rect 18052 29818 18108 29820
rect 18052 29766 18054 29818
rect 18054 29766 18106 29818
rect 18106 29766 18108 29818
rect 18052 29764 18108 29766
rect 18396 29596 18452 29652
rect 20300 30158 20302 30210
rect 20302 30158 20354 30210
rect 20354 30158 20356 30210
rect 20300 30156 20356 30158
rect 20636 30098 20692 30100
rect 20636 30046 20638 30098
rect 20638 30046 20690 30098
rect 20690 30046 20692 30098
rect 20636 30044 20692 30046
rect 19516 29484 19572 29540
rect 18508 29314 18564 29316
rect 18508 29262 18510 29314
rect 18510 29262 18562 29314
rect 18562 29262 18564 29314
rect 18508 29260 18564 29262
rect 18172 29148 18228 29204
rect 16716 27074 16772 27076
rect 16716 27022 16718 27074
rect 16718 27022 16770 27074
rect 16770 27022 16772 27074
rect 16716 27020 16772 27022
rect 19740 29484 19796 29540
rect 20188 29596 20244 29652
rect 19628 29372 19684 29428
rect 19180 29260 19236 29316
rect 20468 29538 20524 29540
rect 20468 29486 20470 29538
rect 20470 29486 20522 29538
rect 20522 29486 20524 29538
rect 20468 29484 20524 29486
rect 20748 29426 20804 29428
rect 20748 29374 20750 29426
rect 20750 29374 20802 29426
rect 20802 29374 20804 29426
rect 20748 29372 20804 29374
rect 19964 29148 20020 29204
rect 20076 28754 20132 28756
rect 20076 28702 20078 28754
rect 20078 28702 20130 28754
rect 20130 28702 20132 28754
rect 20076 28700 20132 28702
rect 21308 30268 21364 30324
rect 22652 30882 22708 30884
rect 22652 30830 22654 30882
rect 22654 30830 22706 30882
rect 22706 30830 22708 30882
rect 22652 30828 22708 30830
rect 22002 30602 22058 30604
rect 22002 30550 22004 30602
rect 22004 30550 22056 30602
rect 22056 30550 22058 30602
rect 22002 30548 22058 30550
rect 22106 30602 22162 30604
rect 22106 30550 22108 30602
rect 22108 30550 22160 30602
rect 22160 30550 22162 30602
rect 22106 30548 22162 30550
rect 22210 30602 22266 30604
rect 22210 30550 22212 30602
rect 22212 30550 22264 30602
rect 22264 30550 22266 30602
rect 22210 30548 22266 30550
rect 21644 30268 21700 30324
rect 22002 29034 22058 29036
rect 22002 28982 22004 29034
rect 22004 28982 22056 29034
rect 22056 28982 22058 29034
rect 22002 28980 22058 28982
rect 22106 29034 22162 29036
rect 22106 28982 22108 29034
rect 22108 28982 22160 29034
rect 22160 28982 22162 29034
rect 22106 28980 22162 28982
rect 22210 29034 22266 29036
rect 22210 28982 22212 29034
rect 22212 28982 22264 29034
rect 22264 28982 22266 29034
rect 22210 28980 22266 28982
rect 24332 30156 24388 30212
rect 23996 30044 24052 30100
rect 22876 29932 22932 29988
rect 22652 29426 22708 29428
rect 22652 29374 22654 29426
rect 22654 29374 22706 29426
rect 22706 29374 22708 29426
rect 23324 29484 23380 29540
rect 22652 29372 22708 29374
rect 22988 29314 23044 29316
rect 22988 29262 22990 29314
rect 22990 29262 23042 29314
rect 23042 29262 23044 29314
rect 22988 29260 23044 29262
rect 21084 28700 21140 28756
rect 17844 28250 17900 28252
rect 17844 28198 17846 28250
rect 17846 28198 17898 28250
rect 17898 28198 17900 28250
rect 17844 28196 17900 28198
rect 17948 28250 18004 28252
rect 17948 28198 17950 28250
rect 17950 28198 18002 28250
rect 18002 28198 18004 28250
rect 17948 28196 18004 28198
rect 18052 28250 18108 28252
rect 18052 28198 18054 28250
rect 18054 28198 18106 28250
rect 18106 28198 18108 28250
rect 18052 28196 18108 28198
rect 17500 27059 17556 27076
rect 17500 27020 17502 27059
rect 17502 27020 17554 27059
rect 17554 27020 17556 27059
rect 14700 25564 14756 25620
rect 15260 25676 15316 25732
rect 14476 25506 14532 25508
rect 14476 25454 14478 25506
rect 14478 25454 14530 25506
rect 14530 25454 14532 25506
rect 14476 25452 14532 25454
rect 14588 25340 14644 25396
rect 15596 25618 15652 25620
rect 15596 25566 15598 25618
rect 15598 25566 15650 25618
rect 15650 25566 15652 25618
rect 15596 25564 15652 25566
rect 15260 25340 15316 25396
rect 15708 25452 15764 25508
rect 14476 25228 14532 25284
rect 13468 24332 13524 24388
rect 13686 24330 13742 24332
rect 13686 24278 13688 24330
rect 13688 24278 13740 24330
rect 13740 24278 13742 24330
rect 13686 24276 13742 24278
rect 13790 24330 13846 24332
rect 13790 24278 13792 24330
rect 13792 24278 13844 24330
rect 13844 24278 13846 24330
rect 13790 24276 13846 24278
rect 13894 24330 13950 24332
rect 13894 24278 13896 24330
rect 13896 24278 13948 24330
rect 13948 24278 13950 24330
rect 13894 24276 13950 24278
rect 13468 23660 13524 23716
rect 13356 23548 13412 23604
rect 13020 22540 13076 22596
rect 13804 23100 13860 23156
rect 13686 22762 13742 22764
rect 13686 22710 13688 22762
rect 13688 22710 13740 22762
rect 13740 22710 13742 22762
rect 13686 22708 13742 22710
rect 13790 22762 13846 22764
rect 13790 22710 13792 22762
rect 13792 22710 13844 22762
rect 13844 22710 13846 22762
rect 13790 22708 13846 22710
rect 13894 22762 13950 22764
rect 13894 22710 13896 22762
rect 13896 22710 13948 22762
rect 13948 22710 13950 22762
rect 13894 22708 13950 22710
rect 13132 21586 13188 21588
rect 13132 21534 13134 21586
rect 13134 21534 13186 21586
rect 13186 21534 13188 21586
rect 13132 21532 13188 21534
rect 14028 22370 14084 22372
rect 14028 22318 14030 22370
rect 14030 22318 14082 22370
rect 14082 22318 14084 22370
rect 14028 22316 14084 22318
rect 13524 22258 13580 22260
rect 13524 22206 13526 22258
rect 13526 22206 13578 22258
rect 13578 22206 13580 22258
rect 13524 22204 13580 22206
rect 14028 21532 14084 21588
rect 12684 20076 12740 20132
rect 13020 20748 13076 20804
rect 12684 19906 12740 19908
rect 12684 19854 12686 19906
rect 12686 19854 12738 19906
rect 12738 19854 12740 19906
rect 12684 19852 12740 19854
rect 9528 18842 9584 18844
rect 9528 18790 9530 18842
rect 9530 18790 9582 18842
rect 9582 18790 9584 18842
rect 9528 18788 9584 18790
rect 9632 18842 9688 18844
rect 9632 18790 9634 18842
rect 9634 18790 9686 18842
rect 9686 18790 9688 18842
rect 9632 18788 9688 18790
rect 9736 18842 9792 18844
rect 9736 18790 9738 18842
rect 9738 18790 9790 18842
rect 9790 18790 9792 18842
rect 9736 18788 9792 18790
rect 9100 18620 9156 18676
rect 8988 18284 9044 18340
rect 11228 18284 11284 18340
rect 13686 21194 13742 21196
rect 13686 21142 13688 21194
rect 13688 21142 13740 21194
rect 13740 21142 13742 21194
rect 13686 21140 13742 21142
rect 13790 21194 13846 21196
rect 13790 21142 13792 21194
rect 13792 21142 13844 21194
rect 13844 21142 13846 21194
rect 13790 21140 13846 21142
rect 13894 21194 13950 21196
rect 13894 21142 13896 21194
rect 13896 21142 13948 21194
rect 13948 21142 13950 21194
rect 13894 21140 13950 21142
rect 13356 20300 13412 20356
rect 13468 20076 13524 20132
rect 13020 19740 13076 19796
rect 12012 18172 12068 18228
rect 12124 18844 12180 18900
rect 12236 18284 12292 18340
rect 12348 18396 12404 18452
rect 12012 17724 12068 17780
rect 11900 17666 11956 17668
rect 10892 17500 10948 17556
rect 11900 17614 11902 17666
rect 11902 17614 11954 17666
rect 11954 17614 11956 17666
rect 11900 17612 11956 17614
rect 8764 17388 8820 17444
rect 9528 17274 9584 17276
rect 9528 17222 9530 17274
rect 9530 17222 9582 17274
rect 9582 17222 9584 17274
rect 9528 17220 9584 17222
rect 9632 17274 9688 17276
rect 9632 17222 9634 17274
rect 9634 17222 9686 17274
rect 9686 17222 9688 17274
rect 9632 17220 9688 17222
rect 9736 17274 9792 17276
rect 9736 17222 9738 17274
rect 9738 17222 9790 17274
rect 9790 17222 9792 17274
rect 9736 17220 9792 17222
rect 6300 16828 6356 16884
rect 5370 16490 5426 16492
rect 5370 16438 5372 16490
rect 5372 16438 5424 16490
rect 5424 16438 5426 16490
rect 5370 16436 5426 16438
rect 5474 16490 5530 16492
rect 5474 16438 5476 16490
rect 5476 16438 5528 16490
rect 5528 16438 5530 16490
rect 5474 16436 5530 16438
rect 5578 16490 5634 16492
rect 5578 16438 5580 16490
rect 5580 16438 5632 16490
rect 5632 16438 5634 16490
rect 5578 16436 5634 16438
rect 4900 16044 4956 16100
rect 5124 16098 5180 16100
rect 5124 16046 5126 16098
rect 5126 16046 5178 16098
rect 5178 16046 5180 16098
rect 5124 16044 5180 16046
rect 5852 16044 5908 16100
rect 5370 14922 5426 14924
rect 5370 14870 5372 14922
rect 5372 14870 5424 14922
rect 5424 14870 5426 14922
rect 5370 14868 5426 14870
rect 5474 14922 5530 14924
rect 5474 14870 5476 14922
rect 5476 14870 5528 14922
rect 5528 14870 5530 14922
rect 5474 14868 5530 14870
rect 5578 14922 5634 14924
rect 5578 14870 5580 14922
rect 5580 14870 5632 14922
rect 5632 14870 5634 14922
rect 5578 14868 5634 14870
rect 3388 14530 3444 14532
rect 3388 14478 3390 14530
rect 3390 14478 3442 14530
rect 3442 14478 3444 14530
rect 3388 14476 3444 14478
rect 2940 13804 2996 13860
rect 3612 13804 3668 13860
rect 3052 13746 3108 13748
rect 3052 13694 3054 13746
rect 3054 13694 3106 13746
rect 3106 13694 3108 13746
rect 4956 13804 5012 13860
rect 3836 13746 3892 13748
rect 3052 13692 3108 13694
rect 2828 13580 2884 13636
rect 2268 13468 2324 13524
rect 3836 13694 3838 13746
rect 3838 13694 3890 13746
rect 3890 13694 3892 13746
rect 3836 13692 3892 13694
rect 4060 13634 4116 13636
rect 4060 13582 4062 13634
rect 4062 13582 4114 13634
rect 4114 13582 4116 13634
rect 4060 13580 4116 13582
rect 2716 12908 2772 12964
rect 3612 13468 3668 13524
rect 4452 13580 4508 13636
rect 2660 12178 2716 12180
rect 2660 12126 2662 12178
rect 2662 12126 2714 12178
rect 2714 12126 2716 12178
rect 2660 12124 2716 12126
rect 2716 11116 2772 11172
rect 3388 12962 3444 12964
rect 3388 12910 3390 12962
rect 3390 12910 3442 12962
rect 3442 12910 3444 12962
rect 3388 12908 3444 12910
rect 3276 12012 3332 12068
rect 3052 11900 3108 11956
rect 4060 12908 4116 12964
rect 4732 12348 4788 12404
rect 3836 12178 3892 12180
rect 3836 12126 3838 12178
rect 3838 12126 3890 12178
rect 3890 12126 3892 12178
rect 3836 12124 3892 12126
rect 4284 12124 4340 12180
rect 3836 11788 3892 11844
rect 3220 11170 3276 11172
rect 3220 11118 3222 11170
rect 3222 11118 3274 11170
rect 3274 11118 3276 11170
rect 3220 11116 3276 11118
rect 3724 11004 3780 11060
rect 3052 10610 3108 10612
rect 3052 10558 3054 10610
rect 3054 10558 3106 10610
rect 3106 10558 3108 10610
rect 3052 10556 3108 10558
rect 3612 10108 3668 10164
rect 2716 9772 2772 9828
rect 3276 9660 3332 9716
rect 3052 9548 3108 9604
rect 2492 8092 2548 8148
rect 2492 5682 2548 5684
rect 2492 5630 2494 5682
rect 2494 5630 2546 5682
rect 2546 5630 2548 5682
rect 2492 5628 2548 5630
rect 2604 7420 2660 7476
rect 3836 10332 3892 10388
rect 4284 11116 4340 11172
rect 4508 12178 4564 12180
rect 4508 12126 4510 12178
rect 4510 12126 4562 12178
rect 4562 12126 4564 12178
rect 4508 12124 4564 12126
rect 5370 13354 5426 13356
rect 5370 13302 5372 13354
rect 5372 13302 5424 13354
rect 5424 13302 5426 13354
rect 5370 13300 5426 13302
rect 5474 13354 5530 13356
rect 5474 13302 5476 13354
rect 5476 13302 5528 13354
rect 5528 13302 5530 13354
rect 5474 13300 5530 13302
rect 5578 13354 5634 13356
rect 5578 13302 5580 13354
rect 5580 13302 5632 13354
rect 5632 13302 5634 13354
rect 5578 13300 5634 13302
rect 5740 13020 5796 13076
rect 5068 12796 5124 12852
rect 8540 16716 8596 16772
rect 10444 16828 10500 16884
rect 9436 16716 9492 16772
rect 11340 16828 11396 16884
rect 7868 16098 7924 16100
rect 7868 16046 7870 16098
rect 7870 16046 7922 16098
rect 7922 16046 7924 16098
rect 7868 16044 7924 16046
rect 8540 16044 8596 16100
rect 7980 15260 8036 15316
rect 6188 14700 6244 14756
rect 6748 14754 6804 14756
rect 6748 14702 6750 14754
rect 6750 14702 6802 14754
rect 6802 14702 6804 14754
rect 6748 14700 6804 14702
rect 7308 14754 7364 14756
rect 7308 14702 7310 14754
rect 7310 14702 7362 14754
rect 7362 14702 7364 14754
rect 7308 14700 7364 14702
rect 7084 13580 7140 13636
rect 5964 12962 6020 12964
rect 5964 12910 5966 12962
rect 5966 12910 6018 12962
rect 6018 12910 6020 12962
rect 5964 12908 6020 12910
rect 6300 12908 6356 12964
rect 6972 12934 7028 12964
rect 5516 12460 5572 12516
rect 3948 9996 4004 10052
rect 3836 9798 3892 9828
rect 3836 9772 3838 9798
rect 3838 9772 3890 9798
rect 3890 9772 3892 9798
rect 3724 9548 3780 9604
rect 3668 9100 3724 9156
rect 3052 8428 3108 8484
rect 3052 8092 3108 8148
rect 3892 8316 3948 8372
rect 4172 8428 4228 8484
rect 4508 11340 4564 11396
rect 4732 11228 4788 11284
rect 4956 11004 5012 11060
rect 5068 11900 5124 11956
rect 5180 11788 5236 11844
rect 5370 11786 5426 11788
rect 5370 11734 5372 11786
rect 5372 11734 5424 11786
rect 5424 11734 5426 11786
rect 5370 11732 5426 11734
rect 5474 11786 5530 11788
rect 5474 11734 5476 11786
rect 5476 11734 5528 11786
rect 5528 11734 5530 11786
rect 5474 11732 5530 11734
rect 5578 11786 5634 11788
rect 5578 11734 5580 11786
rect 5580 11734 5632 11786
rect 5632 11734 5634 11786
rect 5578 11732 5634 11734
rect 5180 10780 5236 10836
rect 4508 10108 4564 10164
rect 4620 10556 4676 10612
rect 5852 10668 5908 10724
rect 5068 10332 5124 10388
rect 6972 12908 6974 12934
rect 6974 12908 7026 12934
rect 7026 12908 7028 12934
rect 5628 10332 5684 10388
rect 6188 11676 6244 11732
rect 5370 10218 5426 10220
rect 5370 10166 5372 10218
rect 5372 10166 5424 10218
rect 5424 10166 5426 10218
rect 5370 10164 5426 10166
rect 5474 10218 5530 10220
rect 5474 10166 5476 10218
rect 5476 10166 5528 10218
rect 5528 10166 5530 10218
rect 5474 10164 5530 10166
rect 5578 10218 5634 10220
rect 5578 10166 5580 10218
rect 5580 10166 5632 10218
rect 5632 10166 5634 10218
rect 5578 10164 5634 10166
rect 4396 9660 4452 9716
rect 4620 9548 4676 9604
rect 4508 8764 4564 8820
rect 4284 8258 4340 8260
rect 4284 8206 4286 8258
rect 4286 8206 4338 8258
rect 4338 8206 4340 8258
rect 4284 8204 4340 8206
rect 4060 8092 4116 8148
rect 2772 6748 2828 6804
rect 3108 6690 3164 6692
rect 3108 6638 3110 6690
rect 3110 6638 3162 6690
rect 3162 6638 3164 6690
rect 3108 6636 3164 6638
rect 3948 6748 4004 6804
rect 4732 8316 4788 8372
rect 4844 9772 4900 9828
rect 3500 6524 3556 6580
rect 2940 5964 2996 6020
rect 3108 6412 3164 6468
rect 3836 6412 3892 6468
rect 4228 6690 4284 6692
rect 4228 6638 4230 6690
rect 4230 6638 4282 6690
rect 4282 6638 4284 6690
rect 4228 6636 4284 6638
rect 4060 6412 4116 6468
rect 3612 6188 3668 6244
rect 3724 6300 3780 6356
rect 3612 5964 3668 6020
rect 2828 5906 2884 5908
rect 2828 5854 2830 5906
rect 2830 5854 2882 5906
rect 2882 5854 2884 5906
rect 2828 5852 2884 5854
rect 3388 5852 3444 5908
rect 1596 4338 1652 4340
rect 1596 4286 1598 4338
rect 1598 4286 1650 4338
rect 1650 4286 1652 4338
rect 1596 4284 1652 4286
rect 2940 5122 2996 5124
rect 2940 5070 2942 5122
rect 2942 5070 2994 5122
rect 2994 5070 2996 5122
rect 2940 5068 2996 5070
rect 3612 5122 3668 5124
rect 3612 5070 3614 5122
rect 3614 5070 3666 5122
rect 3666 5070 3668 5122
rect 3612 5068 3668 5070
rect 4732 6300 4788 6356
rect 4172 5964 4228 6020
rect 5740 9996 5796 10052
rect 4956 9548 5012 9604
rect 5068 9212 5124 9268
rect 4956 7980 5012 8036
rect 5740 9212 5796 9268
rect 5370 8650 5426 8652
rect 5370 8598 5372 8650
rect 5372 8598 5424 8650
rect 5424 8598 5426 8650
rect 5370 8596 5426 8598
rect 5474 8650 5530 8652
rect 5474 8598 5476 8650
rect 5476 8598 5528 8650
rect 5528 8598 5530 8650
rect 5474 8596 5530 8598
rect 5578 8650 5634 8652
rect 5578 8598 5580 8650
rect 5580 8598 5632 8650
rect 5632 8598 5634 8650
rect 5578 8596 5634 8598
rect 6076 9996 6132 10052
rect 5964 9826 6020 9828
rect 5964 9774 5966 9826
rect 5966 9774 6018 9826
rect 6018 9774 6020 9826
rect 5964 9772 6020 9774
rect 6524 12460 6580 12516
rect 6860 12236 6916 12292
rect 6748 11788 6804 11844
rect 6748 9548 6804 9604
rect 6188 9100 6244 9156
rect 6524 9042 6580 9044
rect 6524 8990 6526 9042
rect 6526 8990 6578 9042
rect 6578 8990 6580 9042
rect 6524 8988 6580 8990
rect 6300 8428 6356 8484
rect 6636 8764 6692 8820
rect 5370 7082 5426 7084
rect 5370 7030 5372 7082
rect 5372 7030 5424 7082
rect 5424 7030 5426 7082
rect 5370 7028 5426 7030
rect 5474 7082 5530 7084
rect 5474 7030 5476 7082
rect 5476 7030 5528 7082
rect 5528 7030 5530 7082
rect 5474 7028 5530 7030
rect 5578 7082 5634 7084
rect 5578 7030 5580 7082
rect 5580 7030 5632 7082
rect 5632 7030 5634 7082
rect 5578 7028 5634 7030
rect 5516 6690 5572 6692
rect 5516 6638 5518 6690
rect 5518 6638 5570 6690
rect 5570 6638 5572 6690
rect 5516 6636 5572 6638
rect 4844 6076 4900 6132
rect 3948 5740 4004 5796
rect 4284 5068 4340 5124
rect 4284 4450 4340 4452
rect 4284 4398 4286 4450
rect 4286 4398 4338 4450
rect 4338 4398 4340 4450
rect 4284 4396 4340 4398
rect 3612 4172 3668 4228
rect 5236 6018 5292 6020
rect 5236 5966 5238 6018
rect 5238 5966 5290 6018
rect 5290 5966 5292 6018
rect 5236 5964 5292 5966
rect 4732 5906 4788 5908
rect 4732 5854 4734 5906
rect 4734 5854 4786 5906
rect 4786 5854 4788 5906
rect 4732 5852 4788 5854
rect 5370 5514 5426 5516
rect 5370 5462 5372 5514
rect 5372 5462 5424 5514
rect 5424 5462 5426 5514
rect 5370 5460 5426 5462
rect 5474 5514 5530 5516
rect 5474 5462 5476 5514
rect 5476 5462 5528 5514
rect 5528 5462 5530 5514
rect 5474 5460 5530 5462
rect 5578 5514 5634 5516
rect 5578 5462 5580 5514
rect 5580 5462 5632 5514
rect 5632 5462 5634 5514
rect 5578 5460 5634 5462
rect 4956 5292 5012 5348
rect 4732 5122 4788 5124
rect 4732 5070 4734 5122
rect 4734 5070 4786 5122
rect 4786 5070 4788 5122
rect 4732 5068 4788 5070
rect 4956 5122 5012 5124
rect 4956 5070 4958 5122
rect 4958 5070 5010 5122
rect 5010 5070 5012 5122
rect 4956 5068 5012 5070
rect 4620 4396 4676 4452
rect 5608 4508 5664 4564
rect 5852 7868 5908 7924
rect 6748 8540 6804 8596
rect 6748 8204 6804 8260
rect 6748 6860 6804 6916
rect 5852 6188 5908 6244
rect 6412 5906 6468 5908
rect 6412 5854 6414 5906
rect 6414 5854 6466 5906
rect 6466 5854 6468 5906
rect 6412 5852 6468 5854
rect 6246 5628 6302 5684
rect 6972 11900 7028 11956
rect 7140 11788 7196 11844
rect 8204 14700 8260 14756
rect 7644 12908 7700 12964
rect 7756 13132 7812 13188
rect 7532 12236 7588 12292
rect 7420 11452 7476 11508
rect 7084 11228 7140 11284
rect 7084 9826 7140 9828
rect 7084 9774 7086 9826
rect 7086 9774 7138 9826
rect 7138 9774 7140 9826
rect 7084 9772 7140 9774
rect 7084 9100 7140 9156
rect 7084 8540 7140 8596
rect 7308 9436 7364 9492
rect 7308 9028 7310 9044
rect 7310 9028 7362 9044
rect 7362 9028 7364 9044
rect 7308 8988 7364 9028
rect 8432 12572 8488 12628
rect 11172 15874 11228 15876
rect 11172 15822 11174 15874
rect 11174 15822 11226 15874
rect 11226 15822 11228 15874
rect 11172 15820 11228 15822
rect 9528 15706 9584 15708
rect 9528 15654 9530 15706
rect 9530 15654 9582 15706
rect 9582 15654 9584 15706
rect 9528 15652 9584 15654
rect 9632 15706 9688 15708
rect 9632 15654 9634 15706
rect 9634 15654 9686 15706
rect 9686 15654 9688 15706
rect 9632 15652 9688 15654
rect 9736 15706 9792 15708
rect 9736 15654 9738 15706
rect 9738 15654 9790 15706
rect 9790 15654 9792 15706
rect 9736 15652 9792 15654
rect 8988 15314 9044 15316
rect 8988 15262 8990 15314
rect 8990 15262 9042 15314
rect 9042 15262 9044 15314
rect 8988 15260 9044 15262
rect 9772 15314 9828 15316
rect 9772 15262 9774 15314
rect 9774 15262 9826 15314
rect 9826 15262 9828 15314
rect 9772 15260 9828 15262
rect 12964 19234 13020 19236
rect 12964 19182 12966 19234
rect 12966 19182 13018 19234
rect 13018 19182 13020 19234
rect 12964 19180 13020 19182
rect 13860 20018 13916 20020
rect 13860 19966 13862 20018
rect 13862 19966 13914 20018
rect 13914 19966 13916 20018
rect 13860 19964 13916 19966
rect 14364 23324 14420 23380
rect 16156 25564 16212 25620
rect 16044 25452 16100 25508
rect 15820 24780 15876 24836
rect 15932 25340 15988 25396
rect 17612 26796 17668 26852
rect 18172 26796 18228 26852
rect 17844 26682 17900 26684
rect 17844 26630 17846 26682
rect 17846 26630 17898 26682
rect 17898 26630 17900 26682
rect 17844 26628 17900 26630
rect 17948 26682 18004 26684
rect 17948 26630 17950 26682
rect 17950 26630 18002 26682
rect 18002 26630 18004 26682
rect 17948 26628 18004 26630
rect 18052 26682 18108 26684
rect 18052 26630 18054 26682
rect 18054 26630 18106 26682
rect 18106 26630 18108 26682
rect 18052 26628 18108 26630
rect 17276 26290 17332 26292
rect 17276 26238 17278 26290
rect 17278 26238 17330 26290
rect 17330 26238 17332 26290
rect 17276 26236 17332 26238
rect 16380 25228 16436 25284
rect 16380 24722 16436 24724
rect 16380 24670 16382 24722
rect 16382 24670 16434 24722
rect 16434 24670 16436 24722
rect 16380 24668 16436 24670
rect 18172 25564 18228 25620
rect 19852 26236 19908 26292
rect 17844 25114 17900 25116
rect 17844 25062 17846 25114
rect 17846 25062 17898 25114
rect 17898 25062 17900 25114
rect 17844 25060 17900 25062
rect 17948 25114 18004 25116
rect 17948 25062 17950 25114
rect 17950 25062 18002 25114
rect 18002 25062 18004 25114
rect 17948 25060 18004 25062
rect 18052 25114 18108 25116
rect 18052 25062 18054 25114
rect 18054 25062 18106 25114
rect 18106 25062 18108 25114
rect 18052 25060 18108 25062
rect 16604 24780 16660 24836
rect 17612 24946 17668 24948
rect 17612 24894 17614 24946
rect 17614 24894 17666 24946
rect 17666 24894 17668 24946
rect 17612 24892 17668 24894
rect 17276 24722 17332 24724
rect 17276 24670 17278 24722
rect 17278 24670 17330 24722
rect 17330 24670 17332 24722
rect 17276 24668 17332 24670
rect 16604 23772 16660 23828
rect 16940 23772 16996 23828
rect 16716 23324 16772 23380
rect 14700 22428 14756 22484
rect 14028 20018 14084 20020
rect 14028 19966 14030 20018
rect 14030 19966 14082 20018
rect 14082 19966 14084 20018
rect 14028 19964 14084 19966
rect 13686 19626 13742 19628
rect 13686 19574 13688 19626
rect 13688 19574 13740 19626
rect 13740 19574 13742 19626
rect 13686 19572 13742 19574
rect 13790 19626 13846 19628
rect 13790 19574 13792 19626
rect 13792 19574 13844 19626
rect 13844 19574 13846 19626
rect 13790 19572 13846 19574
rect 13894 19626 13950 19628
rect 13894 19574 13896 19626
rect 13896 19574 13948 19626
rect 13948 19574 13950 19626
rect 13894 19572 13950 19574
rect 14364 19628 14420 19684
rect 13804 19292 13860 19348
rect 13524 19234 13580 19236
rect 13524 19182 13526 19234
rect 13526 19182 13578 19234
rect 13578 19182 13580 19234
rect 13524 19180 13580 19182
rect 13916 19404 13972 19460
rect 14588 19404 14644 19460
rect 15988 21868 16044 21924
rect 16604 21868 16660 21924
rect 17612 23884 17668 23940
rect 18732 25452 18788 25508
rect 18396 24780 18452 24836
rect 18564 24498 18620 24500
rect 18564 24446 18566 24498
rect 18566 24446 18618 24498
rect 18618 24446 18620 24498
rect 18564 24444 18620 24446
rect 19292 25340 19348 25396
rect 19964 25452 20020 25508
rect 18956 24892 19012 24948
rect 19068 24834 19124 24836
rect 19068 24782 19070 24834
rect 19070 24782 19122 24834
rect 19122 24782 19124 24834
rect 19068 24780 19124 24782
rect 20412 27074 20468 27076
rect 20412 27022 20414 27074
rect 20414 27022 20466 27074
rect 20466 27022 20468 27074
rect 20412 27020 20468 27022
rect 20972 26290 21028 26292
rect 20972 26238 20974 26290
rect 20974 26238 21026 26290
rect 21026 26238 21028 26290
rect 20972 26236 21028 26238
rect 20188 25340 20244 25396
rect 20860 25340 20916 25396
rect 19852 24780 19908 24836
rect 19628 24444 19684 24500
rect 19292 24108 19348 24164
rect 17836 23826 17892 23828
rect 17836 23774 17838 23826
rect 17838 23774 17890 23826
rect 17890 23774 17892 23826
rect 17836 23772 17892 23774
rect 17276 23714 17332 23716
rect 17276 23662 17278 23714
rect 17278 23662 17330 23714
rect 17330 23662 17332 23714
rect 17276 23660 17332 23662
rect 17844 23546 17900 23548
rect 17844 23494 17846 23546
rect 17846 23494 17898 23546
rect 17898 23494 17900 23546
rect 17844 23492 17900 23494
rect 17948 23546 18004 23548
rect 17948 23494 17950 23546
rect 17950 23494 18002 23546
rect 18002 23494 18004 23546
rect 17948 23492 18004 23494
rect 18052 23546 18108 23548
rect 18052 23494 18054 23546
rect 18054 23494 18106 23546
rect 18106 23494 18108 23546
rect 18052 23492 18108 23494
rect 18172 23154 18228 23156
rect 18172 23102 18174 23154
rect 18174 23102 18226 23154
rect 18226 23102 18228 23154
rect 18172 23100 18228 23102
rect 17780 22876 17836 22932
rect 18060 22876 18116 22932
rect 16716 21532 16772 21588
rect 16044 20300 16100 20356
rect 13132 18844 13188 18900
rect 14812 19628 14868 19684
rect 12684 18396 12740 18452
rect 12740 18060 12796 18116
rect 12628 17612 12684 17668
rect 12796 17724 12852 17780
rect 13300 18060 13356 18116
rect 14046 18562 14102 18564
rect 14046 18510 14048 18562
rect 14048 18510 14100 18562
rect 14100 18510 14102 18562
rect 14046 18508 14102 18510
rect 13804 18172 13860 18228
rect 15036 19234 15092 19236
rect 15036 19182 15038 19234
rect 15038 19182 15090 19234
rect 15090 19182 15092 19234
rect 15036 19180 15092 19182
rect 13686 18058 13742 18060
rect 13686 18006 13688 18058
rect 13688 18006 13740 18058
rect 13740 18006 13742 18058
rect 13686 18004 13742 18006
rect 13790 18058 13846 18060
rect 13790 18006 13792 18058
rect 13792 18006 13844 18058
rect 13844 18006 13846 18058
rect 13790 18004 13846 18006
rect 13894 18058 13950 18060
rect 13894 18006 13896 18058
rect 13896 18006 13948 18058
rect 13948 18006 13950 18058
rect 14476 18060 14532 18116
rect 13894 18004 13950 18006
rect 14252 17948 14308 18004
rect 13132 17612 13188 17668
rect 13580 17666 13636 17668
rect 13580 17614 13582 17666
rect 13582 17614 13634 17666
rect 13634 17614 13636 17666
rect 16156 20188 16212 20244
rect 16324 19404 16380 19460
rect 18172 22316 18228 22372
rect 17844 21978 17900 21980
rect 17844 21926 17846 21978
rect 17846 21926 17898 21978
rect 17898 21926 17900 21978
rect 17844 21924 17900 21926
rect 17948 21978 18004 21980
rect 17948 21926 17950 21978
rect 17950 21926 18002 21978
rect 18002 21926 18004 21978
rect 17948 21924 18004 21926
rect 18052 21978 18108 21980
rect 18052 21926 18054 21978
rect 18054 21926 18106 21978
rect 18106 21926 18108 21978
rect 18052 21924 18108 21926
rect 17724 21756 17780 21812
rect 16492 19234 16548 19236
rect 16492 19182 16494 19234
rect 16494 19182 16546 19234
rect 16546 19182 16548 19234
rect 16492 19180 16548 19182
rect 16604 19292 16660 19348
rect 15596 18508 15652 18564
rect 17724 21586 17780 21588
rect 17724 21534 17726 21586
rect 17726 21534 17778 21586
rect 17778 21534 17780 21586
rect 17724 21532 17780 21534
rect 18172 21308 18228 21364
rect 17844 20410 17900 20412
rect 17844 20358 17846 20410
rect 17846 20358 17898 20410
rect 17898 20358 17900 20410
rect 17844 20356 17900 20358
rect 17948 20410 18004 20412
rect 17948 20358 17950 20410
rect 17950 20358 18002 20410
rect 18002 20358 18004 20410
rect 17948 20356 18004 20358
rect 18052 20410 18108 20412
rect 18052 20358 18054 20410
rect 18054 20358 18106 20410
rect 18106 20358 18108 20410
rect 18052 20356 18108 20358
rect 17724 20188 17780 20244
rect 16884 19234 16940 19236
rect 16884 19182 16886 19234
rect 16886 19182 16938 19234
rect 16938 19182 16940 19234
rect 16884 19180 16940 19182
rect 16604 18732 16660 18788
rect 14924 18284 14980 18340
rect 15260 18172 15316 18228
rect 14924 17836 14980 17892
rect 13580 17612 13636 17614
rect 12927 16882 12983 16884
rect 12927 16830 12929 16882
rect 12929 16830 12981 16882
rect 12981 16830 12983 16882
rect 12927 16828 12983 16830
rect 14028 16716 14084 16772
rect 13686 16490 13742 16492
rect 13686 16438 13688 16490
rect 13688 16438 13740 16490
rect 13740 16438 13742 16490
rect 13686 16436 13742 16438
rect 13790 16490 13846 16492
rect 13790 16438 13792 16490
rect 13792 16438 13844 16490
rect 13844 16438 13846 16490
rect 13790 16436 13846 16438
rect 13894 16490 13950 16492
rect 13894 16438 13896 16490
rect 13896 16438 13948 16490
rect 13948 16438 13950 16490
rect 13894 16436 13950 16438
rect 12516 15874 12572 15876
rect 12516 15822 12518 15874
rect 12518 15822 12570 15874
rect 12570 15822 12572 15874
rect 12516 15820 12572 15822
rect 11172 15260 11228 15316
rect 9528 14138 9584 14140
rect 9528 14086 9530 14138
rect 9530 14086 9582 14138
rect 9582 14086 9584 14138
rect 9528 14084 9584 14086
rect 9632 14138 9688 14140
rect 9632 14086 9634 14138
rect 9634 14086 9686 14138
rect 9686 14086 9688 14138
rect 9632 14084 9688 14086
rect 9736 14138 9792 14140
rect 9736 14086 9738 14138
rect 9738 14086 9790 14138
rect 9790 14086 9792 14138
rect 9736 14084 9792 14086
rect 9884 13244 9940 13300
rect 11340 13244 11396 13300
rect 9324 13020 9380 13076
rect 8876 12460 8932 12516
rect 7756 12236 7812 12292
rect 7980 12162 7982 12180
rect 7982 12162 8034 12180
rect 8034 12162 8036 12180
rect 7980 12124 8036 12162
rect 8316 12012 8372 12068
rect 8764 12290 8820 12292
rect 8764 12238 8766 12290
rect 8766 12238 8818 12290
rect 8818 12238 8820 12290
rect 8764 12236 8820 12238
rect 7756 11452 7812 11508
rect 7588 9714 7644 9716
rect 7588 9662 7590 9714
rect 7590 9662 7642 9714
rect 7642 9662 7644 9714
rect 7588 9660 7644 9662
rect 7644 9436 7700 9492
rect 7532 9324 7588 9380
rect 7532 8428 7588 8484
rect 7420 8092 7476 8148
rect 6860 5516 6916 5572
rect 8428 9826 8484 9828
rect 8428 9774 8430 9826
rect 8430 9774 8482 9826
rect 8482 9774 8484 9826
rect 8428 9772 8484 9774
rect 8316 8988 8372 9044
rect 7756 8204 7812 8260
rect 7644 7474 7700 7476
rect 7644 7422 7646 7474
rect 7646 7422 7698 7474
rect 7698 7422 7700 7474
rect 7644 7420 7700 7422
rect 7868 7868 7924 7924
rect 7756 7196 7812 7252
rect 7868 7084 7924 7140
rect 6748 5404 6804 5460
rect 6412 5068 6468 5124
rect 7084 6524 7140 6580
rect 7252 5964 7308 6020
rect 7868 6188 7924 6244
rect 8876 11788 8932 11844
rect 8652 11676 8708 11732
rect 9212 11676 9268 11732
rect 9528 12570 9584 12572
rect 9528 12518 9530 12570
rect 9530 12518 9582 12570
rect 9582 12518 9584 12570
rect 9528 12516 9584 12518
rect 9632 12570 9688 12572
rect 9632 12518 9634 12570
rect 9634 12518 9686 12570
rect 9686 12518 9688 12570
rect 9632 12516 9688 12518
rect 9736 12570 9792 12572
rect 9736 12518 9738 12570
rect 9738 12518 9790 12570
rect 9790 12518 9792 12570
rect 9736 12516 9792 12518
rect 10164 13020 10220 13076
rect 9884 11900 9940 11956
rect 10332 11564 10388 11620
rect 10556 12796 10612 12852
rect 10556 12236 10612 12292
rect 9660 11394 9716 11396
rect 9660 11342 9662 11394
rect 9662 11342 9714 11394
rect 9714 11342 9716 11394
rect 9660 11340 9716 11342
rect 9528 11002 9584 11004
rect 9528 10950 9530 11002
rect 9530 10950 9582 11002
rect 9582 10950 9584 11002
rect 9528 10948 9584 10950
rect 9632 11002 9688 11004
rect 9632 10950 9634 11002
rect 9634 10950 9686 11002
rect 9686 10950 9688 11002
rect 9632 10948 9688 10950
rect 9736 11002 9792 11004
rect 9736 10950 9738 11002
rect 9738 10950 9790 11002
rect 9790 10950 9792 11002
rect 9736 10948 9792 10950
rect 10220 11170 10276 11172
rect 10220 11118 10222 11170
rect 10222 11118 10274 11170
rect 10274 11118 10276 11170
rect 10220 11116 10276 11118
rect 10220 10780 10276 10836
rect 11340 13020 11396 13076
rect 10780 12908 10836 12964
rect 10948 12178 11004 12180
rect 10948 12126 10950 12178
rect 10950 12126 11002 12178
rect 11002 12126 11004 12178
rect 10948 12124 11004 12126
rect 11116 11564 11172 11620
rect 11228 12124 11284 12180
rect 11340 12066 11396 12068
rect 11340 12014 11342 12066
rect 11342 12014 11394 12066
rect 11394 12014 11396 12066
rect 11340 12012 11396 12014
rect 12012 12962 12068 12964
rect 12012 12910 12014 12962
rect 12014 12910 12066 12962
rect 12066 12910 12068 12962
rect 12012 12908 12068 12910
rect 12236 12908 12292 12964
rect 12012 12348 12068 12404
rect 11564 11788 11620 11844
rect 9772 10386 9828 10388
rect 9772 10334 9774 10386
rect 9774 10334 9826 10386
rect 9826 10334 9828 10386
rect 9772 10332 9828 10334
rect 10444 10332 10500 10388
rect 9212 10220 9268 10276
rect 9100 9772 9156 9828
rect 8652 9660 8708 9716
rect 9528 9434 9584 9436
rect 9528 9382 9530 9434
rect 9530 9382 9582 9434
rect 9582 9382 9584 9434
rect 9528 9380 9584 9382
rect 9632 9434 9688 9436
rect 9632 9382 9634 9434
rect 9634 9382 9686 9434
rect 9686 9382 9688 9434
rect 9632 9380 9688 9382
rect 9736 9434 9792 9436
rect 9736 9382 9738 9434
rect 9738 9382 9790 9434
rect 9790 9382 9792 9434
rect 9736 9380 9792 9382
rect 10220 9324 10276 9380
rect 10220 9100 10276 9156
rect 9548 8988 9604 9044
rect 8652 8258 8708 8260
rect 8652 8206 8654 8258
rect 8654 8206 8706 8258
rect 8706 8206 8708 8258
rect 8652 8204 8708 8206
rect 8540 7980 8596 8036
rect 9100 7308 9156 7364
rect 10108 8258 10164 8260
rect 8988 7084 9044 7140
rect 8260 6524 8316 6580
rect 8204 6300 8260 6356
rect 6972 5292 7028 5348
rect 6806 5180 6862 5236
rect 7084 5122 7140 5124
rect 7084 5070 7086 5122
rect 7086 5070 7138 5122
rect 7138 5070 7140 5122
rect 7084 5068 7140 5070
rect 5740 4284 5796 4340
rect 5370 3946 5426 3948
rect 5370 3894 5372 3946
rect 5372 3894 5424 3946
rect 5424 3894 5426 3946
rect 5370 3892 5426 3894
rect 5474 3946 5530 3948
rect 5474 3894 5476 3946
rect 5476 3894 5528 3946
rect 5528 3894 5530 3946
rect 5474 3892 5530 3894
rect 5578 3946 5634 3948
rect 5578 3894 5580 3946
rect 5580 3894 5632 3946
rect 5632 3894 5634 3946
rect 5578 3892 5634 3894
rect 8092 5740 8148 5796
rect 8092 5516 8148 5572
rect 8204 4956 8260 5012
rect 8316 6188 8372 6244
rect 10108 8206 10110 8258
rect 10110 8206 10162 8258
rect 10162 8206 10164 8258
rect 10108 8204 10164 8206
rect 9772 8092 9828 8148
rect 9528 7866 9584 7868
rect 9528 7814 9530 7866
rect 9530 7814 9582 7866
rect 9582 7814 9584 7866
rect 9528 7812 9584 7814
rect 9632 7866 9688 7868
rect 9632 7814 9634 7866
rect 9634 7814 9686 7866
rect 9686 7814 9688 7866
rect 9632 7812 9688 7814
rect 9736 7866 9792 7868
rect 9736 7814 9738 7866
rect 9738 7814 9790 7866
rect 9790 7814 9792 7866
rect 9736 7812 9792 7814
rect 9996 7362 10052 7364
rect 9996 7310 9998 7362
rect 9998 7310 10050 7362
rect 10050 7310 10052 7362
rect 9996 7308 10052 7310
rect 9528 6298 9584 6300
rect 9528 6246 9530 6298
rect 9530 6246 9582 6298
rect 9582 6246 9584 6298
rect 9528 6244 9584 6246
rect 9632 6298 9688 6300
rect 9632 6246 9634 6298
rect 9634 6246 9686 6298
rect 9686 6246 9688 6298
rect 9632 6244 9688 6246
rect 9736 6298 9792 6300
rect 9736 6246 9738 6298
rect 9738 6246 9790 6298
rect 9790 6246 9792 6298
rect 9736 6244 9792 6246
rect 9324 6076 9380 6132
rect 9996 6076 10052 6132
rect 8316 4396 8372 4452
rect 8428 5292 8484 5348
rect 8428 5068 8484 5124
rect 9996 5180 10052 5236
rect 10108 5852 10164 5908
rect 10390 6860 10446 6916
rect 10556 7474 10612 7476
rect 10556 7422 10558 7474
rect 10558 7422 10610 7474
rect 10610 7422 10612 7474
rect 10556 7420 10612 7422
rect 10556 6748 10612 6804
rect 10780 6524 10836 6580
rect 10892 9660 10948 9716
rect 10220 5628 10276 5684
rect 11116 11116 11172 11172
rect 11452 11564 11508 11620
rect 11396 9826 11452 9828
rect 11396 9774 11398 9826
rect 11398 9774 11450 9826
rect 11450 9774 11452 9826
rect 11396 9772 11452 9774
rect 11228 9436 11284 9492
rect 11228 9212 11284 9268
rect 11116 7980 11172 8036
rect 11340 8204 11396 8260
rect 11004 7420 11060 7476
rect 11172 6914 11228 6916
rect 11172 6862 11174 6914
rect 11174 6862 11226 6914
rect 11226 6862 11228 6914
rect 11172 6860 11228 6862
rect 11900 12178 11956 12180
rect 11900 12126 11902 12178
rect 11902 12126 11954 12178
rect 11954 12126 11956 12178
rect 11900 12124 11956 12126
rect 14812 17724 14868 17780
rect 14364 16716 14420 16772
rect 14028 15372 14084 15428
rect 15764 17948 15820 18004
rect 15932 17836 15988 17892
rect 15484 17724 15540 17780
rect 16324 18226 16380 18228
rect 16324 18174 16326 18226
rect 16326 18174 16378 18226
rect 16378 18174 16380 18226
rect 16324 18172 16380 18174
rect 16156 17666 16212 17668
rect 16156 17614 16158 17666
rect 16158 17614 16210 17666
rect 16210 17614 16212 17666
rect 16156 17612 16212 17614
rect 14980 17554 15036 17556
rect 14980 17502 14982 17554
rect 14982 17502 15034 17554
rect 15034 17502 15036 17554
rect 14980 17500 15036 17502
rect 14700 16828 14756 16884
rect 14644 15372 14700 15428
rect 15932 15484 15988 15540
rect 14924 15148 14980 15204
rect 13686 14922 13742 14924
rect 13686 14870 13688 14922
rect 13688 14870 13740 14922
rect 13740 14870 13742 14922
rect 13686 14868 13742 14870
rect 13790 14922 13846 14924
rect 13790 14870 13792 14922
rect 13792 14870 13844 14922
rect 13844 14870 13846 14922
rect 13790 14868 13846 14870
rect 13894 14922 13950 14924
rect 13894 14870 13896 14922
rect 13896 14870 13948 14922
rect 13948 14870 13950 14922
rect 13894 14868 13950 14870
rect 15148 13970 15204 13972
rect 15148 13918 15150 13970
rect 15150 13918 15202 13970
rect 15202 13918 15204 13970
rect 15148 13916 15204 13918
rect 14476 13634 14532 13636
rect 14476 13582 14478 13634
rect 14478 13582 14530 13634
rect 14530 13582 14532 13634
rect 14476 13580 14532 13582
rect 13686 13354 13742 13356
rect 13686 13302 13688 13354
rect 13688 13302 13740 13354
rect 13740 13302 13742 13354
rect 13686 13300 13742 13302
rect 13790 13354 13846 13356
rect 13790 13302 13792 13354
rect 13792 13302 13844 13354
rect 13844 13302 13846 13354
rect 13790 13300 13846 13302
rect 13894 13354 13950 13356
rect 13894 13302 13896 13354
rect 13896 13302 13948 13354
rect 13948 13302 13950 13354
rect 13894 13300 13950 13302
rect 14028 13132 14084 13188
rect 12572 12460 12628 12516
rect 12460 12348 12516 12404
rect 12572 11618 12628 11620
rect 12572 11566 12574 11618
rect 12574 11566 12626 11618
rect 12626 11566 12628 11618
rect 12572 11564 12628 11566
rect 13692 12460 13748 12516
rect 14364 13020 14420 13076
rect 14588 12908 14644 12964
rect 14196 12124 14252 12180
rect 15596 12962 15652 12964
rect 15596 12910 15598 12962
rect 15598 12910 15650 12962
rect 15650 12910 15652 12962
rect 15596 12908 15652 12910
rect 13686 11786 13742 11788
rect 13686 11734 13688 11786
rect 13688 11734 13740 11786
rect 13740 11734 13742 11786
rect 13686 11732 13742 11734
rect 13790 11786 13846 11788
rect 13790 11734 13792 11786
rect 13792 11734 13844 11786
rect 13844 11734 13846 11786
rect 13790 11732 13846 11734
rect 13894 11786 13950 11788
rect 13894 11734 13896 11786
rect 13896 11734 13948 11786
rect 13948 11734 13950 11786
rect 14028 11788 14084 11844
rect 13894 11732 13950 11734
rect 14588 11676 14644 11732
rect 15204 12796 15260 12852
rect 13356 11564 13412 11620
rect 15316 12402 15372 12404
rect 15316 12350 15318 12402
rect 15318 12350 15370 12402
rect 15370 12350 15372 12402
rect 15316 12348 15372 12350
rect 14980 11788 15036 11844
rect 14812 11564 14868 11620
rect 12908 11116 12964 11172
rect 12236 10668 12292 10724
rect 12460 10668 12516 10724
rect 12180 10444 12236 10500
rect 11788 9996 11844 10052
rect 12012 10220 12068 10276
rect 11676 9212 11732 9268
rect 11788 9660 11844 9716
rect 11788 8876 11844 8932
rect 11900 9100 11956 9156
rect 11788 8652 11844 8708
rect 11788 8092 11844 8148
rect 11564 7980 11620 8036
rect 12348 9996 12404 10052
rect 12180 9100 12236 9156
rect 12348 8988 12404 9044
rect 12012 8428 12068 8484
rect 12796 10668 12852 10724
rect 13524 11170 13580 11172
rect 13524 11118 13526 11170
rect 13526 11118 13578 11170
rect 13578 11118 13580 11170
rect 13524 11116 13580 11118
rect 13132 10610 13188 10612
rect 13132 10558 13134 10610
rect 13134 10558 13186 10610
rect 13186 10558 13188 10610
rect 13132 10556 13188 10558
rect 14476 11228 14532 11284
rect 14140 10668 14196 10724
rect 13916 10610 13972 10612
rect 13916 10558 13918 10610
rect 13918 10558 13970 10610
rect 13970 10558 13972 10610
rect 13916 10556 13972 10558
rect 13132 10332 13188 10388
rect 13132 9884 13188 9940
rect 13020 9548 13076 9604
rect 12572 9324 12628 9380
rect 12908 9436 12964 9492
rect 12684 9212 12740 9268
rect 12348 8652 12404 8708
rect 12348 8428 12404 8484
rect 12236 8204 12292 8260
rect 12124 8092 12180 8148
rect 12012 7868 12068 7924
rect 11676 6860 11732 6916
rect 11564 6578 11620 6580
rect 11564 6526 11566 6578
rect 11566 6526 11618 6578
rect 11618 6526 11620 6578
rect 11564 6524 11620 6526
rect 10444 6188 10500 6244
rect 10332 5516 10388 5572
rect 9528 4730 9584 4732
rect 9528 4678 9530 4730
rect 9530 4678 9582 4730
rect 9582 4678 9584 4730
rect 9528 4676 9584 4678
rect 9632 4730 9688 4732
rect 9632 4678 9634 4730
rect 9634 4678 9686 4730
rect 9686 4678 9688 4730
rect 9632 4676 9688 4678
rect 9736 4730 9792 4732
rect 9736 4678 9738 4730
rect 9738 4678 9790 4730
rect 9790 4678 9792 4730
rect 9736 4676 9792 4678
rect 9660 4338 9716 4340
rect 9660 4286 9662 4338
rect 9662 4286 9714 4338
rect 9714 4286 9716 4338
rect 9660 4284 9716 4286
rect 10332 5180 10388 5236
rect 10220 4844 10276 4900
rect 10668 6130 10724 6132
rect 10668 6078 10670 6130
rect 10670 6078 10722 6130
rect 10722 6078 10724 6130
rect 10668 6076 10724 6078
rect 10444 5068 10500 5124
rect 11004 5964 11060 6020
rect 11116 5852 11172 5908
rect 10986 4844 11042 4900
rect 11732 6188 11788 6244
rect 11900 6524 11956 6580
rect 11564 5964 11620 6020
rect 11676 5906 11732 5908
rect 11676 5854 11678 5906
rect 11678 5854 11730 5906
rect 11730 5854 11732 5906
rect 11676 5852 11732 5854
rect 11228 5628 11284 5684
rect 11732 5404 11788 5460
rect 11676 4956 11732 5012
rect 11788 4844 11844 4900
rect 12012 6300 12068 6356
rect 12012 6130 12068 6132
rect 12012 6078 12014 6130
rect 12014 6078 12066 6130
rect 12066 6078 12068 6130
rect 12012 6076 12068 6078
rect 12572 8204 12628 8260
rect 12348 7756 12404 7812
rect 12348 7532 12404 7588
rect 12460 7474 12516 7476
rect 12460 7422 12462 7474
rect 12462 7422 12514 7474
rect 12514 7422 12516 7474
rect 12460 7420 12516 7422
rect 12460 6972 12516 7028
rect 13686 10218 13742 10220
rect 13686 10166 13688 10218
rect 13688 10166 13740 10218
rect 13740 10166 13742 10218
rect 13686 10164 13742 10166
rect 13790 10218 13846 10220
rect 13790 10166 13792 10218
rect 13792 10166 13844 10218
rect 13844 10166 13846 10218
rect 13790 10164 13846 10166
rect 13894 10218 13950 10220
rect 13894 10166 13896 10218
rect 13896 10166 13948 10218
rect 13948 10166 13950 10218
rect 13894 10164 13950 10166
rect 13468 9212 13524 9268
rect 13692 9042 13748 9044
rect 13692 8990 13694 9042
rect 13694 8990 13746 9042
rect 13746 8990 13748 9042
rect 13692 8988 13748 8990
rect 14196 9042 14252 9044
rect 14196 8990 14198 9042
rect 14198 8990 14250 9042
rect 14250 8990 14252 9042
rect 14196 8988 14252 8990
rect 14700 11228 14756 11284
rect 16268 15148 16324 15204
rect 15932 12236 15988 12292
rect 16492 15036 16548 15092
rect 17052 17666 17108 17668
rect 17052 17614 17054 17666
rect 17054 17614 17106 17666
rect 17106 17614 17108 17666
rect 17052 17612 17108 17614
rect 16716 16716 16772 16772
rect 16716 15202 16772 15204
rect 16716 15150 16718 15202
rect 16718 15150 16770 15202
rect 16770 15150 16772 15202
rect 16716 15148 16772 15150
rect 16604 13916 16660 13972
rect 16492 13746 16548 13748
rect 16492 13694 16494 13746
rect 16494 13694 16546 13746
rect 16546 13694 16548 13746
rect 16492 13692 16548 13694
rect 16660 13746 16716 13748
rect 16660 13694 16662 13746
rect 16662 13694 16714 13746
rect 16714 13694 16716 13746
rect 16660 13692 16716 13694
rect 16380 13580 16436 13636
rect 16268 13020 16324 13076
rect 16716 13468 16772 13524
rect 16380 12684 16436 12740
rect 16828 12908 16884 12964
rect 16940 13468 16996 13524
rect 15820 11452 15876 11508
rect 16044 11564 16100 11620
rect 15148 11340 15204 11396
rect 15148 10780 15204 10836
rect 14812 10610 14868 10612
rect 14812 10558 14814 10610
rect 14814 10558 14866 10610
rect 14866 10558 14868 10610
rect 14812 10556 14868 10558
rect 15540 11394 15596 11396
rect 15540 11342 15542 11394
rect 15542 11342 15594 11394
rect 15594 11342 15596 11394
rect 15540 11340 15596 11342
rect 14588 8988 14644 9044
rect 15036 8988 15092 9044
rect 13686 8650 13742 8652
rect 13686 8598 13688 8650
rect 13688 8598 13740 8650
rect 13740 8598 13742 8650
rect 13686 8596 13742 8598
rect 13790 8650 13846 8652
rect 13790 8598 13792 8650
rect 13792 8598 13844 8650
rect 13844 8598 13846 8650
rect 13790 8596 13846 8598
rect 13894 8650 13950 8652
rect 13894 8598 13896 8650
rect 13896 8598 13948 8650
rect 13948 8598 13950 8650
rect 13894 8596 13950 8598
rect 12908 7644 12964 7700
rect 12124 5852 12180 5908
rect 12236 6300 12292 6356
rect 13356 7756 13412 7812
rect 12460 6076 12516 6132
rect 13188 6636 13244 6692
rect 13804 7980 13860 8036
rect 13580 7308 13636 7364
rect 13468 7196 13524 7252
rect 14028 7196 14084 7252
rect 13686 7082 13742 7084
rect 13686 7030 13688 7082
rect 13688 7030 13740 7082
rect 13740 7030 13742 7082
rect 13686 7028 13742 7030
rect 13790 7082 13846 7084
rect 13790 7030 13792 7082
rect 13792 7030 13844 7082
rect 13844 7030 13846 7082
rect 13790 7028 13846 7030
rect 13894 7082 13950 7084
rect 13894 7030 13896 7082
rect 13896 7030 13948 7082
rect 13948 7030 13950 7082
rect 13894 7028 13950 7030
rect 13860 6914 13916 6916
rect 13860 6862 13862 6914
rect 13862 6862 13914 6914
rect 13914 6862 13916 6914
rect 13860 6860 13916 6862
rect 14028 6748 14084 6804
rect 13580 6690 13636 6692
rect 13580 6638 13582 6690
rect 13582 6638 13634 6690
rect 13634 6638 13636 6690
rect 13580 6636 13636 6638
rect 13804 6636 13860 6692
rect 13468 6188 13524 6244
rect 12236 5404 12292 5460
rect 12012 5292 12068 5348
rect 13804 5740 13860 5796
rect 13686 5514 13742 5516
rect 13686 5462 13688 5514
rect 13688 5462 13740 5514
rect 13740 5462 13742 5514
rect 13686 5460 13742 5462
rect 13790 5514 13846 5516
rect 13790 5462 13792 5514
rect 13792 5462 13844 5514
rect 13844 5462 13846 5514
rect 13790 5460 13846 5462
rect 13894 5514 13950 5516
rect 13894 5462 13896 5514
rect 13896 5462 13948 5514
rect 13948 5462 13950 5514
rect 13894 5460 13950 5462
rect 14364 6860 14420 6916
rect 14364 6690 14420 6692
rect 14364 6638 14366 6690
rect 14366 6638 14418 6690
rect 14418 6638 14420 6690
rect 14364 6636 14420 6638
rect 14364 6412 14420 6468
rect 14700 7868 14756 7924
rect 14868 7868 14924 7924
rect 14588 7196 14644 7252
rect 15260 8930 15316 8932
rect 15260 8878 15262 8930
rect 15262 8878 15314 8930
rect 15314 8878 15316 8930
rect 15260 8876 15316 8878
rect 15708 10780 15764 10836
rect 15596 9772 15652 9828
rect 16492 12290 16548 12292
rect 16492 12238 16494 12290
rect 16494 12238 16546 12290
rect 16546 12238 16548 12290
rect 16492 12236 16548 12238
rect 16660 12236 16716 12292
rect 16828 12012 16884 12068
rect 15148 8370 15204 8372
rect 15148 8318 15150 8370
rect 15150 8318 15202 8370
rect 15202 8318 15204 8370
rect 15148 8316 15204 8318
rect 14476 5964 14532 6020
rect 13636 5234 13692 5236
rect 13636 5182 13638 5234
rect 13638 5182 13690 5234
rect 13690 5182 13692 5234
rect 13636 5180 13692 5182
rect 13020 4284 13076 4340
rect 14588 5234 14644 5236
rect 14588 5182 14590 5234
rect 14590 5182 14642 5234
rect 14642 5182 14644 5234
rect 14588 5180 14644 5182
rect 4508 3554 4564 3556
rect 4508 3502 4510 3554
rect 4510 3502 4562 3554
rect 4562 3502 4564 3554
rect 4508 3500 4564 3502
rect 13686 3946 13742 3948
rect 13686 3894 13688 3946
rect 13688 3894 13740 3946
rect 13740 3894 13742 3946
rect 13686 3892 13742 3894
rect 13790 3946 13846 3948
rect 13790 3894 13792 3946
rect 13792 3894 13844 3946
rect 13844 3894 13846 3946
rect 13790 3892 13846 3894
rect 13894 3946 13950 3948
rect 13894 3894 13896 3946
rect 13896 3894 13948 3946
rect 13948 3894 13950 3946
rect 13894 3892 13950 3894
rect 11228 3778 11284 3780
rect 11228 3726 11230 3778
rect 11230 3726 11282 3778
rect 11282 3726 11284 3778
rect 11228 3724 11284 3726
rect 5852 3500 5908 3556
rect 4844 3388 4900 3444
rect 6132 3442 6188 3444
rect 6132 3390 6134 3442
rect 6134 3390 6186 3442
rect 6186 3390 6188 3442
rect 6132 3388 6188 3390
rect 15036 6636 15092 6692
rect 14868 6412 14924 6468
rect 14868 5964 14924 6020
rect 15372 7250 15428 7252
rect 15372 7198 15374 7250
rect 15374 7198 15426 7250
rect 15426 7198 15428 7250
rect 15372 7196 15428 7198
rect 15372 6690 15428 6692
rect 15372 6638 15374 6690
rect 15374 6638 15426 6690
rect 15426 6638 15428 6690
rect 15372 6636 15428 6638
rect 15596 7868 15652 7924
rect 16380 11452 16436 11508
rect 15932 8258 15988 8260
rect 15932 8206 15934 8258
rect 15934 8206 15986 8258
rect 15986 8206 15988 8258
rect 15932 8204 15988 8206
rect 15932 7756 15988 7812
rect 15764 7474 15820 7476
rect 15764 7422 15766 7474
rect 15766 7422 15818 7474
rect 15818 7422 15820 7474
rect 15764 7420 15820 7422
rect 18956 23100 19012 23156
rect 19516 23996 19572 24052
rect 20412 24332 20468 24388
rect 18508 22988 18564 23044
rect 19180 22988 19236 23044
rect 20300 23826 20356 23828
rect 20300 23774 20302 23826
rect 20302 23774 20354 23826
rect 20354 23774 20356 23826
rect 20300 23772 20356 23774
rect 22002 27466 22058 27468
rect 22002 27414 22004 27466
rect 22004 27414 22056 27466
rect 22056 27414 22058 27466
rect 22002 27412 22058 27414
rect 22106 27466 22162 27468
rect 22106 27414 22108 27466
rect 22108 27414 22160 27466
rect 22160 27414 22162 27466
rect 22106 27412 22162 27414
rect 22210 27466 22266 27468
rect 22210 27414 22212 27466
rect 22212 27414 22264 27466
rect 22264 27414 22266 27466
rect 22210 27412 22266 27414
rect 21532 27132 21588 27188
rect 21980 27186 22036 27188
rect 21980 27134 21982 27186
rect 21982 27134 22034 27186
rect 22034 27134 22036 27186
rect 21980 27132 22036 27134
rect 23660 29260 23716 29316
rect 24108 29372 24164 29428
rect 23492 27020 23548 27076
rect 21868 26236 21924 26292
rect 22002 25898 22058 25900
rect 22002 25846 22004 25898
rect 22004 25846 22056 25898
rect 22056 25846 22058 25898
rect 22002 25844 22058 25846
rect 22106 25898 22162 25900
rect 22106 25846 22108 25898
rect 22108 25846 22160 25898
rect 22160 25846 22162 25898
rect 22106 25844 22162 25846
rect 22210 25898 22266 25900
rect 22210 25846 22212 25898
rect 22212 25846 22264 25898
rect 22264 25846 22266 25898
rect 22210 25844 22266 25846
rect 21084 24668 21140 24724
rect 21756 24722 21812 24724
rect 21756 24670 21758 24722
rect 21758 24670 21810 24722
rect 21810 24670 21812 24722
rect 21756 24668 21812 24670
rect 22092 25004 22148 25060
rect 22092 24444 22148 24500
rect 22428 24780 22484 24836
rect 22002 24330 22058 24332
rect 22002 24278 22004 24330
rect 22004 24278 22056 24330
rect 22056 24278 22058 24330
rect 22002 24276 22058 24278
rect 22106 24330 22162 24332
rect 22106 24278 22108 24330
rect 22108 24278 22160 24330
rect 22160 24278 22162 24330
rect 22106 24276 22162 24278
rect 22210 24330 22266 24332
rect 22210 24278 22212 24330
rect 22212 24278 22264 24330
rect 22264 24278 22266 24330
rect 22210 24276 22266 24278
rect 22988 24780 23044 24836
rect 22876 24610 22932 24612
rect 22876 24558 22878 24610
rect 22878 24558 22930 24610
rect 22930 24558 22932 24610
rect 22876 24556 22932 24558
rect 22428 23772 22484 23828
rect 20132 23378 20188 23380
rect 20132 23326 20134 23378
rect 20134 23326 20186 23378
rect 20186 23326 20188 23378
rect 20132 23324 20188 23326
rect 19964 22428 20020 22484
rect 19180 22370 19236 22372
rect 19180 22318 19182 22370
rect 19182 22318 19234 22370
rect 19234 22318 19236 22370
rect 19180 22316 19236 22318
rect 18564 21810 18620 21812
rect 18564 21758 18566 21810
rect 18566 21758 18618 21810
rect 18618 21758 18620 21810
rect 18564 21756 18620 21758
rect 18902 21756 18958 21812
rect 19852 21756 19908 21812
rect 18396 21308 18452 21364
rect 17276 17836 17332 17892
rect 17500 17836 17556 17892
rect 17164 15036 17220 15092
rect 17052 11676 17108 11732
rect 16380 9826 16436 9828
rect 16380 9774 16382 9826
rect 16382 9774 16434 9826
rect 16434 9774 16436 9826
rect 16380 9772 16436 9774
rect 17276 14252 17332 14308
rect 17500 13692 17556 13748
rect 17444 13522 17500 13524
rect 17444 13470 17446 13522
rect 17446 13470 17498 13522
rect 17498 13470 17500 13522
rect 17444 13468 17500 13470
rect 18284 19234 18340 19236
rect 18284 19182 18286 19234
rect 18286 19182 18338 19234
rect 18338 19182 18340 19234
rect 18284 19180 18340 19182
rect 18844 20018 18900 20020
rect 18844 19966 18846 20018
rect 18846 19966 18898 20018
rect 18898 19966 18900 20018
rect 18844 19964 18900 19966
rect 18732 19180 18788 19236
rect 19404 19852 19460 19908
rect 17844 18842 17900 18844
rect 17844 18790 17846 18842
rect 17846 18790 17898 18842
rect 17898 18790 17900 18842
rect 17844 18788 17900 18790
rect 17948 18842 18004 18844
rect 17948 18790 17950 18842
rect 17950 18790 18002 18842
rect 18002 18790 18004 18842
rect 17948 18788 18004 18790
rect 18052 18842 18108 18844
rect 18052 18790 18054 18842
rect 18054 18790 18106 18842
rect 18106 18790 18108 18842
rect 18052 18788 18108 18790
rect 17724 18620 17780 18676
rect 18844 18508 18900 18564
rect 17724 18284 17780 18340
rect 17724 18060 17780 18116
rect 17836 17612 17892 17668
rect 18508 17948 18564 18004
rect 19740 19234 19796 19236
rect 19740 19182 19742 19234
rect 19742 19182 19794 19234
rect 19794 19182 19796 19234
rect 19740 19180 19796 19182
rect 19404 18508 19460 18564
rect 19516 18396 19572 18452
rect 19348 17890 19404 17892
rect 19348 17838 19350 17890
rect 19350 17838 19402 17890
rect 19402 17838 19404 17890
rect 19348 17836 19404 17838
rect 18956 17612 19012 17668
rect 17844 17274 17900 17276
rect 17844 17222 17846 17274
rect 17846 17222 17898 17274
rect 17898 17222 17900 17274
rect 17844 17220 17900 17222
rect 17948 17274 18004 17276
rect 17948 17222 17950 17274
rect 17950 17222 18002 17274
rect 18002 17222 18004 17274
rect 17948 17220 18004 17222
rect 18052 17274 18108 17276
rect 18052 17222 18054 17274
rect 18054 17222 18106 17274
rect 18106 17222 18108 17274
rect 18052 17220 18108 17222
rect 17836 17106 17892 17108
rect 17836 17054 17838 17106
rect 17838 17054 17890 17106
rect 17890 17054 17892 17106
rect 17836 17052 17892 17054
rect 18732 17276 18788 17332
rect 18396 16716 18452 16772
rect 17724 16044 17780 16100
rect 17844 15706 17900 15708
rect 17844 15654 17846 15706
rect 17846 15654 17898 15706
rect 17898 15654 17900 15706
rect 17844 15652 17900 15654
rect 17948 15706 18004 15708
rect 17948 15654 17950 15706
rect 17950 15654 18002 15706
rect 18002 15654 18004 15706
rect 17948 15652 18004 15654
rect 18052 15706 18108 15708
rect 18052 15654 18054 15706
rect 18054 15654 18106 15706
rect 18106 15654 18108 15706
rect 18052 15652 18108 15654
rect 17836 15538 17892 15540
rect 17836 15486 17838 15538
rect 17838 15486 17890 15538
rect 17890 15486 17892 15538
rect 17836 15484 17892 15486
rect 19516 17612 19572 17668
rect 21420 21756 21476 21812
rect 22002 22762 22058 22764
rect 22002 22710 22004 22762
rect 22004 22710 22056 22762
rect 22056 22710 22058 22762
rect 22002 22708 22058 22710
rect 22106 22762 22162 22764
rect 22106 22710 22108 22762
rect 22108 22710 22160 22762
rect 22160 22710 22162 22762
rect 22106 22708 22162 22710
rect 22210 22762 22266 22764
rect 22210 22710 22212 22762
rect 22212 22710 22264 22762
rect 22264 22710 22266 22762
rect 22210 22708 22266 22710
rect 21868 21810 21924 21812
rect 21868 21758 21870 21810
rect 21870 21758 21922 21810
rect 21922 21758 21924 21810
rect 21868 21756 21924 21758
rect 20076 20802 20132 20804
rect 20076 20750 20078 20802
rect 20078 20750 20130 20802
rect 20130 20750 20132 20802
rect 20076 20748 20132 20750
rect 20692 20524 20748 20580
rect 19964 19068 20020 19124
rect 20300 18508 20356 18564
rect 21644 20972 21700 21028
rect 21364 20802 21420 20804
rect 21364 20750 21366 20802
rect 21366 20750 21418 20802
rect 21418 20750 21420 20802
rect 21364 20748 21420 20750
rect 22988 24444 23044 24500
rect 25340 30882 25396 30884
rect 25340 30830 25342 30882
rect 25342 30830 25394 30882
rect 25394 30830 25396 30882
rect 25340 30828 25396 30830
rect 24668 30210 24724 30212
rect 24668 30158 24670 30210
rect 24670 30158 24722 30210
rect 24722 30158 24724 30210
rect 24668 30156 24724 30158
rect 25172 30098 25228 30100
rect 25172 30046 25174 30098
rect 25174 30046 25226 30098
rect 25226 30046 25228 30098
rect 25172 30044 25228 30046
rect 24892 29932 24948 29988
rect 25228 29484 25284 29540
rect 25900 29932 25956 29988
rect 25452 29372 25508 29428
rect 24556 28588 24612 28644
rect 24780 28700 24836 28756
rect 25228 28642 25284 28644
rect 25228 28590 25230 28642
rect 25230 28590 25282 28642
rect 25282 28590 25284 28642
rect 25228 28588 25284 28590
rect 26160 29818 26216 29820
rect 26160 29766 26162 29818
rect 26162 29766 26214 29818
rect 26214 29766 26216 29818
rect 26160 29764 26216 29766
rect 26264 29818 26320 29820
rect 26264 29766 26266 29818
rect 26266 29766 26318 29818
rect 26318 29766 26320 29818
rect 26264 29764 26320 29766
rect 26368 29818 26424 29820
rect 26368 29766 26370 29818
rect 26370 29766 26422 29818
rect 26422 29766 26424 29818
rect 26368 29764 26424 29766
rect 30318 30602 30374 30604
rect 30318 30550 30320 30602
rect 30320 30550 30372 30602
rect 30372 30550 30374 30602
rect 30318 30548 30374 30550
rect 30422 30602 30478 30604
rect 30422 30550 30424 30602
rect 30424 30550 30476 30602
rect 30476 30550 30478 30602
rect 30422 30548 30478 30550
rect 30526 30602 30582 30604
rect 30526 30550 30528 30602
rect 30528 30550 30580 30602
rect 30580 30550 30582 30602
rect 30526 30548 30582 30550
rect 26796 29484 26852 29540
rect 26012 28700 26068 28756
rect 26684 28700 26740 28756
rect 26160 28250 26216 28252
rect 26160 28198 26162 28250
rect 26162 28198 26214 28250
rect 26214 28198 26216 28250
rect 26160 28196 26216 28198
rect 26264 28250 26320 28252
rect 26264 28198 26266 28250
rect 26266 28198 26318 28250
rect 26318 28198 26320 28250
rect 26264 28196 26320 28198
rect 26368 28250 26424 28252
rect 26368 28198 26370 28250
rect 26370 28198 26422 28250
rect 26422 28198 26424 28250
rect 26368 28196 26424 28198
rect 27580 29426 27636 29428
rect 27580 29374 27582 29426
rect 27582 29374 27634 29426
rect 27634 29374 27636 29426
rect 27580 29372 27636 29374
rect 29036 29372 29092 29428
rect 27356 28700 27412 28756
rect 27860 28530 27916 28532
rect 27860 28478 27862 28530
rect 27862 28478 27914 28530
rect 27914 28478 27916 28530
rect 27860 28476 27916 28478
rect 28700 28476 28756 28532
rect 23996 25506 24052 25508
rect 23996 25454 23998 25506
rect 23998 25454 24050 25506
rect 24050 25454 24052 25506
rect 23996 25452 24052 25454
rect 24556 25564 24612 25620
rect 23548 25004 23604 25060
rect 23324 24892 23380 24948
rect 23436 24668 23492 24724
rect 23212 24444 23268 24500
rect 22428 21756 22484 21812
rect 21980 21308 22036 21364
rect 22002 21194 22058 21196
rect 22002 21142 22004 21194
rect 22004 21142 22056 21194
rect 22056 21142 22058 21194
rect 22002 21140 22058 21142
rect 22106 21194 22162 21196
rect 22106 21142 22108 21194
rect 22108 21142 22160 21194
rect 22160 21142 22162 21194
rect 22106 21140 22162 21142
rect 22210 21194 22266 21196
rect 22210 21142 22212 21194
rect 22212 21142 22264 21194
rect 22264 21142 22266 21194
rect 22210 21140 22266 21142
rect 22764 22370 22820 22372
rect 22764 22318 22766 22370
rect 22766 22318 22818 22370
rect 22818 22318 22820 22370
rect 22764 22316 22820 22318
rect 22876 21980 22932 22036
rect 23660 24444 23716 24500
rect 24444 25004 24500 25060
rect 24332 24780 24388 24836
rect 23996 24556 24052 24612
rect 24836 24780 24892 24836
rect 26160 26682 26216 26684
rect 26160 26630 26162 26682
rect 26162 26630 26214 26682
rect 26214 26630 26216 26682
rect 26160 26628 26216 26630
rect 26264 26682 26320 26684
rect 26264 26630 26266 26682
rect 26266 26630 26318 26682
rect 26318 26630 26320 26682
rect 26264 26628 26320 26630
rect 26368 26682 26424 26684
rect 26368 26630 26370 26682
rect 26370 26630 26422 26682
rect 26422 26630 26424 26682
rect 26368 26628 26424 26630
rect 27580 28140 27636 28196
rect 28476 28140 28532 28196
rect 28364 27858 28420 27860
rect 28364 27806 28366 27858
rect 28366 27806 28418 27858
rect 28418 27806 28420 27858
rect 28364 27804 28420 27806
rect 27804 27186 27860 27188
rect 27804 27134 27806 27186
rect 27806 27134 27858 27186
rect 27858 27134 27860 27186
rect 27804 27132 27860 27134
rect 27580 26012 27636 26068
rect 28924 27858 28980 27860
rect 28924 27806 28926 27858
rect 28926 27806 28978 27858
rect 28978 27806 28980 27858
rect 28924 27804 28980 27806
rect 28476 27132 28532 27188
rect 28140 26012 28196 26068
rect 28252 26348 28308 26404
rect 26160 25114 26216 25116
rect 26160 25062 26162 25114
rect 26162 25062 26214 25114
rect 26214 25062 26216 25114
rect 26160 25060 26216 25062
rect 26264 25114 26320 25116
rect 26264 25062 26266 25114
rect 26266 25062 26318 25114
rect 26318 25062 26320 25114
rect 26264 25060 26320 25062
rect 26368 25114 26424 25116
rect 26368 25062 26370 25114
rect 26370 25062 26422 25114
rect 26422 25062 26424 25114
rect 26368 25060 26424 25062
rect 26236 24892 26292 24948
rect 25004 24668 25060 24724
rect 23660 23996 23716 24052
rect 24332 24050 24388 24052
rect 24332 23998 24334 24050
rect 24334 23998 24386 24050
rect 24386 23998 24388 24050
rect 24332 23996 24388 23998
rect 25452 23996 25508 24052
rect 27356 24892 27412 24948
rect 27020 24780 27076 24836
rect 26740 24444 26796 24500
rect 26796 23884 26852 23940
rect 26160 23546 26216 23548
rect 26160 23494 26162 23546
rect 26162 23494 26214 23546
rect 26214 23494 26216 23546
rect 26160 23492 26216 23494
rect 26264 23546 26320 23548
rect 26264 23494 26266 23546
rect 26266 23494 26318 23546
rect 26318 23494 26320 23546
rect 26264 23492 26320 23494
rect 26368 23546 26424 23548
rect 26368 23494 26370 23546
rect 26370 23494 26422 23546
rect 26422 23494 26424 23546
rect 26368 23492 26424 23494
rect 28140 25452 28196 25508
rect 28028 25340 28084 25396
rect 28588 26348 28644 26404
rect 29372 26348 29428 26404
rect 27580 24780 27636 24836
rect 27188 24444 27244 24500
rect 27244 23938 27300 23940
rect 27244 23886 27246 23938
rect 27246 23886 27298 23938
rect 27298 23886 27300 23938
rect 27244 23884 27300 23886
rect 27692 24444 27748 24500
rect 28252 24444 28308 24500
rect 28924 26012 28980 26068
rect 29260 25394 29316 25396
rect 29260 25342 29262 25394
rect 29262 25342 29314 25394
rect 29314 25342 29316 25394
rect 29260 25340 29316 25342
rect 28476 23884 28532 23940
rect 29036 23938 29092 23940
rect 29036 23886 29038 23938
rect 29038 23886 29090 23938
rect 29090 23886 29092 23938
rect 29036 23884 29092 23886
rect 23156 21980 23212 22036
rect 22932 21474 22988 21476
rect 22932 21422 22934 21474
rect 22934 21422 22986 21474
rect 22986 21422 22988 21474
rect 22932 21420 22988 21422
rect 23324 21868 23380 21924
rect 22988 21196 23044 21252
rect 22876 20972 22932 21028
rect 22092 20802 22148 20804
rect 21756 20636 21812 20692
rect 22092 20750 22094 20802
rect 22094 20750 22146 20802
rect 22146 20750 22148 20802
rect 22092 20748 22148 20750
rect 22092 20524 22148 20580
rect 21532 19906 21588 19908
rect 21532 19854 21534 19906
rect 21534 19854 21586 19906
rect 21586 19854 21588 19906
rect 21532 19852 21588 19854
rect 20748 18396 20804 18452
rect 19740 17554 19796 17556
rect 19740 17502 19742 17554
rect 19742 17502 19794 17554
rect 19794 17502 19796 17554
rect 19740 17500 19796 17502
rect 20188 17836 20244 17892
rect 19908 17164 19964 17220
rect 20076 17276 20132 17332
rect 19292 16604 19348 16660
rect 19516 16098 19572 16100
rect 19516 16046 19518 16098
rect 19518 16046 19570 16098
rect 19570 16046 19572 16098
rect 19516 16044 19572 16046
rect 18340 15372 18396 15428
rect 18844 15484 18900 15540
rect 17724 14252 17780 14308
rect 18172 14306 18228 14308
rect 18172 14254 18174 14306
rect 18174 14254 18226 14306
rect 18226 14254 18228 14306
rect 18172 14252 18228 14254
rect 17844 14138 17900 14140
rect 17844 14086 17846 14138
rect 17846 14086 17898 14138
rect 17898 14086 17900 14138
rect 17844 14084 17900 14086
rect 17948 14138 18004 14140
rect 17948 14086 17950 14138
rect 17950 14086 18002 14138
rect 18002 14086 18004 14138
rect 17948 14084 18004 14086
rect 18052 14138 18108 14140
rect 18052 14086 18054 14138
rect 18054 14086 18106 14138
rect 18106 14086 18108 14138
rect 18052 14084 18108 14086
rect 17836 13858 17892 13860
rect 17836 13806 17838 13858
rect 17838 13806 17890 13858
rect 17890 13806 17892 13858
rect 17836 13804 17892 13806
rect 18004 13746 18060 13748
rect 18004 13694 18006 13746
rect 18006 13694 18058 13746
rect 18058 13694 18060 13746
rect 18004 13692 18060 13694
rect 17724 13468 17780 13524
rect 17500 12908 17556 12964
rect 17388 12178 17444 12180
rect 17388 12126 17390 12178
rect 17390 12126 17442 12178
rect 17442 12126 17444 12178
rect 17388 12124 17444 12126
rect 17276 9212 17332 9268
rect 17892 12796 17948 12852
rect 18172 12796 18228 12852
rect 18284 12684 18340 12740
rect 17844 12570 17900 12572
rect 17844 12518 17846 12570
rect 17846 12518 17898 12570
rect 17898 12518 17900 12570
rect 17844 12516 17900 12518
rect 17948 12570 18004 12572
rect 17948 12518 17950 12570
rect 17950 12518 18002 12570
rect 18002 12518 18004 12570
rect 17948 12516 18004 12518
rect 18052 12570 18108 12572
rect 18052 12518 18054 12570
rect 18054 12518 18106 12570
rect 18106 12518 18108 12570
rect 18052 12516 18108 12518
rect 18060 12178 18116 12180
rect 18060 12126 18062 12178
rect 18062 12126 18114 12178
rect 18114 12126 18116 12178
rect 18060 12124 18116 12126
rect 17668 11394 17724 11396
rect 17668 11342 17670 11394
rect 17670 11342 17722 11394
rect 17722 11342 17724 11394
rect 17668 11340 17724 11342
rect 17844 11002 17900 11004
rect 17844 10950 17846 11002
rect 17846 10950 17898 11002
rect 17898 10950 17900 11002
rect 17844 10948 17900 10950
rect 17948 11002 18004 11004
rect 17948 10950 17950 11002
rect 17950 10950 18002 11002
rect 18002 10950 18004 11002
rect 17948 10948 18004 10950
rect 18052 11002 18108 11004
rect 18052 10950 18054 11002
rect 18054 10950 18106 11002
rect 18106 10950 18108 11002
rect 18052 10948 18108 10950
rect 18508 13692 18564 13748
rect 18564 13522 18620 13524
rect 18564 13470 18566 13522
rect 18566 13470 18618 13522
rect 18618 13470 18620 13522
rect 18564 13468 18620 13470
rect 20636 17890 20692 17892
rect 20636 17838 20638 17890
rect 20638 17838 20690 17890
rect 20690 17838 20692 17890
rect 20636 17836 20692 17838
rect 20300 17724 20356 17780
rect 21980 19852 22036 19908
rect 22316 20748 22372 20804
rect 22596 20802 22652 20804
rect 22596 20750 22598 20802
rect 22598 20750 22650 20802
rect 22650 20750 22652 20802
rect 22596 20748 22652 20750
rect 22764 20690 22820 20692
rect 22764 20638 22766 20690
rect 22766 20638 22818 20690
rect 22818 20638 22820 20690
rect 22764 20636 22820 20638
rect 22428 20524 22484 20580
rect 22540 20412 22596 20468
rect 22540 19964 22596 20020
rect 22988 20188 23044 20244
rect 25284 22316 25340 22372
rect 23884 21868 23940 21924
rect 23548 21756 23604 21812
rect 23772 21420 23828 21476
rect 34476 29818 34532 29820
rect 34476 29766 34478 29818
rect 34478 29766 34530 29818
rect 34530 29766 34532 29818
rect 34476 29764 34532 29766
rect 34580 29818 34636 29820
rect 34580 29766 34582 29818
rect 34582 29766 34634 29818
rect 34634 29766 34636 29818
rect 34580 29764 34636 29766
rect 34684 29818 34740 29820
rect 34684 29766 34686 29818
rect 34686 29766 34738 29818
rect 34738 29766 34740 29818
rect 34684 29764 34740 29766
rect 30318 29034 30374 29036
rect 30318 28982 30320 29034
rect 30320 28982 30372 29034
rect 30372 28982 30374 29034
rect 30318 28980 30374 28982
rect 30422 29034 30478 29036
rect 30422 28982 30424 29034
rect 30424 28982 30476 29034
rect 30476 28982 30478 29034
rect 30422 28980 30478 28982
rect 30526 29034 30582 29036
rect 30526 28982 30528 29034
rect 30528 28982 30580 29034
rect 30580 28982 30582 29034
rect 30526 28980 30582 28982
rect 34476 28250 34532 28252
rect 34476 28198 34478 28250
rect 34478 28198 34530 28250
rect 34530 28198 34532 28250
rect 34476 28196 34532 28198
rect 34580 28250 34636 28252
rect 34580 28198 34582 28250
rect 34582 28198 34634 28250
rect 34634 28198 34636 28250
rect 34580 28196 34636 28198
rect 34684 28250 34740 28252
rect 34684 28198 34686 28250
rect 34686 28198 34738 28250
rect 34738 28198 34740 28250
rect 34684 28196 34740 28198
rect 30318 27466 30374 27468
rect 30318 27414 30320 27466
rect 30320 27414 30372 27466
rect 30372 27414 30374 27466
rect 30318 27412 30374 27414
rect 30422 27466 30478 27468
rect 30422 27414 30424 27466
rect 30424 27414 30476 27466
rect 30476 27414 30478 27466
rect 30422 27412 30478 27414
rect 30526 27466 30582 27468
rect 30526 27414 30528 27466
rect 30528 27414 30580 27466
rect 30580 27414 30582 27466
rect 30526 27412 30582 27414
rect 34476 26682 34532 26684
rect 34476 26630 34478 26682
rect 34478 26630 34530 26682
rect 34530 26630 34532 26682
rect 34476 26628 34532 26630
rect 34580 26682 34636 26684
rect 34580 26630 34582 26682
rect 34582 26630 34634 26682
rect 34634 26630 34636 26682
rect 34580 26628 34636 26630
rect 34684 26682 34740 26684
rect 34684 26630 34686 26682
rect 34686 26630 34738 26682
rect 34738 26630 34740 26682
rect 34684 26628 34740 26630
rect 29652 26066 29708 26068
rect 29652 26014 29654 26066
rect 29654 26014 29706 26066
rect 29706 26014 29708 26066
rect 29652 26012 29708 26014
rect 30318 25898 30374 25900
rect 30318 25846 30320 25898
rect 30320 25846 30372 25898
rect 30372 25846 30374 25898
rect 30318 25844 30374 25846
rect 30422 25898 30478 25900
rect 30422 25846 30424 25898
rect 30424 25846 30476 25898
rect 30476 25846 30478 25898
rect 30422 25844 30478 25846
rect 30526 25898 30582 25900
rect 30526 25846 30528 25898
rect 30528 25846 30580 25898
rect 30580 25846 30582 25898
rect 30526 25844 30582 25846
rect 29708 25452 29764 25508
rect 31164 25506 31220 25508
rect 31164 25454 31166 25506
rect 31166 25454 31218 25506
rect 31218 25454 31220 25506
rect 31164 25452 31220 25454
rect 30318 24330 30374 24332
rect 30318 24278 30320 24330
rect 30320 24278 30372 24330
rect 30372 24278 30374 24330
rect 30318 24276 30374 24278
rect 30422 24330 30478 24332
rect 30422 24278 30424 24330
rect 30424 24278 30476 24330
rect 30476 24278 30478 24330
rect 30422 24276 30478 24278
rect 30526 24330 30582 24332
rect 30526 24278 30528 24330
rect 30528 24278 30580 24330
rect 30580 24278 30582 24330
rect 30526 24276 30582 24278
rect 30318 22762 30374 22764
rect 30318 22710 30320 22762
rect 30320 22710 30372 22762
rect 30372 22710 30374 22762
rect 30318 22708 30374 22710
rect 30422 22762 30478 22764
rect 30422 22710 30424 22762
rect 30424 22710 30476 22762
rect 30476 22710 30478 22762
rect 30422 22708 30478 22710
rect 30526 22762 30582 22764
rect 30526 22710 30528 22762
rect 30528 22710 30580 22762
rect 30580 22710 30582 22762
rect 30526 22708 30582 22710
rect 26160 21978 26216 21980
rect 26160 21926 26162 21978
rect 26162 21926 26214 21978
rect 26214 21926 26216 21978
rect 26160 21924 26216 21926
rect 26264 21978 26320 21980
rect 26264 21926 26266 21978
rect 26266 21926 26318 21978
rect 26318 21926 26320 21978
rect 26264 21924 26320 21926
rect 26368 21978 26424 21980
rect 26368 21926 26370 21978
rect 26370 21926 26422 21978
rect 26422 21926 26424 21978
rect 26368 21924 26424 21926
rect 25788 21756 25844 21812
rect 26460 21756 26516 21812
rect 25564 21420 25620 21476
rect 23324 20412 23380 20468
rect 23884 20300 23940 20356
rect 26124 20802 26180 20804
rect 26124 20750 26126 20802
rect 26126 20750 26178 20802
rect 26178 20750 26180 20802
rect 26124 20748 26180 20750
rect 29092 20972 29148 21028
rect 26684 20802 26740 20804
rect 26684 20750 26686 20802
rect 26686 20750 26738 20802
rect 26738 20750 26740 20802
rect 26684 20748 26740 20750
rect 27748 20802 27804 20804
rect 27748 20750 27750 20802
rect 27750 20750 27802 20802
rect 27802 20750 27804 20802
rect 27748 20748 27804 20750
rect 24220 20300 24276 20356
rect 26160 20410 26216 20412
rect 26160 20358 26162 20410
rect 26162 20358 26214 20410
rect 26214 20358 26216 20410
rect 26160 20356 26216 20358
rect 26264 20410 26320 20412
rect 26264 20358 26266 20410
rect 26266 20358 26318 20410
rect 26318 20358 26320 20410
rect 26264 20356 26320 20358
rect 26368 20410 26424 20412
rect 26368 20358 26370 20410
rect 26370 20358 26422 20410
rect 26422 20358 26424 20410
rect 26368 20356 26424 20358
rect 22002 19626 22058 19628
rect 22002 19574 22004 19626
rect 22004 19574 22056 19626
rect 22056 19574 22058 19626
rect 22002 19572 22058 19574
rect 22106 19626 22162 19628
rect 22106 19574 22108 19626
rect 22108 19574 22160 19626
rect 22160 19574 22162 19626
rect 22106 19572 22162 19574
rect 22210 19626 22266 19628
rect 22210 19574 22212 19626
rect 22212 19574 22264 19626
rect 22264 19574 22266 19626
rect 22210 19572 22266 19574
rect 20972 19180 21028 19236
rect 21364 19180 21420 19236
rect 22204 19180 22260 19236
rect 20860 17948 20916 18004
rect 22428 18450 22484 18452
rect 22428 18398 22430 18450
rect 22430 18398 22482 18450
rect 22482 18398 22484 18450
rect 22428 18396 22484 18398
rect 21084 17724 21140 17780
rect 22002 18058 22058 18060
rect 22002 18006 22004 18058
rect 22004 18006 22056 18058
rect 22056 18006 22058 18058
rect 22002 18004 22058 18006
rect 22106 18058 22162 18060
rect 22106 18006 22108 18058
rect 22108 18006 22160 18058
rect 22160 18006 22162 18058
rect 22106 18004 22162 18006
rect 22210 18058 22266 18060
rect 22210 18006 22212 18058
rect 22212 18006 22264 18058
rect 22264 18006 22266 18058
rect 22210 18004 22266 18006
rect 20748 16828 20804 16884
rect 19068 15148 19124 15204
rect 18956 13580 19012 13636
rect 18508 12962 18564 12964
rect 18508 12910 18510 12962
rect 18510 12910 18562 12962
rect 18562 12910 18564 12962
rect 18508 12908 18564 12910
rect 18956 13020 19012 13076
rect 18676 12348 18732 12404
rect 18844 12684 18900 12740
rect 18620 12012 18676 12068
rect 18732 12124 18788 12180
rect 18732 11788 18788 11844
rect 18956 12236 19012 12292
rect 18956 11788 19012 11844
rect 17836 9938 17892 9940
rect 17836 9886 17838 9938
rect 17838 9886 17890 9938
rect 17890 9886 17892 9938
rect 17836 9884 17892 9886
rect 17844 9434 17900 9436
rect 17844 9382 17846 9434
rect 17846 9382 17898 9434
rect 17898 9382 17900 9434
rect 17844 9380 17900 9382
rect 17948 9434 18004 9436
rect 17948 9382 17950 9434
rect 17950 9382 18002 9434
rect 18002 9382 18004 9434
rect 17948 9380 18004 9382
rect 18052 9434 18108 9436
rect 18052 9382 18054 9434
rect 18054 9382 18106 9434
rect 18106 9382 18108 9434
rect 18052 9380 18108 9382
rect 18172 9212 18228 9268
rect 16156 7420 16212 7476
rect 15484 6412 15540 6468
rect 15932 6636 15988 6692
rect 17052 8258 17108 8260
rect 17052 8206 17054 8258
rect 17054 8206 17106 8258
rect 17106 8206 17108 8258
rect 17052 8204 17108 8206
rect 16268 6748 16324 6804
rect 16884 6466 16940 6468
rect 16884 6414 16886 6466
rect 16886 6414 16938 6466
rect 16938 6414 16940 6466
rect 16884 6412 16940 6414
rect 16436 6076 16492 6132
rect 17052 5964 17108 6020
rect 16716 5906 16772 5908
rect 16716 5854 16718 5906
rect 16718 5854 16770 5906
rect 16770 5854 16772 5906
rect 16716 5852 16772 5854
rect 15260 5404 15316 5460
rect 16492 5122 16548 5124
rect 16492 5070 16494 5122
rect 16494 5070 16546 5122
rect 16546 5070 16548 5122
rect 16492 5068 16548 5070
rect 17844 7866 17900 7868
rect 17844 7814 17846 7866
rect 17846 7814 17898 7866
rect 17898 7814 17900 7866
rect 17844 7812 17900 7814
rect 17948 7866 18004 7868
rect 17948 7814 17950 7866
rect 17950 7814 18002 7866
rect 18002 7814 18004 7866
rect 17948 7812 18004 7814
rect 18052 7866 18108 7868
rect 18052 7814 18054 7866
rect 18054 7814 18106 7866
rect 18106 7814 18108 7866
rect 18052 7812 18108 7814
rect 17388 6636 17444 6692
rect 18004 6690 18060 6692
rect 18004 6638 18006 6690
rect 18006 6638 18058 6690
rect 18058 6638 18060 6690
rect 18004 6636 18060 6638
rect 17844 6298 17900 6300
rect 17844 6246 17846 6298
rect 17846 6246 17898 6298
rect 17898 6246 17900 6298
rect 17844 6244 17900 6246
rect 17948 6298 18004 6300
rect 17948 6246 17950 6298
rect 17950 6246 18002 6298
rect 18002 6246 18004 6298
rect 17948 6244 18004 6246
rect 18052 6298 18108 6300
rect 18052 6246 18054 6298
rect 18054 6246 18106 6298
rect 18106 6246 18108 6298
rect 18052 6244 18108 6246
rect 17276 6076 17332 6132
rect 18060 5964 18116 6020
rect 17164 5852 17220 5908
rect 17836 5852 17892 5908
rect 18172 5740 18228 5796
rect 18060 5180 18116 5236
rect 17844 4730 17900 4732
rect 17844 4678 17846 4730
rect 17846 4678 17898 4730
rect 17898 4678 17900 4730
rect 17844 4676 17900 4678
rect 17948 4730 18004 4732
rect 17948 4678 17950 4730
rect 17950 4678 18002 4730
rect 18002 4678 18004 4730
rect 17948 4676 18004 4678
rect 18052 4730 18108 4732
rect 18052 4678 18054 4730
rect 18054 4678 18106 4730
rect 18106 4678 18108 4730
rect 18052 4676 18108 4678
rect 14812 4338 14868 4340
rect 14812 4286 14814 4338
rect 14814 4286 14866 4338
rect 14866 4286 14868 4338
rect 14812 4284 14868 4286
rect 16828 4284 16884 4340
rect 17836 4338 17892 4340
rect 17836 4286 17838 4338
rect 17838 4286 17890 4338
rect 17890 4286 17892 4338
rect 17836 4284 17892 4286
rect 18172 4508 18228 4564
rect 21196 17052 21252 17108
rect 21308 17164 21364 17220
rect 22764 19964 22820 20020
rect 23884 19234 23940 19236
rect 23884 19182 23886 19234
rect 23886 19182 23938 19234
rect 23938 19182 23940 19234
rect 23884 19180 23940 19182
rect 27020 20018 27076 20020
rect 27020 19966 27022 20018
rect 27022 19966 27074 20018
rect 27074 19966 27076 20018
rect 27020 19964 27076 19966
rect 26160 18842 26216 18844
rect 26160 18790 26162 18842
rect 26162 18790 26214 18842
rect 26214 18790 26216 18842
rect 26160 18788 26216 18790
rect 26264 18842 26320 18844
rect 26264 18790 26266 18842
rect 26266 18790 26318 18842
rect 26318 18790 26320 18842
rect 26264 18788 26320 18790
rect 26368 18842 26424 18844
rect 26368 18790 26370 18842
rect 26370 18790 26422 18842
rect 26422 18790 26424 18842
rect 26368 18788 26424 18790
rect 22764 17948 22820 18004
rect 22652 17836 22708 17892
rect 22764 17500 22820 17556
rect 22484 17276 22540 17332
rect 27132 18284 27188 18340
rect 21308 16940 21364 16996
rect 22988 17948 23044 18004
rect 23156 17500 23212 17556
rect 21980 16882 22036 16884
rect 21980 16830 21982 16882
rect 21982 16830 22034 16882
rect 22034 16830 22036 16882
rect 21980 16828 22036 16830
rect 21532 16268 21588 16324
rect 22002 16490 22058 16492
rect 22002 16438 22004 16490
rect 22004 16438 22056 16490
rect 22056 16438 22058 16490
rect 22002 16436 22058 16438
rect 22106 16490 22162 16492
rect 22106 16438 22108 16490
rect 22108 16438 22160 16490
rect 22160 16438 22162 16490
rect 22106 16436 22162 16438
rect 22210 16490 22266 16492
rect 22210 16438 22212 16490
rect 22212 16438 22264 16490
rect 22264 16438 22266 16490
rect 22210 16436 22266 16438
rect 22856 16716 22912 16772
rect 25452 17612 25508 17668
rect 23604 16940 23660 16996
rect 23436 16882 23492 16884
rect 23436 16830 23438 16882
rect 23438 16830 23490 16882
rect 23490 16830 23492 16882
rect 23436 16828 23492 16830
rect 23324 16716 23380 16772
rect 24220 16716 24276 16772
rect 22316 16268 22372 16324
rect 21532 15148 21588 15204
rect 22372 15202 22428 15204
rect 22372 15150 22374 15202
rect 22374 15150 22426 15202
rect 22426 15150 22428 15202
rect 22372 15148 22428 15150
rect 22002 14922 22058 14924
rect 22002 14870 22004 14922
rect 22004 14870 22056 14922
rect 22056 14870 22058 14922
rect 22002 14868 22058 14870
rect 22106 14922 22162 14924
rect 22106 14870 22108 14922
rect 22108 14870 22160 14922
rect 22160 14870 22162 14922
rect 22106 14868 22162 14870
rect 22210 14922 22266 14924
rect 22210 14870 22212 14922
rect 22212 14870 22264 14922
rect 22264 14870 22266 14922
rect 22210 14868 22266 14870
rect 22002 13354 22058 13356
rect 22002 13302 22004 13354
rect 22004 13302 22056 13354
rect 22056 13302 22058 13354
rect 22002 13300 22058 13302
rect 22106 13354 22162 13356
rect 22106 13302 22108 13354
rect 22108 13302 22160 13354
rect 22160 13302 22162 13354
rect 22106 13300 22162 13302
rect 22210 13354 22266 13356
rect 22210 13302 22212 13354
rect 22212 13302 22264 13354
rect 22264 13302 22266 13354
rect 22210 13300 22266 13302
rect 21308 13132 21364 13188
rect 20188 12908 20244 12964
rect 19684 12796 19740 12852
rect 19516 12236 19572 12292
rect 21532 12962 21588 12964
rect 21532 12910 21534 12962
rect 21534 12910 21586 12962
rect 21586 12910 21588 12962
rect 21532 12908 21588 12910
rect 22408 12962 22464 12964
rect 22408 12910 22410 12962
rect 22410 12910 22462 12962
rect 22462 12910 22464 12962
rect 22408 12908 22464 12910
rect 19404 11564 19460 11620
rect 19516 8428 19572 8484
rect 22002 11786 22058 11788
rect 22002 11734 22004 11786
rect 22004 11734 22056 11786
rect 22056 11734 22058 11786
rect 22002 11732 22058 11734
rect 22106 11786 22162 11788
rect 22106 11734 22108 11786
rect 22108 11734 22160 11786
rect 22160 11734 22162 11786
rect 22106 11732 22162 11734
rect 22210 11786 22266 11788
rect 22210 11734 22212 11786
rect 22212 11734 22264 11786
rect 22264 11734 22266 11786
rect 22210 11732 22266 11734
rect 21308 9996 21364 10052
rect 25340 16044 25396 16100
rect 23436 15148 23492 15204
rect 22932 13970 22988 13972
rect 22932 13918 22934 13970
rect 22934 13918 22986 13970
rect 22986 13918 22988 13970
rect 22932 13916 22988 13918
rect 23212 13916 23268 13972
rect 23324 13692 23380 13748
rect 23100 13580 23156 13636
rect 22652 13186 22708 13188
rect 22652 13134 22654 13186
rect 22654 13134 22706 13186
rect 22706 13134 22708 13186
rect 22652 13132 22708 13134
rect 24780 15148 24836 15204
rect 25340 14364 25396 14420
rect 23436 13580 23492 13636
rect 22540 10892 22596 10948
rect 24164 13634 24220 13636
rect 24164 13582 24166 13634
rect 24166 13582 24218 13634
rect 24218 13582 24220 13634
rect 24164 13580 24220 13582
rect 25228 13468 25284 13524
rect 23884 13244 23940 13300
rect 23548 12908 23604 12964
rect 24220 12236 24276 12292
rect 26160 17274 26216 17276
rect 26160 17222 26162 17274
rect 26162 17222 26214 17274
rect 26214 17222 26216 17274
rect 26160 17220 26216 17222
rect 26264 17274 26320 17276
rect 26264 17222 26266 17274
rect 26266 17222 26318 17274
rect 26318 17222 26320 17274
rect 26264 17220 26320 17222
rect 26368 17274 26424 17276
rect 26368 17222 26370 17274
rect 26370 17222 26422 17274
rect 26422 17222 26424 17274
rect 26368 17220 26424 17222
rect 27132 17276 27188 17332
rect 27748 20188 27804 20244
rect 29148 20774 29204 20804
rect 29148 20748 29150 20774
rect 29150 20748 29202 20774
rect 29202 20748 29204 20774
rect 28476 20188 28532 20244
rect 28924 20076 28980 20132
rect 28028 19964 28084 20020
rect 27692 18450 27748 18452
rect 27692 18398 27694 18450
rect 27694 18398 27746 18450
rect 27746 18398 27748 18450
rect 27692 18396 27748 18398
rect 27580 17629 27636 17668
rect 27580 17612 27582 17629
rect 27582 17612 27634 17629
rect 27634 17612 27636 17629
rect 27778 17500 27834 17556
rect 27692 17276 27748 17332
rect 26908 16492 26964 16548
rect 26292 16322 26348 16324
rect 26292 16270 26294 16322
rect 26294 16270 26346 16322
rect 26346 16270 26348 16322
rect 26292 16268 26348 16270
rect 26124 16098 26180 16100
rect 26124 16046 26126 16098
rect 26126 16046 26178 16098
rect 26178 16046 26180 16098
rect 26124 16044 26180 16046
rect 26160 15706 26216 15708
rect 26160 15654 26162 15706
rect 26162 15654 26214 15706
rect 26214 15654 26216 15706
rect 26160 15652 26216 15654
rect 26264 15706 26320 15708
rect 26264 15654 26266 15706
rect 26266 15654 26318 15706
rect 26318 15654 26320 15706
rect 26264 15652 26320 15654
rect 26368 15706 26424 15708
rect 26368 15654 26370 15706
rect 26370 15654 26422 15706
rect 26422 15654 26424 15706
rect 26368 15652 26424 15654
rect 26908 15148 26964 15204
rect 27132 16604 27188 16660
rect 27132 16268 27188 16324
rect 27524 15932 27580 15988
rect 27580 15314 27636 15316
rect 27580 15262 27582 15314
rect 27582 15262 27634 15314
rect 27634 15262 27636 15314
rect 27580 15260 27636 15262
rect 27356 15148 27412 15204
rect 28812 19292 28868 19348
rect 29484 21586 29540 21588
rect 29484 21534 29486 21586
rect 29486 21534 29538 21586
rect 29538 21534 29540 21586
rect 29484 21532 29540 21534
rect 29932 21532 29988 21588
rect 30940 21756 30996 21812
rect 34476 25114 34532 25116
rect 34476 25062 34478 25114
rect 34478 25062 34530 25114
rect 34530 25062 34532 25114
rect 34476 25060 34532 25062
rect 34580 25114 34636 25116
rect 34580 25062 34582 25114
rect 34582 25062 34634 25114
rect 34634 25062 34636 25114
rect 34580 25060 34636 25062
rect 34684 25114 34740 25116
rect 34684 25062 34686 25114
rect 34686 25062 34738 25114
rect 34738 25062 34740 25114
rect 34684 25060 34740 25062
rect 34476 23546 34532 23548
rect 34476 23494 34478 23546
rect 34478 23494 34530 23546
rect 34530 23494 34532 23546
rect 34476 23492 34532 23494
rect 34580 23546 34636 23548
rect 34580 23494 34582 23546
rect 34582 23494 34634 23546
rect 34634 23494 34636 23546
rect 34580 23492 34636 23494
rect 34684 23546 34740 23548
rect 34684 23494 34686 23546
rect 34686 23494 34738 23546
rect 34738 23494 34740 23546
rect 34684 23492 34740 23494
rect 34476 21978 34532 21980
rect 34476 21926 34478 21978
rect 34478 21926 34530 21978
rect 34530 21926 34532 21978
rect 34476 21924 34532 21926
rect 34580 21978 34636 21980
rect 34580 21926 34582 21978
rect 34582 21926 34634 21978
rect 34634 21926 34636 21978
rect 34580 21924 34636 21926
rect 34684 21978 34740 21980
rect 34684 21926 34686 21978
rect 34686 21926 34738 21978
rect 34738 21926 34740 21978
rect 34684 21924 34740 21926
rect 30716 21420 30772 21476
rect 30318 21194 30374 21196
rect 30318 21142 30320 21194
rect 30320 21142 30372 21194
rect 30372 21142 30374 21194
rect 30318 21140 30374 21142
rect 30422 21194 30478 21196
rect 30422 21142 30424 21194
rect 30424 21142 30476 21194
rect 30476 21142 30478 21194
rect 30422 21140 30478 21142
rect 30526 21194 30582 21196
rect 30526 21142 30528 21194
rect 30528 21142 30580 21194
rect 30580 21142 30582 21194
rect 30526 21140 30582 21142
rect 30828 20748 30884 20804
rect 29596 19964 29652 20020
rect 29932 20076 29988 20132
rect 29372 19852 29428 19908
rect 29148 19346 29204 19348
rect 29148 19294 29150 19346
rect 29150 19294 29202 19346
rect 29202 19294 29204 19346
rect 29148 19292 29204 19294
rect 28028 16716 28084 16772
rect 28140 17612 28196 17668
rect 28700 18396 28756 18452
rect 28364 17612 28420 17668
rect 28476 17500 28532 17556
rect 28476 16828 28532 16884
rect 28588 17612 28644 17668
rect 29260 18172 29316 18228
rect 28924 16940 28980 16996
rect 28476 16604 28532 16660
rect 27972 16098 28028 16100
rect 27972 16046 27974 16098
rect 27974 16046 28026 16098
rect 28026 16046 28028 16098
rect 27972 16044 28028 16046
rect 27804 15708 27860 15764
rect 28532 15986 28588 15988
rect 28532 15934 28534 15986
rect 28534 15934 28586 15986
rect 28586 15934 28588 15986
rect 28532 15932 28588 15934
rect 28252 15484 28308 15540
rect 28700 15708 28756 15764
rect 27132 14588 27188 14644
rect 26031 14530 26087 14532
rect 26031 14478 26033 14530
rect 26033 14478 26085 14530
rect 26085 14478 26087 14530
rect 26031 14476 26087 14478
rect 25788 14418 25844 14420
rect 25788 14366 25790 14418
rect 25790 14366 25842 14418
rect 25842 14366 25844 14418
rect 25788 14364 25844 14366
rect 26160 14138 26216 14140
rect 26160 14086 26162 14138
rect 26162 14086 26214 14138
rect 26214 14086 26216 14138
rect 26160 14084 26216 14086
rect 26264 14138 26320 14140
rect 26264 14086 26266 14138
rect 26266 14086 26318 14138
rect 26318 14086 26320 14138
rect 26264 14084 26320 14086
rect 26368 14138 26424 14140
rect 26368 14086 26370 14138
rect 26370 14086 26422 14138
rect 26422 14086 26424 14138
rect 26368 14084 26424 14086
rect 26460 13804 26516 13860
rect 23324 10892 23380 10948
rect 22002 10218 22058 10220
rect 22002 10166 22004 10218
rect 22004 10166 22056 10218
rect 22056 10166 22058 10218
rect 22002 10164 22058 10166
rect 22106 10218 22162 10220
rect 22106 10166 22108 10218
rect 22108 10166 22160 10218
rect 22160 10166 22162 10218
rect 22106 10164 22162 10166
rect 22210 10218 22266 10220
rect 22210 10166 22212 10218
rect 22212 10166 22264 10218
rect 22264 10166 22266 10218
rect 22210 10164 22266 10166
rect 21868 9884 21924 9940
rect 21980 9772 22036 9828
rect 21868 8988 21924 9044
rect 22204 8930 22260 8932
rect 22204 8878 22206 8930
rect 22206 8878 22258 8930
rect 22258 8878 22260 8930
rect 22204 8876 22260 8878
rect 22002 8650 22058 8652
rect 22002 8598 22004 8650
rect 22004 8598 22056 8650
rect 22056 8598 22058 8650
rect 22002 8596 22058 8598
rect 22106 8650 22162 8652
rect 22106 8598 22108 8650
rect 22108 8598 22160 8650
rect 22160 8598 22162 8650
rect 22106 8596 22162 8598
rect 22210 8650 22266 8652
rect 22210 8598 22212 8650
rect 22212 8598 22264 8650
rect 22264 8598 22266 8650
rect 22210 8596 22266 8598
rect 22652 9996 22708 10052
rect 22876 10386 22932 10388
rect 22876 10334 22878 10386
rect 22878 10334 22930 10386
rect 22930 10334 22932 10386
rect 22876 10332 22932 10334
rect 23212 9996 23268 10052
rect 23100 9799 23156 9828
rect 23100 9772 23102 9799
rect 23102 9772 23154 9799
rect 23154 9772 23156 9799
rect 24332 11506 24388 11508
rect 24332 11454 24334 11506
rect 24334 11454 24386 11506
rect 24386 11454 24388 11506
rect 24332 11452 24388 11454
rect 23324 9884 23380 9940
rect 23940 9938 23996 9940
rect 23940 9886 23942 9938
rect 23942 9886 23994 9938
rect 23994 9886 23996 9938
rect 23940 9884 23996 9886
rect 24220 9548 24276 9604
rect 22652 8876 22708 8932
rect 22764 9042 22820 9044
rect 22764 8990 22766 9042
rect 22766 8990 22818 9042
rect 22818 8990 22820 9042
rect 22764 8988 22820 8990
rect 22428 8428 22484 8484
rect 22652 8428 22708 8484
rect 18396 6076 18452 6132
rect 19180 6636 19236 6692
rect 19068 6076 19124 6132
rect 18732 5852 18788 5908
rect 18912 5964 18968 6020
rect 18956 5740 19012 5796
rect 19516 6076 19572 6132
rect 19628 5906 19684 5908
rect 19068 5180 19124 5236
rect 18508 5122 18564 5124
rect 18508 5070 18510 5122
rect 18510 5070 18562 5122
rect 18562 5070 18564 5122
rect 18508 5068 18564 5070
rect 19628 5854 19630 5906
rect 19630 5854 19682 5906
rect 19682 5854 19684 5906
rect 19628 5852 19684 5854
rect 19348 5122 19404 5124
rect 19348 5070 19350 5122
rect 19350 5070 19402 5122
rect 19402 5070 19404 5122
rect 19348 5068 19404 5070
rect 19628 5180 19684 5236
rect 19908 6018 19964 6020
rect 19908 5966 19910 6018
rect 19910 5966 19962 6018
rect 19962 5966 19964 6018
rect 19908 5964 19964 5966
rect 22428 7980 22484 8036
rect 22092 7586 22148 7588
rect 22092 7534 22094 7586
rect 22094 7534 22146 7586
rect 22146 7534 22148 7586
rect 22092 7532 22148 7534
rect 22540 7532 22596 7588
rect 22002 7082 22058 7084
rect 22002 7030 22004 7082
rect 22004 7030 22056 7082
rect 22056 7030 22058 7082
rect 22002 7028 22058 7030
rect 22106 7082 22162 7084
rect 22106 7030 22108 7082
rect 22108 7030 22160 7082
rect 22160 7030 22162 7082
rect 22106 7028 22162 7030
rect 22210 7082 22266 7084
rect 22210 7030 22212 7082
rect 22212 7030 22264 7082
rect 22264 7030 22266 7082
rect 22210 7028 22266 7030
rect 21420 6748 21476 6804
rect 21756 6748 21812 6804
rect 21364 5740 21420 5796
rect 21532 5292 21588 5348
rect 22764 8370 22820 8372
rect 22764 8318 22766 8370
rect 22766 8318 22818 8370
rect 22818 8318 22820 8370
rect 22764 8316 22820 8318
rect 23100 8258 23156 8260
rect 23100 8206 23102 8258
rect 23102 8206 23154 8258
rect 23154 8206 23156 8258
rect 23100 8204 23156 8206
rect 22876 7980 22932 8036
rect 23044 7980 23100 8036
rect 22764 7532 22820 7588
rect 22876 7756 22932 7812
rect 23604 8428 23660 8484
rect 25452 11788 25508 11844
rect 25340 11506 25396 11508
rect 25340 11454 25342 11506
rect 25342 11454 25394 11506
rect 25394 11454 25396 11506
rect 25340 11452 25396 11454
rect 24724 11340 24780 11396
rect 25116 11394 25172 11396
rect 25116 11342 25118 11394
rect 25118 11342 25170 11394
rect 25170 11342 25172 11394
rect 25788 13468 25844 13524
rect 26460 13468 26516 13524
rect 26160 12570 26216 12572
rect 26160 12518 26162 12570
rect 26162 12518 26214 12570
rect 26214 12518 26216 12570
rect 26160 12516 26216 12518
rect 26264 12570 26320 12572
rect 26264 12518 26266 12570
rect 26266 12518 26318 12570
rect 26318 12518 26320 12570
rect 26264 12516 26320 12518
rect 26368 12570 26424 12572
rect 26368 12518 26370 12570
rect 26370 12518 26422 12570
rect 26422 12518 26424 12570
rect 26368 12516 26424 12518
rect 26124 11788 26180 11844
rect 26012 11564 26068 11620
rect 25116 11340 25172 11342
rect 25340 10573 25342 10612
rect 25342 10573 25394 10612
rect 25394 10573 25396 10612
rect 25340 10556 25396 10573
rect 24444 10444 24500 10500
rect 25228 10498 25284 10500
rect 25228 10446 25230 10498
rect 25230 10446 25282 10498
rect 25282 10446 25284 10498
rect 25228 10444 25284 10446
rect 25452 10332 25508 10388
rect 24780 9996 24836 10052
rect 25116 9602 25172 9604
rect 25116 9550 25118 9602
rect 25118 9550 25170 9602
rect 25170 9550 25172 9602
rect 25116 9548 25172 9550
rect 25116 8988 25172 9044
rect 23436 8092 23492 8148
rect 23604 7474 23660 7476
rect 23604 7422 23606 7474
rect 23606 7422 23658 7474
rect 23658 7422 23660 7474
rect 23604 7420 23660 7422
rect 23212 7084 23268 7140
rect 23212 6748 23268 6804
rect 22652 5964 22708 6020
rect 22316 5628 22372 5684
rect 22002 5514 22058 5516
rect 22002 5462 22004 5514
rect 22004 5462 22056 5514
rect 22056 5462 22058 5514
rect 22002 5460 22058 5462
rect 22106 5514 22162 5516
rect 22106 5462 22108 5514
rect 22108 5462 22160 5514
rect 22160 5462 22162 5514
rect 22106 5460 22162 5462
rect 22210 5514 22266 5516
rect 22210 5462 22212 5514
rect 22212 5462 22264 5514
rect 22264 5462 22266 5514
rect 22210 5460 22266 5462
rect 22316 5292 22372 5348
rect 22204 5083 22260 5124
rect 22204 5068 22206 5083
rect 22206 5068 22258 5083
rect 22258 5068 22260 5083
rect 18284 4172 18340 4228
rect 14700 3724 14756 3780
rect 11228 3388 11284 3444
rect 9528 3162 9584 3164
rect 9528 3110 9530 3162
rect 9530 3110 9582 3162
rect 9582 3110 9584 3162
rect 9528 3108 9584 3110
rect 9632 3162 9688 3164
rect 9632 3110 9634 3162
rect 9634 3110 9686 3162
rect 9686 3110 9688 3162
rect 9632 3108 9688 3110
rect 9736 3162 9792 3164
rect 9736 3110 9738 3162
rect 9738 3110 9790 3162
rect 9790 3110 9792 3162
rect 9736 3108 9792 3110
rect 17844 3162 17900 3164
rect 17844 3110 17846 3162
rect 17846 3110 17898 3162
rect 17898 3110 17900 3162
rect 17844 3108 17900 3110
rect 17948 3162 18004 3164
rect 17948 3110 17950 3162
rect 17950 3110 18002 3162
rect 18002 3110 18004 3162
rect 17948 3108 18004 3110
rect 18052 3162 18108 3164
rect 18052 3110 18054 3162
rect 18054 3110 18106 3162
rect 18106 3110 18108 3162
rect 18052 3108 18108 3110
rect 21420 3554 21476 3556
rect 21420 3502 21422 3554
rect 21422 3502 21474 3554
rect 21474 3502 21476 3554
rect 21420 3500 21476 3502
rect 22002 3946 22058 3948
rect 22002 3894 22004 3946
rect 22004 3894 22056 3946
rect 22056 3894 22058 3946
rect 22002 3892 22058 3894
rect 22106 3946 22162 3948
rect 22106 3894 22108 3946
rect 22108 3894 22160 3946
rect 22160 3894 22162 3946
rect 22106 3892 22162 3894
rect 22210 3946 22266 3948
rect 22210 3894 22212 3946
rect 22212 3894 22264 3946
rect 22264 3894 22266 3946
rect 22210 3892 22266 3894
rect 23212 6188 23268 6244
rect 24444 8316 24500 8372
rect 24108 7474 24164 7476
rect 24108 7422 24110 7474
rect 24110 7422 24162 7474
rect 24162 7422 24164 7474
rect 24108 7420 24164 7422
rect 24332 7420 24388 7476
rect 24444 6972 24500 7028
rect 25116 8092 25172 8148
rect 23996 6748 24052 6804
rect 23772 6188 23828 6244
rect 23884 6524 23940 6580
rect 23436 6076 23492 6132
rect 23212 5740 23268 5796
rect 23324 5964 23380 6020
rect 23436 5740 23492 5796
rect 24892 6076 24948 6132
rect 23772 5628 23828 5684
rect 23660 5068 23716 5124
rect 24220 5906 24276 5908
rect 24220 5854 24222 5906
rect 24222 5854 24274 5906
rect 24274 5854 24276 5906
rect 24220 5852 24276 5854
rect 24556 5682 24612 5684
rect 24556 5630 24558 5682
rect 24558 5630 24610 5682
rect 24610 5630 24612 5682
rect 24556 5628 24612 5630
rect 23324 4172 23380 4228
rect 21868 3500 21924 3556
rect 24108 4226 24164 4228
rect 24108 4174 24110 4226
rect 24110 4174 24162 4226
rect 24162 4174 24164 4226
rect 24108 4172 24164 4174
rect 25564 9005 25566 9044
rect 25566 9005 25618 9044
rect 25618 9005 25620 9044
rect 25564 8988 25620 9005
rect 25340 8204 25396 8260
rect 25900 11340 25956 11396
rect 26684 13580 26740 13636
rect 26908 13468 26964 13524
rect 26160 11002 26216 11004
rect 26160 10950 26162 11002
rect 26162 10950 26214 11002
rect 26214 10950 26216 11002
rect 26160 10948 26216 10950
rect 26264 11002 26320 11004
rect 26264 10950 26266 11002
rect 26266 10950 26318 11002
rect 26318 10950 26320 11002
rect 26264 10948 26320 10950
rect 26368 11002 26424 11004
rect 26368 10950 26370 11002
rect 26370 10950 26422 11002
rect 26422 10950 26424 11002
rect 26368 10948 26424 10950
rect 27132 11564 27188 11620
rect 26908 11340 26964 11396
rect 27356 14588 27412 14644
rect 27692 14530 27748 14532
rect 27692 14478 27694 14530
rect 27694 14478 27746 14530
rect 27746 14478 27748 14530
rect 27692 14476 27748 14478
rect 28476 15036 28532 15092
rect 28364 14588 28420 14644
rect 28924 15538 28980 15540
rect 28924 15486 28926 15538
rect 28926 15486 28978 15538
rect 28978 15486 28980 15538
rect 28924 15484 28980 15486
rect 29484 18396 29540 18452
rect 30604 20076 30660 20132
rect 31836 21474 31892 21476
rect 31836 21422 31838 21474
rect 31838 21422 31890 21474
rect 31890 21422 31892 21474
rect 31836 21420 31892 21422
rect 32340 21420 32396 21476
rect 31836 20972 31892 21028
rect 32060 20802 32116 20804
rect 32060 20750 32062 20802
rect 32062 20750 32114 20802
rect 32114 20750 32116 20802
rect 32060 20748 32116 20750
rect 34476 20410 34532 20412
rect 34476 20358 34478 20410
rect 34478 20358 34530 20410
rect 34530 20358 34532 20410
rect 34476 20356 34532 20358
rect 34580 20410 34636 20412
rect 34580 20358 34582 20410
rect 34582 20358 34634 20410
rect 34634 20358 34636 20410
rect 34580 20356 34636 20358
rect 34684 20410 34740 20412
rect 34684 20358 34686 20410
rect 34686 20358 34738 20410
rect 34738 20358 34740 20410
rect 34684 20356 34740 20358
rect 30268 19852 30324 19908
rect 30318 19626 30374 19628
rect 30318 19574 30320 19626
rect 30320 19574 30372 19626
rect 30372 19574 30374 19626
rect 30318 19572 30374 19574
rect 30422 19626 30478 19628
rect 30422 19574 30424 19626
rect 30424 19574 30476 19626
rect 30476 19574 30478 19626
rect 30422 19572 30478 19574
rect 30526 19626 30582 19628
rect 30526 19574 30528 19626
rect 30528 19574 30580 19626
rect 30580 19574 30582 19626
rect 30526 19572 30582 19574
rect 31388 19964 31444 20020
rect 30100 19010 30156 19012
rect 30100 18958 30102 19010
rect 30102 18958 30154 19010
rect 30154 18958 30156 19010
rect 30100 18956 30156 18958
rect 30156 18450 30212 18452
rect 30156 18398 30158 18450
rect 30158 18398 30210 18450
rect 30210 18398 30212 18450
rect 30156 18396 30212 18398
rect 31612 19122 31668 19124
rect 31612 19070 31614 19122
rect 31614 19070 31666 19122
rect 31666 19070 31668 19122
rect 31612 19068 31668 19070
rect 31276 18956 31332 19012
rect 31052 18508 31108 18564
rect 30604 18284 30660 18340
rect 29484 17500 29540 17556
rect 29484 16882 29540 16884
rect 29484 16830 29486 16882
rect 29486 16830 29538 16882
rect 29538 16830 29540 16882
rect 29484 16828 29540 16830
rect 29316 16716 29372 16772
rect 29316 16210 29372 16212
rect 29316 16158 29318 16210
rect 29318 16158 29370 16210
rect 29370 16158 29372 16210
rect 29316 16156 29372 16158
rect 29148 15260 29204 15316
rect 29036 14588 29092 14644
rect 29148 15036 29204 15092
rect 28700 13692 28756 13748
rect 28364 12908 28420 12964
rect 30318 18058 30374 18060
rect 30318 18006 30320 18058
rect 30320 18006 30372 18058
rect 30372 18006 30374 18058
rect 30318 18004 30374 18006
rect 30422 18058 30478 18060
rect 30422 18006 30424 18058
rect 30424 18006 30476 18058
rect 30476 18006 30478 18058
rect 30422 18004 30478 18006
rect 30526 18058 30582 18060
rect 30526 18006 30528 18058
rect 30528 18006 30580 18058
rect 30580 18006 30582 18058
rect 30526 18004 30582 18006
rect 30940 18284 30996 18340
rect 31388 18172 31444 18228
rect 31612 18396 31668 18452
rect 31948 18508 32004 18564
rect 32172 19516 32228 19572
rect 32956 19516 33012 19572
rect 32284 19068 32340 19124
rect 33292 19068 33348 19124
rect 30492 17666 30548 17668
rect 30492 17614 30494 17666
rect 30494 17614 30546 17666
rect 30546 17614 30548 17666
rect 30492 17612 30548 17614
rect 30156 16882 30212 16884
rect 30156 16830 30158 16882
rect 30158 16830 30210 16882
rect 30210 16830 30212 16882
rect 30156 16828 30212 16830
rect 30716 17627 30772 17668
rect 30716 17612 30718 17627
rect 30718 17612 30770 17627
rect 30770 17612 30772 17627
rect 30828 16828 30884 16884
rect 31052 16882 31108 16884
rect 31052 16830 31054 16882
rect 31054 16830 31106 16882
rect 31106 16830 31108 16882
rect 31052 16828 31108 16830
rect 30318 16490 30374 16492
rect 30318 16438 30320 16490
rect 30320 16438 30372 16490
rect 30372 16438 30374 16490
rect 30318 16436 30374 16438
rect 30422 16490 30478 16492
rect 30422 16438 30424 16490
rect 30424 16438 30476 16490
rect 30476 16438 30478 16490
rect 30422 16436 30478 16438
rect 30526 16490 30582 16492
rect 30526 16438 30528 16490
rect 30528 16438 30580 16490
rect 30580 16438 30582 16490
rect 30526 16436 30582 16438
rect 31948 18284 32004 18340
rect 31612 17052 31668 17108
rect 31724 18172 31780 18228
rect 31724 17612 31780 17668
rect 30156 15708 30212 15764
rect 30156 15372 30212 15428
rect 30318 14922 30374 14924
rect 30318 14870 30320 14922
rect 30320 14870 30372 14922
rect 30372 14870 30374 14922
rect 30318 14868 30374 14870
rect 30422 14922 30478 14924
rect 30422 14870 30424 14922
rect 30424 14870 30476 14922
rect 30476 14870 30478 14922
rect 30422 14868 30478 14870
rect 30526 14922 30582 14924
rect 30526 14870 30528 14922
rect 30528 14870 30580 14922
rect 30580 14870 30582 14922
rect 30526 14868 30582 14870
rect 29372 14588 29428 14644
rect 29260 13634 29316 13636
rect 29260 13582 29262 13634
rect 29262 13582 29314 13634
rect 29314 13582 29316 13634
rect 29260 13580 29316 13582
rect 29540 14530 29596 14532
rect 29540 14478 29542 14530
rect 29542 14478 29594 14530
rect 29594 14478 29596 14530
rect 29540 14476 29596 14478
rect 29036 12962 29092 12964
rect 29036 12910 29038 12962
rect 29038 12910 29090 12962
rect 29090 12910 29092 12962
rect 29036 12908 29092 12910
rect 28028 11788 28084 11844
rect 27580 11394 27636 11396
rect 27580 11342 27582 11394
rect 27582 11342 27634 11394
rect 27634 11342 27636 11394
rect 27580 11340 27636 11342
rect 26236 9826 26292 9828
rect 26236 9774 26238 9826
rect 26238 9774 26290 9826
rect 26290 9774 26292 9826
rect 26236 9772 26292 9774
rect 26160 9434 26216 9436
rect 26160 9382 26162 9434
rect 26162 9382 26214 9434
rect 26214 9382 26216 9434
rect 26160 9380 26216 9382
rect 26264 9434 26320 9436
rect 26264 9382 26266 9434
rect 26266 9382 26318 9434
rect 26318 9382 26320 9434
rect 26264 9380 26320 9382
rect 26368 9434 26424 9436
rect 26368 9382 26370 9434
rect 26370 9382 26422 9434
rect 26422 9382 26424 9434
rect 26368 9380 26424 9382
rect 26460 7980 26516 8036
rect 26572 8428 26628 8484
rect 27468 9826 27524 9828
rect 27468 9774 27470 9826
rect 27470 9774 27522 9826
rect 27522 9774 27524 9826
rect 27468 9772 27524 9774
rect 28028 9996 28084 10052
rect 28028 9042 28084 9044
rect 28028 8990 28030 9042
rect 28030 8990 28082 9042
rect 28082 8990 28084 9042
rect 28028 8988 28084 8990
rect 26160 7866 26216 7868
rect 26160 7814 26162 7866
rect 26162 7814 26214 7866
rect 26214 7814 26216 7866
rect 26160 7812 26216 7814
rect 26264 7866 26320 7868
rect 26264 7814 26266 7866
rect 26266 7814 26318 7866
rect 26318 7814 26320 7866
rect 26264 7812 26320 7814
rect 26368 7866 26424 7868
rect 26368 7814 26370 7866
rect 26370 7814 26422 7866
rect 26422 7814 26424 7866
rect 26368 7812 26424 7814
rect 25788 7420 25844 7476
rect 27916 8258 27972 8260
rect 27916 8206 27918 8258
rect 27918 8206 27970 8258
rect 27970 8206 27972 8258
rect 27916 8204 27972 8206
rect 30436 14530 30492 14532
rect 30436 14478 30438 14530
rect 30438 14478 30490 14530
rect 30490 14478 30492 14530
rect 30436 14476 30492 14478
rect 30716 13804 30772 13860
rect 31220 16210 31276 16212
rect 31220 16158 31222 16210
rect 31222 16158 31274 16210
rect 31274 16158 31276 16210
rect 31220 16156 31276 16158
rect 31836 16828 31892 16884
rect 34300 18956 34356 19012
rect 33404 18508 33460 18564
rect 33124 18226 33180 18228
rect 33124 18174 33126 18226
rect 33126 18174 33178 18226
rect 33178 18174 33180 18226
rect 33124 18172 33180 18174
rect 32060 17500 32116 17556
rect 32284 17612 32340 17668
rect 31948 16882 32004 16884
rect 31948 16830 31950 16882
rect 31950 16830 32002 16882
rect 32002 16830 32004 16882
rect 31948 16828 32004 16830
rect 33516 17666 33572 17668
rect 33516 17614 33518 17666
rect 33518 17614 33570 17666
rect 33570 17614 33572 17666
rect 33516 17612 33572 17614
rect 34476 18842 34532 18844
rect 34476 18790 34478 18842
rect 34478 18790 34530 18842
rect 34530 18790 34532 18842
rect 34476 18788 34532 18790
rect 34580 18842 34636 18844
rect 34580 18790 34582 18842
rect 34582 18790 34634 18842
rect 34634 18790 34636 18842
rect 34580 18788 34636 18790
rect 34684 18842 34740 18844
rect 34684 18790 34686 18842
rect 34686 18790 34738 18842
rect 34738 18790 34740 18842
rect 34684 18788 34740 18790
rect 34476 17274 34532 17276
rect 34476 17222 34478 17274
rect 34478 17222 34530 17274
rect 34530 17222 34532 17274
rect 34476 17220 34532 17222
rect 34580 17274 34636 17276
rect 34580 17222 34582 17274
rect 34582 17222 34634 17274
rect 34634 17222 34636 17274
rect 34580 17220 34636 17222
rect 34684 17274 34740 17276
rect 34684 17222 34686 17274
rect 34686 17222 34738 17274
rect 34738 17222 34740 17274
rect 34684 17220 34740 17222
rect 34476 15706 34532 15708
rect 34476 15654 34478 15706
rect 34478 15654 34530 15706
rect 34530 15654 34532 15706
rect 34476 15652 34532 15654
rect 34580 15706 34636 15708
rect 34580 15654 34582 15706
rect 34582 15654 34634 15706
rect 34634 15654 34636 15706
rect 34580 15652 34636 15654
rect 34684 15706 34740 15708
rect 34684 15654 34686 15706
rect 34686 15654 34738 15706
rect 34738 15654 34740 15706
rect 34684 15652 34740 15654
rect 32956 15372 33012 15428
rect 31836 14812 31892 14868
rect 32060 14700 32116 14756
rect 30940 14364 30996 14420
rect 31612 14418 31668 14420
rect 31612 14366 31614 14418
rect 31614 14366 31666 14418
rect 31666 14366 31668 14418
rect 31612 14364 31668 14366
rect 30318 13354 30374 13356
rect 30318 13302 30320 13354
rect 30320 13302 30372 13354
rect 30372 13302 30374 13354
rect 30318 13300 30374 13302
rect 30422 13354 30478 13356
rect 30422 13302 30424 13354
rect 30424 13302 30476 13354
rect 30476 13302 30478 13354
rect 30422 13300 30478 13302
rect 30526 13354 30582 13356
rect 30526 13302 30528 13354
rect 30528 13302 30580 13354
rect 30580 13302 30582 13354
rect 30526 13300 30582 13302
rect 29932 12962 29988 12964
rect 29932 12910 29934 12962
rect 29934 12910 29986 12962
rect 29986 12910 29988 12962
rect 29932 12908 29988 12910
rect 30268 12796 30324 12852
rect 29708 12236 29764 12292
rect 31164 12962 31220 12964
rect 31164 12910 31166 12962
rect 31166 12910 31218 12962
rect 31218 12910 31220 12962
rect 31164 12908 31220 12910
rect 31276 12796 31332 12852
rect 29372 12124 29428 12180
rect 31164 12178 31220 12180
rect 31164 12126 31166 12178
rect 31166 12126 31218 12178
rect 31218 12126 31220 12178
rect 31164 12124 31220 12126
rect 29316 11788 29372 11844
rect 31724 13356 31780 13412
rect 32284 13356 32340 13412
rect 31388 12124 31444 12180
rect 31612 12684 31668 12740
rect 31836 12178 31892 12180
rect 31836 12126 31838 12178
rect 31838 12126 31890 12178
rect 31890 12126 31892 12178
rect 31836 12124 31892 12126
rect 30318 11786 30374 11788
rect 30318 11734 30320 11786
rect 30320 11734 30372 11786
rect 30372 11734 30374 11786
rect 30318 11732 30374 11734
rect 30422 11786 30478 11788
rect 30422 11734 30424 11786
rect 30424 11734 30476 11786
rect 30476 11734 30478 11786
rect 30422 11732 30478 11734
rect 30526 11786 30582 11788
rect 30526 11734 30528 11786
rect 30528 11734 30580 11786
rect 30580 11734 30582 11786
rect 30526 11732 30582 11734
rect 31276 11788 31332 11844
rect 29764 11340 29820 11396
rect 28588 9772 28644 9828
rect 28476 9660 28532 9716
rect 28588 9548 28644 9604
rect 28364 9212 28420 9268
rect 28252 8764 28308 8820
rect 28924 8764 28980 8820
rect 29596 10444 29652 10500
rect 29260 9996 29316 10052
rect 29596 9884 29652 9940
rect 29372 9660 29428 9716
rect 29260 9212 29316 9268
rect 29148 9042 29204 9044
rect 29148 8990 29150 9042
rect 29150 8990 29202 9042
rect 29202 8990 29204 9042
rect 29148 8988 29204 8990
rect 28140 8258 28196 8260
rect 28140 8206 28142 8258
rect 28142 8206 28194 8258
rect 28194 8206 28196 8258
rect 28140 8204 28196 8206
rect 29036 8258 29092 8260
rect 29036 8206 29038 8258
rect 29038 8206 29090 8258
rect 29090 8206 29092 8258
rect 29036 8204 29092 8206
rect 27580 8034 27636 8036
rect 27580 7982 27582 8034
rect 27582 7982 27634 8034
rect 27634 7982 27636 8034
rect 27580 7980 27636 7982
rect 28252 7980 28308 8036
rect 25284 6130 25340 6132
rect 25284 6078 25286 6130
rect 25286 6078 25338 6130
rect 25338 6078 25340 6130
rect 25284 6076 25340 6078
rect 26160 6298 26216 6300
rect 26160 6246 26162 6298
rect 26162 6246 26214 6298
rect 26214 6246 26216 6298
rect 26160 6244 26216 6246
rect 26264 6298 26320 6300
rect 26264 6246 26266 6298
rect 26266 6246 26318 6298
rect 26318 6246 26320 6298
rect 26264 6244 26320 6246
rect 26368 6298 26424 6300
rect 26368 6246 26370 6298
rect 26370 6246 26422 6298
rect 26422 6246 26424 6298
rect 26368 6244 26424 6246
rect 26348 5346 26404 5348
rect 26348 5294 26350 5346
rect 26350 5294 26402 5346
rect 26402 5294 26404 5346
rect 26348 5292 26404 5294
rect 25676 5122 25732 5124
rect 25676 5070 25678 5122
rect 25678 5070 25730 5122
rect 25730 5070 25732 5122
rect 25676 5068 25732 5070
rect 26160 4730 26216 4732
rect 26160 4678 26162 4730
rect 26162 4678 26214 4730
rect 26214 4678 26216 4730
rect 26160 4676 26216 4678
rect 26264 4730 26320 4732
rect 26264 4678 26266 4730
rect 26266 4678 26318 4730
rect 26318 4678 26320 4730
rect 26264 4676 26320 4678
rect 26368 4730 26424 4732
rect 26368 4678 26370 4730
rect 26370 4678 26422 4730
rect 26422 4678 26424 4730
rect 26368 4676 26424 4678
rect 26908 7474 26964 7476
rect 26908 7422 26910 7474
rect 26910 7422 26962 7474
rect 26962 7422 26964 7474
rect 26908 7420 26964 7422
rect 27468 6188 27524 6244
rect 27244 5516 27300 5572
rect 26908 5122 26964 5124
rect 26908 5070 26910 5122
rect 26910 5070 26962 5122
rect 26962 5070 26964 5122
rect 26908 5068 26964 5070
rect 27356 5068 27412 5124
rect 27804 5180 27860 5236
rect 28252 6748 28308 6804
rect 28140 6524 28196 6580
rect 28140 5852 28196 5908
rect 28476 5964 28532 6020
rect 28700 5852 28756 5908
rect 28252 5180 28308 5236
rect 26572 4508 26628 4564
rect 26348 4338 26404 4340
rect 26348 4286 26350 4338
rect 26350 4286 26402 4338
rect 26402 4286 26404 4338
rect 26348 4284 26404 4286
rect 28364 4284 28420 4340
rect 26012 4226 26068 4228
rect 26012 4174 26014 4226
rect 26014 4174 26066 4226
rect 26066 4174 26068 4226
rect 26012 4172 26068 4174
rect 27244 4226 27300 4228
rect 27244 4174 27246 4226
rect 27246 4174 27298 4226
rect 27298 4174 27300 4226
rect 27244 4172 27300 4174
rect 25116 3612 25172 3668
rect 26348 3666 26404 3668
rect 26348 3614 26350 3666
rect 26350 3614 26402 3666
rect 26402 3614 26404 3666
rect 26348 3612 26404 3614
rect 28644 3500 28700 3556
rect 29932 10556 29988 10612
rect 30940 10573 30942 10612
rect 30942 10573 30994 10612
rect 30994 10573 30996 10612
rect 30940 10556 30996 10573
rect 34300 14530 34356 14532
rect 34300 14478 34302 14530
rect 34302 14478 34354 14530
rect 34354 14478 34356 14530
rect 34300 14476 34356 14478
rect 34476 14138 34532 14140
rect 34476 14086 34478 14138
rect 34478 14086 34530 14138
rect 34530 14086 34532 14138
rect 34476 14084 34532 14086
rect 34580 14138 34636 14140
rect 34580 14086 34582 14138
rect 34582 14086 34634 14138
rect 34634 14086 34636 14138
rect 34580 14084 34636 14086
rect 34684 14138 34740 14140
rect 34684 14086 34686 14138
rect 34686 14086 34738 14138
rect 34738 14086 34740 14138
rect 34684 14084 34740 14086
rect 33068 13356 33124 13412
rect 33852 13356 33908 13412
rect 32396 12908 32452 12964
rect 32284 11788 32340 11844
rect 33628 12947 33684 12964
rect 33628 12908 33630 12947
rect 33630 12908 33682 12947
rect 33682 12908 33684 12947
rect 30828 10498 30884 10500
rect 30828 10446 30830 10498
rect 30830 10446 30882 10498
rect 30882 10446 30884 10498
rect 30828 10444 30884 10446
rect 29820 9772 29876 9828
rect 29932 9548 29988 9604
rect 30318 10218 30374 10220
rect 30318 10166 30320 10218
rect 30320 10166 30372 10218
rect 30372 10166 30374 10218
rect 30318 10164 30374 10166
rect 30422 10218 30478 10220
rect 30422 10166 30424 10218
rect 30424 10166 30476 10218
rect 30476 10166 30478 10218
rect 30422 10164 30478 10166
rect 30526 10218 30582 10220
rect 30526 10166 30528 10218
rect 30528 10166 30580 10218
rect 30580 10166 30582 10218
rect 30526 10164 30582 10166
rect 30380 9938 30436 9940
rect 30380 9886 30382 9938
rect 30382 9886 30434 9938
rect 30434 9886 30436 9938
rect 30380 9884 30436 9886
rect 30716 9826 30772 9828
rect 30716 9774 30718 9826
rect 30718 9774 30770 9826
rect 30770 9774 30772 9826
rect 30716 9772 30772 9774
rect 30492 9212 30548 9268
rect 31724 9548 31780 9604
rect 29372 8930 29428 8932
rect 29372 8878 29374 8930
rect 29374 8878 29426 8930
rect 29426 8878 29428 8930
rect 29372 8876 29428 8878
rect 29932 8764 29988 8820
rect 29764 7586 29820 7588
rect 29764 7534 29766 7586
rect 29766 7534 29818 7586
rect 29818 7534 29820 7586
rect 29764 7532 29820 7534
rect 29484 7474 29540 7476
rect 29484 7422 29486 7474
rect 29486 7422 29538 7474
rect 29538 7422 29540 7474
rect 29484 7420 29540 7422
rect 29764 7084 29820 7140
rect 30156 8988 30212 9044
rect 30492 8930 30548 8932
rect 30492 8878 30494 8930
rect 30494 8878 30546 8930
rect 30546 8878 30548 8930
rect 30492 8876 30548 8878
rect 30318 8650 30374 8652
rect 30318 8598 30320 8650
rect 30320 8598 30372 8650
rect 30372 8598 30374 8650
rect 30318 8596 30374 8598
rect 30422 8650 30478 8652
rect 30422 8598 30424 8650
rect 30424 8598 30476 8650
rect 30476 8598 30478 8650
rect 30422 8596 30478 8598
rect 30526 8650 30582 8652
rect 30526 8598 30528 8650
rect 30528 8598 30580 8650
rect 30580 8598 30582 8650
rect 30526 8596 30582 8598
rect 29932 7084 29988 7140
rect 29596 6636 29652 6692
rect 30318 7082 30374 7084
rect 30318 7030 30320 7082
rect 30320 7030 30372 7082
rect 30372 7030 30374 7082
rect 30318 7028 30374 7030
rect 30422 7082 30478 7084
rect 30422 7030 30424 7082
rect 30424 7030 30476 7082
rect 30476 7030 30478 7082
rect 30422 7028 30478 7030
rect 30526 7082 30582 7084
rect 30526 7030 30528 7082
rect 30528 7030 30580 7082
rect 30580 7030 30582 7082
rect 30526 7028 30582 7030
rect 29596 5964 29652 6020
rect 29484 5906 29540 5908
rect 29484 5854 29486 5906
rect 29486 5854 29538 5906
rect 29538 5854 29540 5906
rect 29484 5852 29540 5854
rect 29484 5122 29540 5124
rect 29484 5070 29486 5122
rect 29486 5070 29538 5122
rect 29538 5070 29540 5122
rect 29484 5068 29540 5070
rect 30156 6300 30212 6356
rect 30044 5964 30100 6020
rect 29820 5628 29876 5684
rect 31612 7474 31668 7476
rect 31612 7422 31614 7474
rect 31614 7422 31666 7474
rect 31666 7422 31668 7474
rect 31612 7420 31668 7422
rect 30604 6188 30660 6244
rect 30380 6076 30436 6132
rect 30380 5740 30436 5796
rect 30268 5628 30324 5684
rect 30716 5628 30772 5684
rect 30318 5514 30374 5516
rect 30318 5462 30320 5514
rect 30320 5462 30372 5514
rect 30372 5462 30374 5514
rect 30318 5460 30374 5462
rect 30422 5514 30478 5516
rect 30422 5462 30424 5514
rect 30424 5462 30476 5514
rect 30476 5462 30478 5514
rect 30422 5460 30478 5462
rect 30526 5514 30582 5516
rect 30526 5462 30528 5514
rect 30528 5462 30580 5514
rect 30580 5462 30582 5514
rect 30526 5460 30582 5462
rect 30380 5122 30436 5124
rect 30380 5070 30382 5122
rect 30382 5070 30434 5122
rect 30434 5070 30436 5122
rect 30380 5068 30436 5070
rect 30604 4844 30660 4900
rect 29764 4562 29820 4564
rect 29764 4510 29766 4562
rect 29766 4510 29818 4562
rect 29818 4510 29820 4562
rect 29764 4508 29820 4510
rect 30318 3946 30374 3948
rect 30318 3894 30320 3946
rect 30320 3894 30372 3946
rect 30372 3894 30374 3946
rect 30318 3892 30374 3894
rect 30422 3946 30478 3948
rect 30422 3894 30424 3946
rect 30424 3894 30476 3946
rect 30476 3894 30478 3946
rect 30422 3892 30478 3894
rect 30526 3946 30582 3948
rect 30526 3894 30528 3946
rect 30528 3894 30580 3946
rect 30580 3894 30582 3946
rect 30526 3892 30582 3894
rect 30996 5628 31052 5684
rect 31276 5740 31332 5796
rect 30940 5180 30996 5236
rect 30940 4844 30996 4900
rect 31052 3836 31108 3892
rect 31052 3539 31108 3556
rect 31052 3500 31054 3539
rect 31054 3500 31106 3539
rect 31106 3500 31108 3539
rect 31388 5628 31444 5684
rect 32956 10610 33012 10612
rect 32956 10558 32958 10610
rect 32958 10558 33010 10610
rect 33010 10558 33012 10610
rect 32956 10556 33012 10558
rect 33180 10780 33236 10836
rect 33628 12684 33684 12740
rect 34476 12570 34532 12572
rect 34476 12518 34478 12570
rect 34478 12518 34530 12570
rect 34530 12518 34532 12570
rect 34476 12516 34532 12518
rect 34580 12570 34636 12572
rect 34580 12518 34582 12570
rect 34582 12518 34634 12570
rect 34634 12518 34636 12570
rect 34580 12516 34636 12518
rect 34684 12570 34740 12572
rect 34684 12518 34686 12570
rect 34686 12518 34738 12570
rect 34738 12518 34740 12570
rect 34684 12516 34740 12518
rect 34476 11002 34532 11004
rect 34476 10950 34478 11002
rect 34478 10950 34530 11002
rect 34530 10950 34532 11002
rect 34476 10948 34532 10950
rect 34580 11002 34636 11004
rect 34580 10950 34582 11002
rect 34582 10950 34634 11002
rect 34634 10950 34636 11002
rect 34580 10948 34636 10950
rect 34684 11002 34740 11004
rect 34684 10950 34686 11002
rect 34686 10950 34738 11002
rect 34738 10950 34740 11002
rect 34684 10948 34740 10950
rect 34076 10556 34132 10612
rect 33292 9660 33348 9716
rect 34476 9434 34532 9436
rect 34476 9382 34478 9434
rect 34478 9382 34530 9434
rect 34530 9382 34532 9434
rect 34476 9380 34532 9382
rect 34580 9434 34636 9436
rect 34580 9382 34582 9434
rect 34582 9382 34634 9434
rect 34634 9382 34636 9434
rect 34580 9380 34636 9382
rect 34684 9434 34740 9436
rect 34684 9382 34686 9434
rect 34686 9382 34738 9434
rect 34738 9382 34740 9434
rect 34684 9380 34740 9382
rect 31892 8988 31948 9044
rect 34476 7866 34532 7868
rect 34476 7814 34478 7866
rect 34478 7814 34530 7866
rect 34530 7814 34532 7866
rect 34476 7812 34532 7814
rect 34580 7866 34636 7868
rect 34580 7814 34582 7866
rect 34582 7814 34634 7866
rect 34634 7814 34636 7866
rect 34580 7812 34636 7814
rect 34684 7866 34740 7868
rect 34684 7814 34686 7866
rect 34686 7814 34738 7866
rect 34738 7814 34740 7866
rect 34684 7812 34740 7814
rect 31836 7308 31892 7364
rect 32060 7362 32116 7364
rect 32060 7310 32062 7362
rect 32062 7310 32114 7362
rect 32114 7310 32116 7362
rect 32060 7308 32116 7310
rect 33628 7420 33684 7476
rect 32172 6802 32228 6804
rect 32172 6750 32174 6802
rect 32174 6750 32226 6802
rect 32226 6750 32228 6802
rect 32172 6748 32228 6750
rect 31948 5852 32004 5908
rect 31612 5068 31668 5124
rect 32172 6076 32228 6132
rect 33292 6748 33348 6804
rect 33124 6076 33180 6132
rect 33404 5906 33460 5908
rect 33404 5854 33406 5906
rect 33406 5854 33458 5906
rect 33458 5854 33460 5906
rect 33404 5852 33460 5854
rect 34076 7420 34132 7476
rect 34476 6298 34532 6300
rect 34476 6246 34478 6298
rect 34478 6246 34530 6298
rect 34530 6246 34532 6298
rect 34476 6244 34532 6246
rect 34580 6298 34636 6300
rect 34580 6246 34582 6298
rect 34582 6246 34634 6298
rect 34634 6246 34636 6298
rect 34580 6244 34636 6246
rect 34684 6298 34740 6300
rect 34684 6246 34686 6298
rect 34686 6246 34738 6298
rect 34738 6246 34740 6298
rect 34684 6244 34740 6246
rect 34076 5740 34132 5796
rect 31948 5180 32004 5236
rect 31500 4114 31556 4116
rect 31500 4062 31502 4114
rect 31502 4062 31554 4114
rect 31554 4062 31556 4114
rect 31500 4060 31556 4062
rect 32396 5292 32452 5348
rect 31948 3724 32004 3780
rect 32172 4060 32228 4116
rect 34476 4730 34532 4732
rect 34476 4678 34478 4730
rect 34478 4678 34530 4730
rect 34530 4678 34532 4730
rect 34476 4676 34532 4678
rect 34580 4730 34636 4732
rect 34580 4678 34582 4730
rect 34582 4678 34634 4730
rect 34634 4678 34636 4730
rect 34580 4676 34636 4678
rect 34684 4730 34740 4732
rect 34684 4678 34686 4730
rect 34686 4678 34738 4730
rect 34738 4678 34740 4730
rect 34684 4676 34740 4678
rect 26160 3162 26216 3164
rect 26160 3110 26162 3162
rect 26162 3110 26214 3162
rect 26214 3110 26216 3162
rect 26160 3108 26216 3110
rect 26264 3162 26320 3164
rect 26264 3110 26266 3162
rect 26266 3110 26318 3162
rect 26318 3110 26320 3162
rect 26264 3108 26320 3110
rect 26368 3162 26424 3164
rect 26368 3110 26370 3162
rect 26370 3110 26422 3162
rect 26422 3110 26424 3162
rect 26368 3108 26424 3110
rect 32844 3836 32900 3892
rect 32564 3778 32620 3780
rect 32564 3726 32566 3778
rect 32566 3726 32618 3778
rect 32618 3726 32620 3778
rect 32564 3724 32620 3726
rect 32284 3554 32340 3556
rect 32284 3502 32286 3554
rect 32286 3502 32338 3554
rect 32338 3502 32340 3554
rect 32284 3500 32340 3502
rect 34476 3162 34532 3164
rect 34476 3110 34478 3162
rect 34478 3110 34530 3162
rect 34530 3110 34532 3162
rect 34476 3108 34532 3110
rect 34580 3162 34636 3164
rect 34580 3110 34582 3162
rect 34582 3110 34634 3162
rect 34634 3110 34636 3162
rect 34580 3108 34636 3110
rect 34684 3162 34740 3164
rect 34684 3110 34686 3162
rect 34686 3110 34738 3162
rect 34738 3110 34740 3162
rect 34684 3108 34740 3110
<< metal3 >>
rect 5360 32116 5370 32172
rect 5426 32116 5474 32172
rect 5530 32116 5578 32172
rect 5634 32116 5644 32172
rect 13676 32116 13686 32172
rect 13742 32116 13790 32172
rect 13846 32116 13894 32172
rect 13950 32116 13960 32172
rect 21992 32116 22002 32172
rect 22058 32116 22106 32172
rect 22162 32116 22210 32172
rect 22266 32116 22276 32172
rect 30308 32116 30318 32172
rect 30374 32116 30422 32172
rect 30478 32116 30526 32172
rect 30582 32116 30592 32172
rect 19618 31836 19628 31892
rect 19684 31836 20524 31892
rect 20580 31836 20590 31892
rect 14802 31500 14812 31556
rect 14868 31500 15820 31556
rect 15876 31500 15886 31556
rect 9518 31332 9528 31388
rect 9584 31332 9632 31388
rect 9688 31332 9736 31388
rect 9792 31332 9802 31388
rect 17834 31332 17844 31388
rect 17900 31332 17948 31388
rect 18004 31332 18052 31388
rect 18108 31332 18118 31388
rect 26150 31332 26160 31388
rect 26216 31332 26264 31388
rect 26320 31332 26368 31388
rect 26424 31332 26434 31388
rect 34466 31332 34476 31388
rect 34532 31332 34580 31388
rect 34636 31332 34684 31388
rect 34740 31332 34750 31388
rect 22642 30828 22652 30884
rect 22708 30828 25340 30884
rect 25396 30828 25406 30884
rect 5360 30548 5370 30604
rect 5426 30548 5474 30604
rect 5530 30548 5578 30604
rect 5634 30548 5644 30604
rect 13676 30548 13686 30604
rect 13742 30548 13790 30604
rect 13846 30548 13894 30604
rect 13950 30548 13960 30604
rect 21992 30548 22002 30604
rect 22058 30548 22106 30604
rect 22162 30548 22210 30604
rect 22266 30548 22276 30604
rect 30308 30548 30318 30604
rect 30374 30548 30422 30604
rect 30478 30548 30526 30604
rect 30582 30548 30592 30604
rect 20850 30268 20860 30324
rect 20916 30268 21308 30324
rect 21364 30268 21644 30324
rect 21700 30268 21710 30324
rect 10434 30156 10444 30212
rect 10500 30156 11676 30212
rect 11732 30156 11742 30212
rect 16818 30156 16828 30212
rect 16884 30156 17724 30212
rect 17780 30156 17790 30212
rect 18050 30156 18060 30212
rect 18116 30156 18620 30212
rect 18676 30156 18686 30212
rect 18946 30156 18956 30212
rect 19012 30156 20300 30212
rect 20356 30156 20366 30212
rect 24322 30156 24332 30212
rect 24388 30156 24668 30212
rect 24724 30156 24734 30212
rect 11554 30044 11564 30100
rect 11620 30044 14700 30100
rect 14756 30044 14766 30100
rect 20132 30044 20636 30100
rect 20692 30044 20702 30100
rect 23986 30044 23996 30100
rect 24052 30044 25172 30100
rect 25228 30044 25238 30100
rect 20132 29988 20188 30044
rect 11778 29932 11788 29988
rect 11844 29932 13692 29988
rect 13748 29932 15708 29988
rect 15764 29932 18508 29988
rect 18564 29932 20188 29988
rect 22866 29932 22876 29988
rect 22932 29932 24892 29988
rect 24948 29932 25900 29988
rect 25956 29932 25966 29988
rect 9518 29764 9528 29820
rect 9584 29764 9632 29820
rect 9688 29764 9736 29820
rect 9792 29764 9802 29820
rect 17834 29764 17844 29820
rect 17900 29764 17948 29820
rect 18004 29764 18052 29820
rect 18108 29764 18118 29820
rect 26150 29764 26160 29820
rect 26216 29764 26264 29820
rect 26320 29764 26368 29820
rect 26424 29764 26434 29820
rect 34466 29764 34476 29820
rect 34532 29764 34580 29820
rect 34636 29764 34684 29820
rect 34740 29764 34750 29820
rect 16370 29596 16380 29652
rect 16436 29596 17332 29652
rect 17388 29596 18396 29652
rect 18452 29596 20188 29652
rect 20244 29596 20254 29652
rect 14634 29484 14644 29540
rect 14700 29484 15932 29540
rect 15988 29484 17052 29540
rect 17108 29484 17118 29540
rect 19506 29484 19516 29540
rect 19572 29484 19740 29540
rect 19796 29484 20468 29540
rect 20524 29484 20534 29540
rect 23314 29484 23324 29540
rect 23380 29484 25228 29540
rect 25284 29484 26796 29540
rect 26852 29484 26862 29540
rect 12674 29372 12684 29428
rect 12740 29372 13468 29428
rect 13524 29372 13534 29428
rect 14242 29372 14252 29428
rect 14308 29372 15428 29428
rect 15484 29372 15494 29428
rect 16258 29372 16268 29428
rect 16324 29372 16828 29428
rect 16884 29372 16894 29428
rect 19618 29372 19628 29428
rect 19684 29372 20748 29428
rect 20804 29372 20814 29428
rect 22642 29372 22652 29428
rect 22708 29372 24108 29428
rect 24164 29372 24174 29428
rect 25442 29372 25452 29428
rect 25508 29372 27580 29428
rect 27636 29372 29036 29428
rect 29092 29372 29102 29428
rect 12114 29260 12124 29316
rect 12180 29260 12348 29316
rect 12404 29260 12908 29316
rect 12964 29260 13356 29316
rect 13412 29260 13422 29316
rect 18498 29260 18508 29316
rect 18564 29260 19180 29316
rect 19236 29260 19246 29316
rect 22978 29260 22988 29316
rect 23044 29260 23660 29316
rect 23716 29260 23726 29316
rect 13234 29148 13244 29204
rect 13300 29148 13748 29204
rect 13804 29148 14364 29204
rect 14420 29148 14430 29204
rect 14802 29148 14812 29204
rect 14868 29148 14878 29204
rect 18162 29148 18172 29204
rect 18228 29148 19964 29204
rect 20020 29148 20030 29204
rect 5360 28980 5370 29036
rect 5426 28980 5474 29036
rect 5530 28980 5578 29036
rect 5634 28980 5644 29036
rect 13676 28980 13686 29036
rect 13742 28980 13790 29036
rect 13846 28980 13894 29036
rect 13950 28980 13960 29036
rect 14812 28868 14868 29148
rect 21992 28980 22002 29036
rect 22058 28980 22106 29036
rect 22162 28980 22210 29036
rect 22266 28980 22276 29036
rect 30308 28980 30318 29036
rect 30374 28980 30422 29036
rect 30478 28980 30526 29036
rect 30582 28980 30592 29036
rect 13906 28812 13916 28868
rect 13972 28812 15708 28868
rect 15764 28812 15774 28868
rect 14354 28700 14364 28756
rect 14420 28700 15428 28756
rect 15484 28700 15494 28756
rect 20066 28700 20076 28756
rect 20132 28700 21084 28756
rect 21140 28700 21150 28756
rect 24770 28700 24780 28756
rect 24836 28700 26012 28756
rect 26068 28700 26684 28756
rect 26740 28700 27356 28756
rect 27412 28700 27422 28756
rect 13346 28588 13356 28644
rect 13412 28588 13636 28644
rect 13692 28588 13702 28644
rect 13804 28588 15820 28644
rect 15876 28588 16716 28644
rect 16772 28588 16782 28644
rect 24546 28588 24556 28644
rect 24612 28588 25228 28644
rect 25284 28588 25294 28644
rect 13804 28532 13860 28588
rect 13458 28476 13468 28532
rect 13524 28476 13860 28532
rect 27850 28476 27860 28532
rect 27916 28476 28700 28532
rect 28756 28476 28766 28532
rect 9518 28196 9528 28252
rect 9584 28196 9632 28252
rect 9688 28196 9736 28252
rect 9792 28196 9802 28252
rect 17834 28196 17844 28252
rect 17900 28196 17948 28252
rect 18004 28196 18052 28252
rect 18108 28196 18118 28252
rect 26150 28196 26160 28252
rect 26216 28196 26264 28252
rect 26320 28196 26368 28252
rect 26424 28196 26434 28252
rect 34466 28196 34476 28252
rect 34532 28196 34580 28252
rect 34636 28196 34684 28252
rect 34740 28196 34750 28252
rect 27570 28140 27580 28196
rect 27636 28140 28476 28196
rect 28532 28140 28542 28196
rect 11442 27804 11452 27860
rect 11508 27804 12348 27860
rect 12404 27804 12414 27860
rect 12898 27804 12908 27860
rect 12964 27804 13244 27860
rect 13300 27804 13310 27860
rect 28354 27804 28364 27860
rect 28420 27804 28924 27860
rect 28980 27804 28990 27860
rect 5360 27412 5370 27468
rect 5426 27412 5474 27468
rect 5530 27412 5578 27468
rect 5634 27412 5644 27468
rect 13676 27412 13686 27468
rect 13742 27412 13790 27468
rect 13846 27412 13894 27468
rect 13950 27412 13960 27468
rect 21992 27412 22002 27468
rect 22058 27412 22106 27468
rect 22162 27412 22210 27468
rect 22266 27412 22276 27468
rect 30308 27412 30318 27468
rect 30374 27412 30422 27468
rect 30478 27412 30526 27468
rect 30582 27412 30592 27468
rect 21522 27132 21532 27188
rect 21588 27132 21980 27188
rect 22036 27132 22046 27188
rect 27794 27132 27804 27188
rect 27860 27132 28476 27188
rect 28532 27132 28542 27188
rect 12674 27020 12684 27076
rect 12740 27020 14028 27076
rect 14084 27020 14094 27076
rect 14466 27020 14476 27076
rect 14532 27020 16716 27076
rect 16772 27020 17500 27076
rect 17556 27020 17566 27076
rect 20402 27020 20412 27076
rect 20468 27020 23492 27076
rect 23548 27020 23558 27076
rect 6066 26908 6076 26964
rect 6132 26908 6972 26964
rect 7028 26908 7038 26964
rect 5786 26796 5796 26852
rect 5852 26796 7532 26852
rect 7588 26796 7598 26852
rect 17602 26796 17612 26852
rect 17668 26796 18172 26852
rect 18228 26796 18238 26852
rect 9518 26628 9528 26684
rect 9584 26628 9632 26684
rect 9688 26628 9736 26684
rect 9792 26628 9802 26684
rect 17834 26628 17844 26684
rect 17900 26628 17948 26684
rect 18004 26628 18052 26684
rect 18108 26628 18118 26684
rect 26150 26628 26160 26684
rect 26216 26628 26264 26684
rect 26320 26628 26368 26684
rect 26424 26628 26434 26684
rect 34466 26628 34476 26684
rect 34532 26628 34580 26684
rect 34636 26628 34684 26684
rect 34740 26628 34750 26684
rect 28242 26348 28252 26404
rect 28308 26348 28588 26404
rect 28644 26348 29372 26404
rect 29428 26348 29438 26404
rect 4610 26236 4620 26292
rect 4676 26236 5292 26292
rect 5348 26236 5796 26292
rect 5852 26236 5862 26292
rect 7970 26236 7980 26292
rect 8036 26236 8876 26292
rect 8932 26236 9660 26292
rect 9716 26236 9726 26292
rect 12114 26236 12124 26292
rect 12180 26236 12684 26292
rect 12740 26236 12750 26292
rect 14242 26236 14252 26292
rect 14308 26236 17276 26292
rect 17332 26236 17342 26292
rect 19842 26236 19852 26292
rect 19908 26236 20972 26292
rect 21028 26236 21868 26292
rect 21924 26236 21934 26292
rect 3042 26124 3052 26180
rect 3108 26124 4844 26180
rect 4900 26124 4910 26180
rect 10490 26124 10500 26180
rect 10556 26124 10892 26180
rect 10948 26124 13188 26180
rect 13244 26124 13254 26180
rect 8194 26012 8204 26068
rect 8260 26012 12292 26068
rect 12348 26012 12358 26068
rect 27570 26012 27580 26068
rect 27636 26012 28140 26068
rect 28196 26012 28924 26068
rect 28980 26012 29652 26068
rect 29708 26012 29718 26068
rect 5360 25844 5370 25900
rect 5426 25844 5474 25900
rect 5530 25844 5578 25900
rect 5634 25844 5644 25900
rect 13676 25844 13686 25900
rect 13742 25844 13790 25900
rect 13846 25844 13894 25900
rect 13950 25844 13960 25900
rect 21992 25844 22002 25900
rect 22058 25844 22106 25900
rect 22162 25844 22210 25900
rect 22266 25844 22276 25900
rect 30308 25844 30318 25900
rect 30374 25844 30422 25900
rect 30478 25844 30526 25900
rect 30582 25844 30592 25900
rect 6738 25788 6748 25844
rect 6804 25788 8652 25844
rect 8708 25788 10220 25844
rect 10276 25788 10286 25844
rect 7410 25676 7420 25732
rect 7476 25676 7812 25732
rect 7868 25676 7878 25732
rect 8754 25676 8764 25732
rect 8820 25676 15260 25732
rect 15316 25676 15326 25732
rect 8764 25620 8820 25676
rect 6514 25564 6524 25620
rect 6580 25564 6860 25620
rect 6916 25564 8820 25620
rect 13682 25564 13692 25620
rect 13748 25564 14700 25620
rect 14756 25564 15596 25620
rect 15652 25564 16156 25620
rect 16212 25564 16222 25620
rect 18162 25564 18172 25620
rect 18228 25564 24556 25620
rect 24612 25564 24622 25620
rect 7522 25452 7532 25508
rect 7588 25452 8764 25508
rect 8820 25452 9828 25508
rect 9884 25452 9894 25508
rect 9986 25452 9996 25508
rect 10052 25452 13524 25508
rect 13580 25452 13590 25508
rect 14466 25452 14476 25508
rect 14532 25452 15708 25508
rect 15764 25452 15774 25508
rect 16034 25452 16044 25508
rect 16100 25452 18732 25508
rect 18788 25452 19964 25508
rect 20020 25452 20030 25508
rect 23986 25452 23996 25508
rect 24052 25452 28140 25508
rect 28196 25452 28206 25508
rect 29698 25452 29708 25508
rect 29764 25452 31164 25508
rect 31220 25452 31230 25508
rect 11004 25396 11060 25452
rect 10994 25340 11004 25396
rect 11060 25340 11070 25396
rect 12562 25340 12572 25396
rect 12628 25340 14588 25396
rect 14644 25340 14654 25396
rect 15250 25340 15260 25396
rect 15316 25340 15932 25396
rect 15988 25340 15998 25396
rect 19282 25340 19292 25396
rect 19348 25340 20188 25396
rect 20244 25340 20860 25396
rect 20916 25340 20926 25396
rect 28018 25340 28028 25396
rect 28084 25340 29260 25396
rect 29316 25340 29326 25396
rect 1586 25228 1596 25284
rect 1652 25228 2268 25284
rect 2324 25228 4620 25284
rect 4676 25228 4686 25284
rect 7298 25228 7308 25284
rect 7364 25228 7374 25284
rect 7942 25228 7980 25284
rect 8036 25228 8046 25284
rect 8362 25228 8372 25284
rect 8428 25228 14476 25284
rect 14532 25228 14542 25284
rect 15092 25228 16380 25284
rect 16436 25228 16446 25284
rect 7308 25172 7364 25228
rect 15092 25172 15148 25228
rect 6738 25116 6748 25172
rect 6804 25116 7364 25172
rect 13458 25116 13468 25172
rect 13524 25116 14140 25172
rect 14196 25116 15148 25172
rect 9518 25060 9528 25116
rect 9584 25060 9632 25116
rect 9688 25060 9736 25116
rect 9792 25060 9802 25116
rect 17834 25060 17844 25116
rect 17900 25060 17948 25116
rect 18004 25060 18052 25116
rect 18108 25060 18118 25116
rect 26150 25060 26160 25116
rect 26216 25060 26264 25116
rect 26320 25060 26368 25116
rect 26424 25060 26434 25116
rect 34466 25060 34476 25116
rect 34532 25060 34580 25116
rect 34636 25060 34684 25116
rect 34740 25060 34750 25116
rect 5058 25004 5068 25060
rect 5124 25004 9380 25060
rect 9324 24948 9380 25004
rect 10892 25004 13692 25060
rect 13748 25004 13758 25060
rect 22082 25004 22092 25060
rect 22148 25004 23548 25060
rect 23604 25004 23614 25060
rect 24434 25004 24444 25060
rect 24500 25004 24510 25060
rect 10892 24948 10948 25004
rect 24444 24948 24500 25004
rect 5170 24892 5180 24948
rect 5236 24892 6524 24948
rect 6580 24892 6590 24948
rect 9324 24892 10948 24948
rect 11106 24892 11116 24948
rect 11172 24892 12740 24948
rect 12796 24892 12806 24948
rect 17602 24892 17612 24948
rect 17668 24892 18956 24948
rect 19012 24892 19022 24948
rect 23314 24892 23324 24948
rect 23380 24892 26236 24948
rect 26292 24892 27356 24948
rect 27412 24892 27422 24948
rect 4386 24780 4396 24836
rect 4452 24780 5068 24836
rect 5124 24780 5134 24836
rect 6234 24780 6244 24836
rect 6300 24780 7532 24836
rect 7588 24780 7598 24836
rect 7690 24780 7700 24836
rect 7756 24780 8428 24836
rect 8484 24780 8494 24836
rect 12002 24780 12012 24836
rect 12068 24780 12908 24836
rect 12964 24780 13244 24836
rect 13300 24780 15820 24836
rect 15876 24780 15886 24836
rect 16594 24780 16604 24836
rect 16660 24780 18396 24836
rect 18452 24780 19068 24836
rect 19124 24780 19852 24836
rect 19908 24780 19918 24836
rect 22418 24780 22428 24836
rect 22484 24780 22988 24836
rect 23044 24780 23054 24836
rect 24322 24780 24332 24836
rect 24388 24780 24836 24836
rect 24892 24780 27020 24836
rect 27076 24780 27580 24836
rect 27636 24780 27646 24836
rect 4946 24668 4956 24724
rect 5012 24668 6636 24724
rect 6692 24668 6702 24724
rect 7970 24668 7980 24724
rect 8036 24668 8260 24724
rect 8316 24668 8326 24724
rect 11666 24668 11676 24724
rect 11732 24668 12460 24724
rect 12516 24668 12526 24724
rect 16370 24668 16380 24724
rect 16436 24668 17276 24724
rect 17332 24668 17342 24724
rect 21074 24668 21084 24724
rect 21140 24668 21756 24724
rect 21812 24668 23436 24724
rect 23492 24668 25004 24724
rect 25060 24668 25070 24724
rect 6300 24612 6356 24668
rect 6290 24556 6300 24612
rect 6356 24556 6366 24612
rect 22866 24556 22876 24612
rect 22932 24556 23996 24612
rect 24052 24556 24062 24612
rect 18554 24444 18564 24500
rect 18620 24444 19628 24500
rect 19684 24444 19694 24500
rect 20132 24444 22092 24500
rect 22148 24444 22158 24500
rect 22978 24444 22988 24500
rect 23044 24444 23212 24500
rect 23268 24444 23660 24500
rect 23716 24444 26740 24500
rect 26796 24444 27188 24500
rect 27244 24444 27692 24500
rect 27748 24444 28252 24500
rect 28308 24444 28318 24500
rect 20132 24388 20188 24444
rect 7196 24332 13468 24388
rect 13524 24332 13534 24388
rect 20132 24332 20412 24388
rect 20468 24332 20478 24388
rect 5360 24276 5370 24332
rect 5426 24276 5474 24332
rect 5530 24276 5578 24332
rect 5634 24276 5644 24332
rect 7130 24220 7140 24276
rect 7196 24220 7252 24332
rect 13676 24276 13686 24332
rect 13742 24276 13790 24332
rect 13846 24276 13894 24332
rect 13950 24276 13960 24332
rect 9202 24220 9212 24276
rect 9268 24220 12236 24276
rect 12292 24220 12302 24276
rect 20132 24164 20188 24332
rect 21992 24276 22002 24332
rect 22058 24276 22106 24332
rect 22162 24276 22210 24332
rect 22266 24276 22276 24332
rect 30308 24276 30318 24332
rect 30374 24276 30422 24332
rect 30478 24276 30526 24332
rect 30582 24276 30592 24332
rect 3042 24108 3052 24164
rect 3108 24108 4340 24164
rect 4396 24108 4406 24164
rect 8306 24108 8316 24164
rect 8372 24108 9324 24164
rect 9380 24108 9390 24164
rect 19282 24108 19292 24164
rect 19348 24108 20188 24164
rect 4890 23996 4900 24052
rect 4956 23996 7140 24052
rect 7196 23996 7206 24052
rect 8194 23996 8204 24052
rect 8260 23996 10220 24052
rect 10276 23996 10892 24052
rect 10948 23996 10958 24052
rect 11834 23996 11844 24052
rect 11900 23996 12348 24052
rect 12404 23996 12414 24052
rect 19506 23996 19516 24052
rect 19572 23996 23660 24052
rect 23716 23996 23726 24052
rect 24322 23996 24332 24052
rect 24388 23996 25452 24052
rect 25508 23996 25518 24052
rect 4610 23884 4620 23940
rect 4676 23884 5796 23940
rect 5852 23884 5862 23940
rect 6850 23884 6860 23940
rect 6916 23884 9828 23940
rect 9884 23884 9894 23940
rect 11218 23884 11228 23940
rect 11284 23884 11564 23940
rect 11620 23884 12236 23940
rect 12292 23884 17612 23940
rect 17668 23884 17678 23940
rect 26786 23884 26796 23940
rect 26852 23884 27244 23940
rect 27300 23884 27310 23940
rect 28466 23884 28476 23940
rect 28532 23884 29036 23940
rect 29092 23884 29102 23940
rect 4386 23772 4396 23828
rect 4452 23772 4732 23828
rect 4788 23772 4798 23828
rect 6290 23772 6300 23828
rect 6356 23772 7868 23828
rect 7924 23772 7934 23828
rect 8866 23772 8876 23828
rect 8932 23772 9548 23828
rect 9604 23772 16604 23828
rect 16660 23772 16940 23828
rect 16996 23772 17836 23828
rect 17892 23772 17902 23828
rect 20132 23772 20300 23828
rect 20356 23772 22428 23828
rect 22484 23772 22494 23828
rect 20132 23716 20188 23772
rect 6066 23660 6076 23716
rect 6132 23660 6860 23716
rect 6916 23660 6926 23716
rect 8530 23660 8540 23716
rect 8596 23660 10052 23716
rect 13458 23660 13468 23716
rect 13524 23660 17276 23716
rect 17332 23660 20188 23716
rect 9996 23604 10052 23660
rect 3938 23548 3948 23604
rect 4004 23548 4732 23604
rect 4788 23548 5180 23604
rect 5236 23548 6300 23604
rect 6356 23548 6366 23604
rect 9996 23548 13356 23604
rect 13412 23548 13422 23604
rect 9518 23492 9528 23548
rect 9584 23492 9632 23548
rect 9688 23492 9736 23548
rect 9792 23492 9802 23548
rect 17834 23492 17844 23548
rect 17900 23492 17948 23548
rect 18004 23492 18052 23548
rect 18108 23492 18118 23548
rect 26150 23492 26160 23548
rect 26216 23492 26264 23548
rect 26320 23492 26368 23548
rect 26424 23492 26434 23548
rect 34466 23492 34476 23548
rect 34532 23492 34580 23548
rect 34636 23492 34684 23548
rect 34740 23492 34750 23548
rect 3602 23436 3612 23492
rect 3668 23436 3836 23492
rect 3892 23436 3902 23492
rect 12392 23324 12402 23380
rect 12458 23324 12684 23380
rect 12740 23324 14364 23380
rect 14420 23324 14430 23380
rect 16706 23324 16716 23380
rect 16772 23324 20132 23380
rect 20188 23324 20198 23380
rect 4274 23212 4284 23268
rect 4340 23212 5608 23268
rect 5664 23212 6636 23268
rect 6692 23212 6702 23268
rect 4172 23100 4844 23156
rect 4900 23100 4910 23156
rect 6402 23100 6412 23156
rect 6468 23100 7532 23156
rect 7588 23100 7598 23156
rect 12786 23100 12796 23156
rect 12852 23100 13804 23156
rect 13860 23100 13870 23156
rect 18162 23100 18172 23156
rect 18228 23100 18956 23156
rect 19012 23100 19022 23156
rect 4172 23044 4228 23100
rect 4162 22988 4172 23044
rect 4228 22988 4238 23044
rect 6738 22988 6748 23044
rect 6804 22988 8484 23044
rect 8540 22988 8550 23044
rect 18498 22988 18508 23044
rect 18564 22988 19180 23044
rect 19236 22988 19246 23044
rect 5842 22876 5852 22932
rect 5908 22876 7532 22932
rect 7588 22876 7598 22932
rect 7914 22876 7924 22932
rect 7980 22876 9324 22932
rect 9380 22876 9390 22932
rect 12460 22876 14140 22932
rect 14196 22876 17780 22932
rect 17836 22876 18060 22932
rect 18116 22876 18126 22932
rect 8418 22764 8428 22820
rect 8484 22764 8988 22820
rect 9044 22764 9054 22820
rect 5360 22708 5370 22764
rect 5426 22708 5474 22764
rect 5530 22708 5578 22764
rect 5634 22708 5644 22764
rect 12460 22708 12516 22876
rect 13676 22708 13686 22764
rect 13742 22708 13790 22764
rect 13846 22708 13894 22764
rect 13950 22708 13960 22764
rect 21992 22708 22002 22764
rect 22058 22708 22106 22764
rect 22162 22708 22210 22764
rect 22266 22708 22276 22764
rect 30308 22708 30318 22764
rect 30374 22708 30422 22764
rect 30478 22708 30526 22764
rect 30582 22708 30592 22764
rect 8642 22652 8652 22708
rect 8708 22652 12460 22708
rect 12516 22652 12526 22708
rect 6850 22540 6860 22596
rect 6916 22540 9884 22596
rect 9940 22540 9950 22596
rect 12058 22540 12068 22596
rect 12124 22540 13020 22596
rect 13076 22540 13086 22596
rect 3378 22428 3388 22484
rect 3444 22428 4060 22484
rect 4116 22428 4126 22484
rect 7858 22428 7868 22484
rect 7924 22428 8876 22484
rect 8932 22428 8942 22484
rect 12226 22428 12236 22484
rect 12292 22428 12796 22484
rect 12852 22428 12862 22484
rect 14690 22428 14700 22484
rect 14756 22428 19964 22484
rect 20020 22428 20030 22484
rect 3042 22316 3052 22372
rect 3108 22316 4452 22372
rect 4508 22316 4518 22372
rect 8082 22316 8092 22372
rect 8148 22316 8540 22372
rect 8596 22316 8606 22372
rect 14018 22316 14028 22372
rect 14084 22316 14252 22372
rect 14308 22316 14318 22372
rect 18162 22316 18172 22372
rect 18228 22316 19180 22372
rect 19236 22316 19246 22372
rect 22754 22316 22764 22372
rect 22820 22316 25284 22372
rect 25340 22316 25350 22372
rect 8866 22204 8876 22260
rect 8932 22204 11788 22260
rect 11844 22204 11854 22260
rect 12114 22204 12124 22260
rect 12180 22204 13524 22260
rect 13580 22204 13590 22260
rect 8642 22092 8652 22148
rect 8708 22092 9548 22148
rect 9604 22092 9614 22148
rect 10938 22092 10948 22148
rect 11004 22092 11564 22148
rect 11620 22092 11630 22148
rect 22866 21980 22876 22036
rect 22932 21980 23156 22036
rect 23212 21980 23222 22036
rect 9518 21924 9528 21980
rect 9584 21924 9632 21980
rect 9688 21924 9736 21980
rect 9792 21924 9802 21980
rect 17834 21924 17844 21980
rect 17900 21924 17948 21980
rect 18004 21924 18052 21980
rect 18108 21924 18118 21980
rect 26150 21924 26160 21980
rect 26216 21924 26264 21980
rect 26320 21924 26368 21980
rect 26424 21924 26434 21980
rect 34466 21924 34476 21980
rect 34532 21924 34580 21980
rect 34636 21924 34684 21980
rect 34740 21924 34750 21980
rect 15978 21868 15988 21924
rect 16044 21868 16604 21924
rect 16660 21868 16670 21924
rect 23314 21868 23324 21924
rect 23380 21868 23884 21924
rect 23940 21868 23950 21924
rect 17714 21756 17724 21812
rect 17780 21756 18564 21812
rect 18620 21756 18630 21812
rect 18732 21756 18902 21812
rect 18958 21756 19852 21812
rect 19908 21756 19918 21812
rect 21410 21756 21420 21812
rect 21476 21756 21868 21812
rect 21924 21756 22428 21812
rect 22484 21756 22494 21812
rect 23538 21756 23548 21812
rect 23604 21756 25788 21812
rect 25844 21756 26460 21812
rect 26516 21756 26526 21812
rect 30930 21756 30940 21812
rect 30996 21756 31948 21812
rect 18732 21588 18788 21756
rect 31892 21588 31948 21756
rect 3602 21532 3612 21588
rect 3668 21532 4060 21588
rect 4116 21532 4844 21588
rect 4900 21532 8316 21588
rect 8372 21532 8764 21588
rect 8820 21532 8830 21588
rect 12786 21532 12796 21588
rect 12852 21532 13132 21588
rect 13188 21532 14028 21588
rect 14084 21532 14094 21588
rect 16706 21532 16716 21588
rect 16772 21532 17724 21588
rect 17780 21532 18788 21588
rect 29474 21532 29484 21588
rect 29540 21532 29932 21588
rect 29988 21532 29998 21588
rect 31892 21532 32340 21588
rect 8418 21420 8428 21476
rect 8484 21420 9044 21476
rect 9100 21420 11564 21476
rect 11620 21420 22932 21476
rect 22988 21420 23772 21476
rect 23828 21420 25564 21476
rect 25620 21420 25630 21476
rect 30706 21420 30716 21476
rect 30772 21420 31836 21476
rect 31892 21420 31902 21476
rect 32284 21420 32340 21532
rect 32396 21420 32406 21476
rect 18162 21308 18172 21364
rect 18228 21308 18396 21364
rect 18452 21308 18462 21364
rect 21970 21308 21980 21364
rect 22036 21308 22484 21364
rect 22428 21252 22484 21308
rect 22428 21196 22988 21252
rect 23044 21196 23054 21252
rect 5360 21140 5370 21196
rect 5426 21140 5474 21196
rect 5530 21140 5578 21196
rect 5634 21140 5644 21196
rect 13676 21140 13686 21196
rect 13742 21140 13790 21196
rect 13846 21140 13894 21196
rect 13950 21140 13960 21196
rect 21992 21140 22002 21196
rect 22058 21140 22106 21196
rect 22162 21140 22210 21196
rect 22266 21140 22276 21196
rect 30308 21140 30318 21196
rect 30374 21140 30422 21196
rect 30478 21140 30526 21196
rect 30582 21140 30592 21196
rect 5002 20972 5012 21028
rect 5068 20972 5628 21028
rect 5684 20972 5694 21028
rect 21634 20972 21644 21028
rect 21700 20972 22876 21028
rect 22932 20972 22942 21028
rect 29082 20972 29092 21028
rect 29148 20972 31836 21028
rect 31892 20972 31902 21028
rect 3658 20860 3668 20916
rect 3724 20860 4172 20916
rect 4228 20860 7196 20916
rect 7252 20860 7262 20916
rect 5954 20748 5964 20804
rect 6020 20748 9212 20804
rect 9268 20748 9278 20804
rect 11778 20748 11788 20804
rect 11844 20748 13020 20804
rect 13076 20748 13086 20804
rect 20066 20748 20076 20804
rect 20132 20748 21364 20804
rect 21420 20748 21430 20804
rect 22082 20748 22092 20804
rect 22148 20748 22316 20804
rect 22372 20748 22382 20804
rect 22586 20748 22596 20804
rect 22652 20748 26124 20804
rect 26180 20748 26684 20804
rect 26740 20748 26750 20804
rect 27738 20748 27748 20804
rect 27804 20748 29148 20804
rect 29204 20748 29214 20804
rect 30818 20748 30828 20804
rect 30884 20748 32060 20804
rect 32116 20748 32126 20804
rect 3938 20636 3948 20692
rect 4004 20636 4014 20692
rect 21746 20636 21756 20692
rect 21812 20636 22764 20692
rect 22820 20636 22830 20692
rect 3948 20132 4004 20636
rect 20682 20524 20692 20580
rect 20748 20524 22092 20580
rect 22148 20524 22428 20580
rect 22484 20524 22494 20580
rect 12506 20412 12516 20468
rect 12572 20412 12796 20468
rect 12852 20412 12862 20468
rect 22530 20412 22540 20468
rect 22596 20412 23324 20468
rect 23380 20412 23390 20468
rect 9518 20356 9528 20412
rect 9584 20356 9632 20412
rect 9688 20356 9736 20412
rect 9792 20356 9802 20412
rect 17834 20356 17844 20412
rect 17900 20356 17948 20412
rect 18004 20356 18052 20412
rect 18108 20356 18118 20412
rect 26150 20356 26160 20412
rect 26216 20356 26264 20412
rect 26320 20356 26368 20412
rect 26424 20356 26434 20412
rect 34466 20356 34476 20412
rect 34532 20356 34580 20412
rect 34636 20356 34684 20412
rect 34740 20356 34750 20412
rect 4498 20300 4508 20356
rect 4564 20300 5796 20356
rect 5852 20300 5862 20356
rect 13346 20300 13356 20356
rect 13412 20300 16044 20356
rect 16100 20300 16110 20356
rect 23874 20300 23884 20356
rect 23940 20300 24220 20356
rect 24276 20300 24286 20356
rect 16146 20188 16156 20244
rect 16212 20188 17724 20244
rect 17780 20188 17790 20244
rect 22978 20188 22988 20244
rect 23044 20188 23548 20244
rect 23604 20188 27748 20244
rect 27804 20188 27814 20244
rect 28466 20188 28476 20244
rect 28532 20188 28542 20244
rect 28476 20132 28532 20188
rect 2818 20076 2828 20132
rect 2884 20076 3612 20132
rect 3668 20076 4004 20132
rect 5506 20076 5516 20132
rect 5572 20076 7084 20132
rect 7140 20076 7150 20132
rect 12674 20076 12684 20132
rect 12740 20076 13468 20132
rect 13524 20076 13534 20132
rect 28476 20076 28924 20132
rect 28980 20076 28990 20132
rect 29922 20076 29932 20132
rect 29988 20076 30604 20132
rect 30660 20076 30670 20132
rect 3956 19964 3966 20020
rect 4022 19964 4284 20020
rect 4340 19964 4350 20020
rect 4722 19964 4732 20020
rect 4788 19964 5852 20020
rect 5908 19964 5918 20020
rect 7522 19964 7532 20020
rect 7588 19964 8820 20020
rect 8876 19964 8886 20020
rect 9426 19964 9436 20020
rect 9492 19964 10332 20020
rect 10388 19964 13860 20020
rect 13916 19964 13926 20020
rect 14018 19964 14028 20020
rect 14084 19964 18844 20020
rect 18900 19964 18910 20020
rect 22530 19964 22540 20020
rect 22596 19964 22764 20020
rect 22820 19964 22830 20020
rect 27010 19964 27020 20020
rect 27076 19964 28028 20020
rect 28084 19964 29596 20020
rect 29652 19964 31388 20020
rect 31444 19964 31454 20020
rect 3714 19852 3724 19908
rect 3780 19852 4508 19908
rect 4564 19852 4574 19908
rect 11554 19852 11564 19908
rect 11620 19852 12684 19908
rect 12740 19852 12750 19908
rect 19394 19852 19404 19908
rect 19460 19852 21532 19908
rect 21588 19852 21980 19908
rect 22036 19852 22046 19908
rect 29362 19852 29372 19908
rect 29428 19852 30268 19908
rect 30324 19852 30334 19908
rect 13010 19740 13020 19796
rect 13076 19740 14420 19796
rect 14364 19684 14420 19740
rect 14354 19628 14364 19684
rect 14420 19628 14812 19684
rect 14868 19628 14878 19684
rect 5360 19572 5370 19628
rect 5426 19572 5474 19628
rect 5530 19572 5578 19628
rect 5634 19572 5644 19628
rect 13676 19572 13686 19628
rect 13742 19572 13790 19628
rect 13846 19572 13894 19628
rect 13950 19572 13960 19628
rect 21992 19572 22002 19628
rect 22058 19572 22106 19628
rect 22162 19572 22210 19628
rect 22266 19572 22276 19628
rect 30308 19572 30318 19628
rect 30374 19572 30422 19628
rect 30478 19572 30526 19628
rect 30582 19572 30592 19628
rect 14028 19516 14140 19572
rect 14196 19516 14206 19572
rect 32162 19516 32172 19572
rect 32228 19516 32956 19572
rect 33012 19516 33022 19572
rect 14028 19460 14084 19516
rect 13906 19404 13916 19460
rect 13972 19404 14084 19460
rect 14578 19404 14588 19460
rect 14644 19404 15596 19460
rect 15652 19404 16324 19460
rect 16380 19404 16390 19460
rect 7186 19292 7196 19348
rect 7252 19292 8540 19348
rect 8596 19292 8606 19348
rect 13794 19292 13804 19348
rect 13860 19292 16604 19348
rect 16660 19292 16670 19348
rect 28802 19292 28812 19348
rect 28868 19292 29148 19348
rect 29204 19292 29214 19348
rect 4946 19180 4956 19236
rect 5012 19180 7308 19236
rect 7364 19180 7374 19236
rect 12954 19180 12964 19236
rect 13020 19180 13524 19236
rect 13580 19180 13590 19236
rect 15026 19180 15036 19236
rect 15092 19180 16492 19236
rect 16548 19180 16558 19236
rect 16874 19180 16884 19236
rect 16940 19180 18284 19236
rect 18340 19180 18732 19236
rect 18788 19180 18798 19236
rect 19730 19180 19740 19236
rect 19796 19180 20972 19236
rect 21028 19180 21364 19236
rect 21420 19180 21430 19236
rect 22194 19180 22204 19236
rect 22260 19180 23884 19236
rect 23940 19180 23950 19236
rect 18732 19124 18788 19180
rect 18732 19068 19964 19124
rect 20020 19068 20030 19124
rect 31602 19068 31612 19124
rect 31668 19068 32284 19124
rect 32340 19068 33292 19124
rect 33348 19068 33358 19124
rect 30090 18956 30100 19012
rect 30156 18956 31276 19012
rect 31332 18956 34300 19012
rect 34356 18956 34366 19012
rect 3266 18844 3276 18900
rect 3332 18844 3948 18900
rect 4004 18844 6416 18900
rect 6472 18844 8428 18900
rect 8484 18844 8494 18900
rect 12114 18844 12124 18900
rect 12180 18844 13132 18900
rect 13188 18844 13198 18900
rect 9518 18788 9528 18844
rect 9584 18788 9632 18844
rect 9688 18788 9736 18844
rect 9792 18788 9802 18844
rect 17834 18788 17844 18844
rect 17900 18788 17948 18844
rect 18004 18788 18052 18844
rect 18108 18788 18118 18844
rect 26150 18788 26160 18844
rect 26216 18788 26264 18844
rect 26320 18788 26368 18844
rect 26424 18788 26434 18844
rect 34466 18788 34476 18844
rect 34532 18788 34580 18844
rect 34636 18788 34684 18844
rect 34740 18788 34750 18844
rect 3826 18732 3836 18788
rect 3892 18732 4900 18788
rect 4956 18732 7196 18788
rect 7252 18732 7262 18788
rect 16566 18732 16604 18788
rect 16660 18732 16670 18788
rect 6402 18620 6412 18676
rect 6468 18620 8540 18676
rect 8596 18620 9100 18676
rect 9156 18620 9166 18676
rect 17714 18620 17724 18676
rect 17780 18620 20188 18676
rect 20132 18564 20188 18620
rect 6290 18508 6300 18564
rect 6356 18508 7084 18564
rect 7140 18508 7150 18564
rect 14036 18508 14046 18564
rect 14102 18508 15596 18564
rect 15652 18508 15662 18564
rect 18834 18508 18844 18564
rect 18900 18508 19404 18564
rect 19460 18508 19470 18564
rect 20132 18508 20300 18564
rect 20356 18508 20366 18564
rect 31042 18508 31052 18564
rect 31108 18508 31948 18564
rect 32004 18508 33404 18564
rect 33460 18508 33470 18564
rect 2594 18396 2604 18452
rect 2660 18396 4060 18452
rect 4116 18396 4126 18452
rect 7746 18396 7756 18452
rect 7812 18396 8428 18452
rect 8484 18396 8494 18452
rect 12338 18396 12348 18452
rect 12404 18396 12684 18452
rect 12740 18396 19516 18452
rect 19572 18396 19582 18452
rect 20738 18396 20748 18452
rect 20804 18396 22428 18452
rect 22484 18396 22494 18452
rect 27682 18396 27692 18452
rect 27748 18396 28700 18452
rect 28756 18396 29484 18452
rect 29540 18396 29550 18452
rect 30146 18396 30156 18452
rect 30212 18396 31612 18452
rect 31668 18396 31678 18452
rect 3378 18284 3388 18340
rect 3444 18284 4508 18340
rect 4564 18284 5292 18340
rect 5348 18284 5740 18340
rect 5796 18284 5806 18340
rect 7988 18284 7998 18340
rect 8054 18284 8988 18340
rect 9044 18284 9054 18340
rect 11218 18284 11228 18340
rect 11284 18284 12236 18340
rect 12292 18284 14924 18340
rect 14980 18284 17724 18340
rect 17780 18284 17790 18340
rect 27122 18284 27132 18340
rect 27188 18284 30604 18340
rect 30660 18284 30670 18340
rect 30930 18284 30940 18340
rect 30996 18284 31948 18340
rect 32004 18284 32014 18340
rect 4050 18172 4060 18228
rect 4116 18172 7644 18228
rect 7700 18172 7710 18228
rect 12002 18172 12012 18228
rect 12068 18172 13804 18228
rect 13860 18172 13870 18228
rect 15250 18172 15260 18228
rect 15316 18172 16324 18228
rect 16380 18172 16390 18228
rect 29250 18172 29260 18228
rect 29316 18172 31388 18228
rect 31444 18172 31454 18228
rect 31714 18172 31724 18228
rect 31780 18172 33124 18228
rect 33180 18172 33190 18228
rect 12730 18060 12740 18116
rect 12796 18060 13300 18116
rect 13356 18060 13366 18116
rect 14466 18060 14476 18116
rect 14532 18060 17724 18116
rect 17780 18060 17790 18116
rect 5360 18004 5370 18060
rect 5426 18004 5474 18060
rect 5530 18004 5578 18060
rect 5634 18004 5644 18060
rect 13676 18004 13686 18060
rect 13742 18004 13790 18060
rect 13846 18004 13894 18060
rect 13950 18004 13960 18060
rect 21992 18004 22002 18060
rect 22058 18004 22106 18060
rect 22162 18004 22210 18060
rect 22266 18004 22276 18060
rect 30308 18004 30318 18060
rect 30374 18004 30422 18060
rect 30478 18004 30526 18060
rect 30582 18004 30592 18060
rect 14242 17948 14252 18004
rect 14308 17948 15596 18004
rect 15652 17948 15662 18004
rect 15754 17948 15764 18004
rect 15820 17948 18508 18004
rect 18564 17948 18574 18004
rect 18722 17948 18732 18004
rect 18788 17948 20860 18004
rect 20916 17948 20926 18004
rect 22754 17948 22764 18004
rect 22820 17948 22988 18004
rect 23044 17948 23054 18004
rect 3602 17836 3612 17892
rect 3668 17836 4060 17892
rect 4116 17836 4396 17892
rect 4452 17836 5964 17892
rect 6020 17836 6030 17892
rect 14914 17836 14924 17892
rect 14980 17836 15932 17892
rect 15988 17836 15998 17892
rect 17266 17836 17276 17892
rect 17332 17836 17500 17892
rect 17556 17836 19348 17892
rect 19404 17836 19414 17892
rect 20178 17836 20188 17892
rect 20244 17836 20636 17892
rect 20692 17836 22652 17892
rect 22708 17836 22718 17892
rect 7634 17724 7644 17780
rect 7700 17724 8092 17780
rect 8148 17724 8316 17780
rect 8372 17724 8382 17780
rect 12002 17724 12012 17780
rect 12068 17724 12796 17780
rect 12852 17724 12862 17780
rect 14242 17724 14252 17780
rect 14308 17724 14812 17780
rect 14868 17724 15484 17780
rect 15540 17724 18732 17780
rect 18788 17724 18798 17780
rect 18956 17724 20300 17780
rect 20356 17724 21084 17780
rect 21140 17724 21150 17780
rect 18956 17668 19012 17724
rect 4274 17612 4284 17668
rect 4340 17612 5740 17668
rect 5796 17612 6300 17668
rect 6356 17612 6366 17668
rect 7746 17612 7756 17668
rect 7812 17612 7822 17668
rect 11890 17612 11900 17668
rect 11956 17612 12628 17668
rect 12684 17612 12694 17668
rect 13122 17612 13132 17668
rect 13188 17612 13580 17668
rect 13636 17612 16156 17668
rect 16212 17612 17052 17668
rect 17108 17612 17118 17668
rect 17826 17612 17836 17668
rect 17892 17612 18956 17668
rect 19012 17612 19022 17668
rect 19506 17612 19516 17668
rect 19572 17612 23548 17668
rect 23604 17612 25452 17668
rect 25508 17612 25518 17668
rect 27570 17612 27580 17668
rect 27636 17612 28140 17668
rect 28196 17612 28364 17668
rect 28420 17612 28430 17668
rect 28578 17612 28588 17668
rect 28644 17612 30492 17668
rect 30548 17612 30558 17668
rect 30706 17612 30716 17668
rect 30772 17612 31724 17668
rect 31780 17612 31790 17668
rect 32274 17612 32284 17668
rect 32340 17612 33516 17668
rect 33572 17612 33582 17668
rect 7756 17556 7812 17612
rect 4162 17500 4172 17556
rect 4228 17500 4956 17556
rect 5012 17500 6972 17556
rect 7028 17500 7812 17556
rect 10882 17500 10892 17556
rect 10948 17500 14980 17556
rect 15036 17500 15046 17556
rect 19730 17500 19740 17556
rect 19796 17500 22764 17556
rect 22820 17500 23156 17556
rect 23212 17500 23222 17556
rect 27768 17500 27778 17556
rect 27834 17500 28476 17556
rect 28532 17500 28542 17556
rect 29474 17500 29484 17556
rect 29540 17500 32060 17556
rect 32116 17500 32126 17556
rect 7298 17388 7308 17444
rect 7364 17388 7812 17444
rect 7868 17388 8764 17444
rect 8820 17388 8830 17444
rect 3938 17276 3948 17332
rect 4004 17276 4228 17332
rect 18722 17276 18732 17332
rect 18788 17276 20076 17332
rect 20132 17276 22484 17332
rect 22540 17276 22550 17332
rect 27122 17276 27132 17332
rect 27188 17276 27692 17332
rect 27748 17276 27758 17332
rect 4172 16884 4228 17276
rect 9518 17220 9528 17276
rect 9584 17220 9632 17276
rect 9688 17220 9736 17276
rect 9792 17220 9802 17276
rect 17834 17220 17844 17276
rect 17900 17220 17948 17276
rect 18004 17220 18052 17276
rect 18108 17220 18118 17276
rect 26150 17220 26160 17276
rect 26216 17220 26264 17276
rect 26320 17220 26368 17276
rect 26424 17220 26434 17276
rect 34466 17220 34476 17276
rect 34532 17220 34580 17276
rect 34636 17220 34684 17276
rect 34740 17220 34750 17276
rect 19898 17164 19908 17220
rect 19964 17164 21308 17220
rect 21364 17164 21374 17220
rect 17826 17052 17836 17108
rect 17892 17052 21196 17108
rect 21252 17052 21262 17108
rect 31602 17052 31612 17108
rect 31668 17052 31678 17108
rect 21298 16940 21308 16996
rect 21364 16940 23604 16996
rect 23660 16940 23670 16996
rect 26908 16940 28924 16996
rect 28980 16940 28990 16996
rect 4162 16828 4172 16884
rect 4228 16828 4238 16884
rect 4498 16828 4508 16884
rect 4564 16828 6300 16884
rect 6356 16828 6366 16884
rect 10434 16828 10444 16884
rect 10500 16828 11340 16884
rect 11396 16828 12927 16884
rect 12983 16828 14700 16884
rect 14756 16828 14766 16884
rect 19292 16828 20748 16884
rect 20804 16828 20814 16884
rect 21970 16828 21980 16884
rect 22036 16828 23436 16884
rect 23492 16828 23502 16884
rect 8530 16716 8540 16772
rect 8596 16716 9436 16772
rect 9492 16716 9502 16772
rect 14018 16716 14028 16772
rect 14084 16716 14364 16772
rect 14420 16716 14430 16772
rect 16706 16716 16716 16772
rect 16772 16716 18396 16772
rect 18452 16716 18462 16772
rect 19292 16660 19348 16828
rect 22846 16716 22856 16772
rect 22912 16716 23324 16772
rect 23380 16716 24220 16772
rect 24276 16716 24286 16772
rect 19282 16604 19292 16660
rect 19348 16604 19358 16660
rect 26908 16548 26964 16940
rect 31612 16884 31668 17052
rect 28466 16828 28476 16884
rect 28532 16828 29484 16884
rect 29540 16828 29550 16884
rect 30146 16828 30156 16884
rect 30212 16828 30828 16884
rect 30884 16828 30894 16884
rect 31042 16828 31052 16884
rect 31108 16828 31668 16884
rect 31826 16828 31836 16884
rect 31892 16828 31948 16884
rect 32004 16828 32014 16884
rect 28018 16716 28028 16772
rect 28084 16716 29316 16772
rect 29372 16716 29382 16772
rect 27122 16604 27132 16660
rect 27188 16604 28476 16660
rect 28532 16604 28542 16660
rect 26898 16492 26908 16548
rect 26964 16492 26974 16548
rect 5360 16436 5370 16492
rect 5426 16436 5474 16492
rect 5530 16436 5578 16492
rect 5634 16436 5644 16492
rect 13676 16436 13686 16492
rect 13742 16436 13790 16492
rect 13846 16436 13894 16492
rect 13950 16436 13960 16492
rect 21992 16436 22002 16492
rect 22058 16436 22106 16492
rect 22162 16436 22210 16492
rect 22266 16436 22276 16492
rect 30308 16436 30318 16492
rect 30374 16436 30422 16492
rect 30478 16436 30526 16492
rect 30582 16436 30592 16492
rect 21522 16268 21532 16324
rect 21588 16268 22316 16324
rect 22372 16268 22382 16324
rect 26282 16268 26292 16324
rect 26348 16268 27132 16324
rect 27188 16268 27198 16324
rect 29306 16156 29316 16212
rect 29372 16156 31220 16212
rect 31276 16156 31286 16212
rect 1810 16044 1820 16100
rect 1876 16044 4900 16100
rect 4956 16044 5124 16100
rect 5180 16044 5852 16100
rect 5908 16044 7868 16100
rect 7924 16044 8540 16100
rect 8596 16044 8606 16100
rect 17714 16044 17724 16100
rect 17780 16044 19516 16100
rect 19572 16044 19582 16100
rect 25330 16044 25340 16100
rect 25396 16044 26124 16100
rect 26180 16044 27972 16100
rect 28028 16044 28038 16100
rect 27514 15932 27524 15988
rect 27580 15932 28532 15988
rect 28588 15932 28598 15988
rect 11162 15820 11172 15876
rect 11228 15820 12516 15876
rect 12572 15820 12582 15876
rect 27794 15708 27804 15764
rect 27860 15708 28700 15764
rect 28756 15708 30156 15764
rect 30212 15708 30222 15764
rect 9518 15652 9528 15708
rect 9584 15652 9632 15708
rect 9688 15652 9736 15708
rect 9792 15652 9802 15708
rect 17834 15652 17844 15708
rect 17900 15652 17948 15708
rect 18004 15652 18052 15708
rect 18108 15652 18118 15708
rect 26150 15652 26160 15708
rect 26216 15652 26264 15708
rect 26320 15652 26368 15708
rect 26424 15652 26434 15708
rect 34466 15652 34476 15708
rect 34532 15652 34580 15708
rect 34636 15652 34684 15708
rect 34740 15652 34750 15708
rect 15922 15484 15932 15540
rect 15988 15484 17836 15540
rect 17892 15484 18844 15540
rect 18900 15484 18910 15540
rect 28242 15484 28252 15540
rect 28308 15484 28924 15540
rect 28980 15484 28990 15540
rect 14018 15372 14028 15428
rect 14084 15372 14644 15428
rect 14700 15372 18340 15428
rect 18396 15372 18406 15428
rect 30146 15372 30156 15428
rect 30212 15372 32956 15428
rect 33012 15372 33022 15428
rect 7970 15260 7980 15316
rect 8036 15260 8988 15316
rect 9044 15260 9772 15316
rect 9828 15260 11172 15316
rect 11228 15260 11238 15316
rect 27570 15260 27580 15316
rect 27636 15260 29148 15316
rect 29204 15260 29214 15316
rect 14914 15148 14924 15204
rect 14980 15148 16268 15204
rect 16324 15148 16716 15204
rect 16772 15148 16782 15204
rect 19058 15148 19068 15204
rect 19124 15148 21532 15204
rect 21588 15148 22372 15204
rect 22428 15148 23436 15204
rect 23492 15148 24780 15204
rect 24836 15148 24846 15204
rect 26898 15148 26908 15204
rect 26964 15148 27356 15204
rect 27412 15148 27422 15204
rect 16482 15036 16492 15092
rect 16548 15036 17164 15092
rect 17220 15036 17230 15092
rect 28466 15036 28476 15092
rect 28532 15036 29148 15092
rect 29204 15036 29214 15092
rect 5360 14868 5370 14924
rect 5426 14868 5474 14924
rect 5530 14868 5578 14924
rect 5634 14868 5644 14924
rect 13676 14868 13686 14924
rect 13742 14868 13790 14924
rect 13846 14868 13894 14924
rect 13950 14868 13960 14924
rect 21992 14868 22002 14924
rect 22058 14868 22106 14924
rect 22162 14868 22210 14924
rect 22266 14868 22276 14924
rect 30308 14868 30318 14924
rect 30374 14868 30422 14924
rect 30478 14868 30526 14924
rect 30582 14868 30592 14924
rect 31826 14812 31836 14868
rect 31892 14756 31948 14868
rect 6178 14700 6188 14756
rect 6244 14700 6748 14756
rect 6804 14700 6814 14756
rect 7298 14700 7308 14756
rect 7364 14700 8204 14756
rect 8260 14700 8270 14756
rect 31892 14700 32060 14756
rect 32116 14700 32126 14756
rect 27122 14588 27132 14644
rect 27188 14588 27356 14644
rect 27412 14588 27422 14644
rect 28354 14588 28364 14644
rect 28420 14588 29036 14644
rect 29092 14588 29372 14644
rect 29428 14588 29438 14644
rect 3350 14476 3388 14532
rect 3444 14476 3454 14532
rect 26021 14476 26031 14532
rect 26087 14476 27692 14532
rect 27748 14476 29540 14532
rect 29596 14476 29606 14532
rect 30426 14476 30436 14532
rect 30492 14476 34300 14532
rect 34356 14476 34366 14532
rect 25330 14364 25340 14420
rect 25396 14364 25788 14420
rect 25844 14364 25854 14420
rect 30930 14364 30940 14420
rect 30996 14364 31612 14420
rect 31668 14364 31678 14420
rect 17266 14252 17276 14308
rect 17332 14252 17724 14308
rect 17780 14252 18172 14308
rect 18228 14252 18238 14308
rect 9518 14084 9528 14140
rect 9584 14084 9632 14140
rect 9688 14084 9736 14140
rect 9792 14084 9802 14140
rect 17834 14084 17844 14140
rect 17900 14084 17948 14140
rect 18004 14084 18052 14140
rect 18108 14084 18118 14140
rect 26150 14084 26160 14140
rect 26216 14084 26264 14140
rect 26320 14084 26368 14140
rect 26424 14084 26434 14140
rect 34466 14084 34476 14140
rect 34532 14084 34580 14140
rect 34636 14084 34684 14140
rect 34740 14084 34750 14140
rect 15138 13916 15148 13972
rect 15204 13916 16604 13972
rect 16660 13916 22932 13972
rect 22988 13916 23212 13972
rect 23268 13916 23278 13972
rect 2930 13804 2940 13860
rect 2996 13804 3612 13860
rect 3668 13804 4956 13860
rect 5012 13804 5022 13860
rect 16492 13804 17836 13860
rect 17892 13804 17902 13860
rect 26450 13804 26460 13860
rect 26516 13804 30716 13860
rect 30772 13804 30782 13860
rect 16492 13748 16548 13804
rect 3042 13692 3052 13748
rect 3108 13692 3836 13748
rect 3892 13692 3902 13748
rect 16370 13692 16380 13748
rect 16436 13692 16492 13748
rect 16548 13692 16558 13748
rect 16650 13692 16660 13748
rect 16716 13692 17500 13748
rect 17556 13692 18004 13748
rect 18060 13692 18070 13748
rect 18498 13692 18508 13748
rect 18564 13692 18844 13748
rect 18900 13692 18910 13748
rect 23314 13692 23324 13748
rect 23380 13692 28700 13748
rect 28756 13692 28766 13748
rect 2818 13580 2828 13636
rect 2884 13580 4060 13636
rect 4116 13580 4126 13636
rect 4442 13580 4452 13636
rect 4508 13580 7084 13636
rect 7140 13580 7150 13636
rect 14466 13580 14476 13636
rect 14532 13580 15148 13636
rect 16370 13580 16380 13636
rect 16436 13580 17780 13636
rect 18610 13580 18620 13636
rect 18676 13580 18956 13636
rect 19012 13580 19022 13636
rect 23090 13580 23100 13636
rect 23156 13580 23436 13636
rect 23492 13580 24164 13636
rect 24220 13580 24230 13636
rect 26674 13580 26684 13636
rect 26740 13580 29260 13636
rect 29316 13580 29326 13636
rect 15092 13524 15148 13580
rect 17724 13524 17780 13580
rect 2258 13468 2268 13524
rect 2324 13468 3612 13524
rect 3668 13468 3678 13524
rect 15092 13468 16716 13524
rect 16772 13468 16782 13524
rect 16930 13468 16940 13524
rect 16996 13468 17444 13524
rect 17500 13468 17510 13524
rect 17714 13468 17724 13524
rect 17780 13468 18564 13524
rect 18620 13468 18630 13524
rect 23884 13468 25228 13524
rect 25284 13468 25294 13524
rect 25778 13468 25788 13524
rect 25844 13468 26460 13524
rect 26516 13468 26908 13524
rect 26964 13468 26974 13524
rect 5360 13300 5370 13356
rect 5426 13300 5474 13356
rect 5530 13300 5578 13356
rect 5634 13300 5644 13356
rect 13676 13300 13686 13356
rect 13742 13300 13790 13356
rect 13846 13300 13894 13356
rect 13950 13300 13960 13356
rect 21992 13300 22002 13356
rect 22058 13300 22106 13356
rect 22162 13300 22210 13356
rect 22266 13300 22276 13356
rect 23884 13300 23940 13468
rect 31714 13356 31724 13412
rect 31780 13356 32284 13412
rect 32340 13356 33068 13412
rect 33124 13356 33852 13412
rect 33908 13356 33918 13412
rect 30308 13300 30318 13356
rect 30374 13300 30422 13356
rect 30478 13300 30526 13356
rect 30582 13300 30592 13356
rect 9874 13244 9884 13300
rect 9940 13244 11340 13300
rect 11396 13244 11406 13300
rect 23874 13244 23884 13300
rect 23940 13244 23950 13300
rect 7746 13132 7756 13188
rect 7812 13132 14028 13188
rect 14084 13132 14094 13188
rect 21298 13132 21308 13188
rect 21364 13132 22652 13188
rect 22708 13132 22718 13188
rect 5730 13020 5740 13076
rect 5796 13020 9324 13076
rect 9380 13020 10164 13076
rect 10220 13020 10836 13076
rect 11330 13020 11340 13076
rect 11396 13020 14364 13076
rect 14420 13020 15148 13076
rect 16258 13020 16268 13076
rect 16324 13020 18956 13076
rect 19012 13020 19022 13076
rect 10780 12964 10836 13020
rect 15092 12964 15148 13020
rect 2706 12908 2716 12964
rect 2772 12908 3388 12964
rect 3444 12908 3454 12964
rect 4050 12908 4060 12964
rect 4116 12908 5964 12964
rect 6020 12908 6300 12964
rect 6356 12908 6366 12964
rect 6962 12908 6972 12964
rect 7028 12908 7644 12964
rect 7700 12908 7710 12964
rect 10770 12908 10780 12964
rect 10836 12908 10846 12964
rect 12002 12908 12012 12964
rect 12068 12908 12236 12964
rect 12292 12908 14588 12964
rect 14644 12908 14654 12964
rect 15092 12908 15596 12964
rect 15652 12908 16828 12964
rect 16884 12908 16894 12964
rect 17490 12908 17500 12964
rect 17556 12908 18508 12964
rect 18564 12908 18574 12964
rect 20178 12908 20188 12964
rect 20244 12908 21532 12964
rect 21588 12908 21598 12964
rect 22398 12908 22408 12964
rect 22464 12908 23548 12964
rect 23604 12908 23614 12964
rect 28354 12908 28364 12964
rect 28420 12908 29036 12964
rect 29092 12908 29102 12964
rect 29922 12908 29932 12964
rect 29988 12908 31164 12964
rect 31220 12908 31230 12964
rect 32386 12908 32396 12964
rect 32452 12908 33628 12964
rect 33684 12908 33694 12964
rect 5058 12796 5068 12852
rect 5124 12796 10556 12852
rect 10612 12796 10622 12852
rect 15194 12796 15204 12852
rect 15260 12796 17892 12852
rect 17948 12740 18004 12852
rect 18162 12796 18172 12852
rect 18228 12796 19684 12852
rect 19740 12796 19750 12852
rect 30258 12796 30268 12852
rect 30324 12796 31276 12852
rect 31332 12796 31342 12852
rect 16342 12684 16380 12740
rect 16436 12684 16446 12740
rect 17948 12684 18284 12740
rect 18340 12684 18350 12740
rect 18806 12684 18844 12740
rect 18900 12684 18910 12740
rect 31602 12684 31612 12740
rect 31668 12684 33628 12740
rect 33684 12684 33694 12740
rect 8422 12572 8432 12628
rect 8488 12572 8498 12628
rect 8428 12516 8484 12572
rect 9518 12516 9528 12572
rect 9584 12516 9632 12572
rect 9688 12516 9736 12572
rect 9792 12516 9802 12572
rect 17834 12516 17844 12572
rect 17900 12516 17948 12572
rect 18004 12516 18052 12572
rect 18108 12516 18118 12572
rect 26150 12516 26160 12572
rect 26216 12516 26264 12572
rect 26320 12516 26368 12572
rect 26424 12516 26434 12572
rect 34466 12516 34476 12572
rect 34532 12516 34580 12572
rect 34636 12516 34684 12572
rect 34740 12516 34750 12572
rect 4284 12460 5516 12516
rect 5572 12460 5582 12516
rect 6514 12460 6524 12516
rect 6580 12460 8876 12516
rect 8932 12460 8942 12516
rect 12012 12460 12572 12516
rect 12628 12460 13692 12516
rect 13748 12460 13758 12516
rect 4284 12180 4340 12460
rect 12012 12404 12068 12460
rect 4508 12348 4732 12404
rect 4788 12348 12012 12404
rect 12068 12348 12078 12404
rect 12450 12348 12460 12404
rect 12516 12348 15316 12404
rect 15372 12348 15382 12404
rect 4508 12180 4564 12348
rect 18620 12292 18676 12404
rect 18732 12348 18742 12404
rect 6850 12236 6860 12292
rect 6916 12236 7532 12292
rect 7588 12236 7598 12292
rect 7746 12236 7756 12292
rect 7812 12236 8764 12292
rect 8820 12236 8830 12292
rect 10546 12236 10556 12292
rect 10612 12236 12516 12292
rect 15922 12236 15932 12292
rect 15988 12236 16492 12292
rect 16548 12236 16558 12292
rect 16650 12236 16660 12292
rect 16716 12236 18956 12292
rect 19012 12236 19516 12292
rect 19572 12236 19582 12292
rect 24210 12236 24220 12292
rect 24276 12236 29708 12292
rect 29764 12236 29774 12292
rect 12460 12180 12516 12236
rect 2650 12124 2660 12180
rect 2716 12124 3836 12180
rect 3892 12124 4284 12180
rect 4340 12124 4350 12180
rect 4498 12124 4508 12180
rect 4564 12124 4574 12180
rect 7970 12124 7980 12180
rect 8036 12124 8428 12180
rect 8484 12124 8494 12180
rect 10938 12124 10948 12180
rect 11004 12124 11228 12180
rect 11284 12124 11900 12180
rect 11956 12124 11966 12180
rect 12460 12124 14196 12180
rect 14252 12124 17388 12180
rect 17444 12124 17454 12180
rect 18050 12124 18060 12180
rect 18116 12124 18732 12180
rect 18788 12124 18798 12180
rect 29362 12124 29372 12180
rect 29428 12124 31164 12180
rect 31220 12124 31230 12180
rect 31378 12124 31388 12180
rect 31444 12124 31836 12180
rect 31892 12124 31902 12180
rect 3266 12012 3276 12068
rect 3332 12012 8316 12068
rect 8372 12012 11340 12068
rect 11396 12012 11406 12068
rect 16818 12012 16828 12068
rect 16884 12012 18620 12068
rect 18676 12012 18686 12068
rect 3042 11900 3052 11956
rect 3108 11900 5068 11956
rect 5124 11900 5134 11956
rect 6962 11900 6972 11956
rect 7028 11900 9884 11956
rect 9940 11900 9950 11956
rect 3826 11788 3836 11844
rect 3892 11788 5180 11844
rect 5236 11788 5246 11844
rect 6738 11788 6748 11844
rect 6804 11788 7140 11844
rect 7196 11788 7206 11844
rect 8372 11788 8876 11844
rect 8932 11788 11564 11844
rect 11620 11788 11630 11844
rect 14018 11788 14028 11844
rect 14084 11788 14980 11844
rect 15036 11788 15046 11844
rect 18722 11788 18732 11844
rect 18788 11788 18956 11844
rect 19012 11788 19022 11844
rect 25442 11788 25452 11844
rect 25508 11788 26124 11844
rect 26180 11788 28028 11844
rect 28084 11788 29316 11844
rect 29372 11788 29382 11844
rect 31266 11788 31276 11844
rect 31332 11788 32284 11844
rect 32340 11788 32350 11844
rect 5360 11732 5370 11788
rect 5426 11732 5474 11788
rect 5530 11732 5578 11788
rect 5634 11732 5644 11788
rect 8372 11732 8428 11788
rect 13676 11732 13686 11788
rect 13742 11732 13790 11788
rect 13846 11732 13894 11788
rect 13950 11732 13960 11788
rect 21992 11732 22002 11788
rect 22058 11732 22106 11788
rect 22162 11732 22210 11788
rect 22266 11732 22276 11788
rect 30308 11732 30318 11788
rect 30374 11732 30422 11788
rect 30478 11732 30526 11788
rect 30582 11732 30592 11788
rect 6178 11676 6188 11732
rect 6244 11676 8428 11732
rect 8642 11676 8652 11732
rect 8708 11676 9212 11732
rect 9268 11676 9278 11732
rect 14578 11676 14588 11732
rect 14644 11676 17052 11732
rect 17108 11676 17118 11732
rect 10322 11564 10332 11620
rect 10388 11564 11116 11620
rect 11172 11564 11452 11620
rect 11508 11564 12572 11620
rect 12628 11564 13356 11620
rect 13412 11564 13422 11620
rect 14802 11564 14812 11620
rect 14868 11564 16044 11620
rect 16100 11564 16110 11620
rect 19394 11564 19404 11620
rect 19460 11564 19470 11620
rect 26002 11564 26012 11620
rect 26068 11564 27132 11620
rect 27188 11564 27198 11620
rect 7410 11452 7420 11508
rect 7476 11452 7756 11508
rect 7812 11452 7822 11508
rect 15810 11452 15820 11508
rect 15876 11452 16380 11508
rect 16436 11452 16446 11508
rect 4498 11340 4508 11396
rect 4564 11340 9660 11396
rect 9716 11340 15148 11396
rect 15204 11340 15214 11396
rect 15530 11340 15540 11396
rect 15596 11340 17668 11396
rect 17724 11340 17734 11396
rect 4722 11228 4732 11284
rect 4788 11228 7084 11284
rect 7140 11228 7150 11284
rect 14466 11228 14476 11284
rect 14532 11228 14700 11284
rect 14756 11228 15148 11284
rect 15092 11172 15148 11228
rect 19404 11172 19460 11564
rect 24322 11452 24332 11508
rect 24388 11452 25340 11508
rect 25396 11452 25406 11508
rect 24714 11340 24724 11396
rect 24780 11340 25116 11396
rect 25172 11340 25900 11396
rect 25956 11340 26908 11396
rect 26964 11340 27580 11396
rect 27636 11340 29764 11396
rect 29820 11340 29830 11396
rect 2706 11116 2716 11172
rect 2772 11116 3220 11172
rect 3276 11116 4284 11172
rect 4340 11116 4350 11172
rect 10210 11116 10220 11172
rect 10276 11116 11116 11172
rect 11172 11116 11182 11172
rect 12898 11116 12908 11172
rect 12964 11116 13524 11172
rect 13580 11116 13590 11172
rect 15092 11116 19460 11172
rect 3714 11004 3724 11060
rect 3780 11004 4956 11060
rect 5012 11004 5022 11060
rect 9518 10948 9528 11004
rect 9584 10948 9632 11004
rect 9688 10948 9736 11004
rect 9792 10948 9802 11004
rect 17834 10948 17844 11004
rect 17900 10948 17948 11004
rect 18004 10948 18052 11004
rect 18108 10948 18118 11004
rect 26150 10948 26160 11004
rect 26216 10948 26264 11004
rect 26320 10948 26368 11004
rect 26424 10948 26434 11004
rect 34466 10948 34476 11004
rect 34532 10948 34580 11004
rect 34636 10948 34684 11004
rect 34740 10948 34750 11004
rect 22530 10892 22540 10948
rect 22596 10892 23324 10948
rect 23380 10892 23390 10948
rect 5170 10780 5180 10836
rect 5236 10780 8428 10836
rect 8484 10780 10220 10836
rect 10276 10780 10286 10836
rect 15138 10780 15148 10836
rect 15204 10780 15708 10836
rect 15764 10780 15774 10836
rect 33170 10780 33180 10836
rect 33236 10780 33246 10836
rect 5842 10668 5852 10724
rect 5908 10668 8428 10724
rect 12226 10668 12236 10724
rect 12292 10668 12460 10724
rect 12516 10668 12796 10724
rect 12852 10668 14140 10724
rect 14196 10668 14206 10724
rect 3042 10556 3052 10612
rect 3108 10556 4620 10612
rect 4676 10556 4686 10612
rect 8372 10500 8428 10668
rect 33180 10612 33236 10780
rect 13122 10556 13132 10612
rect 13188 10556 13916 10612
rect 13972 10556 14812 10612
rect 14868 10556 14878 10612
rect 25330 10556 25340 10612
rect 25396 10556 29932 10612
rect 29988 10556 29998 10612
rect 30930 10556 30940 10612
rect 30996 10556 32956 10612
rect 33012 10556 34076 10612
rect 34132 10556 34142 10612
rect 8372 10444 12180 10500
rect 12236 10444 13188 10500
rect 24434 10444 24444 10500
rect 24500 10444 25228 10500
rect 25284 10444 25294 10500
rect 29586 10444 29596 10500
rect 29652 10444 30828 10500
rect 30884 10444 30894 10500
rect 13132 10388 13188 10444
rect 3826 10332 3836 10388
rect 3892 10332 5068 10388
rect 5124 10332 5628 10388
rect 5684 10332 9772 10388
rect 9828 10332 10444 10388
rect 10500 10332 10510 10388
rect 13122 10332 13132 10388
rect 13188 10332 13198 10388
rect 22866 10332 22876 10388
rect 22932 10332 25452 10388
rect 25508 10332 25518 10388
rect 9202 10220 9212 10276
rect 9268 10220 12012 10276
rect 12068 10220 12078 10276
rect 5360 10164 5370 10220
rect 5426 10164 5474 10220
rect 5530 10164 5578 10220
rect 5634 10164 5644 10220
rect 13676 10164 13686 10220
rect 13742 10164 13790 10220
rect 13846 10164 13894 10220
rect 13950 10164 13960 10220
rect 21992 10164 22002 10220
rect 22058 10164 22106 10220
rect 22162 10164 22210 10220
rect 22266 10164 22276 10220
rect 30308 10164 30318 10220
rect 30374 10164 30422 10220
rect 30478 10164 30526 10220
rect 30582 10164 30592 10220
rect 3602 10108 3612 10164
rect 3668 10108 4284 10164
rect 4340 10108 4350 10164
rect 4498 10108 4508 10164
rect 4564 10108 4602 10164
rect 3938 9996 3948 10052
rect 4004 9996 5740 10052
rect 5796 9996 6076 10052
rect 6132 9996 6142 10052
rect 11778 9996 11788 10052
rect 11844 9996 12348 10052
rect 12404 9996 12414 10052
rect 21298 9996 21308 10052
rect 21364 9996 22652 10052
rect 22708 9996 22718 10052
rect 23100 9996 23212 10052
rect 23268 9996 24780 10052
rect 24836 9996 24846 10052
rect 28018 9996 28028 10052
rect 28084 9996 29260 10052
rect 29316 9996 29326 10052
rect 23100 9940 23156 9996
rect 13122 9884 13132 9940
rect 13188 9884 17836 9940
rect 17892 9884 17902 9940
rect 21858 9884 21868 9940
rect 21924 9884 23156 9940
rect 23314 9884 23324 9940
rect 23380 9884 23940 9940
rect 23996 9884 24006 9940
rect 29586 9884 29596 9940
rect 29652 9884 30380 9940
rect 30436 9884 30446 9940
rect 2706 9772 2716 9828
rect 2772 9772 3836 9828
rect 3892 9772 3902 9828
rect 4834 9772 4844 9828
rect 4900 9772 5964 9828
rect 6020 9772 7084 9828
rect 7140 9772 7150 9828
rect 8418 9772 8428 9828
rect 8484 9772 9100 9828
rect 9156 9772 11396 9828
rect 11452 9772 11462 9828
rect 15586 9772 15596 9828
rect 15652 9772 16380 9828
rect 16436 9772 16446 9828
rect 21970 9772 21980 9828
rect 22036 9772 23100 9828
rect 23156 9772 26236 9828
rect 26292 9772 26302 9828
rect 27458 9772 27468 9828
rect 27524 9772 28588 9828
rect 28644 9772 29820 9828
rect 29876 9772 30716 9828
rect 30772 9772 30782 9828
rect 3266 9660 3276 9716
rect 3332 9660 4396 9716
rect 4452 9660 4462 9716
rect 7578 9660 7588 9716
rect 7644 9660 8652 9716
rect 8708 9660 8718 9716
rect 10882 9660 10892 9716
rect 10948 9660 11788 9716
rect 11844 9660 11854 9716
rect 28466 9660 28476 9716
rect 28532 9660 29372 9716
rect 29428 9660 33292 9716
rect 33348 9660 33358 9716
rect 3042 9548 3052 9604
rect 3108 9548 3724 9604
rect 3780 9548 3790 9604
rect 4610 9548 4620 9604
rect 4676 9548 4956 9604
rect 5012 9548 5022 9604
rect 6738 9548 6748 9604
rect 6804 9548 6916 9604
rect 6860 9380 6916 9548
rect 8372 9548 13020 9604
rect 13076 9548 13086 9604
rect 24210 9548 24220 9604
rect 24276 9548 25116 9604
rect 25172 9548 25182 9604
rect 28578 9548 28588 9604
rect 28644 9548 29932 9604
rect 29988 9548 31724 9604
rect 31780 9548 31790 9604
rect 8372 9492 8428 9548
rect 7298 9436 7308 9492
rect 7364 9436 7644 9492
rect 7700 9436 8428 9492
rect 11218 9436 11228 9492
rect 11284 9436 12908 9492
rect 12964 9436 12974 9492
rect 9518 9380 9528 9436
rect 9584 9380 9632 9436
rect 9688 9380 9736 9436
rect 9792 9380 9802 9436
rect 17834 9380 17844 9436
rect 17900 9380 17948 9436
rect 18004 9380 18052 9436
rect 18108 9380 18118 9436
rect 26150 9380 26160 9436
rect 26216 9380 26264 9436
rect 26320 9380 26368 9436
rect 26424 9380 26434 9436
rect 34466 9380 34476 9436
rect 34532 9380 34580 9436
rect 34636 9380 34684 9436
rect 34740 9380 34750 9436
rect 6860 9324 7532 9380
rect 7588 9324 7598 9380
rect 10210 9324 10220 9380
rect 10276 9324 12572 9380
rect 12628 9324 12638 9380
rect 5058 9212 5068 9268
rect 5124 9212 5740 9268
rect 5796 9212 11228 9268
rect 11284 9212 11294 9268
rect 11666 9212 11676 9268
rect 11732 9212 12684 9268
rect 12740 9212 13468 9268
rect 13524 9212 13534 9268
rect 17266 9212 17276 9268
rect 17332 9212 18172 9268
rect 18228 9212 18238 9268
rect 28354 9212 28364 9268
rect 28420 9212 29260 9268
rect 29316 9212 30492 9268
rect 30548 9212 30558 9268
rect 3658 9100 3668 9156
rect 3724 9100 6188 9156
rect 6244 9100 6254 9156
rect 7074 9100 7084 9156
rect 7140 9100 10220 9156
rect 10276 9100 10286 9156
rect 11890 9100 11900 9156
rect 11956 9100 12180 9156
rect 12236 9100 12246 9156
rect 6514 8988 6524 9044
rect 6580 8988 7308 9044
rect 7364 8988 7374 9044
rect 8306 8988 8316 9044
rect 8372 8988 9548 9044
rect 9604 8988 9614 9044
rect 12338 8988 12348 9044
rect 12404 8988 13692 9044
rect 13748 8988 13758 9044
rect 14186 8988 14196 9044
rect 14252 8988 14588 9044
rect 14644 8988 15036 9044
rect 15092 8988 15102 9044
rect 21858 8988 21868 9044
rect 21924 8988 22764 9044
rect 22820 8988 22830 9044
rect 25106 8988 25116 9044
rect 25172 8988 25564 9044
rect 25620 8988 25630 9044
rect 28018 8988 28028 9044
rect 28084 8988 29148 9044
rect 29204 8988 30156 9044
rect 30212 8988 31892 9044
rect 31948 8988 31958 9044
rect 11778 8876 11788 8932
rect 11844 8876 15260 8932
rect 15316 8876 15326 8932
rect 22194 8876 22204 8932
rect 22260 8876 22652 8932
rect 22708 8876 22718 8932
rect 29362 8876 29372 8932
rect 29428 8876 30492 8932
rect 30548 8876 30558 8932
rect 4498 8764 4508 8820
rect 4564 8764 6636 8820
rect 6692 8764 6702 8820
rect 28242 8764 28252 8820
rect 28308 8764 28924 8820
rect 28980 8764 29932 8820
rect 29988 8764 29998 8820
rect 11778 8652 11788 8708
rect 11844 8652 12348 8708
rect 12404 8652 12414 8708
rect 5360 8596 5370 8652
rect 5426 8596 5474 8652
rect 5530 8596 5578 8652
rect 5634 8596 5644 8652
rect 13676 8596 13686 8652
rect 13742 8596 13790 8652
rect 13846 8596 13894 8652
rect 13950 8596 13960 8652
rect 21992 8596 22002 8652
rect 22058 8596 22106 8652
rect 22162 8596 22210 8652
rect 22266 8596 22276 8652
rect 30308 8596 30318 8652
rect 30374 8596 30422 8652
rect 30478 8596 30526 8652
rect 30582 8596 30592 8652
rect 6738 8540 6748 8596
rect 6804 8540 7084 8596
rect 7140 8540 7150 8596
rect 3042 8428 3052 8484
rect 3108 8428 4172 8484
rect 4228 8428 4238 8484
rect 6290 8428 6300 8484
rect 6356 8428 7532 8484
rect 7588 8428 7598 8484
rect 12002 8428 12012 8484
rect 12068 8428 12348 8484
rect 12404 8428 12414 8484
rect 19506 8428 19516 8484
rect 19572 8428 22428 8484
rect 22484 8428 22652 8484
rect 22708 8428 23604 8484
rect 23660 8428 26572 8484
rect 26628 8428 26638 8484
rect 3882 8316 3892 8372
rect 3948 8316 4732 8372
rect 4788 8316 15148 8372
rect 15204 8316 15214 8372
rect 22754 8316 22764 8372
rect 22820 8316 24444 8372
rect 24500 8316 24510 8372
rect 4246 8204 4284 8260
rect 4340 8204 6748 8260
rect 6804 8204 6814 8260
rect 7746 8204 7756 8260
rect 7812 8204 8652 8260
rect 8708 8204 8718 8260
rect 10098 8204 10108 8260
rect 10164 8204 11340 8260
rect 11396 8204 12236 8260
rect 12292 8204 12572 8260
rect 12628 8204 12638 8260
rect 15922 8204 15932 8260
rect 15988 8204 17052 8260
rect 17108 8204 17118 8260
rect 23090 8204 23100 8260
rect 23156 8204 25340 8260
rect 25396 8204 25406 8260
rect 27906 8204 27916 8260
rect 27972 8204 28140 8260
rect 28196 8204 29036 8260
rect 29092 8204 29102 8260
rect 2482 8092 2492 8148
rect 2548 8092 3052 8148
rect 3108 8092 4060 8148
rect 4116 8092 4126 8148
rect 7410 8092 7420 8148
rect 7476 8092 9772 8148
rect 9828 8092 9838 8148
rect 11778 8092 11788 8148
rect 11844 8092 12124 8148
rect 12180 8092 12190 8148
rect 8540 8036 8596 8092
rect 4946 7980 4956 8036
rect 5012 7980 8428 8036
rect 8530 7980 8540 8036
rect 8596 7980 8606 8036
rect 9324 7980 11116 8036
rect 11172 7980 11182 8036
rect 11554 7980 11564 8036
rect 11620 7980 13804 8036
rect 13860 7980 13870 8036
rect 22418 7980 22428 8036
rect 22484 7980 22876 8036
rect 22932 7980 23044 8036
rect 23100 7980 23110 8036
rect 8372 7924 8428 7980
rect 9324 7924 9380 7980
rect 5842 7868 5852 7924
rect 5908 7868 7868 7924
rect 7924 7868 7934 7924
rect 8372 7868 9380 7924
rect 11116 7924 11172 7980
rect 11116 7868 12012 7924
rect 12068 7868 14700 7924
rect 14756 7868 14766 7924
rect 14858 7868 14868 7924
rect 14924 7868 15596 7924
rect 15652 7868 15662 7924
rect 9518 7812 9528 7868
rect 9584 7812 9632 7868
rect 9688 7812 9736 7868
rect 9792 7812 9802 7868
rect 14700 7812 14756 7868
rect 17834 7812 17844 7868
rect 17900 7812 17948 7868
rect 18004 7812 18052 7868
rect 18108 7812 18118 7868
rect 23212 7812 23268 8204
rect 23426 8092 23436 8148
rect 23492 8092 25116 8148
rect 25172 8092 25182 8148
rect 26450 7980 26460 8036
rect 26516 7980 26908 8036
rect 27570 7980 27580 8036
rect 27636 7980 28252 8036
rect 28308 7980 28318 8036
rect 26150 7812 26160 7868
rect 26216 7812 26264 7868
rect 26320 7812 26368 7868
rect 26424 7812 26434 7868
rect 12338 7756 12348 7812
rect 12404 7756 13356 7812
rect 13412 7756 13422 7812
rect 14700 7756 15932 7812
rect 15988 7756 15998 7812
rect 22866 7756 22876 7812
rect 22932 7756 23268 7812
rect 12898 7644 12908 7700
rect 12964 7644 12974 7700
rect 12908 7588 12964 7644
rect 26852 7588 26908 7980
rect 34466 7812 34476 7868
rect 34532 7812 34580 7868
rect 34636 7812 34684 7868
rect 34740 7812 34750 7868
rect 12338 7532 12348 7588
rect 12404 7532 12964 7588
rect 22082 7532 22092 7588
rect 22148 7532 22540 7588
rect 22596 7532 22764 7588
rect 22820 7532 22830 7588
rect 26852 7532 29764 7588
rect 29820 7532 29830 7588
rect 2594 7420 2604 7476
rect 2660 7420 7644 7476
rect 7700 7420 7710 7476
rect 10546 7420 10556 7476
rect 10612 7420 11004 7476
rect 11060 7420 11070 7476
rect 12450 7420 12460 7476
rect 12516 7420 15764 7476
rect 15820 7420 16156 7476
rect 16212 7420 16222 7476
rect 23594 7420 23604 7476
rect 23660 7420 24108 7476
rect 24164 7420 24174 7476
rect 24322 7420 24332 7476
rect 24388 7420 25788 7476
rect 25844 7420 26908 7476
rect 26964 7420 26974 7476
rect 29474 7420 29484 7476
rect 29540 7420 31612 7476
rect 31668 7420 33628 7476
rect 33684 7420 34076 7476
rect 34132 7420 34142 7476
rect 9090 7308 9100 7364
rect 9156 7308 9996 7364
rect 10052 7308 10062 7364
rect 13020 7308 13580 7364
rect 13636 7308 13646 7364
rect 31826 7308 31836 7364
rect 31892 7308 32060 7364
rect 32116 7308 32126 7364
rect 7746 7196 7756 7252
rect 7812 7196 10948 7252
rect 10892 7140 10948 7196
rect 13020 7140 13076 7308
rect 13458 7196 13468 7252
rect 13524 7196 14028 7252
rect 14084 7196 14094 7252
rect 14578 7196 14588 7252
rect 14644 7196 15372 7252
rect 15428 7196 15438 7252
rect 7858 7084 7868 7140
rect 7924 7084 8988 7140
rect 9044 7084 9054 7140
rect 10892 7084 13076 7140
rect 23202 7084 23212 7140
rect 23268 7084 26908 7140
rect 5360 7028 5370 7084
rect 5426 7028 5474 7084
rect 5530 7028 5578 7084
rect 5634 7028 5644 7084
rect 8988 7028 9044 7084
rect 13676 7028 13686 7084
rect 13742 7028 13790 7084
rect 13846 7028 13894 7084
rect 13950 7028 13960 7084
rect 21992 7028 22002 7084
rect 22058 7028 22106 7084
rect 22162 7028 22210 7084
rect 22266 7028 22276 7084
rect 8988 6972 12460 7028
rect 12516 6972 12526 7028
rect 24434 6972 24444 7028
rect 24500 6972 24510 7028
rect 6738 6860 6748 6916
rect 6804 6860 6814 6916
rect 10380 6860 10390 6916
rect 10446 6860 11172 6916
rect 11228 6860 11676 6916
rect 11732 6860 11742 6916
rect 13850 6860 13860 6916
rect 13916 6860 14364 6916
rect 14420 6860 14430 6916
rect 6748 6804 6804 6860
rect 24444 6804 24500 6972
rect 2762 6748 2772 6804
rect 2828 6748 3948 6804
rect 4004 6748 4014 6804
rect 6748 6748 8092 6804
rect 8148 6748 10556 6804
rect 10612 6748 10622 6804
rect 14018 6748 14028 6804
rect 14084 6748 16268 6804
rect 16324 6748 16334 6804
rect 21410 6748 21420 6804
rect 21476 6748 21756 6804
rect 21812 6748 23212 6804
rect 23268 6748 23278 6804
rect 23986 6748 23996 6804
rect 24052 6748 24500 6804
rect 26852 6804 26908 7084
rect 29708 6804 29764 7140
rect 29820 7084 29830 7140
rect 29922 7084 29932 7140
rect 29988 7084 29998 7140
rect 26852 6748 28252 6804
rect 28308 6748 28318 6804
rect 29596 6748 29764 6804
rect 29596 6692 29652 6748
rect 3098 6636 3108 6692
rect 3164 6636 3388 6692
rect 3444 6636 3454 6692
rect 3612 6636 4228 6692
rect 4284 6636 5516 6692
rect 5572 6636 5582 6692
rect 13178 6636 13188 6692
rect 13244 6636 13580 6692
rect 13636 6636 13646 6692
rect 13794 6636 13804 6692
rect 13860 6636 14364 6692
rect 14420 6636 14430 6692
rect 15026 6636 15036 6692
rect 15092 6636 15372 6692
rect 15428 6636 15932 6692
rect 15988 6636 17388 6692
rect 17444 6636 17454 6692
rect 17994 6636 18004 6692
rect 18060 6636 19180 6692
rect 19236 6636 19246 6692
rect 29586 6636 29596 6692
rect 29652 6636 29662 6692
rect 3612 6580 3668 6636
rect 3490 6524 3500 6580
rect 3556 6524 3668 6580
rect 7074 6524 7084 6580
rect 7140 6524 8260 6580
rect 8316 6524 8326 6580
rect 10770 6524 10780 6580
rect 10836 6524 11564 6580
rect 11620 6524 11630 6580
rect 11890 6524 11900 6580
rect 11956 6524 15148 6580
rect 23874 6524 23884 6580
rect 23940 6524 28140 6580
rect 28196 6524 28206 6580
rect 15092 6468 15148 6524
rect 3098 6412 3108 6468
rect 3164 6412 3836 6468
rect 3892 6412 3902 6468
rect 4050 6412 4060 6468
rect 4116 6412 13524 6468
rect 14354 6412 14364 6468
rect 14420 6412 14868 6468
rect 14924 6412 14934 6468
rect 15092 6412 15484 6468
rect 15540 6412 16884 6468
rect 16940 6412 16950 6468
rect 3714 6300 3724 6356
rect 3780 6300 4732 6356
rect 4788 6300 8204 6356
rect 8260 6300 8270 6356
rect 12002 6300 12012 6356
rect 12068 6300 12236 6356
rect 12292 6300 12302 6356
rect 9518 6244 9528 6300
rect 9584 6244 9632 6300
rect 9688 6244 9736 6300
rect 9792 6244 9802 6300
rect 13468 6244 13524 6412
rect 29932 6356 29988 7084
rect 30308 7028 30318 7084
rect 30374 7028 30422 7084
rect 30478 7028 30526 7084
rect 30582 7028 30592 7084
rect 32162 6748 32172 6804
rect 32228 6748 33292 6804
rect 33348 6748 33358 6804
rect 29932 6300 30156 6356
rect 30212 6300 30222 6356
rect 17834 6244 17844 6300
rect 17900 6244 17948 6300
rect 18004 6244 18052 6300
rect 18108 6244 18118 6300
rect 26150 6244 26160 6300
rect 26216 6244 26264 6300
rect 26320 6244 26368 6300
rect 26424 6244 26434 6300
rect 34466 6244 34476 6300
rect 34532 6244 34580 6300
rect 34636 6244 34684 6300
rect 34740 6244 34750 6300
rect 3602 6188 3612 6244
rect 3668 6188 5852 6244
rect 5908 6188 5918 6244
rect 7858 6188 7868 6244
rect 7924 6188 8316 6244
rect 8372 6188 8382 6244
rect 10434 6188 10444 6244
rect 10500 6188 11732 6244
rect 11788 6188 11798 6244
rect 13458 6188 13468 6244
rect 13524 6188 13534 6244
rect 23202 6188 23212 6244
rect 23268 6188 23772 6244
rect 23828 6188 23838 6244
rect 27458 6188 27468 6244
rect 27524 6188 30604 6244
rect 30660 6188 30670 6244
rect 4834 6076 4844 6132
rect 4900 6076 4910 6132
rect 9314 6076 9324 6132
rect 9380 6076 9996 6132
rect 10052 6076 10668 6132
rect 10724 6076 10734 6132
rect 12002 6076 12012 6132
rect 12068 6076 12460 6132
rect 12516 6076 12526 6132
rect 16426 6076 16436 6132
rect 16492 6076 17276 6132
rect 17332 6076 17342 6132
rect 18386 6076 18396 6132
rect 18452 6076 19068 6132
rect 19124 6076 19516 6132
rect 19572 6076 19582 6132
rect 23426 6076 23436 6132
rect 23492 6076 24892 6132
rect 24948 6076 25284 6132
rect 25340 6076 25350 6132
rect 30370 6076 30380 6132
rect 30436 6076 32172 6132
rect 32228 6076 33124 6132
rect 33180 6076 33190 6132
rect 4844 6020 4900 6076
rect 2930 5964 2940 6020
rect 2996 5964 3612 6020
rect 3668 5964 3678 6020
rect 4162 5964 4172 6020
rect 4228 5964 4900 6020
rect 4956 5964 5236 6020
rect 5292 5964 7252 6020
rect 7308 5964 7318 6020
rect 10994 5964 11004 6020
rect 11060 5964 11564 6020
rect 11620 5964 14476 6020
rect 14532 5964 14868 6020
rect 14924 5964 14934 6020
rect 17042 5964 17052 6020
rect 17108 5964 18060 6020
rect 18116 5964 18126 6020
rect 18902 5964 18912 6020
rect 18968 5964 19908 6020
rect 19964 5964 19974 6020
rect 22642 5964 22652 6020
rect 22708 5964 23324 6020
rect 23380 5964 23390 6020
rect 28466 5964 28476 6020
rect 28532 5964 29596 6020
rect 29652 5964 30044 6020
rect 30100 5964 30110 6020
rect 2818 5852 2828 5908
rect 2884 5852 3388 5908
rect 3444 5852 3454 5908
rect 4498 5852 4508 5908
rect 4564 5852 4732 5908
rect 4788 5852 4798 5908
rect 4956 5796 5012 5964
rect 6402 5852 6412 5908
rect 6468 5852 10108 5908
rect 10164 5852 10174 5908
rect 11106 5852 11116 5908
rect 11172 5852 11676 5908
rect 11732 5852 12124 5908
rect 12180 5852 12190 5908
rect 16706 5852 16716 5908
rect 16772 5852 17164 5908
rect 17220 5852 17230 5908
rect 17826 5852 17836 5908
rect 17892 5852 18732 5908
rect 18788 5852 19628 5908
rect 19684 5852 19694 5908
rect 23436 5852 24220 5908
rect 24276 5852 24286 5908
rect 28130 5852 28140 5908
rect 28196 5852 28700 5908
rect 28756 5852 29484 5908
rect 29540 5852 29550 5908
rect 31938 5852 31948 5908
rect 32004 5852 33404 5908
rect 33460 5852 33470 5908
rect 23436 5796 23492 5852
rect 3938 5740 3948 5796
rect 4004 5740 5012 5796
rect 8054 5740 8092 5796
rect 8148 5740 8158 5796
rect 8372 5740 13804 5796
rect 13860 5740 13870 5796
rect 18162 5740 18172 5796
rect 18228 5740 18956 5796
rect 19012 5740 19022 5796
rect 21354 5740 21364 5796
rect 21420 5740 23212 5796
rect 23268 5740 23278 5796
rect 23426 5740 23436 5796
rect 23492 5740 23502 5796
rect 27244 5740 30380 5796
rect 30436 5740 31276 5796
rect 31332 5740 34076 5796
rect 34132 5740 34142 5796
rect 8372 5684 8428 5740
rect 2482 5628 2492 5684
rect 2548 5628 6246 5684
rect 6302 5628 8428 5684
rect 10210 5628 10220 5684
rect 10276 5628 11228 5684
rect 11284 5628 11294 5684
rect 22306 5628 22316 5684
rect 6850 5516 6860 5572
rect 6916 5516 8092 5572
rect 8148 5516 10332 5572
rect 10388 5516 10398 5572
rect 5360 5460 5370 5516
rect 5426 5460 5474 5516
rect 5530 5460 5578 5516
rect 5634 5460 5644 5516
rect 13676 5460 13686 5516
rect 13742 5460 13790 5516
rect 13846 5460 13894 5516
rect 13950 5460 13960 5516
rect 21992 5460 22002 5516
rect 22058 5460 22106 5516
rect 22162 5460 22210 5516
rect 22266 5460 22276 5516
rect 6738 5404 6748 5460
rect 6804 5404 11732 5460
rect 11788 5404 12236 5460
rect 12292 5404 12302 5460
rect 15092 5404 15260 5460
rect 15316 5404 15326 5460
rect 4946 5292 4956 5348
rect 5012 5292 6972 5348
rect 7028 5292 7038 5348
rect 8418 5292 8428 5348
rect 8484 5292 12012 5348
rect 12068 5292 12078 5348
rect 6796 5180 6806 5236
rect 6862 5180 9996 5236
rect 10052 5180 10062 5236
rect 10322 5180 10332 5236
rect 10388 5180 11732 5236
rect 13626 5180 13636 5236
rect 13692 5180 14588 5236
rect 14644 5180 14654 5236
rect 11676 5124 11732 5180
rect 15092 5124 15148 5404
rect 21522 5292 21532 5348
rect 21588 5292 22316 5348
rect 22372 5292 22428 5684
rect 23762 5628 23772 5684
rect 23828 5628 24556 5684
rect 24612 5628 24622 5684
rect 27244 5572 27300 5740
rect 29810 5628 29820 5684
rect 29876 5628 30268 5684
rect 30324 5628 30716 5684
rect 30772 5628 30996 5684
rect 31052 5628 31388 5684
rect 31444 5628 31454 5684
rect 27234 5516 27244 5572
rect 27300 5516 27310 5572
rect 30308 5460 30318 5516
rect 30374 5460 30422 5516
rect 30478 5460 30526 5516
rect 30582 5460 30592 5516
rect 26338 5292 26348 5348
rect 26404 5292 32396 5348
rect 32452 5292 32462 5348
rect 18050 5180 18060 5236
rect 18116 5180 19068 5236
rect 19124 5180 19628 5236
rect 19684 5180 19694 5236
rect 27794 5180 27804 5236
rect 27860 5180 28252 5236
rect 28308 5180 28318 5236
rect 30930 5180 30940 5236
rect 30996 5180 31948 5236
rect 32004 5180 32014 5236
rect 2930 5068 2940 5124
rect 2996 5068 3612 5124
rect 3668 5068 3678 5124
rect 4274 5068 4284 5124
rect 4340 5068 4732 5124
rect 4788 5068 4798 5124
rect 4946 5068 4956 5124
rect 5012 5068 6412 5124
rect 6468 5068 6478 5124
rect 7074 5068 7084 5124
rect 7140 5068 8428 5124
rect 8484 5068 8494 5124
rect 8764 5068 10444 5124
rect 10500 5068 10510 5124
rect 11676 5068 15148 5124
rect 16482 5068 16492 5124
rect 16548 5068 18508 5124
rect 18564 5068 19348 5124
rect 19404 5068 19414 5124
rect 22194 5068 22204 5124
rect 22260 5068 23660 5124
rect 23716 5068 23726 5124
rect 25666 5068 25676 5124
rect 25732 5068 26908 5124
rect 26964 5068 26974 5124
rect 27346 5068 27356 5124
rect 27412 5068 29484 5124
rect 29540 5068 29550 5124
rect 30370 5068 30380 5124
rect 30436 5068 31612 5124
rect 31668 5068 31678 5124
rect 8764 5012 8820 5068
rect 11676 5012 11732 5068
rect 8194 4956 8204 5012
rect 8260 4956 8820 5012
rect 11666 4956 11676 5012
rect 11732 4956 11742 5012
rect 10210 4844 10220 4900
rect 10276 4844 10986 4900
rect 11042 4844 11788 4900
rect 11844 4844 11854 4900
rect 30594 4844 30604 4900
rect 30660 4844 30940 4900
rect 30996 4844 31006 4900
rect 9518 4676 9528 4732
rect 9584 4676 9632 4732
rect 9688 4676 9736 4732
rect 9792 4676 9802 4732
rect 17834 4676 17844 4732
rect 17900 4676 17948 4732
rect 18004 4676 18052 4732
rect 18108 4676 18118 4732
rect 26150 4676 26160 4732
rect 26216 4676 26264 4732
rect 26320 4676 26368 4732
rect 26424 4676 26434 4732
rect 34466 4676 34476 4732
rect 34532 4676 34580 4732
rect 34636 4676 34684 4732
rect 34740 4676 34750 4732
rect 5598 4508 5608 4564
rect 5664 4508 18172 4564
rect 18228 4508 18238 4564
rect 26562 4508 26572 4564
rect 26628 4508 29764 4564
rect 29820 4508 29830 4564
rect 4274 4396 4284 4452
rect 4340 4396 4620 4452
rect 4676 4396 4686 4452
rect 8306 4396 8316 4452
rect 8372 4396 9716 4452
rect 9660 4340 9716 4396
rect 1586 4284 1596 4340
rect 1652 4284 5740 4340
rect 5796 4284 5806 4340
rect 9650 4284 9660 4340
rect 9716 4284 13020 4340
rect 13076 4284 14812 4340
rect 14868 4284 14878 4340
rect 16818 4284 16828 4340
rect 16884 4284 17836 4340
rect 17892 4284 17902 4340
rect 26338 4284 26348 4340
rect 26404 4284 28364 4340
rect 28420 4284 28430 4340
rect 3602 4172 3612 4228
rect 3668 4172 18284 4228
rect 18340 4172 18350 4228
rect 23314 4172 23324 4228
rect 23380 4172 24108 4228
rect 24164 4172 24174 4228
rect 26002 4172 26012 4228
rect 26068 4172 27244 4228
rect 27300 4172 27310 4228
rect 31490 4060 31500 4116
rect 31556 4060 32172 4116
rect 32228 4060 32238 4116
rect 5360 3892 5370 3948
rect 5426 3892 5474 3948
rect 5530 3892 5578 3948
rect 5634 3892 5644 3948
rect 13676 3892 13686 3948
rect 13742 3892 13790 3948
rect 13846 3892 13894 3948
rect 13950 3892 13960 3948
rect 21992 3892 22002 3948
rect 22058 3892 22106 3948
rect 22162 3892 22210 3948
rect 22266 3892 22276 3948
rect 30308 3892 30318 3948
rect 30374 3892 30422 3948
rect 30478 3892 30526 3948
rect 30582 3892 30592 3948
rect 31042 3836 31052 3892
rect 31108 3836 32844 3892
rect 32900 3836 32910 3892
rect 11218 3724 11228 3780
rect 11284 3724 14700 3780
rect 14756 3724 14766 3780
rect 31938 3724 31948 3780
rect 32004 3724 32564 3780
rect 32620 3724 32630 3780
rect 25106 3612 25116 3668
rect 25172 3612 26348 3668
rect 26404 3612 26414 3668
rect 4498 3500 4508 3556
rect 4564 3500 5852 3556
rect 5908 3500 5918 3556
rect 21410 3500 21420 3556
rect 21476 3500 21868 3556
rect 21924 3500 21934 3556
rect 28634 3500 28644 3556
rect 28700 3500 31052 3556
rect 31108 3500 32284 3556
rect 32340 3500 32350 3556
rect 4834 3388 4844 3444
rect 4900 3388 6132 3444
rect 6188 3388 11228 3444
rect 11284 3388 11294 3444
rect 9518 3108 9528 3164
rect 9584 3108 9632 3164
rect 9688 3108 9736 3164
rect 9792 3108 9802 3164
rect 17834 3108 17844 3164
rect 17900 3108 17948 3164
rect 18004 3108 18052 3164
rect 18108 3108 18118 3164
rect 26150 3108 26160 3164
rect 26216 3108 26264 3164
rect 26320 3108 26368 3164
rect 26424 3108 26434 3164
rect 34466 3108 34476 3164
rect 34532 3108 34580 3164
rect 34636 3108 34684 3164
rect 34740 3108 34750 3164
<< via3 >>
rect 5370 32116 5426 32172
rect 5474 32116 5530 32172
rect 5578 32116 5634 32172
rect 13686 32116 13742 32172
rect 13790 32116 13846 32172
rect 13894 32116 13950 32172
rect 22002 32116 22058 32172
rect 22106 32116 22162 32172
rect 22210 32116 22266 32172
rect 30318 32116 30374 32172
rect 30422 32116 30478 32172
rect 30526 32116 30582 32172
rect 9528 31332 9584 31388
rect 9632 31332 9688 31388
rect 9736 31332 9792 31388
rect 17844 31332 17900 31388
rect 17948 31332 18004 31388
rect 18052 31332 18108 31388
rect 26160 31332 26216 31388
rect 26264 31332 26320 31388
rect 26368 31332 26424 31388
rect 34476 31332 34532 31388
rect 34580 31332 34636 31388
rect 34684 31332 34740 31388
rect 5370 30548 5426 30604
rect 5474 30548 5530 30604
rect 5578 30548 5634 30604
rect 13686 30548 13742 30604
rect 13790 30548 13846 30604
rect 13894 30548 13950 30604
rect 22002 30548 22058 30604
rect 22106 30548 22162 30604
rect 22210 30548 22266 30604
rect 30318 30548 30374 30604
rect 30422 30548 30478 30604
rect 30526 30548 30582 30604
rect 9528 29764 9584 29820
rect 9632 29764 9688 29820
rect 9736 29764 9792 29820
rect 17844 29764 17900 29820
rect 17948 29764 18004 29820
rect 18052 29764 18108 29820
rect 26160 29764 26216 29820
rect 26264 29764 26320 29820
rect 26368 29764 26424 29820
rect 34476 29764 34532 29820
rect 34580 29764 34636 29820
rect 34684 29764 34740 29820
rect 5370 28980 5426 29036
rect 5474 28980 5530 29036
rect 5578 28980 5634 29036
rect 13686 28980 13742 29036
rect 13790 28980 13846 29036
rect 13894 28980 13950 29036
rect 22002 28980 22058 29036
rect 22106 28980 22162 29036
rect 22210 28980 22266 29036
rect 30318 28980 30374 29036
rect 30422 28980 30478 29036
rect 30526 28980 30582 29036
rect 9528 28196 9584 28252
rect 9632 28196 9688 28252
rect 9736 28196 9792 28252
rect 17844 28196 17900 28252
rect 17948 28196 18004 28252
rect 18052 28196 18108 28252
rect 26160 28196 26216 28252
rect 26264 28196 26320 28252
rect 26368 28196 26424 28252
rect 34476 28196 34532 28252
rect 34580 28196 34636 28252
rect 34684 28196 34740 28252
rect 5370 27412 5426 27468
rect 5474 27412 5530 27468
rect 5578 27412 5634 27468
rect 13686 27412 13742 27468
rect 13790 27412 13846 27468
rect 13894 27412 13950 27468
rect 22002 27412 22058 27468
rect 22106 27412 22162 27468
rect 22210 27412 22266 27468
rect 30318 27412 30374 27468
rect 30422 27412 30478 27468
rect 30526 27412 30582 27468
rect 9528 26628 9584 26684
rect 9632 26628 9688 26684
rect 9736 26628 9792 26684
rect 17844 26628 17900 26684
rect 17948 26628 18004 26684
rect 18052 26628 18108 26684
rect 26160 26628 26216 26684
rect 26264 26628 26320 26684
rect 26368 26628 26424 26684
rect 34476 26628 34532 26684
rect 34580 26628 34636 26684
rect 34684 26628 34740 26684
rect 5370 25844 5426 25900
rect 5474 25844 5530 25900
rect 5578 25844 5634 25900
rect 13686 25844 13742 25900
rect 13790 25844 13846 25900
rect 13894 25844 13950 25900
rect 22002 25844 22058 25900
rect 22106 25844 22162 25900
rect 22210 25844 22266 25900
rect 30318 25844 30374 25900
rect 30422 25844 30478 25900
rect 30526 25844 30582 25900
rect 7980 25228 8036 25284
rect 9528 25060 9584 25116
rect 9632 25060 9688 25116
rect 9736 25060 9792 25116
rect 17844 25060 17900 25116
rect 17948 25060 18004 25116
rect 18052 25060 18108 25116
rect 26160 25060 26216 25116
rect 26264 25060 26320 25116
rect 26368 25060 26424 25116
rect 34476 25060 34532 25116
rect 34580 25060 34636 25116
rect 34684 25060 34740 25116
rect 7980 24668 8036 24724
rect 5370 24276 5426 24332
rect 5474 24276 5530 24332
rect 5578 24276 5634 24332
rect 13686 24276 13742 24332
rect 13790 24276 13846 24332
rect 13894 24276 13950 24332
rect 22002 24276 22058 24332
rect 22106 24276 22162 24332
rect 22210 24276 22266 24332
rect 30318 24276 30374 24332
rect 30422 24276 30478 24332
rect 30526 24276 30582 24332
rect 9528 23492 9584 23548
rect 9632 23492 9688 23548
rect 9736 23492 9792 23548
rect 17844 23492 17900 23548
rect 17948 23492 18004 23548
rect 18052 23492 18108 23548
rect 26160 23492 26216 23548
rect 26264 23492 26320 23548
rect 26368 23492 26424 23548
rect 34476 23492 34532 23548
rect 34580 23492 34636 23548
rect 34684 23492 34740 23548
rect 14140 22876 14196 22932
rect 5370 22708 5426 22764
rect 5474 22708 5530 22764
rect 5578 22708 5634 22764
rect 13686 22708 13742 22764
rect 13790 22708 13846 22764
rect 13894 22708 13950 22764
rect 22002 22708 22058 22764
rect 22106 22708 22162 22764
rect 22210 22708 22266 22764
rect 30318 22708 30374 22764
rect 30422 22708 30478 22764
rect 30526 22708 30582 22764
rect 14252 22316 14308 22372
rect 9528 21924 9584 21980
rect 9632 21924 9688 21980
rect 9736 21924 9792 21980
rect 17844 21924 17900 21980
rect 17948 21924 18004 21980
rect 18052 21924 18108 21980
rect 26160 21924 26216 21980
rect 26264 21924 26320 21980
rect 26368 21924 26424 21980
rect 34476 21924 34532 21980
rect 34580 21924 34636 21980
rect 34684 21924 34740 21980
rect 16604 21868 16660 21924
rect 5370 21140 5426 21196
rect 5474 21140 5530 21196
rect 5578 21140 5634 21196
rect 13686 21140 13742 21196
rect 13790 21140 13846 21196
rect 13894 21140 13950 21196
rect 22002 21140 22058 21196
rect 22106 21140 22162 21196
rect 22210 21140 22266 21196
rect 30318 21140 30374 21196
rect 30422 21140 30478 21196
rect 30526 21140 30582 21196
rect 9528 20356 9584 20412
rect 9632 20356 9688 20412
rect 9736 20356 9792 20412
rect 17844 20356 17900 20412
rect 17948 20356 18004 20412
rect 18052 20356 18108 20412
rect 26160 20356 26216 20412
rect 26264 20356 26320 20412
rect 26368 20356 26424 20412
rect 34476 20356 34532 20412
rect 34580 20356 34636 20412
rect 34684 20356 34740 20412
rect 23548 20188 23604 20244
rect 5370 19572 5426 19628
rect 5474 19572 5530 19628
rect 5578 19572 5634 19628
rect 13686 19572 13742 19628
rect 13790 19572 13846 19628
rect 13894 19572 13950 19628
rect 22002 19572 22058 19628
rect 22106 19572 22162 19628
rect 22210 19572 22266 19628
rect 30318 19572 30374 19628
rect 30422 19572 30478 19628
rect 30526 19572 30582 19628
rect 14140 19516 14196 19572
rect 15596 19404 15652 19460
rect 9528 18788 9584 18844
rect 9632 18788 9688 18844
rect 9736 18788 9792 18844
rect 17844 18788 17900 18844
rect 17948 18788 18004 18844
rect 18052 18788 18108 18844
rect 26160 18788 26216 18844
rect 26264 18788 26320 18844
rect 26368 18788 26424 18844
rect 34476 18788 34532 18844
rect 34580 18788 34636 18844
rect 34684 18788 34740 18844
rect 16604 18732 16660 18788
rect 5370 18004 5426 18060
rect 5474 18004 5530 18060
rect 5578 18004 5634 18060
rect 13686 18004 13742 18060
rect 13790 18004 13846 18060
rect 13894 18004 13950 18060
rect 22002 18004 22058 18060
rect 22106 18004 22162 18060
rect 22210 18004 22266 18060
rect 30318 18004 30374 18060
rect 30422 18004 30478 18060
rect 30526 18004 30582 18060
rect 15596 17948 15652 18004
rect 18732 17948 18788 18004
rect 14252 17724 14308 17780
rect 18732 17724 18788 17780
rect 23548 17612 23604 17668
rect 9528 17220 9584 17276
rect 9632 17220 9688 17276
rect 9736 17220 9792 17276
rect 17844 17220 17900 17276
rect 17948 17220 18004 17276
rect 18052 17220 18108 17276
rect 26160 17220 26216 17276
rect 26264 17220 26320 17276
rect 26368 17220 26424 17276
rect 34476 17220 34532 17276
rect 34580 17220 34636 17276
rect 34684 17220 34740 17276
rect 5370 16436 5426 16492
rect 5474 16436 5530 16492
rect 5578 16436 5634 16492
rect 13686 16436 13742 16492
rect 13790 16436 13846 16492
rect 13894 16436 13950 16492
rect 22002 16436 22058 16492
rect 22106 16436 22162 16492
rect 22210 16436 22266 16492
rect 30318 16436 30374 16492
rect 30422 16436 30478 16492
rect 30526 16436 30582 16492
rect 9528 15652 9584 15708
rect 9632 15652 9688 15708
rect 9736 15652 9792 15708
rect 17844 15652 17900 15708
rect 17948 15652 18004 15708
rect 18052 15652 18108 15708
rect 26160 15652 26216 15708
rect 26264 15652 26320 15708
rect 26368 15652 26424 15708
rect 34476 15652 34532 15708
rect 34580 15652 34636 15708
rect 34684 15652 34740 15708
rect 5370 14868 5426 14924
rect 5474 14868 5530 14924
rect 5578 14868 5634 14924
rect 13686 14868 13742 14924
rect 13790 14868 13846 14924
rect 13894 14868 13950 14924
rect 22002 14868 22058 14924
rect 22106 14868 22162 14924
rect 22210 14868 22266 14924
rect 30318 14868 30374 14924
rect 30422 14868 30478 14924
rect 30526 14868 30582 14924
rect 3388 14476 3444 14532
rect 9528 14084 9584 14140
rect 9632 14084 9688 14140
rect 9736 14084 9792 14140
rect 17844 14084 17900 14140
rect 17948 14084 18004 14140
rect 18052 14084 18108 14140
rect 26160 14084 26216 14140
rect 26264 14084 26320 14140
rect 26368 14084 26424 14140
rect 34476 14084 34532 14140
rect 34580 14084 34636 14140
rect 34684 14084 34740 14140
rect 16380 13692 16436 13748
rect 18844 13692 18900 13748
rect 18620 13580 18676 13636
rect 5370 13300 5426 13356
rect 5474 13300 5530 13356
rect 5578 13300 5634 13356
rect 13686 13300 13742 13356
rect 13790 13300 13846 13356
rect 13894 13300 13950 13356
rect 22002 13300 22058 13356
rect 22106 13300 22162 13356
rect 22210 13300 22266 13356
rect 30318 13300 30374 13356
rect 30422 13300 30478 13356
rect 30526 13300 30582 13356
rect 16380 12684 16436 12740
rect 18844 12684 18900 12740
rect 9528 12516 9584 12572
rect 9632 12516 9688 12572
rect 9736 12516 9792 12572
rect 17844 12516 17900 12572
rect 17948 12516 18004 12572
rect 18052 12516 18108 12572
rect 26160 12516 26216 12572
rect 26264 12516 26320 12572
rect 26368 12516 26424 12572
rect 34476 12516 34532 12572
rect 34580 12516 34636 12572
rect 34684 12516 34740 12572
rect 8428 12124 8484 12180
rect 18620 12012 18676 12068
rect 5370 11732 5426 11788
rect 5474 11732 5530 11788
rect 5578 11732 5634 11788
rect 13686 11732 13742 11788
rect 13790 11732 13846 11788
rect 13894 11732 13950 11788
rect 22002 11732 22058 11788
rect 22106 11732 22162 11788
rect 22210 11732 22266 11788
rect 30318 11732 30374 11788
rect 30422 11732 30478 11788
rect 30526 11732 30582 11788
rect 9528 10948 9584 11004
rect 9632 10948 9688 11004
rect 9736 10948 9792 11004
rect 17844 10948 17900 11004
rect 17948 10948 18004 11004
rect 18052 10948 18108 11004
rect 26160 10948 26216 11004
rect 26264 10948 26320 11004
rect 26368 10948 26424 11004
rect 34476 10948 34532 11004
rect 34580 10948 34636 11004
rect 34684 10948 34740 11004
rect 8428 10780 8484 10836
rect 5370 10164 5426 10220
rect 5474 10164 5530 10220
rect 5578 10164 5634 10220
rect 13686 10164 13742 10220
rect 13790 10164 13846 10220
rect 13894 10164 13950 10220
rect 22002 10164 22058 10220
rect 22106 10164 22162 10220
rect 22210 10164 22266 10220
rect 30318 10164 30374 10220
rect 30422 10164 30478 10220
rect 30526 10164 30582 10220
rect 4284 10108 4340 10164
rect 4508 10108 4564 10164
rect 9528 9380 9584 9436
rect 9632 9380 9688 9436
rect 9736 9380 9792 9436
rect 17844 9380 17900 9436
rect 17948 9380 18004 9436
rect 18052 9380 18108 9436
rect 26160 9380 26216 9436
rect 26264 9380 26320 9436
rect 26368 9380 26424 9436
rect 34476 9380 34532 9436
rect 34580 9380 34636 9436
rect 34684 9380 34740 9436
rect 5370 8596 5426 8652
rect 5474 8596 5530 8652
rect 5578 8596 5634 8652
rect 13686 8596 13742 8652
rect 13790 8596 13846 8652
rect 13894 8596 13950 8652
rect 22002 8596 22058 8652
rect 22106 8596 22162 8652
rect 22210 8596 22266 8652
rect 30318 8596 30374 8652
rect 30422 8596 30478 8652
rect 30526 8596 30582 8652
rect 4284 8204 4340 8260
rect 9528 7812 9584 7868
rect 9632 7812 9688 7868
rect 9736 7812 9792 7868
rect 17844 7812 17900 7868
rect 17948 7812 18004 7868
rect 18052 7812 18108 7868
rect 26160 7812 26216 7868
rect 26264 7812 26320 7868
rect 26368 7812 26424 7868
rect 34476 7812 34532 7868
rect 34580 7812 34636 7868
rect 34684 7812 34740 7868
rect 5370 7028 5426 7084
rect 5474 7028 5530 7084
rect 5578 7028 5634 7084
rect 13686 7028 13742 7084
rect 13790 7028 13846 7084
rect 13894 7028 13950 7084
rect 22002 7028 22058 7084
rect 22106 7028 22162 7084
rect 22210 7028 22266 7084
rect 8092 6748 8148 6804
rect 3388 6636 3444 6692
rect 9528 6244 9584 6300
rect 9632 6244 9688 6300
rect 9736 6244 9792 6300
rect 30318 7028 30374 7084
rect 30422 7028 30478 7084
rect 30526 7028 30582 7084
rect 17844 6244 17900 6300
rect 17948 6244 18004 6300
rect 18052 6244 18108 6300
rect 26160 6244 26216 6300
rect 26264 6244 26320 6300
rect 26368 6244 26424 6300
rect 34476 6244 34532 6300
rect 34580 6244 34636 6300
rect 34684 6244 34740 6300
rect 4508 5852 4564 5908
rect 8092 5740 8148 5796
rect 5370 5460 5426 5516
rect 5474 5460 5530 5516
rect 5578 5460 5634 5516
rect 13686 5460 13742 5516
rect 13790 5460 13846 5516
rect 13894 5460 13950 5516
rect 22002 5460 22058 5516
rect 22106 5460 22162 5516
rect 22210 5460 22266 5516
rect 30318 5460 30374 5516
rect 30422 5460 30478 5516
rect 30526 5460 30582 5516
rect 9528 4676 9584 4732
rect 9632 4676 9688 4732
rect 9736 4676 9792 4732
rect 17844 4676 17900 4732
rect 17948 4676 18004 4732
rect 18052 4676 18108 4732
rect 26160 4676 26216 4732
rect 26264 4676 26320 4732
rect 26368 4676 26424 4732
rect 34476 4676 34532 4732
rect 34580 4676 34636 4732
rect 34684 4676 34740 4732
rect 5370 3892 5426 3948
rect 5474 3892 5530 3948
rect 5578 3892 5634 3948
rect 13686 3892 13742 3948
rect 13790 3892 13846 3948
rect 13894 3892 13950 3948
rect 22002 3892 22058 3948
rect 22106 3892 22162 3948
rect 22210 3892 22266 3948
rect 30318 3892 30374 3948
rect 30422 3892 30478 3948
rect 30526 3892 30582 3948
rect 9528 3108 9584 3164
rect 9632 3108 9688 3164
rect 9736 3108 9792 3164
rect 17844 3108 17900 3164
rect 17948 3108 18004 3164
rect 18052 3108 18108 3164
rect 26160 3108 26216 3164
rect 26264 3108 26320 3164
rect 26368 3108 26424 3164
rect 34476 3108 34532 3164
rect 34580 3108 34636 3164
rect 34684 3108 34740 3164
<< metal4 >>
rect 5342 32172 5662 32204
rect 5342 32116 5370 32172
rect 5426 32116 5474 32172
rect 5530 32116 5578 32172
rect 5634 32116 5662 32172
rect 5342 30604 5662 32116
rect 5342 30548 5370 30604
rect 5426 30548 5474 30604
rect 5530 30548 5578 30604
rect 5634 30548 5662 30604
rect 5342 29036 5662 30548
rect 5342 28980 5370 29036
rect 5426 28980 5474 29036
rect 5530 28980 5578 29036
rect 5634 28980 5662 29036
rect 5342 27468 5662 28980
rect 5342 27412 5370 27468
rect 5426 27412 5474 27468
rect 5530 27412 5578 27468
rect 5634 27412 5662 27468
rect 5342 25900 5662 27412
rect 5342 25844 5370 25900
rect 5426 25844 5474 25900
rect 5530 25844 5578 25900
rect 5634 25844 5662 25900
rect 5342 24332 5662 25844
rect 9500 31388 9820 32204
rect 9500 31332 9528 31388
rect 9584 31332 9632 31388
rect 9688 31332 9736 31388
rect 9792 31332 9820 31388
rect 9500 29820 9820 31332
rect 9500 29764 9528 29820
rect 9584 29764 9632 29820
rect 9688 29764 9736 29820
rect 9792 29764 9820 29820
rect 9500 28252 9820 29764
rect 9500 28196 9528 28252
rect 9584 28196 9632 28252
rect 9688 28196 9736 28252
rect 9792 28196 9820 28252
rect 9500 26684 9820 28196
rect 9500 26628 9528 26684
rect 9584 26628 9632 26684
rect 9688 26628 9736 26684
rect 9792 26628 9820 26684
rect 7980 25284 8036 25294
rect 7980 24724 8036 25228
rect 7980 24658 8036 24668
rect 9500 25116 9820 26628
rect 9500 25060 9528 25116
rect 9584 25060 9632 25116
rect 9688 25060 9736 25116
rect 9792 25060 9820 25116
rect 5342 24276 5370 24332
rect 5426 24276 5474 24332
rect 5530 24276 5578 24332
rect 5634 24276 5662 24332
rect 5342 22764 5662 24276
rect 5342 22708 5370 22764
rect 5426 22708 5474 22764
rect 5530 22708 5578 22764
rect 5634 22708 5662 22764
rect 5342 21196 5662 22708
rect 5342 21140 5370 21196
rect 5426 21140 5474 21196
rect 5530 21140 5578 21196
rect 5634 21140 5662 21196
rect 5342 19628 5662 21140
rect 5342 19572 5370 19628
rect 5426 19572 5474 19628
rect 5530 19572 5578 19628
rect 5634 19572 5662 19628
rect 5342 18060 5662 19572
rect 5342 18004 5370 18060
rect 5426 18004 5474 18060
rect 5530 18004 5578 18060
rect 5634 18004 5662 18060
rect 5342 16492 5662 18004
rect 5342 16436 5370 16492
rect 5426 16436 5474 16492
rect 5530 16436 5578 16492
rect 5634 16436 5662 16492
rect 5342 14924 5662 16436
rect 5342 14868 5370 14924
rect 5426 14868 5474 14924
rect 5530 14868 5578 14924
rect 5634 14868 5662 14924
rect 3388 14532 3444 14542
rect 3388 6692 3444 14476
rect 5342 13356 5662 14868
rect 5342 13300 5370 13356
rect 5426 13300 5474 13356
rect 5530 13300 5578 13356
rect 5634 13300 5662 13356
rect 5342 11788 5662 13300
rect 9500 23548 9820 25060
rect 9500 23492 9528 23548
rect 9584 23492 9632 23548
rect 9688 23492 9736 23548
rect 9792 23492 9820 23548
rect 9500 21980 9820 23492
rect 9500 21924 9528 21980
rect 9584 21924 9632 21980
rect 9688 21924 9736 21980
rect 9792 21924 9820 21980
rect 9500 20412 9820 21924
rect 9500 20356 9528 20412
rect 9584 20356 9632 20412
rect 9688 20356 9736 20412
rect 9792 20356 9820 20412
rect 9500 18844 9820 20356
rect 9500 18788 9528 18844
rect 9584 18788 9632 18844
rect 9688 18788 9736 18844
rect 9792 18788 9820 18844
rect 9500 17276 9820 18788
rect 9500 17220 9528 17276
rect 9584 17220 9632 17276
rect 9688 17220 9736 17276
rect 9792 17220 9820 17276
rect 9500 15708 9820 17220
rect 9500 15652 9528 15708
rect 9584 15652 9632 15708
rect 9688 15652 9736 15708
rect 9792 15652 9820 15708
rect 9500 14140 9820 15652
rect 9500 14084 9528 14140
rect 9584 14084 9632 14140
rect 9688 14084 9736 14140
rect 9792 14084 9820 14140
rect 9500 12572 9820 14084
rect 9500 12516 9528 12572
rect 9584 12516 9632 12572
rect 9688 12516 9736 12572
rect 9792 12516 9820 12572
rect 5342 11732 5370 11788
rect 5426 11732 5474 11788
rect 5530 11732 5578 11788
rect 5634 11732 5662 11788
rect 5342 10220 5662 11732
rect 8428 12180 8484 12190
rect 8428 10836 8484 12124
rect 8428 10770 8484 10780
rect 9500 11004 9820 12516
rect 9500 10948 9528 11004
rect 9584 10948 9632 11004
rect 9688 10948 9736 11004
rect 9792 10948 9820 11004
rect 4284 10164 4340 10174
rect 4284 8260 4340 10108
rect 4284 8194 4340 8204
rect 4508 10164 4564 10174
rect 3388 6626 3444 6636
rect 4508 5908 4564 10108
rect 4508 5842 4564 5852
rect 5342 10164 5370 10220
rect 5426 10164 5474 10220
rect 5530 10164 5578 10220
rect 5634 10164 5662 10220
rect 5342 8652 5662 10164
rect 5342 8596 5370 8652
rect 5426 8596 5474 8652
rect 5530 8596 5578 8652
rect 5634 8596 5662 8652
rect 5342 7084 5662 8596
rect 5342 7028 5370 7084
rect 5426 7028 5474 7084
rect 5530 7028 5578 7084
rect 5634 7028 5662 7084
rect 5342 5516 5662 7028
rect 9500 9436 9820 10948
rect 9500 9380 9528 9436
rect 9584 9380 9632 9436
rect 9688 9380 9736 9436
rect 9792 9380 9820 9436
rect 9500 7868 9820 9380
rect 9500 7812 9528 7868
rect 9584 7812 9632 7868
rect 9688 7812 9736 7868
rect 9792 7812 9820 7868
rect 8092 6804 8148 6814
rect 8092 5796 8148 6748
rect 8092 5730 8148 5740
rect 9500 6300 9820 7812
rect 9500 6244 9528 6300
rect 9584 6244 9632 6300
rect 9688 6244 9736 6300
rect 9792 6244 9820 6300
rect 5342 5460 5370 5516
rect 5426 5460 5474 5516
rect 5530 5460 5578 5516
rect 5634 5460 5662 5516
rect 5342 3948 5662 5460
rect 5342 3892 5370 3948
rect 5426 3892 5474 3948
rect 5530 3892 5578 3948
rect 5634 3892 5662 3948
rect 5342 3076 5662 3892
rect 9500 4732 9820 6244
rect 9500 4676 9528 4732
rect 9584 4676 9632 4732
rect 9688 4676 9736 4732
rect 9792 4676 9820 4732
rect 9500 3164 9820 4676
rect 9500 3108 9528 3164
rect 9584 3108 9632 3164
rect 9688 3108 9736 3164
rect 9792 3108 9820 3164
rect 9500 3076 9820 3108
rect 13658 32172 13978 32204
rect 13658 32116 13686 32172
rect 13742 32116 13790 32172
rect 13846 32116 13894 32172
rect 13950 32116 13978 32172
rect 13658 30604 13978 32116
rect 13658 30548 13686 30604
rect 13742 30548 13790 30604
rect 13846 30548 13894 30604
rect 13950 30548 13978 30604
rect 13658 29036 13978 30548
rect 13658 28980 13686 29036
rect 13742 28980 13790 29036
rect 13846 28980 13894 29036
rect 13950 28980 13978 29036
rect 13658 27468 13978 28980
rect 13658 27412 13686 27468
rect 13742 27412 13790 27468
rect 13846 27412 13894 27468
rect 13950 27412 13978 27468
rect 13658 25900 13978 27412
rect 13658 25844 13686 25900
rect 13742 25844 13790 25900
rect 13846 25844 13894 25900
rect 13950 25844 13978 25900
rect 13658 24332 13978 25844
rect 13658 24276 13686 24332
rect 13742 24276 13790 24332
rect 13846 24276 13894 24332
rect 13950 24276 13978 24332
rect 13658 22764 13978 24276
rect 17816 31388 18136 32204
rect 17816 31332 17844 31388
rect 17900 31332 17948 31388
rect 18004 31332 18052 31388
rect 18108 31332 18136 31388
rect 17816 29820 18136 31332
rect 17816 29764 17844 29820
rect 17900 29764 17948 29820
rect 18004 29764 18052 29820
rect 18108 29764 18136 29820
rect 17816 28252 18136 29764
rect 17816 28196 17844 28252
rect 17900 28196 17948 28252
rect 18004 28196 18052 28252
rect 18108 28196 18136 28252
rect 17816 26684 18136 28196
rect 17816 26628 17844 26684
rect 17900 26628 17948 26684
rect 18004 26628 18052 26684
rect 18108 26628 18136 26684
rect 17816 25116 18136 26628
rect 17816 25060 17844 25116
rect 17900 25060 17948 25116
rect 18004 25060 18052 25116
rect 18108 25060 18136 25116
rect 17816 23548 18136 25060
rect 17816 23492 17844 23548
rect 17900 23492 17948 23548
rect 18004 23492 18052 23548
rect 18108 23492 18136 23548
rect 13658 22708 13686 22764
rect 13742 22708 13790 22764
rect 13846 22708 13894 22764
rect 13950 22708 13978 22764
rect 13658 21196 13978 22708
rect 13658 21140 13686 21196
rect 13742 21140 13790 21196
rect 13846 21140 13894 21196
rect 13950 21140 13978 21196
rect 13658 19628 13978 21140
rect 13658 19572 13686 19628
rect 13742 19572 13790 19628
rect 13846 19572 13894 19628
rect 13950 19572 13978 19628
rect 13658 18060 13978 19572
rect 14140 22932 14196 22942
rect 14140 19572 14196 22876
rect 14140 19506 14196 19516
rect 14252 22372 14308 22382
rect 13658 18004 13686 18060
rect 13742 18004 13790 18060
rect 13846 18004 13894 18060
rect 13950 18004 13978 18060
rect 13658 16492 13978 18004
rect 14252 17780 14308 22316
rect 17816 21980 18136 23492
rect 16604 21924 16660 21934
rect 15596 19460 15652 19470
rect 15596 18004 15652 19404
rect 16604 18788 16660 21868
rect 16604 18722 16660 18732
rect 17816 21924 17844 21980
rect 17900 21924 17948 21980
rect 18004 21924 18052 21980
rect 18108 21924 18136 21980
rect 17816 20412 18136 21924
rect 17816 20356 17844 20412
rect 17900 20356 17948 20412
rect 18004 20356 18052 20412
rect 18108 20356 18136 20412
rect 17816 18844 18136 20356
rect 17816 18788 17844 18844
rect 17900 18788 17948 18844
rect 18004 18788 18052 18844
rect 18108 18788 18136 18844
rect 15596 17938 15652 17948
rect 14252 17714 14308 17724
rect 13658 16436 13686 16492
rect 13742 16436 13790 16492
rect 13846 16436 13894 16492
rect 13950 16436 13978 16492
rect 13658 14924 13978 16436
rect 13658 14868 13686 14924
rect 13742 14868 13790 14924
rect 13846 14868 13894 14924
rect 13950 14868 13978 14924
rect 13658 13356 13978 14868
rect 17816 17276 18136 18788
rect 21974 32172 22294 32204
rect 21974 32116 22002 32172
rect 22058 32116 22106 32172
rect 22162 32116 22210 32172
rect 22266 32116 22294 32172
rect 21974 30604 22294 32116
rect 21974 30548 22002 30604
rect 22058 30548 22106 30604
rect 22162 30548 22210 30604
rect 22266 30548 22294 30604
rect 21974 29036 22294 30548
rect 21974 28980 22002 29036
rect 22058 28980 22106 29036
rect 22162 28980 22210 29036
rect 22266 28980 22294 29036
rect 21974 27468 22294 28980
rect 21974 27412 22002 27468
rect 22058 27412 22106 27468
rect 22162 27412 22210 27468
rect 22266 27412 22294 27468
rect 21974 25900 22294 27412
rect 21974 25844 22002 25900
rect 22058 25844 22106 25900
rect 22162 25844 22210 25900
rect 22266 25844 22294 25900
rect 21974 24332 22294 25844
rect 21974 24276 22002 24332
rect 22058 24276 22106 24332
rect 22162 24276 22210 24332
rect 22266 24276 22294 24332
rect 21974 22764 22294 24276
rect 21974 22708 22002 22764
rect 22058 22708 22106 22764
rect 22162 22708 22210 22764
rect 22266 22708 22294 22764
rect 21974 21196 22294 22708
rect 21974 21140 22002 21196
rect 22058 21140 22106 21196
rect 22162 21140 22210 21196
rect 22266 21140 22294 21196
rect 21974 19628 22294 21140
rect 26132 31388 26452 32204
rect 26132 31332 26160 31388
rect 26216 31332 26264 31388
rect 26320 31332 26368 31388
rect 26424 31332 26452 31388
rect 26132 29820 26452 31332
rect 26132 29764 26160 29820
rect 26216 29764 26264 29820
rect 26320 29764 26368 29820
rect 26424 29764 26452 29820
rect 26132 28252 26452 29764
rect 26132 28196 26160 28252
rect 26216 28196 26264 28252
rect 26320 28196 26368 28252
rect 26424 28196 26452 28252
rect 26132 26684 26452 28196
rect 26132 26628 26160 26684
rect 26216 26628 26264 26684
rect 26320 26628 26368 26684
rect 26424 26628 26452 26684
rect 26132 25116 26452 26628
rect 26132 25060 26160 25116
rect 26216 25060 26264 25116
rect 26320 25060 26368 25116
rect 26424 25060 26452 25116
rect 26132 23548 26452 25060
rect 26132 23492 26160 23548
rect 26216 23492 26264 23548
rect 26320 23492 26368 23548
rect 26424 23492 26452 23548
rect 26132 21980 26452 23492
rect 26132 21924 26160 21980
rect 26216 21924 26264 21980
rect 26320 21924 26368 21980
rect 26424 21924 26452 21980
rect 26132 20412 26452 21924
rect 26132 20356 26160 20412
rect 26216 20356 26264 20412
rect 26320 20356 26368 20412
rect 26424 20356 26452 20412
rect 21974 19572 22002 19628
rect 22058 19572 22106 19628
rect 22162 19572 22210 19628
rect 22266 19572 22294 19628
rect 21974 18060 22294 19572
rect 18732 18004 18788 18014
rect 18732 17780 18788 17948
rect 18732 17714 18788 17724
rect 21974 18004 22002 18060
rect 22058 18004 22106 18060
rect 22162 18004 22210 18060
rect 22266 18004 22294 18060
rect 17816 17220 17844 17276
rect 17900 17220 17948 17276
rect 18004 17220 18052 17276
rect 18108 17220 18136 17276
rect 17816 15708 18136 17220
rect 17816 15652 17844 15708
rect 17900 15652 17948 15708
rect 18004 15652 18052 15708
rect 18108 15652 18136 15708
rect 17816 14140 18136 15652
rect 17816 14084 17844 14140
rect 17900 14084 17948 14140
rect 18004 14084 18052 14140
rect 18108 14084 18136 14140
rect 13658 13300 13686 13356
rect 13742 13300 13790 13356
rect 13846 13300 13894 13356
rect 13950 13300 13978 13356
rect 13658 11788 13978 13300
rect 16380 13748 16436 13758
rect 16380 12740 16436 13692
rect 16380 12674 16436 12684
rect 13658 11732 13686 11788
rect 13742 11732 13790 11788
rect 13846 11732 13894 11788
rect 13950 11732 13978 11788
rect 13658 10220 13978 11732
rect 13658 10164 13686 10220
rect 13742 10164 13790 10220
rect 13846 10164 13894 10220
rect 13950 10164 13978 10220
rect 13658 8652 13978 10164
rect 13658 8596 13686 8652
rect 13742 8596 13790 8652
rect 13846 8596 13894 8652
rect 13950 8596 13978 8652
rect 13658 7084 13978 8596
rect 13658 7028 13686 7084
rect 13742 7028 13790 7084
rect 13846 7028 13894 7084
rect 13950 7028 13978 7084
rect 13658 5516 13978 7028
rect 13658 5460 13686 5516
rect 13742 5460 13790 5516
rect 13846 5460 13894 5516
rect 13950 5460 13978 5516
rect 13658 3948 13978 5460
rect 13658 3892 13686 3948
rect 13742 3892 13790 3948
rect 13846 3892 13894 3948
rect 13950 3892 13978 3948
rect 13658 3076 13978 3892
rect 17816 12572 18136 14084
rect 21974 16492 22294 18004
rect 23548 20244 23604 20254
rect 23548 17668 23604 20188
rect 23548 17602 23604 17612
rect 26132 18844 26452 20356
rect 26132 18788 26160 18844
rect 26216 18788 26264 18844
rect 26320 18788 26368 18844
rect 26424 18788 26452 18844
rect 21974 16436 22002 16492
rect 22058 16436 22106 16492
rect 22162 16436 22210 16492
rect 22266 16436 22294 16492
rect 21974 14924 22294 16436
rect 21974 14868 22002 14924
rect 22058 14868 22106 14924
rect 22162 14868 22210 14924
rect 22266 14868 22294 14924
rect 18844 13748 18900 13758
rect 17816 12516 17844 12572
rect 17900 12516 17948 12572
rect 18004 12516 18052 12572
rect 18108 12516 18136 12572
rect 17816 11004 18136 12516
rect 18620 13636 18676 13646
rect 18620 12068 18676 13580
rect 18844 12740 18900 13692
rect 18844 12674 18900 12684
rect 21974 13356 22294 14868
rect 21974 13300 22002 13356
rect 22058 13300 22106 13356
rect 22162 13300 22210 13356
rect 22266 13300 22294 13356
rect 18620 12002 18676 12012
rect 17816 10948 17844 11004
rect 17900 10948 17948 11004
rect 18004 10948 18052 11004
rect 18108 10948 18136 11004
rect 17816 9436 18136 10948
rect 17816 9380 17844 9436
rect 17900 9380 17948 9436
rect 18004 9380 18052 9436
rect 18108 9380 18136 9436
rect 17816 7868 18136 9380
rect 17816 7812 17844 7868
rect 17900 7812 17948 7868
rect 18004 7812 18052 7868
rect 18108 7812 18136 7868
rect 17816 6300 18136 7812
rect 17816 6244 17844 6300
rect 17900 6244 17948 6300
rect 18004 6244 18052 6300
rect 18108 6244 18136 6300
rect 17816 4732 18136 6244
rect 17816 4676 17844 4732
rect 17900 4676 17948 4732
rect 18004 4676 18052 4732
rect 18108 4676 18136 4732
rect 17816 3164 18136 4676
rect 17816 3108 17844 3164
rect 17900 3108 17948 3164
rect 18004 3108 18052 3164
rect 18108 3108 18136 3164
rect 17816 3076 18136 3108
rect 21974 11788 22294 13300
rect 21974 11732 22002 11788
rect 22058 11732 22106 11788
rect 22162 11732 22210 11788
rect 22266 11732 22294 11788
rect 21974 10220 22294 11732
rect 21974 10164 22002 10220
rect 22058 10164 22106 10220
rect 22162 10164 22210 10220
rect 22266 10164 22294 10220
rect 21974 8652 22294 10164
rect 21974 8596 22002 8652
rect 22058 8596 22106 8652
rect 22162 8596 22210 8652
rect 22266 8596 22294 8652
rect 21974 7084 22294 8596
rect 21974 7028 22002 7084
rect 22058 7028 22106 7084
rect 22162 7028 22210 7084
rect 22266 7028 22294 7084
rect 21974 5516 22294 7028
rect 21974 5460 22002 5516
rect 22058 5460 22106 5516
rect 22162 5460 22210 5516
rect 22266 5460 22294 5516
rect 21974 3948 22294 5460
rect 21974 3892 22002 3948
rect 22058 3892 22106 3948
rect 22162 3892 22210 3948
rect 22266 3892 22294 3948
rect 21974 3076 22294 3892
rect 26132 17276 26452 18788
rect 26132 17220 26160 17276
rect 26216 17220 26264 17276
rect 26320 17220 26368 17276
rect 26424 17220 26452 17276
rect 26132 15708 26452 17220
rect 26132 15652 26160 15708
rect 26216 15652 26264 15708
rect 26320 15652 26368 15708
rect 26424 15652 26452 15708
rect 26132 14140 26452 15652
rect 26132 14084 26160 14140
rect 26216 14084 26264 14140
rect 26320 14084 26368 14140
rect 26424 14084 26452 14140
rect 26132 12572 26452 14084
rect 26132 12516 26160 12572
rect 26216 12516 26264 12572
rect 26320 12516 26368 12572
rect 26424 12516 26452 12572
rect 26132 11004 26452 12516
rect 26132 10948 26160 11004
rect 26216 10948 26264 11004
rect 26320 10948 26368 11004
rect 26424 10948 26452 11004
rect 26132 9436 26452 10948
rect 26132 9380 26160 9436
rect 26216 9380 26264 9436
rect 26320 9380 26368 9436
rect 26424 9380 26452 9436
rect 26132 7868 26452 9380
rect 26132 7812 26160 7868
rect 26216 7812 26264 7868
rect 26320 7812 26368 7868
rect 26424 7812 26452 7868
rect 26132 6300 26452 7812
rect 26132 6244 26160 6300
rect 26216 6244 26264 6300
rect 26320 6244 26368 6300
rect 26424 6244 26452 6300
rect 26132 4732 26452 6244
rect 26132 4676 26160 4732
rect 26216 4676 26264 4732
rect 26320 4676 26368 4732
rect 26424 4676 26452 4732
rect 26132 3164 26452 4676
rect 26132 3108 26160 3164
rect 26216 3108 26264 3164
rect 26320 3108 26368 3164
rect 26424 3108 26452 3164
rect 26132 3076 26452 3108
rect 30290 32172 30610 32204
rect 30290 32116 30318 32172
rect 30374 32116 30422 32172
rect 30478 32116 30526 32172
rect 30582 32116 30610 32172
rect 30290 30604 30610 32116
rect 30290 30548 30318 30604
rect 30374 30548 30422 30604
rect 30478 30548 30526 30604
rect 30582 30548 30610 30604
rect 30290 29036 30610 30548
rect 30290 28980 30318 29036
rect 30374 28980 30422 29036
rect 30478 28980 30526 29036
rect 30582 28980 30610 29036
rect 30290 27468 30610 28980
rect 30290 27412 30318 27468
rect 30374 27412 30422 27468
rect 30478 27412 30526 27468
rect 30582 27412 30610 27468
rect 30290 25900 30610 27412
rect 30290 25844 30318 25900
rect 30374 25844 30422 25900
rect 30478 25844 30526 25900
rect 30582 25844 30610 25900
rect 30290 24332 30610 25844
rect 30290 24276 30318 24332
rect 30374 24276 30422 24332
rect 30478 24276 30526 24332
rect 30582 24276 30610 24332
rect 30290 22764 30610 24276
rect 30290 22708 30318 22764
rect 30374 22708 30422 22764
rect 30478 22708 30526 22764
rect 30582 22708 30610 22764
rect 30290 21196 30610 22708
rect 30290 21140 30318 21196
rect 30374 21140 30422 21196
rect 30478 21140 30526 21196
rect 30582 21140 30610 21196
rect 30290 19628 30610 21140
rect 30290 19572 30318 19628
rect 30374 19572 30422 19628
rect 30478 19572 30526 19628
rect 30582 19572 30610 19628
rect 30290 18060 30610 19572
rect 30290 18004 30318 18060
rect 30374 18004 30422 18060
rect 30478 18004 30526 18060
rect 30582 18004 30610 18060
rect 30290 16492 30610 18004
rect 30290 16436 30318 16492
rect 30374 16436 30422 16492
rect 30478 16436 30526 16492
rect 30582 16436 30610 16492
rect 30290 14924 30610 16436
rect 30290 14868 30318 14924
rect 30374 14868 30422 14924
rect 30478 14868 30526 14924
rect 30582 14868 30610 14924
rect 30290 13356 30610 14868
rect 30290 13300 30318 13356
rect 30374 13300 30422 13356
rect 30478 13300 30526 13356
rect 30582 13300 30610 13356
rect 30290 11788 30610 13300
rect 30290 11732 30318 11788
rect 30374 11732 30422 11788
rect 30478 11732 30526 11788
rect 30582 11732 30610 11788
rect 30290 10220 30610 11732
rect 30290 10164 30318 10220
rect 30374 10164 30422 10220
rect 30478 10164 30526 10220
rect 30582 10164 30610 10220
rect 30290 8652 30610 10164
rect 30290 8596 30318 8652
rect 30374 8596 30422 8652
rect 30478 8596 30526 8652
rect 30582 8596 30610 8652
rect 30290 7084 30610 8596
rect 30290 7028 30318 7084
rect 30374 7028 30422 7084
rect 30478 7028 30526 7084
rect 30582 7028 30610 7084
rect 30290 5516 30610 7028
rect 30290 5460 30318 5516
rect 30374 5460 30422 5516
rect 30478 5460 30526 5516
rect 30582 5460 30610 5516
rect 30290 3948 30610 5460
rect 30290 3892 30318 3948
rect 30374 3892 30422 3948
rect 30478 3892 30526 3948
rect 30582 3892 30610 3948
rect 30290 3076 30610 3892
rect 34448 31388 34768 32204
rect 34448 31332 34476 31388
rect 34532 31332 34580 31388
rect 34636 31332 34684 31388
rect 34740 31332 34768 31388
rect 34448 29820 34768 31332
rect 34448 29764 34476 29820
rect 34532 29764 34580 29820
rect 34636 29764 34684 29820
rect 34740 29764 34768 29820
rect 34448 28252 34768 29764
rect 34448 28196 34476 28252
rect 34532 28196 34580 28252
rect 34636 28196 34684 28252
rect 34740 28196 34768 28252
rect 34448 26684 34768 28196
rect 34448 26628 34476 26684
rect 34532 26628 34580 26684
rect 34636 26628 34684 26684
rect 34740 26628 34768 26684
rect 34448 25116 34768 26628
rect 34448 25060 34476 25116
rect 34532 25060 34580 25116
rect 34636 25060 34684 25116
rect 34740 25060 34768 25116
rect 34448 23548 34768 25060
rect 34448 23492 34476 23548
rect 34532 23492 34580 23548
rect 34636 23492 34684 23548
rect 34740 23492 34768 23548
rect 34448 21980 34768 23492
rect 34448 21924 34476 21980
rect 34532 21924 34580 21980
rect 34636 21924 34684 21980
rect 34740 21924 34768 21980
rect 34448 20412 34768 21924
rect 34448 20356 34476 20412
rect 34532 20356 34580 20412
rect 34636 20356 34684 20412
rect 34740 20356 34768 20412
rect 34448 18844 34768 20356
rect 34448 18788 34476 18844
rect 34532 18788 34580 18844
rect 34636 18788 34684 18844
rect 34740 18788 34768 18844
rect 34448 17276 34768 18788
rect 34448 17220 34476 17276
rect 34532 17220 34580 17276
rect 34636 17220 34684 17276
rect 34740 17220 34768 17276
rect 34448 15708 34768 17220
rect 34448 15652 34476 15708
rect 34532 15652 34580 15708
rect 34636 15652 34684 15708
rect 34740 15652 34768 15708
rect 34448 14140 34768 15652
rect 34448 14084 34476 14140
rect 34532 14084 34580 14140
rect 34636 14084 34684 14140
rect 34740 14084 34768 14140
rect 34448 12572 34768 14084
rect 34448 12516 34476 12572
rect 34532 12516 34580 12572
rect 34636 12516 34684 12572
rect 34740 12516 34768 12572
rect 34448 11004 34768 12516
rect 34448 10948 34476 11004
rect 34532 10948 34580 11004
rect 34636 10948 34684 11004
rect 34740 10948 34768 11004
rect 34448 9436 34768 10948
rect 34448 9380 34476 9436
rect 34532 9380 34580 9436
rect 34636 9380 34684 9436
rect 34740 9380 34768 9436
rect 34448 7868 34768 9380
rect 34448 7812 34476 7868
rect 34532 7812 34580 7868
rect 34636 7812 34684 7868
rect 34740 7812 34768 7868
rect 34448 6300 34768 7812
rect 34448 6244 34476 6300
rect 34532 6244 34580 6300
rect 34636 6244 34684 6300
rect 34740 6244 34768 6300
rect 34448 4732 34768 6244
rect 34448 4676 34476 4732
rect 34532 4676 34580 4732
rect 34636 4676 34684 4732
rect 34740 4676 34768 4732
rect 34448 3164 34768 4676
rect 34448 3108 34476 3164
rect 34532 3108 34580 3164
rect 34636 3108 34684 3164
rect 34740 3108 34768 3164
rect 34448 3076 34768 3108
use gf180mcu_as_sc_mcu7t3v3__inv_2  _0481_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751532043
transform 1 0 23408 0 -1 17248
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _0482_
timestamp 1751532043
transform -1 0 23408 0 1 17248
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _0483_
timestamp 1751532043
transform -1 0 21616 0 1 18816
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _0484_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751740063
transform -1 0 19936 0 1 18816
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _0485_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1753960525
transform -1 0 20272 0 1 17248
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0486_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751534193
transform 1 0 17472 0 -1 15680
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _0487_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751531619
transform 1 0 17584 0 1 29792
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _0488_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751889808
transform -1 0 17920 0 1 28224
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _0489_
timestamp 1751740063
transform -1 0 13216 0 -1 29792
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0490_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751889408
transform -1 0 16016 0 1 28224
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _0491_
timestamp 1751531619
transform 1 0 13888 0 1 26656
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _0492_
timestamp 1751889808
transform -1 0 17024 0 1 26656
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _0493_
timestamp 1751532043
transform 1 0 18368 0 -1 25088
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__nand4_2  _0494_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1753172561
transform 1 0 23632 0 1 28224
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__nand4_2  _0495_
timestamp 1753172561
transform -1 0 28560 0 1 25088
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _0496_
timestamp 1751889808
transform -1 0 24304 0 1 25088
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _0497_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1753371985
transform -1 0 19824 0 1 23520
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _0498_
timestamp 1751740063
transform -1 0 24416 0 -1 26656
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _0499_
timestamp 1751531619
transform -1 0 19824 0 -1 23520
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0500_
timestamp 1751534193
transform 1 0 17696 0 -1 21952
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _0501_
timestamp 1753371985
transform -1 0 18816 0 -1 23520
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _0502_
timestamp 1751532043
transform -1 0 16240 0 1 20384
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _0503_
timestamp 1751740063
transform 1 0 12096 0 1 20384
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _0504_
timestamp 1753960525
transform 1 0 16016 0 1 18816
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _0505_
timestamp 1751532043
transform -1 0 18816 0 -1 21952
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _0506_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1753182340
transform 1 0 17024 0 1 21952
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0507_
timestamp 1751534193
transform 1 0 16352 0 -1 15680
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0508_
timestamp 1751889408
transform -1 0 19152 0 -1 14112
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand4_2  _0509_
timestamp 1753172561
transform 1 0 15456 0 1 12544
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _0510_
timestamp 1753960525
transform -1 0 17024 0 -1 14112
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__nand3_2  _0511_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1752345181
transform 1 0 15008 0 -1 9408
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _0512_
timestamp 1751532043
transform 1 0 11200 0 -1 6272
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0513_
timestamp 1751534193
transform -1 0 11536 0 -1 4704
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0514_
timestamp 1751534193
transform 1 0 11648 0 -1 6272
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0515_
timestamp 1751534193
transform 1 0 12096 0 1 4704
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _0516_
timestamp 1751532043
transform 1 0 15008 0 1 12544
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _0517_
timestamp 1753960525
transform -1 0 18368 0 -1 14112
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0518_
timestamp 1751534193
transform -1 0 19152 0 1 10976
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _0519_
timestamp 1753960525
transform -1 0 17024 0 -1 12544
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__nand2b_2  _0520_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751905124
transform -1 0 17024 0 1 10976
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0521_
timestamp 1751534193
transform -1 0 14000 0 -1 10976
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _0522_
timestamp 1751532043
transform -1 0 14448 0 1 12544
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _0523_
timestamp 1751740063
transform 1 0 17024 0 1 26656
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _0524_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1753441877
transform -1 0 19376 0 1 21952
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__nand4_2  _0525_
timestamp 1753172561
transform 1 0 17136 0 1 18816
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _0526_
timestamp 1751531619
transform 1 0 18480 0 -1 12544
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _0527_
timestamp 1753182340
transform 1 0 17248 0 -1 12544
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _0528_
timestamp 1751889808
transform -1 0 17024 0 -1 6272
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0529_
timestamp 1751534193
transform 1 0 17808 0 -1 4704
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0530_
timestamp 1751534193
transform 1 0 17248 0 -1 6272
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0531_
timestamp 1751534193
transform 1 0 17808 0 1 14112
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _0532_
timestamp 1753371985
transform -1 0 19040 0 1 6272
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _0533_
timestamp 1751531619
transform 1 0 17136 0 1 6272
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _0534_
timestamp 1751532043
transform -1 0 15120 0 -1 6272
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0535_
timestamp 1751534193
transform -1 0 11088 0 -1 6272
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0536_
timestamp 1751534193
transform -1 0 10080 0 -1 4704
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0537_
timestamp 1751534193
transform -1 0 16016 0 -1 6272
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _0538_
timestamp 1751532043
transform 1 0 19488 0 1 12544
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _0539_
timestamp 1753441877
transform -1 0 18368 0 1 12544
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _0540_
timestamp 1753960525
transform 1 0 18368 0 1 12544
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0541_
timestamp 1751534193
transform -1 0 14560 0 1 10976
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _0542_
timestamp 1751740063
transform -1 0 13328 0 -1 10976
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _0543_
timestamp 1751532043
transform -1 0 13776 0 1 10976
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0544_
timestamp 1751889408
transform -1 0 12768 0 1 9408
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _0545_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751914308
transform -1 0 12096 0 1 4704
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _0546_
timestamp 1753960525
transform 1 0 19040 0 -1 6272
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _0547_
timestamp 1753441877
transform -1 0 19824 0 1 4704
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__nand2b_2  _0548_
timestamp 1751905124
transform -1 0 19040 0 -1 6272
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _0549_
timestamp 1751532043
transform -1 0 17136 0 1 6272
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _0550_
timestamp 1753441877
transform 1 0 11536 0 -1 4704
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _0551_
timestamp 1753960525
transform 1 0 12432 0 -1 6272
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__nand3_2  _0552_
timestamp 1752345181
transform -1 0 18704 0 1 4704
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _0553_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1753277515
transform 1 0 4592 0 -1 4704
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _0554_
timestamp 1751531619
transform -1 0 5040 0 1 3136
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0555_
timestamp 1751534193
transform -1 0 3696 0 1 4704
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0556_
timestamp 1751534193
transform -1 0 2912 0 -1 6272
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0557_
timestamp 1751534193
transform 1 0 15344 0 1 6272
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nand3_2  _0558_
timestamp 1752345181
transform -1 0 16576 0 1 9408
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0559_
timestamp 1751889408
transform -1 0 15008 0 -1 10976
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0560_
timestamp 1751534193
transform 1 0 14336 0 -1 9408
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0561_
timestamp 1751534193
transform -1 0 16688 0 1 6272
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _0562_
timestamp 1753441877
transform -1 0 16240 0 -1 7840
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0563_
timestamp 1751889408
transform 1 0 14336 0 1 6272
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0564_
timestamp 1751534193
transform -1 0 12992 0 1 10976
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0565_
timestamp 1751534193
transform -1 0 12320 0 1 10976
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _0566_
timestamp 1753371985
transform 1 0 9968 0 -1 12544
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0567_
timestamp 1751889408
transform -1 0 11984 0 1 9408
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _0568_
timestamp 1753182340
transform -1 0 9968 0 1 10976
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _0569_
timestamp 1751532043
transform 1 0 11984 0 -1 10976
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _0570_
timestamp 1753960525
transform 1 0 12320 0 -1 7840
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _0571_
timestamp 1751889808
transform 1 0 13328 0 1 6272
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0572_
timestamp 1751534193
transform 1 0 5488 0 1 6272
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0573_
timestamp 1751534193
transform -1 0 10864 0 -1 4704
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _0574_
timestamp 1751889808
transform -1 0 12768 0 -1 9408
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _0575_
timestamp 1753960525
transform -1 0 12096 0 1 6272
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _0576_
timestamp 1751531619
transform -1 0 11648 0 1 12544
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0577_
timestamp 1751534193
transform -1 0 10640 0 1 10976
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _0578_
timestamp 1751532043
transform 1 0 11088 0 -1 9408
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _0579_
timestamp 1753182340
transform -1 0 12320 0 -1 7840
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _0580_
timestamp 1751740063
transform 1 0 13328 0 1 7840
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _0581_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1753868718
transform 1 0 13888 0 -1 7840
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0582_
timestamp 1751534193
transform 1 0 15568 0 1 7840
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _0583_
timestamp 1751889808
transform -1 0 11536 0 1 10976
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _0584_
timestamp 1753441877
transform -1 0 8400 0 1 4704
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _0585_
timestamp 1751531619
transform 1 0 3696 0 1 4704
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _0586_
timestamp 1751889808
transform 1 0 4704 0 -1 6272
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0587_
timestamp 1751534193
transform -1 0 9072 0 1 6272
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _0588_
timestamp 1751914308
transform 1 0 6944 0 -1 6272
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _0589_
timestamp 1753441877
transform -1 0 13888 0 -1 9408
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _0590_
timestamp 1751531619
transform 1 0 5488 0 1 9408
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0591_
timestamp 1751534193
transform -1 0 7504 0 1 7840
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _0592_
timestamp 1753371985
transform 1 0 5712 0 -1 9408
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _0593_
timestamp 1753371985
transform 1 0 7056 0 -1 9408
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _0594_
timestamp 1751531619
transform -1 0 11200 0 1 9408
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0595_
timestamp 1751534193
transform -1 0 10192 0 -1 10976
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _0596_
timestamp 1753441877
transform -1 0 10864 0 -1 7840
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__aoi22_2  _0597_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1753579406
transform 1 0 7728 0 1 7840
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _0598_
timestamp 1751889808
transform 1 0 7056 0 1 9408
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _0599_
timestamp 1753277515
transform -1 0 8624 0 -1 4704
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _0600_
timestamp 1753371985
transform 1 0 7280 0 1 6272
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _0601_
timestamp 1751531619
transform -1 0 8960 0 -1 9408
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand3_2  _0602_
timestamp 1752345181
transform 1 0 9296 0 1 7840
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _0603_
timestamp 1751889808
transform -1 0 8624 0 1 9408
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _0604_
timestamp 1753441877
transform -1 0 10640 0 1 12544
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0605_
timestamp 1751534193
transform -1 0 15568 0 1 7840
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _0606_
timestamp 1751531619
transform 1 0 4144 0 1 9408
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__aoi31_2  _0607_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1753891287
transform -1 0 6160 0 -1 10976
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0608_
timestamp 1751534193
transform 1 0 13328 0 1 12544
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _0609_
timestamp 1753441877
transform -1 0 12208 0 -1 12544
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__aoi31_2  _0610_
timestamp 1753891287
transform 1 0 7392 0 -1 12544
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _0611_
timestamp 1751532043
transform -1 0 3024 0 1 4704
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0612_
timestamp 1751889408
transform -1 0 7952 0 -1 7840
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _0613_
timestamp 1753868718
transform 1 0 6832 0 1 10976
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _0614_
timestamp 1753960525
transform -1 0 8512 0 -1 10976
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0615_
timestamp 1751534193
transform -1 0 7728 0 1 14112
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0616_
timestamp 1751534193
transform -1 0 3136 0 -1 10976
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _0617_
timestamp 1751889808
transform -1 0 3920 0 -1 10976
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _0618_
timestamp 1751740063
transform -1 0 4704 0 -1 9408
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _0619_
timestamp 1753868718
transform -1 0 4144 0 1 9408
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0620_
timestamp 1751534193
transform -1 0 4592 0 -1 10976
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _0621_
timestamp 1753371985
transform -1 0 3696 0 -1 12544
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _0622_
timestamp 1751531619
transform -1 0 4816 0 1 7840
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _0623_
timestamp 1751889808
transform -1 0 3248 0 -1 14112
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _0624_
timestamp 1753371985
transform 1 0 3248 0 -1 14112
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _0625_
timestamp 1751531619
transform 1 0 2128 0 1 12544
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _0626_
timestamp 1751531619
transform -1 0 5264 0 1 12544
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _0627_
timestamp 1751531619
transform -1 0 5824 0 -1 12544
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _0628_
timestamp 1753960525
transform -1 0 4480 0 1 10976
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _0629_
timestamp 1751914308
transform 1 0 3696 0 -1 12544
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _0630_
timestamp 1751740063
transform -1 0 6272 0 1 12544
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _0631_
timestamp 1753371985
transform -1 0 5488 0 -1 14112
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__aoi22_2  _0632_
timestamp 1753579406
transform 1 0 2912 0 1 12544
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _0633_
timestamp 1753371985
transform -1 0 5264 0 1 6272
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_4  _0634_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1753432499
transform 1 0 10976 0 1 7840
box -86 -86 2214 870
use gf180mcu_as_sc_mcu7t3v3__nor2b_2  _0635_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1752061876
transform -1 0 3920 0 -1 7840
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _0636_
timestamp 1753868718
transform -1 0 4144 0 -1 6272
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _0637_
timestamp 1753441877
transform -1 0 7280 0 1 4704
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _0638_
timestamp 1751531619
transform -1 0 10752 0 1 4704
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _0639_
timestamp 1753441877
transform -1 0 6720 0 -1 6272
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _0640_
timestamp 1753371985
transform 1 0 2688 0 -1 9408
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _0641_
timestamp 1753371985
transform 1 0 2912 0 1 7840
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _0642_
timestamp 1753868718
transform -1 0 4144 0 1 6272
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0643_
timestamp 1751534193
transform -1 0 3472 0 1 14112
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _0644_
timestamp 1751531619
transform 1 0 4480 0 1 4704
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _0645_
timestamp 1751889808
transform -1 0 18256 0 1 10976
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _0646_
timestamp 1753960525
transform -1 0 15904 0 1 10976
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__nand2b_2  _0647_
timestamp 1751905124
transform -1 0 8624 0 1 12544
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _0648_
timestamp 1753371985
transform 1 0 6160 0 -1 12544
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _0649_
timestamp 1753868718
transform -1 0 7504 0 1 12544
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0650_
timestamp 1751534193
transform 1 0 6384 0 1 14112
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0651_
timestamp 1751889408
transform 1 0 26432 0 1 20384
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0652_
timestamp 1751534193
transform -1 0 26768 0 1 4704
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0653_
timestamp 1751534193
transform -1 0 22624 0 1 6272
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0654_
timestamp 1751534193
transform 1 0 14784 0 -1 14112
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _0655_
timestamp 1751532043
transform -1 0 21616 0 1 4704
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _0656_
timestamp 1751889808
transform -1 0 30352 0 -1 18816
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _0657_
timestamp 1751532043
transform -1 0 33376 0 -1 18816
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _0658_
timestamp 1751532043
transform 1 0 26096 0 1 15680
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__nand4_2  _0659_
timestamp 1753172561
transform -1 0 31360 0 1 17248
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _0660_
timestamp 1753182340
transform 1 0 29344 0 -1 17248
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _0661_
timestamp 1751740063
transform 1 0 25088 0 -1 9408
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0662_
timestamp 1751889408
transform 1 0 26432 0 1 12544
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _0663_
timestamp 1751740063
transform -1 0 22400 0 1 9408
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0664_
timestamp 1751889408
transform 1 0 29232 0 -1 7840
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand4_2  _0665_
timestamp 1753172561
transform 1 0 25424 0 1 9408
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _0666_
timestamp 1751532043
transform -1 0 32144 0 1 7840
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _0667_
timestamp 1751740063
transform -1 0 31472 0 -1 10976
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _0668_
timestamp 1751740063
transform 1 0 26768 0 1 4704
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0669_
timestamp 1751889408
transform -1 0 29792 0 1 4704
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand4_2  _0670_
timestamp 1753172561
transform -1 0 30464 0 -1 10976
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _0671_
timestamp 1751740063
transform -1 0 25872 0 -1 10976
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand3_2  _0672_
timestamp 1752345181
transform 1 0 23632 0 -1 12544
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _0673_
timestamp 1751531619
transform 1 0 23072 0 -1 14112
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0674_
timestamp 1751534193
transform -1 0 28784 0 1 12544
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0675_
timestamp 1751534193
transform -1 0 28000 0 1 7840
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _0676_
timestamp 1751740063
transform -1 0 21952 0 1 7840
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0677_
timestamp 1751534193
transform 1 0 19488 0 1 15680
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0678_
timestamp 1751534193
transform 1 0 22624 0 1 23520
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0679_
timestamp 1751889408
transform 1 0 22512 0 -1 9408
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _0680_
timestamp 1753182340
transform -1 0 23632 0 1 9408
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0681_
timestamp 1751534193
transform -1 0 21392 0 -1 10976
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0682_
timestamp 1751534193
transform 1 0 30128 0 -1 15680
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0683_
timestamp 1751534193
transform -1 0 26544 0 -1 14112
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _0684_
timestamp 1753277515
transform -1 0 24192 0 -1 10976
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _0685_
timestamp 1751740063
transform -1 0 25984 0 1 10976
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand4_2  _0686_
timestamp 1753172561
transform 1 0 22288 0 1 7840
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _0687_
timestamp 1753960525
transform 1 0 22736 0 -1 7840
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _0688_
timestamp 1751531619
transform -1 0 24640 0 -1 7840
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _0689_
timestamp 1751740063
transform -1 0 24640 0 1 7840
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _0690_
timestamp 1751532043
transform -1 0 25536 0 -1 6272
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _0691_
timestamp 1751740063
transform -1 0 24752 0 -1 4704
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0692_
timestamp 1751889408
transform -1 0 24080 0 1 3136
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _0693_
timestamp 1753182340
transform 1 0 22736 0 -1 4704
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0694_
timestamp 1751534193
transform 1 0 24192 0 -1 6272
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _0695_
timestamp 1753182340
transform 1 0 22960 0 -1 6272
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _0696_
timestamp 1751740063
transform 1 0 22176 0 -1 6272
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _0697_
timestamp 1753182340
transform 1 0 21616 0 1 4704
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0698_
timestamp 1751534193
transform -1 0 21504 0 1 3136
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _0699_
timestamp 1751740063
transform -1 0 28672 0 1 6272
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0700_
timestamp 1751889408
transform -1 0 29232 0 1 3136
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _0701_
timestamp 1753182340
transform 1 0 27552 0 1 4704
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0702_
timestamp 1751534193
transform -1 0 26432 0 -1 4704
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0703_
timestamp 1751534193
transform 1 0 28112 0 1 7840
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _0704_
timestamp 1751740063
transform -1 0 31584 0 1 3136
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0705_
timestamp 1751889408
transform 1 0 32032 0 1 3136
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _0706_
timestamp 1753182340
transform 1 0 30128 0 1 4704
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0707_
timestamp 1751534193
transform 1 0 32816 0 1 3136
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _0708_
timestamp 1751740063
transform 1 0 31472 0 -1 7840
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0709_
timestamp 1751889408
transform -1 0 33712 0 -1 6272
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _0710_
timestamp 1753182340
transform 1 0 31360 0 -1 6272
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0711_
timestamp 1751534193
transform 1 0 32928 0 -1 7840
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _0712_
timestamp 1753277515
transform 1 0 29344 0 1 6272
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _0713_
timestamp 1751740063
transform 1 0 26768 0 -1 7840
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand4_2  _0714_
timestamp 1753172561
transform -1 0 30688 0 -1 6272
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _0715_
timestamp 1751740063
transform 1 0 27776 0 -1 9408
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _0716_
timestamp 1751889808
transform 1 0 29008 0 1 7840
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _0717_
timestamp 1753371985
transform 1 0 28560 0 -1 9408
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _0718_
timestamp 1751740063
transform -1 0 31024 0 1 9408
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _0719_
timestamp 1751532043
transform -1 0 27552 0 1 9408
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _0720_
timestamp 1753182340
transform 1 0 27552 0 1 9408
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _0721_
timestamp 1753182340
transform -1 0 30240 0 1 9408
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0722_
timestamp 1751534193
transform -1 0 27552 0 1 10976
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _0723_
timestamp 1751740063
transform -1 0 33376 0 1 10976
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0724_
timestamp 1751889408
transform 1 0 32928 0 -1 10976
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _0725_
timestamp 1753182340
transform 1 0 31472 0 -1 10976
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0726_
timestamp 1751534193
transform 1 0 32928 0 -1 9408
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0727_
timestamp 1751534193
transform 1 0 29008 0 1 12544
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _0728_
timestamp 1751740063
transform -1 0 34160 0 1 12544
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0729_
timestamp 1751889408
transform -1 0 32592 0 1 10976
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _0730_
timestamp 1753182340
transform 1 0 31024 0 -1 12544
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0731_
timestamp 1751534193
transform -1 0 30352 0 1 12544
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nand3_2  _0732_
timestamp 1752345181
transform 1 0 31472 0 -1 14112
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _0733_
timestamp 1751740063
transform 1 0 30688 0 -1 14112
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _0734_
timestamp 1751740063
transform 1 0 30576 0 1 14112
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0735_
timestamp 1751889408
transform 1 0 31472 0 -1 15680
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0736_
timestamp 1751534193
transform 1 0 32928 0 -1 14112
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _0737_
timestamp 1751532043
transform -1 0 31136 0 -1 17248
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _0738_
timestamp 1751740063
transform 1 0 30464 0 -1 18816
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _0739_
timestamp 1751889808
transform 1 0 32928 0 -1 17248
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _0740_
timestamp 1753371985
transform 1 0 31472 0 1 15680
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _0741_
timestamp 1751740063
transform -1 0 32480 0 -1 20384
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _0742_
timestamp 1753182340
transform 1 0 31136 0 -1 17248
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _0743_
timestamp 1753182340
transform 1 0 31248 0 -1 18816
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0744_
timestamp 1751534193
transform 1 0 32928 0 -1 20384
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _0745_
timestamp 1751740063
transform -1 0 29792 0 1 18816
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0746_
timestamp 1751889408
transform -1 0 29792 0 1 17248
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0747_
timestamp 1751534193
transform -1 0 29344 0 -1 15680
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _0748_
timestamp 1753182340
transform -1 0 29344 0 -1 18816
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0749_
timestamp 1751534193
transform -1 0 28560 0 1 20384
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _0750_
timestamp 1751740063
transform -1 0 28672 0 -1 15680
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0751_
timestamp 1751889408
transform 1 0 29008 0 1 14112
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _0752_
timestamp 1753182340
transform -1 0 28560 0 1 14112
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0753_
timestamp 1751534193
transform -1 0 28112 0 1 12544
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _0754_
timestamp 1753277515
transform -1 0 27104 0 1 14112
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _0755_
timestamp 1751740063
transform -1 0 25872 0 -1 14112
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _0756_
timestamp 1751531619
transform 1 0 27104 0 -1 15680
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _0757_
timestamp 1753960525
transform 1 0 27664 0 1 15680
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _0758_
timestamp 1753371985
transform 1 0 26544 0 1 15680
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__aoi31_2  _0759_
timestamp 1753891287
transform 1 0 26544 0 1 17248
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _0760_
timestamp 1751532043
transform -1 0 28560 0 1 17248
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _0761_
timestamp 1753182340
transform 1 0 28112 0 -1 17248
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _0762_
timestamp 1753182340
transform 1 0 26880 0 -1 18816
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0763_
timestamp 1751534193
transform -1 0 26992 0 -1 20384
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _0764_
timestamp 1751889808
transform -1 0 29680 0 -1 21952
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _0765_
timestamp 1753371985
transform 1 0 30016 0 -1 20384
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0766_
timestamp 1751889408
transform 1 0 31808 0 1 20384
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0767_
timestamp 1751534193
transform -1 0 31024 0 -1 23520
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0768_
timestamp 1751534193
transform 1 0 20272 0 -1 23520
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0769_
timestamp 1751534193
transform 1 0 21504 0 -1 21952
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0770_
timestamp 1751889408
transform -1 0 18480 0 -1 20384
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0771_
timestamp 1751534193
transform 1 0 19936 0 1 18816
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _0772_
timestamp 1751531619
transform 1 0 17248 0 -1 18816
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0773_
timestamp 1751534193
transform 1 0 20272 0 1 17248
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _0774_
timestamp 1751740063
transform 1 0 18704 0 1 15680
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0775_
timestamp 1751889408
transform 1 0 20160 0 1 20384
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _0776_
timestamp 1753960525
transform 1 0 22288 0 1 20384
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0777_
timestamp 1751534193
transform 1 0 23520 0 -1 20384
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0778_
timestamp 1751534193
transform -1 0 18256 0 1 23520
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _0779_
timestamp 1751740063
transform 1 0 6160 0 -1 23520
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _0780_
timestamp 1751532043
transform 1 0 13328 0 1 25088
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _0781_
timestamp 1751740063
transform -1 0 10192 0 -1 26656
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _0782_
timestamp 1753182340
transform -1 0 8736 0 1 23520
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _0783_
timestamp 1753960525
transform -1 0 8848 0 -1 23520
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0784_
timestamp 1751889408
transform -1 0 9632 0 1 23520
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _0785_
timestamp 1751889808
transform -1 0 25872 0 -1 23520
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _0786_
timestamp 1751531619
transform 1 0 22288 0 1 21952
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _0787_
timestamp 1753371985
transform -1 0 24192 0 -1 21952
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0788_
timestamp 1751534193
transform -1 0 8736 0 -1 21952
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _0789_
timestamp 1751889808
transform -1 0 4368 0 1 17248
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0790_
timestamp 1751889408
transform -1 0 4256 0 1 20384
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0791_
timestamp 1751534193
transform -1 0 3584 0 1 17248
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0792_
timestamp 1751534193
transform 1 0 4368 0 1 17248
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _0793_
timestamp 1751889808
transform -1 0 5488 0 -1 18816
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0794_
timestamp 1751534193
transform -1 0 4592 0 -1 17248
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0795_
timestamp 1751534193
transform 1 0 4592 0 -1 17248
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__aoi22_2  _0796_
timestamp 1753579406
transform 1 0 3136 0 -1 18816
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__nand3_2  _0797_
timestamp 1752345181
transform -1 0 4368 0 1 18816
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _0798_
timestamp 1751889808
transform -1 0 4144 0 1 23520
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0799_
timestamp 1751889408
transform -1 0 16912 0 1 23520
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0800_
timestamp 1751534193
transform -1 0 14560 0 1 25088
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0801_
timestamp 1751889408
transform -1 0 16688 0 -1 25088
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0802_
timestamp 1751534193
transform 1 0 15232 0 1 25088
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0803_
timestamp 1751889408
transform -1 0 4704 0 -1 25088
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _0804_
timestamp 1753960525
transform 1 0 3584 0 1 21952
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0805_
timestamp 1751534193
transform -1 0 3136 0 1 21952
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _0806_
timestamp 1751532043
transform 1 0 4816 0 -1 21952
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _0807_
timestamp 1751531619
transform 1 0 2352 0 1 18816
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _0808_
timestamp 1751914308
transform 1 0 2912 0 -1 20384
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _0809_
timestamp 1751889808
transform -1 0 4816 0 -1 21952
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0810_
timestamp 1751534193
transform 1 0 9520 0 1 21952
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _0811_
timestamp 1751889808
transform -1 0 6384 0 1 23520
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0812_
timestamp 1751889408
transform -1 0 5488 0 -1 25088
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _0813_
timestamp 1753960525
transform -1 0 5264 0 1 23520
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0814_
timestamp 1751534193
transform -1 0 3136 0 -1 25088
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _0815_
timestamp 1751531619
transform 1 0 4368 0 1 18816
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _0816_
timestamp 1751889808
transform 1 0 8288 0 -1 20384
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _0817_
timestamp 1751532043
transform 1 0 7616 0 1 17248
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _0818_
timestamp 1751531619
transform 1 0 6832 0 1 17248
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _0819_
timestamp 1751531619
transform -1 0 8624 0 1 18816
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand4_2  _0820_
timestamp 1753172561
transform 1 0 6720 0 -1 20384
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _0821_
timestamp 1751889808
transform -1 0 10416 0 1 23520
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0822_
timestamp 1751889408
transform 1 0 6608 0 -1 25088
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _0823_
timestamp 1753960525
transform -1 0 7504 0 1 23520
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0824_
timestamp 1751534193
transform -1 0 5264 0 1 25088
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0825_
timestamp 1751534193
transform -1 0 21504 0 -1 21952
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0826_
timestamp 1751534193
transform 1 0 12432 0 1 21952
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _0827_
timestamp 1751532043
transform 1 0 13104 0 -1 21952
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0828_
timestamp 1751534193
transform 1 0 16912 0 1 23520
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0829_
timestamp 1751534193
transform 1 0 17248 0 -1 25088
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _0830_
timestamp 1751531619
transform 1 0 5488 0 1 17248
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _0831_
timestamp 1751914308
transform 1 0 6944 0 -1 18816
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _0832_
timestamp 1753868718
transform 1 0 11088 0 1 21952
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _0833_
timestamp 1753960525
transform 1 0 12880 0 -1 23520
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0834_
timestamp 1751889408
transform -1 0 14112 0 1 21952
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0835_
timestamp 1751534193
transform -1 0 12208 0 -1 21952
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nand2b_2  _0836_
timestamp 1751905124
transform -1 0 6608 0 1 18816
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _0837_
timestamp 1751889808
transform -1 0 5040 0 -1 20384
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _0838_
timestamp 1751740063
transform 1 0 8288 0 -1 18816
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _0839_
timestamp 1751531619
transform 1 0 8624 0 1 18816
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand3_2  _0840_
timestamp 1752345181
transform 1 0 5040 0 -1 20384
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _0841_
timestamp 1753960525
transform 1 0 5488 0 1 20384
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _0842_
timestamp 1751889808
transform -1 0 7616 0 1 25088
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0843_
timestamp 1751889408
transform -1 0 6832 0 1 25088
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _0844_
timestamp 1753960525
transform 1 0 7392 0 -1 25088
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0845_
timestamp 1751534193
transform 1 0 8064 0 -1 28224
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0846_
timestamp 1751889408
transform 1 0 6160 0 -1 18816
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _0847_
timestamp 1753960525
transform 1 0 6720 0 1 18816
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _0848_
timestamp 1751531619
transform 1 0 7056 0 1 20384
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _0849_
timestamp 1751889808
transform -1 0 12880 0 -1 26656
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0850_
timestamp 1751889408
transform -1 0 9072 0 -1 26656
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _0851_
timestamp 1753960525
transform -1 0 8736 0 1 25088
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0852_
timestamp 1751534193
transform -1 0 7392 0 1 26656
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _0853_
timestamp 1753277515
transform 1 0 4592 0 -1 23520
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _0854_
timestamp 1753371985
transform 1 0 7280 0 1 21952
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _0855_
timestamp 1753960525
transform 1 0 8400 0 1 21952
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0856_
timestamp 1751534193
transform -1 0 18256 0 -1 17248
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0857_
timestamp 1751534193
transform -1 0 14784 0 1 21952
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _0858_
timestamp 1753371985
transform 1 0 10864 0 1 23520
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0859_
timestamp 1751889408
transform 1 0 12208 0 -1 25088
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0860_
timestamp 1751534193
transform -1 0 11648 0 -1 26656
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao22_2  _0861_
timestamp 1753868718
transform 1 0 15904 0 1 25088
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0862_
timestamp 1751534193
transform 1 0 17136 0 1 25088
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _0863_
timestamp 1751740063
transform -1 0 23520 0 -1 25088
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0864_
timestamp 1751889408
transform 1 0 24304 0 1 25088
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _0865_
timestamp 1753182340
transform 1 0 23520 0 -1 25088
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0866_
timestamp 1751534193
transform 1 0 25088 0 -1 25088
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _0867_
timestamp 1751740063
transform -1 0 27552 0 1 23520
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0868_
timestamp 1751889408
transform 1 0 27328 0 -1 25088
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _0869_
timestamp 1753182340
transform 1 0 27552 0 1 23520
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0870_
timestamp 1751534193
transform 1 0 29008 0 1 23520
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _0871_
timestamp 1751740063
transform -1 0 29120 0 -1 26656
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0872_
timestamp 1751889408
transform 1 0 29120 0 -1 26656
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _0873_
timestamp 1753182340
transform 1 0 28112 0 -1 25088
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0874_
timestamp 1751534193
transform 1 0 29344 0 -1 25088
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0875_
timestamp 1751534193
transform 1 0 22848 0 -1 26656
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _0876_
timestamp 1751740063
transform -1 0 28112 0 -1 26656
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0877_
timestamp 1751889408
transform -1 0 28672 0 -1 28224
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _0878_
timestamp 1753182340
transform 1 0 26656 0 -1 28224
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0879_
timestamp 1751534193
transform -1 0 26992 0 -1 26656
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _0880_
timestamp 1751740063
transform 1 0 26544 0 1 28224
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0881_
timestamp 1751889408
transform 1 0 27328 0 1 28224
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0882_
timestamp 1751889408
transform 1 0 28672 0 -1 28224
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _0883_
timestamp 1753182340
transform 1 0 26768 0 -1 29792
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0884_
timestamp 1751534193
transform 1 0 27216 0 -1 31360
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _0885_
timestamp 1751740063
transform 1 0 25088 0 -1 28224
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0886_
timestamp 1751889408
transform 1 0 25200 0 1 28224
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _0887_
timestamp 1753182340
transform 1 0 25088 0 -1 29792
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0888_
timestamp 1751534193
transform -1 0 25760 0 -1 31360
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _0889_
timestamp 1751740063
transform 1 0 22400 0 -1 29792
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0890_
timestamp 1751889408
transform 1 0 24640 0 1 29792
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _0891_
timestamp 1753182340
transform 1 0 23184 0 -1 29792
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0892_
timestamp 1751534193
transform -1 0 23408 0 1 28224
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _0893_
timestamp 1751889808
transform -1 0 24080 0 -1 28224
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0894_
timestamp 1751889408
transform 1 0 20160 0 1 26656
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _0895_
timestamp 1751531619
transform -1 0 22624 0 -1 25088
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0896_
timestamp 1751889408
transform 1 0 20720 0 -1 26656
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0897_
timestamp 1751534193
transform 1 0 21168 0 -1 28224
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _0898_
timestamp 1753960525
transform 1 0 19824 0 1 23520
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _0899_
timestamp 1753371985
transform 1 0 19600 0 1 25088
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0900_
timestamp 1751534193
transform -1 0 17472 0 1 17248
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0901_
timestamp 1751534193
transform -1 0 16240 0 1 17248
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _0902_
timestamp 1751889808
transform -1 0 12096 0 1 20384
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _0903_
timestamp 1751532043
transform -1 0 12880 0 1 17248
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _0904_
timestamp 1751914308
transform 1 0 11088 0 1 17248
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _0905_
timestamp 1753371985
transform -1 0 13552 0 -1 20384
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0906_
timestamp 1751889408
transform -1 0 11872 0 1 18816
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0907_
timestamp 1751534193
transform -1 0 11088 0 1 18816
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__inv_2  _0908_
timestamp 1751532043
transform -1 0 18592 0 -1 15680
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _0909_
timestamp 1753277515
transform -1 0 14000 0 -1 17248
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0910_
timestamp 1751889408
transform 1 0 12208 0 -1 18816
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _0911_
timestamp 1751914308
transform 1 0 12992 0 -1 18816
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _0912_
timestamp 1753960525
transform 1 0 15456 0 -1 18816
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0913_
timestamp 1751889408
transform -1 0 15568 0 1 17248
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0914_
timestamp 1751534193
transform -1 0 10976 0 1 17248
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _0915_
timestamp 1751740063
transform 1 0 13888 0 1 20384
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _0916_
timestamp 1751914308
transform 1 0 14224 0 1 18816
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _0917_
timestamp 1753960525
transform 1 0 14336 0 -1 18816
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _0918_
timestamp 1751740063
transform -1 0 15680 0 1 20384
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__or2_2  _0919_
timestamp 1751889808
transform -1 0 14112 0 1 18816
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _0920_
timestamp 1753371985
transform 1 0 11984 0 1 18816
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__mux2_2  _0921_
timestamp 1751914308
transform 1 0 13440 0 1 17248
box -86 -86 1430 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _0922_
timestamp 1753960525
transform 1 0 14336 0 -1 15680
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0923_
timestamp 1751889408
transform 1 0 14560 0 -1 17248
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0924_
timestamp 1751534193
transform 1 0 15344 0 -1 17248
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _0925_
timestamp 1753441877
transform -1 0 22960 0 1 17248
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _0926_
timestamp 1753371985
transform 1 0 20720 0 -1 17248
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _0927_
timestamp 1751531619
transform 1 0 18368 0 1 17248
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _0928_
timestamp 1753441877
transform 1 0 18256 0 -1 17248
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _0929_
timestamp 1753371985
transform -1 0 20496 0 -1 17248
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0930_
timestamp 1751889408
transform 1 0 21840 0 -1 20384
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _0931_
timestamp 1753960525
transform -1 0 22288 0 1 20384
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0932_
timestamp 1751534193
transform -1 0 20160 0 1 20384
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _0933_
timestamp 1753277515
transform 1 0 21840 0 -1 17248
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _0934_
timestamp 1753441877
transform 1 0 20832 0 -1 18816
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__aoi21_2  _0935_
timestamp 1753371985
transform -1 0 23072 0 -1 18816
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__ao21_2  _0936_
timestamp 1753441877
transform 1 0 11984 0 1 23520
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0937_
timestamp 1751534193
transform 1 0 14560 0 1 25088
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _0938_
timestamp 1753277515
transform 1 0 21392 0 1 12544
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0939_
timestamp 1751889408
transform 1 0 21056 0 -1 14112
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0940_
timestamp 1751534193
transform 1 0 21840 0 -1 14112
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _0941_
timestamp 1751531619
transform -1 0 19488 0 1 25088
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0942_
timestamp 1751534193
transform 1 0 20272 0 1 29792
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _0943_
timestamp 1751740063
transform -1 0 12320 0 -1 29792
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0944_
timestamp 1751889408
transform 1 0 13216 0 -1 29792
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _0945_
timestamp 1753182340
transform 1 0 12096 0 -1 28224
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0946_
timestamp 1751534193
transform -1 0 11536 0 -1 28224
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _0947_
timestamp 1753277515
transform -1 0 14896 0 1 29792
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _0948_
timestamp 1751740063
transform -1 0 13776 0 1 31360
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0949_
timestamp 1751889408
transform 1 0 14112 0 -1 29792
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__ao31_2  _0950_
timestamp 1753960525
transform 1 0 13328 0 1 28224
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__nand2_2  _0951_
timestamp 1751531619
transform 1 0 14448 0 1 28224
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _0952_
timestamp 1751740063
transform -1 0 15456 0 1 26656
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _0953_
timestamp 1751740063
transform -1 0 16464 0 -1 29792
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0954_
timestamp 1751889408
transform 1 0 16800 0 1 29792
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _0955_
timestamp 1753182340
transform 1 0 15568 0 1 29792
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0956_
timestamp 1751534193
transform -1 0 16240 0 1 31360
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _0957_
timestamp 1751740063
transform 1 0 17920 0 -1 29792
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__and2_2  _0958_
timestamp 1751889408
transform 1 0 19936 0 -1 29792
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__nor3_2  _0959_
timestamp 1753182340
transform 1 0 18704 0 -1 29792
box -86 -86 1318 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _0960_
timestamp 1751534193
transform 1 0 20720 0 -1 29792
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__xnor2_2  _0961_
timestamp 1753277515
transform 1 0 18704 0 1 29792
box -86 -86 1654 870
use gf180mcu_as_sc_mcu7t3v3__nor2_2  _0962_
timestamp 1751740063
transform 1 0 19040 0 1 31360
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _0963_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751632746
transform 1 0 16240 0 1 7840
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _0964_
timestamp 1751632746
transform 1 0 7840 0 1 15680
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _0965_
timestamp 1751632746
transform -1 0 9072 0 -1 15680
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _0966_
timestamp 1751632746
transform 1 0 1792 0 1 15680
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _0967_
timestamp 1751632746
transform 1 0 1568 0 -1 15680
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _0968_
timestamp 1751632746
transform 1 0 5376 0 -1 17248
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _0969_
timestamp 1751632746
transform 1 0 19376 0 -1 7840
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _0970_
timestamp 1751632746
transform 1 0 19488 0 -1 9408
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _0971_
timestamp 1751632746
transform -1 0 25200 0 1 10976
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _0972_
timestamp 1751632746
transform 1 0 23072 0 1 6272
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _0973_
timestamp 1751632746
transform 1 0 22960 0 1 4704
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _0974_
timestamp 1751632746
transform 1 0 19600 0 -1 4704
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _0975_
timestamp 1751632746
transform 1 0 26432 0 -1 4704
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _0976_
timestamp 1751632746
transform 1 0 31360 0 1 4704
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _0977_
timestamp 1751632746
transform 1 0 31360 0 1 6272
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _0978_
timestamp 1751632746
transform 1 0 26096 0 -1 6272
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _0979_
timestamp 1751632746
transform 1 0 29680 0 -1 9408
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _0980_
timestamp 1751632746
transform 1 0 25872 0 -1 10976
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _0981_
timestamp 1751632746
transform 1 0 31360 0 1 9408
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _0982_
timestamp 1751632746
transform 1 0 30352 0 1 12544
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _0983_
timestamp 1751632746
transform -1 0 34384 0 1 14112
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _0984_
timestamp 1751632746
transform -1 0 34384 0 1 17248
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _0985_
timestamp 1751632746
transform -1 0 34384 0 1 18816
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _0986_
timestamp 1751632746
transform 1 0 26992 0 -1 20384
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _0987_
timestamp 1751632746
transform 1 0 26544 0 -1 14112
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _0988_
timestamp 1751632746
transform 1 0 23072 0 1 12544
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _0989_
timestamp 1751632746
transform -1 0 28112 0 -1 17248
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _0990_
timestamp 1751632746
transform 1 0 25088 0 1 18816
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _0991_
timestamp 1751632746
transform -1 0 32704 0 -1 21952
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _0992_
timestamp 1751632746
transform 1 0 17024 0 1 9408
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _0993_
timestamp 1751632746
transform 1 0 11760 0 -1 14112
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _0994_
timestamp 1751632746
transform -1 0 12320 0 1 14112
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _0995_
timestamp 1751632746
transform 1 0 14000 0 -1 4704
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _0996_
timestamp 1751632746
transform 1 0 13776 0 1 4704
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _0997_
timestamp 1751632746
transform 1 0 1568 0 -1 4704
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _0998_
timestamp 1751632746
transform 1 0 23408 0 1 20384
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _0999_
timestamp 1751632746
transform 1 0 23072 0 1 21952
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1000_
timestamp 1751632746
transform 1 0 1568 0 -1 23520
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1001_
timestamp 1751632746
transform 1 0 1568 0 1 25088
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1002_
timestamp 1751632746
transform 1 0 2240 0 -1 26656
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1003_
timestamp 1751632746
transform -1 0 12880 0 -1 23520
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1004_
timestamp 1751632746
transform 1 0 7504 0 1 26656
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1005_
timestamp 1751632746
transform 1 0 5264 0 -1 26656
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1006_
timestamp 1751632746
transform 1 0 10080 0 1 25088
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1007_
timestamp 1751632746
transform 1 0 17248 0 -1 26656
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1008_
timestamp 1751632746
transform 1 0 23520 0 1 23520
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1009_
timestamp 1751632746
transform -1 0 29568 0 -1 23520
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1010_
timestamp 1751632746
transform -1 0 32032 0 1 25088
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1011_
timestamp 1751632746
transform 1 0 25088 0 1 26656
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1012_
timestamp 1751632746
transform -1 0 28784 0 1 29792
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1013_
timestamp 1751632746
transform 1 0 21840 0 -1 31360
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1014_
timestamp 1751632746
transform 1 0 21616 0 1 29792
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1015_
timestamp 1751632746
transform 1 0 21168 0 1 26656
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1016_
timestamp 1751632746
transform -1 0 21840 0 -1 25088
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1017_
timestamp 1751632746
transform 1 0 9408 0 -1 20384
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1018_
timestamp 1751632746
transform 1 0 9408 0 -1 17248
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1019_
timestamp 1751632746
transform 1 0 14000 0 -1 20384
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1020_
timestamp 1751632746
transform -1 0 17024 0 1 15680
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1021_
timestamp 1751632746
transform 1 0 21504 0 1 15680
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1022_
timestamp 1751632746
transform 1 0 19040 0 -1 15680
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1023_
timestamp 1751632746
transform 1 0 18816 0 -1 20384
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1024_
timestamp 1751632746
transform -1 0 24752 0 1 18816
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1025_
timestamp 1751632746
transform 1 0 14000 0 -1 23520
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1026_
timestamp 1751632746
transform -1 0 22736 0 -1 12544
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1027_
timestamp 1751632746
transform 1 0 9632 0 1 29792
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1028_
timestamp 1751632746
transform 1 0 9632 0 1 28224
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1029_
timestamp 1751632746
transform -1 0 14000 0 -1 31360
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1030_
timestamp 1751632746
transform 1 0 14000 0 -1 28224
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1031_
timestamp 1751632746
transform 1 0 14000 0 -1 31360
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1032_
timestamp 1751632746
transform -1 0 20944 0 1 28224
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__dfxtp_2  _1033_
timestamp 1751632746
transform -1 0 21392 0 -1 31360
box -86 -86 3110 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1034_
timestamp 1751534193
transform -1 0 20496 0 1 4704
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1035_
timestamp 1751534193
transform 1 0 25088 0 -1 4704
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  _1036_
timestamp 1751534193
transform 1 0 32928 0 -1 4704
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0511__A dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751532392
transform 1 0 14112 0 -1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0516__A
timestamp 1751532392
transform 1 0 14784 0 1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0554__A
timestamp 1751532392
transform -1 0 6272 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0619__B
timestamp 1751532392
transform -1 0 2912 0 1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0628__D
timestamp 1751532392
transform 1 0 3136 0 1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0642__A
timestamp 1751532392
transform -1 0 2912 0 1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0654__A
timestamp 1751532392
transform -1 0 14784 0 1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0673__A
timestamp 1751532392
transform 1 0 22848 0 -1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0680__A
timestamp 1751532392
transform -1 0 24080 0 1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0768__A
timestamp 1751532392
transform 1 0 20048 0 -1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0785__B
timestamp 1751532392
transform 1 0 26096 0 -1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0787__B
timestamp 1751532392
transform -1 0 23072 0 -1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0799__A
timestamp 1751532392
transform 1 0 15904 0 1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0801__A
timestamp 1751532392
transform -1 0 16576 0 -1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0832__C
timestamp 1751532392
transform 1 0 10864 0 1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0854__C
timestamp 1751532392
transform -1 0 9184 0 -1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0865__A
timestamp 1751532392
transform -1 0 23520 0 1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0869__A
timestamp 1751532392
transform 1 0 27104 0 -1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0873__A
timestamp 1751532392
transform 1 0 26656 0 -1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0964__CLK
timestamp 1751532392
transform 1 0 11088 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0965__CLK
timestamp 1751532392
transform 1 0 9632 0 -1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0966__CLK
timestamp 1751532392
transform 1 0 5040 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0967__CLK
timestamp 1751532392
transform 1 0 4816 0 -1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0968__CLK
timestamp 1751532392
transform -1 0 8848 0 -1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0969__CLK
timestamp 1751532392
transform 1 0 22848 0 1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0970__CLK
timestamp 1751532392
transform 1 0 23520 0 -1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0971__CLK
timestamp 1751532392
transform 1 0 24640 0 -1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0972__CLK
timestamp 1751532392
transform 1 0 26320 0 1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0973__CLK
timestamp 1751532392
transform 1 0 25872 0 -1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0974__CLK
timestamp 1751532392
transform -1 0 22848 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0975__CLK
timestamp 1751532392
transform 1 0 29680 0 -1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0976__CLK
timestamp 1751532392
transform -1 0 30800 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0977__CLK
timestamp 1751532392
transform 1 0 31136 0 1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0978__CLK
timestamp 1751532392
transform 1 0 30912 0 -1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0979__CLK
timestamp 1751532392
transform 1 0 30016 0 1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0980__CLK
timestamp 1751532392
transform 1 0 30128 0 1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0981__CLK
timestamp 1751532392
transform 1 0 31136 0 1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0982__CLK
timestamp 1751532392
transform 1 0 30240 0 -1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0983__CLK
timestamp 1751532392
transform 1 0 30352 0 1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0984__CLK
timestamp 1751532392
transform -1 0 31360 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0985__CLK
timestamp 1751532392
transform 1 0 31136 0 1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0986__CLK
timestamp 1751532392
transform 1 0 30016 0 1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0987__CLK
timestamp 1751532392
transform 1 0 29792 0 -1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0988__CLK
timestamp 1751532392
transform 1 0 26656 0 1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0989__CLK
timestamp 1751532392
transform -1 0 29456 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0991__CLK
timestamp 1751532392
transform 1 0 33152 0 -1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0996__D
timestamp 1751532392
transform -1 0 13776 0 1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__0997__CLK
timestamp 1751532392
transform -1 0 5824 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1000__CLK
timestamp 1751532392
transform 1 0 4928 0 1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1001__CLK
timestamp 1751532392
transform 1 0 5712 0 1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1002__CLK
timestamp 1751532392
transform 1 0 5712 0 1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1004__CLK
timestamp 1751532392
transform 1 0 10752 0 1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1005__CLK
timestamp 1751532392
transform 1 0 10416 0 -1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1006__CLK
timestamp 1751532392
transform 1 0 13104 0 -1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1009__CLK
timestamp 1751532392
transform 1 0 29792 0 -1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1010__CLK
timestamp 1751532392
transform 1 0 32256 0 1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1012__CLK
timestamp 1751532392
transform 1 0 29232 0 1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1017__CLK
timestamp 1751532392
transform 1 0 13776 0 -1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1018__CLK
timestamp 1751532392
transform 1 0 12432 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1021__CLK
timestamp 1751532392
transform 1 0 24752 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1022__CLK
timestamp 1751532392
transform 1 0 22288 0 -1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1026__CLK
timestamp 1751532392
transform 1 0 21952 0 1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1027__CLK
timestamp 1751532392
transform 1 0 12880 0 1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA__1028__CLK
timestamp 1751532392
transform 1 0 12880 0 1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_clkbuf_0_wb_clk_i_A
timestamp 1751532392
transform 1 0 17808 0 1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_clkbuf_3_0__f_wb_clk_i_A
timestamp 1751532392
transform 1 0 12432 0 -1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_clkbuf_3_1__f_wb_clk_i_A
timestamp 1751532392
transform 1 0 15232 0 -1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_clkbuf_3_2__f_wb_clk_i_A
timestamp 1751532392
transform -1 0 12096 0 -1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_clkbuf_3_3__f_wb_clk_i_A
timestamp 1751532392
transform -1 0 16128 0 -1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_clkbuf_3_4__f_wb_clk_i_A
timestamp 1751532392
transform -1 0 26432 0 1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_clkbuf_3_5__f_wb_clk_i_A
timestamp 1751532392
transform -1 0 29456 0 1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_clkbuf_3_6__f_wb_clk_i_A
timestamp 1751532392
transform 1 0 21840 0 -1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_clkbuf_3_7__f_wb_clk_i_A
timestamp 1751532392
transform 1 0 27664 0 1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_clkload0_A
timestamp 1751532392
transform 1 0 8960 0 -1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_clkload2_A
timestamp 1751532392
transform 1 0 9744 0 1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_clkload4_A
timestamp 1751532392
transform 1 0 24080 0 -1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_clkload5_A
timestamp 1751532392
transform 1 0 29680 0 1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_clkload6_A
timestamp 1751532392
transform 1 0 32032 0 1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__diode_2  ANTENNA_input1_A
timestamp 1751532392
transform -1 0 10864 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkbuf_0_wb_clk_i dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751661108
transform 1 0 18032 0 -1 18816
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkbuf_3_0__f_wb_clk_i
timestamp 1751661108
transform -1 0 12208 0 -1 15680
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkbuf_3_1__f_wb_clk_i
timestamp 1751661108
transform 1 0 12208 0 -1 12544
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkbuf_3_2__f_wb_clk_i
timestamp 1751661108
transform -1 0 12208 0 -1 25088
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkbuf_3_3__f_wb_clk_i
timestamp 1751661108
transform 1 0 13104 0 -1 25088
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkbuf_3_4__f_wb_clk_i
timestamp 1751661108
transform 1 0 25088 0 -1 12544
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkbuf_3_5__f_wb_clk_i
timestamp 1751661108
transform 1 0 27888 0 -1 12544
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkbuf_3_6__f_wb_clk_i
timestamp 1751661108
transform 1 0 22064 0 -1 23520
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkbuf_3_7__f_wb_clk_i
timestamp 1751661108
transform 1 0 29008 0 1 20384
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__inv_6  clkload0 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751896485
transform 1 0 7840 0 1 14112
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__inv_6  clkload1
timestamp 1751896485
transform 1 0 11984 0 1 12544
box -86 -86 1206 870
use gf180mcu_as_sc_mcu7t3v3__inv_4  clkload2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751633659
transform 1 0 8736 0 1 25088
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkload3
timestamp 1751661108
transform 1 0 13328 0 1 23520
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__inv_4  clkload4
timestamp 1751633659
transform 1 0 22848 0 -1 12544
box -86 -86 870 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_4  clkload5 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751558652
transform 1 0 27552 0 1 10976
box -86 -86 1094 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  clkload6
timestamp 1751661108
transform 1 0 29008 0 1 21952
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  fanout5
timestamp 1751534193
transform 1 0 24752 0 1 9408
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_0_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751532351
transform 1 0 1568 0 1 3136
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_0_18 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751532312
transform 1 0 3360 0 1 3136
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_0_33 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751532423
transform 1 0 5040 0 1 3136
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_0_36 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751532440
transform 1 0 5376 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_0_40
timestamp 1751532440
transform 1 0 5824 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_0_44
timestamp 1751532351
transform 1 0 6272 0 1 3136
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_0_60
timestamp 1751532312
transform 1 0 8064 0 1 3136
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_0_70
timestamp 1751532312
transform 1 0 9184 0 1 3136
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_0_78 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751532246
transform 1 0 10080 0 1 3136
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_0_82
timestamp 1751532423
transform 1 0 10528 0 1 3136
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_0_91
timestamp 1751532312
transform 1 0 11536 0 1 3136
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_0_99
timestamp 1751532440
transform 1 0 12432 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_0_101
timestamp 1751532423
transform 1 0 12656 0 1 3136
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_0_104
timestamp 1751532351
transform 1 0 12992 0 1 3136
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_0_120
timestamp 1751532351
transform 1 0 14784 0 1 3136
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_0_138
timestamp 1751532246
transform 1 0 16800 0 1 3136
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_0_142
timestamp 1751532440
transform 1 0 17248 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_0_144
timestamp 1751532423
transform 1 0 17472 0 1 3136
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_0_172
timestamp 1751532440
transform 1 0 20608 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_0_180
timestamp 1751532312
transform 1 0 21504 0 1 3136
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_0_188
timestamp 1751532440
transform 1 0 22400 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_0_192
timestamp 1751532246
transform 1 0 22848 0 1 3136
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_0_203
timestamp 1751532423
transform 1 0 24080 0 1 3136
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_0_206
timestamp 1751532246
transform 1 0 24416 0 1 3136
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_0_210
timestamp 1751532440
transform 1 0 24864 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_0_212
timestamp 1751532423
transform 1 0 25088 0 1 3136
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_0_240
timestamp 1751532440
transform 1 0 28224 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_0_249
timestamp 1751532312
transform 1 0 29232 0 1 3136
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_0_257
timestamp 1751532246
transform 1 0 30128 0 1 3136
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_0_270
timestamp 1751532440
transform 1 0 31584 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_0_287
timestamp 1751532312
transform 1 0 33488 0 1 3136
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_1_43
timestamp 1751532312
transform 1 0 6160 0 -1 4704
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_1_65
timestamp 1751532246
transform 1 0 8624 0 -1 4704
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_1_69
timestamp 1751532423
transform 1 0 9072 0 -1 4704
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_1_78
timestamp 1751532423
transform 1 0 10080 0 -1 4704
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_1_101
timestamp 1751532312
transform 1 0 12656 0 -1 4704
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_1_109
timestamp 1751532246
transform 1 0 13552 0 -1 4704
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_1_142
timestamp 1751532246
transform 1 0 17248 0 -1 4704
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_1_146
timestamp 1751532423
transform 1 0 17696 0 -1 4704
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_1_153
timestamp 1751532312
transform 1 0 18480 0 -1 4704
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_1_161
timestamp 1751532440
transform 1 0 19376 0 -1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_1_190
timestamp 1751532423
transform 1 0 22624 0 -1 4704
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_1_209
timestamp 1751532423
transform 1 0 24752 0 -1 4704
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_1_251
timestamp 1751532440
transform 1 0 29456 0 -1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_1_288
timestamp 1751532246
transform 1 0 33600 0 -1 4704
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_1_292
timestamp 1751532440
transform 1 0 34048 0 -1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_1_294
timestamp 1751532423
transform 1 0 34272 0 -1 4704
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_2_2
timestamp 1751532312
transform 1 0 1568 0 1 4704
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_2_10
timestamp 1751532423
transform 1 0 2464 0 1 4704
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_2_37
timestamp 1751532246
transform 1 0 5488 0 1 4704
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_2_41
timestamp 1751532440
transform 1 0 5936 0 1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_2_63
timestamp 1751532312
transform 1 0 8400 0 1 4704
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_2_71
timestamp 1751532246
transform 1 0 9296 0 1 4704
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_2_75
timestamp 1751532440
transform 1 0 9744 0 1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_2_102
timestamp 1751532440
transform 1 0 12768 0 1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_2_104
timestamp 1751532423
transform 1 0 12992 0 1 4704
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_2_107
timestamp 1751532440
transform 1 0 13328 0 1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_2_138
timestamp 1751532246
transform 1 0 16800 0 1 4704
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_2_142
timestamp 1751532440
transform 1 0 17248 0 1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_2_171
timestamp 1751532246
transform 1 0 20496 0 1 4704
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_2_192
timestamp 1751532423
transform 1 0 22848 0 1 4704
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_2_220
timestamp 1751532423
transform 1 0 25984 0 1 4704
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_2_254
timestamp 1751532440
transform 1 0 29792 0 1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_2_256
timestamp 1751532423
transform 1 0 30016 0 1 4704
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_3_2
timestamp 1751532246
transform 1 0 1568 0 -1 6272
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_3_6
timestamp 1751532440
transform 1 0 2016 0 -1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_3_25
timestamp 1751532246
transform 1 0 4144 0 -1 6272
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_3_29
timestamp 1751532423
transform 1 0 4592 0 -1 6272
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_3_37
timestamp 1751532423
transform 1 0 5488 0 -1 6272
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_3_48
timestamp 1751532440
transform 1 0 6720 0 -1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_3_62
timestamp 1751532312
transform 1 0 8288 0 -1 6272
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_3_72
timestamp 1751532312
transform 1 0 9408 0 -1 6272
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_3_80
timestamp 1751532423
transform 1 0 10304 0 -1 6272
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_3_87
timestamp 1751532423
transform 1 0 11088 0 -1 6272
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_3_98
timestamp 1751532423
transform 1 0 12320 0 -1 6272
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_3_109
timestamp 1751532312
transform 1 0 13552 0 -1 6272
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_3_117
timestamp 1751532440
transform 1 0 14448 0 -1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_3_123
timestamp 1751532440
transform 1 0 15120 0 -1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_3_131
timestamp 1751532440
transform 1 0 16016 0 -1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_3_168
timestamp 1751532351
transform 1 0 20160 0 -1 6272
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_3_184
timestamp 1751532440
transform 1 0 21952 0 -1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_3_216
timestamp 1751532440
transform 1 0 25536 0 -1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_3_218
timestamp 1751532423
transform 1 0 25760 0 -1 6272
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_3_262
timestamp 1751532440
transform 1 0 30688 0 -1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_3_266
timestamp 1751532440
transform 1 0 31136 0 -1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_3_279
timestamp 1751532423
transform 1 0 32592 0 -1 6272
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_3_289
timestamp 1751532246
transform 1 0 33712 0 -1 6272
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_3_293
timestamp 1751532440
transform 1 0 34160 0 -1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_4_2
timestamp 1751532312
transform 1 0 1568 0 1 6272
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_4_10
timestamp 1751532440
transform 1 0 2464 0 1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_4_43
timestamp 1751532312
transform 1 0 6160 0 1 6272
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_4_51
timestamp 1751532440
transform 1 0 7056 0 1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_4_69
timestamp 1751532351
transform 1 0 9072 0 1 6272
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_4_85
timestamp 1751532423
transform 1 0 10864 0 1 6272
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_4_96
timestamp 1751532312
transform 1 0 12096 0 1 6272
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_4_104
timestamp 1751532423
transform 1 0 12992 0 1 6272
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_4_114
timestamp 1751532440
transform 1 0 14112 0 1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_4_123
timestamp 1751532440
transform 1 0 15120 0 1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_4_158
timestamp 1751532351
transform 1 0 19040 0 1 6272
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_4_174
timestamp 1751532423
transform 1 0 20832 0 1 6272
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_4_177
timestamp 1751532246
transform 1 0 21168 0 1 6272
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_4_181
timestamp 1751532440
transform 1 0 21616 0 1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_4_183
timestamp 1751532423
transform 1 0 21840 0 1 6272
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_4_190
timestamp 1751532440
transform 1 0 22624 0 1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_4_221
timestamp 1751532440
transform 1 0 26096 0 1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_4_225
timestamp 1751532312
transform 1 0 26544 0 1 6272
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_4_233
timestamp 1751532246
transform 1 0 27440 0 1 6272
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_4_244
timestamp 1751532423
transform 1 0 28672 0 1 6272
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_4_247
timestamp 1751532440
transform 1 0 29008 0 1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_4_249
timestamp 1751532423
transform 1 0 29232 0 1 6272
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_4_264
timestamp 1751532440
transform 1 0 30912 0 1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_5_2
timestamp 1751532312
transform 1 0 1568 0 -1 7840
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_5_10
timestamp 1751532440
transform 1 0 2464 0 -1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_5_12
timestamp 1751532423
transform 1 0 2688 0 -1 7840
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_5_23
timestamp 1751532351
transform 1 0 3920 0 -1 7840
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_5_39
timestamp 1751532312
transform 1 0 5712 0 -1 7840
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_5_47
timestamp 1751532246
transform 1 0 6608 0 -1 7840
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_5_51
timestamp 1751532423
transform 1 0 7056 0 -1 7840
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_5_59
timestamp 1751532312
transform 1 0 7952 0 -1 7840
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_5_67
timestamp 1751532440
transform 1 0 8848 0 -1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_5_69
timestamp 1751532423
transform 1 0 9072 0 -1 7840
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_5_72
timestamp 1751532440
transform 1 0 9408 0 -1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_5_74
timestamp 1751532423
transform 1 0 9632 0 -1 7840
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_5_85
timestamp 1751532440
transform 1 0 10864 0 -1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_5_108
timestamp 1751532246
transform 1 0 13440 0 -1 7840
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_5_133
timestamp 1751532246
transform 1 0 16240 0 -1 7840
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_5_137
timestamp 1751532440
transform 1 0 16688 0 -1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_5_139
timestamp 1751532423
transform 1 0 16912 0 -1 7840
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_5_142
timestamp 1751532351
transform 1 0 17248 0 -1 7840
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_5_158
timestamp 1751532440
transform 1 0 19040 0 -1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_5_160
timestamp 1751532423
transform 1 0 19264 0 -1 7840
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_5_188
timestamp 1751532440
transform 1 0 22400 0 -1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_5_190
timestamp 1751532423
transform 1 0 22624 0 -1 7840
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_5_208
timestamp 1751532440
transform 1 0 24640 0 -1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_5_212
timestamp 1751532312
transform 1 0 25088 0 -1 7840
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_5_220
timestamp 1751532246
transform 1 0 25984 0 -1 7840
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_5_224
timestamp 1751532440
transform 1 0 26432 0 -1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_5_226
timestamp 1751532423
transform 1 0 26656 0 -1 7840
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_5_234
timestamp 1751532312
transform 1 0 27552 0 -1 7840
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_5_242
timestamp 1751532246
transform 1 0 28448 0 -1 7840
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_5_246
timestamp 1751532440
transform 1 0 28896 0 -1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_5_248
timestamp 1751532423
transform 1 0 29120 0 -1 7840
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_5_256
timestamp 1751532312
transform 1 0 30016 0 -1 7840
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_5_264
timestamp 1751532246
transform 1 0 30912 0 -1 7840
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_5_268
timestamp 1751532423
transform 1 0 31360 0 -1 7840
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_5_276
timestamp 1751532246
transform 1 0 32256 0 -1 7840
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_5_288
timestamp 1751532246
transform 1 0 33600 0 -1 7840
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_5_292
timestamp 1751532440
transform 1 0 34048 0 -1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_5_294
timestamp 1751532423
transform 1 0 34272 0 -1 7840
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_6_2
timestamp 1751532312
transform 1 0 1568 0 1 7840
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_6_10
timestamp 1751532246
transform 1 0 2464 0 1 7840
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_6_31
timestamp 1751532246
transform 1 0 4816 0 1 7840
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_6_37
timestamp 1751532312
transform 1 0 5488 0 1 7840
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_6_45
timestamp 1751532246
transform 1 0 6384 0 1 7840
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_6_55
timestamp 1751532440
transform 1 0 7504 0 1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_6_82
timestamp 1751532246
transform 1 0 10528 0 1 7840
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_6_114
timestamp 1751532246
transform 1 0 14112 0 1 7840
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_6_118
timestamp 1751532440
transform 1 0 14560 0 1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_6_120
timestamp 1751532423
transform 1 0 14784 0 1 7840
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_6_160
timestamp 1751532312
transform 1 0 19264 0 1 7840
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_6_168
timestamp 1751532246
transform 1 0 20160 0 1 7840
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_6_172
timestamp 1751532440
transform 1 0 20608 0 1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_6_174
timestamp 1751532423
transform 1 0 20832 0 1 7840
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_6_184
timestamp 1751532440
transform 1 0 21952 0 1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_6_186
timestamp 1751532423
transform 1 0 22176 0 1 7840
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_6_208
timestamp 1751532351
transform 1 0 24640 0 1 7840
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_6_224
timestamp 1751532312
transform 1 0 26432 0 1 7840
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_6_238
timestamp 1751532423
transform 1 0 28000 0 1 7840
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_6_254
timestamp 1751532440
transform 1 0 29792 0 1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_6_258
timestamp 1751532312
transform 1 0 30240 0 1 7840
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_6_268
timestamp 1751532440
transform 1 0 31360 0 1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_6_270
timestamp 1751532423
transform 1 0 31584 0 1 7840
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_6_275
timestamp 1751532351
transform 1 0 32144 0 1 7840
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_6_291
timestamp 1751532246
transform 1 0 33936 0 1 7840
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_7_2
timestamp 1751532312
transform 1 0 1568 0 -1 9408
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_7_10
timestamp 1751532440
transform 1 0 2464 0 -1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_7_22
timestamp 1751532423
transform 1 0 3808 0 -1 9408
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_7_30
timestamp 1751532312
transform 1 0 4704 0 -1 9408
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_7_38
timestamp 1751532423
transform 1 0 5600 0 -1 9408
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_7_49
timestamp 1751532440
transform 1 0 6832 0 -1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_7_68
timestamp 1751532440
transform 1 0 8960 0 -1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_7_72
timestamp 1751532312
transform 1 0 9408 0 -1 9408
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_7_80
timestamp 1751532246
transform 1 0 10304 0 -1 9408
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_7_84
timestamp 1751532440
transform 1 0 10752 0 -1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_7_86
timestamp 1751532423
transform 1 0 10976 0 -1 9408
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_7_91
timestamp 1751532246
transform 1 0 11536 0 -1 9408
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_7_112
timestamp 1751532440
transform 1 0 13888 0 -1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_7_133
timestamp 1751532246
transform 1 0 16240 0 -1 9408
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_7_137
timestamp 1751532440
transform 1 0 16688 0 -1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_7_139
timestamp 1751532423
transform 1 0 16912 0 -1 9408
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_7_142
timestamp 1751532351
transform 1 0 17248 0 -1 9408
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_7_158
timestamp 1751532246
transform 1 0 19040 0 -1 9408
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_7_196
timestamp 1751532440
transform 1 0 23296 0 -1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_7_200
timestamp 1751532312
transform 1 0 23744 0 -1 9408
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_7_208
timestamp 1751532440
transform 1 0 24640 0 -1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_7_219
timestamp 1751532351
transform 1 0 25872 0 -1 9408
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_7_235
timestamp 1751532423
transform 1 0 27664 0 -1 9408
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_7_288
timestamp 1751532246
transform 1 0 33600 0 -1 9408
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_7_292
timestamp 1751532440
transform 1 0 34048 0 -1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_7_294
timestamp 1751532423
transform 1 0 34272 0 -1 9408
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_8_2
timestamp 1751532312
transform 1 0 1568 0 1 9408
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_8_10
timestamp 1751532440
transform 1 0 2464 0 1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_8_32
timestamp 1751532440
transform 1 0 4928 0 1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_8_34
timestamp 1751532423
transform 1 0 5152 0 1 9408
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_8_44
timestamp 1751532246
transform 1 0 6272 0 1 9408
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_8_48
timestamp 1751532440
transform 1 0 6720 0 1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_8_50
timestamp 1751532423
transform 1 0 6944 0 1 9408
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_8_65
timestamp 1751532351
transform 1 0 8624 0 1 9408
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_8_102
timestamp 1751532440
transform 1 0 12768 0 1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_8_104
timestamp 1751532423
transform 1 0 12992 0 1 9408
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_8_107
timestamp 1751532351
transform 1 0 13328 0 1 9408
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_8_123
timestamp 1751532440
transform 1 0 15120 0 1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_8_136
timestamp 1751532246
transform 1 0 16576 0 1 9408
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_8_167
timestamp 1751532312
transform 1 0 20048 0 1 9408
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_8_177
timestamp 1751532246
transform 1 0 21168 0 1 9408
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_8_199
timestamp 1751532440
transform 1 0 23632 0 1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_8_203
timestamp 1751532246
transform 1 0 24080 0 1 9408
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_8_207
timestamp 1751532440
transform 1 0 24528 0 1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_8_229
timestamp 1751532423
transform 1 0 26992 0 1 9408
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_8_265
timestamp 1751532440
transform 1 0 31024 0 1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_8_267
timestamp 1751532423
transform 1 0 31248 0 1 9408
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_9_2
timestamp 1751532312
transform 1 0 1568 0 -1 10976
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_9_43
timestamp 1751532312
transform 1 0 6160 0 -1 10976
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_9_51
timestamp 1751532440
transform 1 0 7056 0 -1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_9_53
timestamp 1751532423
transform 1 0 7280 0 -1 10976
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_9_64
timestamp 1751532246
transform 1 0 8512 0 -1 10976
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_9_68
timestamp 1751532440
transform 1 0 8960 0 -1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_9_72
timestamp 1751532423
transform 1 0 9408 0 -1 10976
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_9_79
timestamp 1751532351
transform 1 0 10192 0 -1 10976
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_9_99
timestamp 1751532423
transform 1 0 12432 0 -1 10976
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_9_113
timestamp 1751532440
transform 1 0 14000 0 -1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_9_122
timestamp 1751532351
transform 1 0 15008 0 -1 10976
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_9_138
timestamp 1751532440
transform 1 0 16800 0 -1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_9_142
timestamp 1751532351
transform 1 0 17248 0 -1 10976
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_9_158
timestamp 1751532312
transform 1 0 19040 0 -1 10976
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_9_166
timestamp 1751532246
transform 1 0 19936 0 -1 10976
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_9_170
timestamp 1751532440
transform 1 0 20384 0 -1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_9_172
timestamp 1751532423
transform 1 0 20608 0 -1 10976
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_9_179
timestamp 1751532312
transform 1 0 21392 0 -1 10976
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_9_187
timestamp 1751532440
transform 1 0 22288 0 -1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_9_189
timestamp 1751532423
transform 1 0 22512 0 -1 10976
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_9_204
timestamp 1751532246
transform 1 0 24192 0 -1 10976
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_9_260
timestamp 1751532440
transform 1 0 30464 0 -1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_9_289
timestamp 1751532246
transform 1 0 33712 0 -1 10976
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_9_293
timestamp 1751532440
transform 1 0 34160 0 -1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_10_2
timestamp 1751532312
transform 1 0 1568 0 1 10976
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_10_10
timestamp 1751532246
transform 1 0 2464 0 1 10976
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_10_14
timestamp 1751532440
transform 1 0 2912 0 1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_10_28
timestamp 1751532246
transform 1 0 4480 0 1 10976
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_10_32
timestamp 1751532440
transform 1 0 4928 0 1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_10_34
timestamp 1751532423
transform 1 0 5152 0 1 10976
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_10_37
timestamp 1751532312
transform 1 0 5488 0 1 10976
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_10_45
timestamp 1751532246
transform 1 0 6384 0 1 10976
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_10_60
timestamp 1751532246
transform 1 0 8064 0 1 10976
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_10_64
timestamp 1751532440
transform 1 0 8512 0 1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_10_83
timestamp 1751532423
transform 1 0 10640 0 1 10976
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_10_91
timestamp 1751532423
transform 1 0 11536 0 1 10976
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_10_104
timestamp 1751532423
transform 1 0 12992 0 1 10976
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_10_111
timestamp 1751532423
transform 1 0 13776 0 1 10976
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_10_118
timestamp 1751532440
transform 1 0 14560 0 1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_10_140
timestamp 1751532246
transform 1 0 17024 0 1 10976
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_10_151
timestamp 1751532440
transform 1 0 18256 0 1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_10_159
timestamp 1751532351
transform 1 0 19152 0 1 10976
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_10_177
timestamp 1751532246
transform 1 0 21168 0 1 10976
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_10_181
timestamp 1751532440
transform 1 0 21616 0 1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_10_183
timestamp 1751532423
transform 1 0 21840 0 1 10976
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_10_220
timestamp 1751532440
transform 1 0 25984 0 1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_10_224
timestamp 1751532440
transform 1 0 26432 0 1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_10_243
timestamp 1751532440
transform 1 0 28560 0 1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_10_247
timestamp 1751532440
transform 1 0 29008 0 1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_10_251
timestamp 1751532440
transform 1 0 29456 0 1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_10_255
timestamp 1751532440
transform 1 0 29904 0 1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_10_259
timestamp 1751532312
transform 1 0 30352 0 1 10976
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_10_267
timestamp 1751532246
transform 1 0 31248 0 1 10976
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_10_271
timestamp 1751532423
transform 1 0 31696 0 1 10976
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_10_286
timestamp 1751532312
transform 1 0 33376 0 1 10976
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_10_294
timestamp 1751532423
transform 1 0 34272 0 1 10976
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_11_2
timestamp 1751532312
transform 1 0 1568 0 -1 12544
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_11_10
timestamp 1751532423
transform 1 0 2464 0 -1 12544
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_11_40
timestamp 1751532440
transform 1 0 5824 0 -1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_11_42
timestamp 1751532423
transform 1 0 6048 0 -1 12544
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_11_53
timestamp 1751532423
transform 1 0 7280 0 -1 12544
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_11_68
timestamp 1751532440
transform 1 0 8960 0 -1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_11_72
timestamp 1751532246
transform 1 0 9408 0 -1 12544
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_11_76
timestamp 1751532423
transform 1 0 9856 0 -1 12544
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_11_122
timestamp 1751532440
transform 1 0 15008 0 -1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_11_126
timestamp 1751532246
transform 1 0 15456 0 -1 12544
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_11_160
timestamp 1751532246
transform 1 0 19264 0 -1 12544
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_11_191
timestamp 1751532423
transform 1 0 22736 0 -1 12544
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_11_262
timestamp 1751532440
transform 1 0 30688 0 -1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_11_264
timestamp 1751532423
transform 1 0 30912 0 -1 12544
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_11_276
timestamp 1751532246
transform 1 0 32256 0 -1 12544
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_11_282
timestamp 1751532312
transform 1 0 32928 0 -1 12544
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_11_290
timestamp 1751532246
transform 1 0 33824 0 -1 12544
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_11_294
timestamp 1751532423
transform 1 0 34272 0 -1 12544
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_12_2
timestamp 1751532246
transform 1 0 1568 0 1 12544
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_12_6
timestamp 1751532423
transform 1 0 2016 0 1 12544
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_12_65
timestamp 1751532312
transform 1 0 8624 0 1 12544
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_12_83
timestamp 1751532440
transform 1 0 10640 0 1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_12_92
timestamp 1751532440
transform 1 0 11648 0 1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_12_94
timestamp 1751532423
transform 1 0 11872 0 1 12544
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_12_117
timestamp 1751532440
transform 1 0 14448 0 1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_12_119
timestamp 1751532423
transform 1 0 14672 0 1 12544
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_12_140
timestamp 1751532440
transform 1 0 17024 0 1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_12_166
timestamp 1751532312
transform 1 0 19936 0 1 12544
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_12_174
timestamp 1751532423
transform 1 0 20832 0 1 12544
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_12_177
timestamp 1751532440
transform 1 0 21168 0 1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_12_193
timestamp 1751532423
transform 1 0 22960 0 1 12544
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_12_221
timestamp 1751532440
transform 1 0 26096 0 1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_12_223
timestamp 1751532423
transform 1 0 26320 0 1 12544
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_12_231
timestamp 1751532440
transform 1 0 27216 0 1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_12_293
timestamp 1751532440
transform 1 0 34160 0 1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_13_2
timestamp 1751532312
transform 1 0 1568 0 -1 14112
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_13_37
timestamp 1751532351
transform 1 0 5488 0 -1 14112
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_13_53
timestamp 1751532312
transform 1 0 7280 0 -1 14112
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_13_61
timestamp 1751532246
transform 1 0 8176 0 -1 14112
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_13_65
timestamp 1751532440
transform 1 0 8624 0 -1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_13_67
timestamp 1751532423
transform 1 0 8848 0 -1 14112
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_13_72
timestamp 1751532440
transform 1 0 9408 0 -1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_13_76
timestamp 1751532351
transform 1 0 9856 0 -1 14112
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_13_92
timestamp 1751532423
transform 1 0 11648 0 -1 14112
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_13_126
timestamp 1751532246
transform 1 0 15456 0 -1 14112
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_13_159
timestamp 1751532351
transform 1 0 19152 0 -1 14112
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_13_175
timestamp 1751532423
transform 1 0 20944 0 -1 14112
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_13_189
timestamp 1751532440
transform 1 0 22512 0 -1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_13_191
timestamp 1751532423
transform 1 0 22736 0 -1 14112
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_13_201
timestamp 1751532440
transform 1 0 23856 0 -1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_13_205
timestamp 1751532246
transform 1 0 24304 0 -1 14112
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_13_209
timestamp 1751532423
transform 1 0 24752 0 -1 14112
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_13_252
timestamp 1751532440
transform 1 0 29568 0 -1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_13_256
timestamp 1751532440
transform 1 0 30016 0 -1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_13_260
timestamp 1751532440
transform 1 0 30464 0 -1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_13_288
timestamp 1751532246
transform 1 0 33600 0 -1 14112
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_13_292
timestamp 1751532440
transform 1 0 34048 0 -1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_13_294
timestamp 1751532423
transform 1 0 34272 0 -1 14112
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_14_2
timestamp 1751532312
transform 1 0 1568 0 1 14112
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_14_10
timestamp 1751532440
transform 1 0 2464 0 1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_14_12
timestamp 1751532423
transform 1 0 2688 0 1 14112
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_14_19
timestamp 1751532351
transform 1 0 3472 0 1 14112
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_14_37
timestamp 1751532312
transform 1 0 5488 0 1 14112
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_14_57
timestamp 1751532423
transform 1 0 7728 0 1 14112
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_14_68
timestamp 1751532440
transform 1 0 8960 0 1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_14_70
timestamp 1751532423
transform 1 0 9184 0 1 14112
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_14_98
timestamp 1751532246
transform 1 0 12320 0 1 14112
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_14_102
timestamp 1751532440
transform 1 0 12768 0 1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_14_104
timestamp 1751532423
transform 1 0 12992 0 1 14112
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_14_107
timestamp 1751532312
transform 1 0 13328 0 1 14112
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_14_115
timestamp 1751532440
transform 1 0 14224 0 1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_14_117
timestamp 1751532423
transform 1 0 14448 0 1 14112
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_14_120
timestamp 1751532351
transform 1 0 14784 0 1 14112
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_14_136
timestamp 1751532312
transform 1 0 16576 0 1 14112
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_14_144
timestamp 1751532440
transform 1 0 17472 0 1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_14_146
timestamp 1751532423
transform 1 0 17696 0 1 14112
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_14_153
timestamp 1751532351
transform 1 0 18480 0 1 14112
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_14_169
timestamp 1751532246
transform 1 0 20272 0 1 14112
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_14_173
timestamp 1751532440
transform 1 0 20720 0 1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_14_177
timestamp 1751532351
transform 1 0 21168 0 1 14112
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_14_193
timestamp 1751532351
transform 1 0 22960 0 1 14112
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_14_209
timestamp 1751532246
transform 1 0 24752 0 1 14112
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_14_213
timestamp 1751532440
transform 1 0 25200 0 1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_14_215
timestamp 1751532423
transform 1 0 25424 0 1 14112
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_14_230
timestamp 1751532440
transform 1 0 27104 0 1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_14_243
timestamp 1751532440
transform 1 0 28560 0 1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_14_254
timestamp 1751532246
transform 1 0 29792 0 1 14112
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_14_258
timestamp 1751532423
transform 1 0 30240 0 1 14112
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_15_29
timestamp 1751532440
transform 1 0 4592 0 -1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_15_33
timestamp 1751532312
transform 1 0 5040 0 -1 15680
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_15_41
timestamp 1751532423
transform 1 0 5936 0 -1 15680
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_15_69
timestamp 1751532423
transform 1 0 9072 0 -1 15680
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_15_97
timestamp 1751532440
transform 1 0 12208 0 -1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_15_101
timestamp 1751532312
transform 1 0 12656 0 -1 15680
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_15_109
timestamp 1751532246
transform 1 0 13552 0 -1 15680
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_15_113
timestamp 1751532440
transform 1 0 14000 0 -1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_15_115
timestamp 1751532423
transform 1 0 14224 0 -1 15680
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_15_126
timestamp 1751532312
transform 1 0 15456 0 -1 15680
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_15_142
timestamp 1751532440
transform 1 0 17248 0 -1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_15_154
timestamp 1751532246
transform 1 0 18592 0 -1 15680
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_15_185
timestamp 1751532440
transform 1 0 22064 0 -1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_15_189
timestamp 1751532351
transform 1 0 22512 0 -1 15680
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_15_205
timestamp 1751532246
transform 1 0 24304 0 -1 15680
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_15_209
timestamp 1751532423
transform 1 0 24752 0 -1 15680
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_15_212
timestamp 1751532351
transform 1 0 25088 0 -1 15680
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_15_228
timestamp 1751532440
transform 1 0 26880 0 -1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_15_250
timestamp 1751532246
transform 1 0 29344 0 -1 15680
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_15_254
timestamp 1751532440
transform 1 0 29792 0 -1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_15_256
timestamp 1751532423
transform 1 0 30016 0 -1 15680
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_15_263
timestamp 1751532246
transform 1 0 30800 0 -1 15680
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_15_267
timestamp 1751532440
transform 1 0 31248 0 -1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_15_276
timestamp 1751532246
transform 1 0 32256 0 -1 15680
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_15_282
timestamp 1751532312
transform 1 0 32928 0 -1 15680
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_15_290
timestamp 1751532246
transform 1 0 33824 0 -1 15680
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_15_294
timestamp 1751532423
transform 1 0 34272 0 -1 15680
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_16_2
timestamp 1751532440
transform 1 0 1568 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_16_31
timestamp 1751532440
transform 1 0 4816 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_16_37
timestamp 1751532351
transform 1 0 5488 0 1 15680
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_16_53
timestamp 1751532246
transform 1 0 7280 0 1 15680
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_16_57
timestamp 1751532423
transform 1 0 7728 0 1 15680
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_16_85
timestamp 1751532440
transform 1 0 10864 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_16_89
timestamp 1751532312
transform 1 0 11312 0 1 15680
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_16_97
timestamp 1751532440
transform 1 0 12208 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_16_101
timestamp 1751532246
transform 1 0 12656 0 1 15680
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_16_107
timestamp 1751532246
transform 1 0 13328 0 1 15680
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_16_111
timestamp 1751532440
transform 1 0 13776 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_16_140
timestamp 1751532312
transform 1 0 17024 0 1 15680
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_16_148
timestamp 1751532246
transform 1 0 17920 0 1 15680
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_16_152
timestamp 1751532440
transform 1 0 18368 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_16_154
timestamp 1751532423
transform 1 0 18592 0 1 15680
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_16_168
timestamp 1751532246
transform 1 0 20160 0 1 15680
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_16_172
timestamp 1751532440
transform 1 0 20608 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_16_174
timestamp 1751532423
transform 1 0 20832 0 1 15680
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_16_177
timestamp 1751532440
transform 1 0 21168 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_16_179
timestamp 1751532423
transform 1 0 21392 0 1 15680
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_16_207
timestamp 1751532440
transform 1 0 24528 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_16_211
timestamp 1751532312
transform 1 0 24976 0 1 15680
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_16_219
timestamp 1751532440
transform 1 0 25872 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_16_247
timestamp 1751532440
transform 1 0 29008 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_16_251
timestamp 1751532312
transform 1 0 29456 0 1 15680
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_16_259
timestamp 1751532246
transform 1 0 30352 0 1 15680
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_16_263
timestamp 1751532440
transform 1 0 30800 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_16_265
timestamp 1751532423
transform 1 0 31024 0 1 15680
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_16_268
timestamp 1751532423
transform 1 0 31360 0 1 15680
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_16_279
timestamp 1751532351
transform 1 0 32592 0 1 15680
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_17_2
timestamp 1751532351
transform 1 0 1568 0 -1 17248
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_17_18
timestamp 1751532246
transform 1 0 3360 0 -1 17248
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_17_22
timestamp 1751532423
transform 1 0 3808 0 -1 17248
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_17_35
timestamp 1751532423
transform 1 0 5264 0 -1 17248
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_17_63
timestamp 1751532440
transform 1 0 8400 0 -1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_17_67
timestamp 1751532440
transform 1 0 8848 0 -1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_17_69
timestamp 1751532423
transform 1 0 9072 0 -1 17248
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_17_113
timestamp 1751532246
transform 1 0 14000 0 -1 17248
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_17_117
timestamp 1751532423
transform 1 0 14448 0 -1 17248
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_17_131
timestamp 1751532312
transform 1 0 16016 0 -1 17248
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_17_139
timestamp 1751532423
transform 1 0 16912 0 -1 17248
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_17_142
timestamp 1751532440
transform 1 0 17248 0 -1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_17_144
timestamp 1751532423
transform 1 0 17472 0 -1 17248
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_17_171
timestamp 1751532440
transform 1 0 20496 0 -1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_17_201
timestamp 1751532312
transform 1 0 23856 0 -1 17248
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_17_209
timestamp 1751532423
transform 1 0 24752 0 -1 17248
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_17_261
timestamp 1751532423
transform 1 0 30576 0 -1 17248
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_17_277
timestamp 1751532440
transform 1 0 32368 0 -1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_17_279
timestamp 1751532423
transform 1 0 32592 0 -1 17248
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_17_289
timestamp 1751532246
transform 1 0 33712 0 -1 17248
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_17_293
timestamp 1751532440
transform 1 0 34160 0 -1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_18_2
timestamp 1751532312
transform 1 0 1568 0 1 17248
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_18_10
timestamp 1751532246
transform 1 0 2464 0 1 17248
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_18_33
timestamp 1751532440
transform 1 0 5040 0 1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_18_44
timestamp 1751532246
transform 1 0 6272 0 1 17248
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_18_48
timestamp 1751532423
transform 1 0 6720 0 1 17248
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_18_60
timestamp 1751532351
transform 1 0 8064 0 1 17248
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_18_76
timestamp 1751532246
transform 1 0 9856 0 1 17248
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_18_86
timestamp 1751532423
transform 1 0 10976 0 1 17248
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_18_103
timestamp 1751532440
transform 1 0 12880 0 1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_18_107
timestamp 1751532423
transform 1 0 13328 0 1 17248
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_18_133
timestamp 1751532246
transform 1 0 16240 0 1 17248
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_18_137
timestamp 1751532423
transform 1 0 16688 0 1 17248
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_18_144
timestamp 1751532440
transform 1 0 17472 0 1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_18_146
timestamp 1751532423
transform 1 0 17696 0 1 17248
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_18_149
timestamp 1751532440
transform 1 0 18032 0 1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_18_151
timestamp 1751532423
transform 1 0 18256 0 1 17248
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_18_177
timestamp 1751532246
transform 1 0 21168 0 1 17248
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_18_181
timestamp 1751532440
transform 1 0 21616 0 1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_18_197
timestamp 1751532351
transform 1 0 23408 0 1 17248
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_18_213
timestamp 1751532312
transform 1 0 25200 0 1 17248
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_18_221
timestamp 1751532246
transform 1 0 26096 0 1 17248
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_18_243
timestamp 1751532440
transform 1 0 28560 0 1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_19_2
timestamp 1751532312
transform 1 0 1568 0 -1 18816
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_19_10
timestamp 1751532246
transform 1 0 2464 0 -1 18816
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_19_14
timestamp 1751532440
transform 1 0 2912 0 -1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_19_37
timestamp 1751532246
transform 1 0 5488 0 -1 18816
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_19_41
timestamp 1751532440
transform 1 0 5936 0 -1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_19_69
timestamp 1751532423
transform 1 0 9072 0 -1 18816
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_19_72
timestamp 1751532351
transform 1 0 9408 0 -1 18816
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_19_88
timestamp 1751532312
transform 1 0 11200 0 -1 18816
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_19_96
timestamp 1751532423
transform 1 0 12096 0 -1 18816
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_19_136
timestamp 1751532246
transform 1 0 16576 0 -1 18816
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_19_194
timestamp 1751532351
transform 1 0 23072 0 -1 18816
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_19_212
timestamp 1751532351
transform 1 0 25088 0 -1 18816
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_19_250
timestamp 1751532440
transform 1 0 29344 0 -1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_19_259
timestamp 1751532423
transform 1 0 30352 0 -1 18816
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_19_278
timestamp 1751532440
transform 1 0 32480 0 -1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_19_286
timestamp 1751532312
transform 1 0 33376 0 -1 18816
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_19_294
timestamp 1751532423
transform 1 0 34272 0 -1 18816
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_20_2
timestamp 1751532246
transform 1 0 1568 0 1 18816
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_20_6
timestamp 1751532440
transform 1 0 2016 0 1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_20_8
timestamp 1751532423
transform 1 0 2240 0 1 18816
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_20_34
timestamp 1751532423
transform 1 0 5152 0 1 18816
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_20_47
timestamp 1751532423
transform 1 0 6608 0 1 18816
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_20_72
timestamp 1751532312
transform 1 0 9408 0 1 18816
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_20_80
timestamp 1751532423
transform 1 0 10304 0 1 18816
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_20_94
timestamp 1751532423
transform 1 0 11872 0 1 18816
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_20_114
timestamp 1751532423
transform 1 0 14112 0 1 18816
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_20_127
timestamp 1751532246
transform 1 0 15568 0 1 18816
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_20_155
timestamp 1751532246
transform 1 0 18704 0 1 18816
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_20_172
timestamp 1751532440
transform 1 0 20608 0 1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_20_174
timestamp 1751532423
transform 1 0 20832 0 1 18816
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_20_181
timestamp 1751532423
transform 1 0 21616 0 1 18816
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_20_209
timestamp 1751532440
transform 1 0 24752 0 1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_20_211
timestamp 1751532423
transform 1 0 24976 0 1 18816
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_20_239
timestamp 1751532246
transform 1 0 28112 0 1 18816
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_20_243
timestamp 1751532440
transform 1 0 28560 0 1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_20_254
timestamp 1751532440
transform 1 0 29792 0 1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_20_258
timestamp 1751532312
transform 1 0 30240 0 1 18816
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_21_2
timestamp 1751532312
transform 1 0 1568 0 -1 20384
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_21_10
timestamp 1751532246
transform 1 0 2464 0 -1 20384
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_21_44
timestamp 1751532246
transform 1 0 6272 0 -1 20384
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_21_69
timestamp 1751532423
transform 1 0 9072 0 -1 20384
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_21_109
timestamp 1751532440
transform 1 0 13552 0 -1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_21_142
timestamp 1751532246
transform 1 0 17248 0 -1 20384
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_21_153
timestamp 1751532440
transform 1 0 18480 0 -1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_21_155
timestamp 1751532423
transform 1 0 18704 0 -1 20384
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_21_190
timestamp 1751532312
transform 1 0 22624 0 -1 20384
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_21_204
timestamp 1751532246
transform 1 0 24192 0 -1 20384
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_21_208
timestamp 1751532440
transform 1 0 24640 0 -1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_21_212
timestamp 1751532312
transform 1 0 25088 0 -1 20384
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_21_220
timestamp 1751532440
transform 1 0 25984 0 -1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_21_222
timestamp 1751532423
transform 1 0 26208 0 -1 20384
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_21_266
timestamp 1751532246
transform 1 0 31136 0 -1 20384
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_21_270
timestamp 1751532423
transform 1 0 31584 0 -1 20384
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_21_278
timestamp 1751532440
transform 1 0 32480 0 -1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_21_288
timestamp 1751532246
transform 1 0 33600 0 -1 20384
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_21_292
timestamp 1751532440
transform 1 0 34048 0 -1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_21_294
timestamp 1751532423
transform 1 0 34272 0 -1 20384
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_22_2
timestamp 1751532351
transform 1 0 1568 0 1 20384
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_22_18
timestamp 1751532423
transform 1 0 3360 0 1 20384
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_22_26
timestamp 1751532312
transform 1 0 4256 0 1 20384
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_22_34
timestamp 1751532423
transform 1 0 5152 0 1 20384
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_22_47
timestamp 1751532246
transform 1 0 6608 0 1 20384
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_22_58
timestamp 1751532351
transform 1 0 7840 0 1 20384
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_22_74
timestamp 1751532312
transform 1 0 9632 0 1 20384
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_22_82
timestamp 1751532246
transform 1 0 10528 0 1 20384
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_22_86
timestamp 1751532440
transform 1 0 10976 0 1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_22_88
timestamp 1751532423
transform 1 0 11200 0 1 20384
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_22_103
timestamp 1751532440
transform 1 0 12880 0 1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_22_107
timestamp 1751532246
transform 1 0 13328 0 1 20384
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_22_111
timestamp 1751532423
transform 1 0 13776 0 1 20384
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_22_119
timestamp 1751532440
transform 1 0 14672 0 1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_22_128
timestamp 1751532423
transform 1 0 15680 0 1 20384
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_22_133
timestamp 1751532351
transform 1 0 16240 0 1 20384
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_22_149
timestamp 1751532312
transform 1 0 18032 0 1 20384
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_22_157
timestamp 1751532246
transform 1 0 18928 0 1 20384
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_22_161
timestamp 1751532423
transform 1 0 19376 0 1 20384
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_22_231
timestamp 1751532246
transform 1 0 27216 0 1 20384
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_22_243
timestamp 1751532440
transform 1 0 28560 0 1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_22_279
timestamp 1751532351
transform 1 0 32592 0 1 20384
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_23_2
timestamp 1751532351
transform 1 0 1568 0 -1 21952
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_23_18
timestamp 1751532246
transform 1 0 3360 0 -1 21952
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_23_22
timestamp 1751532440
transform 1 0 3808 0 -1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_23_35
timestamp 1751532351
transform 1 0 5264 0 -1 21952
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_23_51
timestamp 1751532312
transform 1 0 7056 0 -1 21952
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_23_59
timestamp 1751532423
transform 1 0 7952 0 -1 21952
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_23_66
timestamp 1751532440
transform 1 0 8736 0 -1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_23_72
timestamp 1751532351
transform 1 0 9408 0 -1 21952
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_23_88
timestamp 1751532440
transform 1 0 11200 0 -1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_23_90
timestamp 1751532423
transform 1 0 11424 0 -1 21952
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_23_97
timestamp 1751532312
transform 1 0 12208 0 -1 21952
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_23_109
timestamp 1751532351
transform 1 0 13552 0 -1 21952
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_23_125
timestamp 1751532312
transform 1 0 15344 0 -1 21952
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_23_133
timestamp 1751532246
transform 1 0 16240 0 -1 21952
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_23_137
timestamp 1751532440
transform 1 0 16688 0 -1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_23_139
timestamp 1751532423
transform 1 0 16912 0 -1 21952
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_23_142
timestamp 1751532246
transform 1 0 17248 0 -1 21952
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_23_156
timestamp 1751532351
transform 1 0 18816 0 -1 21952
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_23_172
timestamp 1751532440
transform 1 0 20608 0 -1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_23_186
timestamp 1751532246
transform 1 0 22176 0 -1 21952
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_23_190
timestamp 1751532440
transform 1 0 22624 0 -1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_23_204
timestamp 1751532246
transform 1 0 24192 0 -1 21952
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_23_208
timestamp 1751532440
transform 1 0 24640 0 -1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_23_212
timestamp 1751532351
transform 1 0 25088 0 -1 21952
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_23_228
timestamp 1751532351
transform 1 0 26880 0 -1 21952
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_23_244
timestamp 1751532440
transform 1 0 28672 0 -1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_23_282
timestamp 1751532440
transform 1 0 32928 0 -1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_23_286
timestamp 1751532312
transform 1 0 33376 0 -1 21952
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_23_294
timestamp 1751532423
transform 1 0 34272 0 -1 21952
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_24_2
timestamp 1751532312
transform 1 0 1568 0 1 21952
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_24_16
timestamp 1751532246
transform 1 0 3136 0 1 21952
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_24_30
timestamp 1751532440
transform 1 0 4704 0 1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_24_34
timestamp 1751532423
transform 1 0 5152 0 1 21952
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_24_37
timestamp 1751532351
transform 1 0 5488 0 1 21952
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_24_79
timestamp 1751532246
transform 1 0 10192 0 1 21952
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_24_83
timestamp 1751532440
transform 1 0 10640 0 1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_24_98
timestamp 1751532423
transform 1 0 12320 0 1 21952
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_24_120
timestamp 1751532312
transform 1 0 14784 0 1 21952
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_24_128
timestamp 1751532440
transform 1 0 15680 0 1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_24_132
timestamp 1751532312
transform 1 0 16128 0 1 21952
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_24_161
timestamp 1751532312
transform 1 0 19376 0 1 21952
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_24_169
timestamp 1751532246
transform 1 0 20272 0 1 21952
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_24_173
timestamp 1751532440
transform 1 0 20720 0 1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_24_177
timestamp 1751532312
transform 1 0 21168 0 1 21952
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_24_185
timestamp 1751532440
transform 1 0 22064 0 1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_24_221
timestamp 1751532351
transform 1 0 26096 0 1 21952
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_24_237
timestamp 1751532312
transform 1 0 27888 0 1 21952
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_24_272
timestamp 1751532440
transform 1 0 31808 0 1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_24_276
timestamp 1751532351
transform 1 0 32256 0 1 21952
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_24_292
timestamp 1751532440
transform 1 0 34048 0 1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_24_294
timestamp 1751532423
transform 1 0 34272 0 1 21952
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_25_50
timestamp 1751532246
transform 1 0 6944 0 -1 23520
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_25_54
timestamp 1751532440
transform 1 0 7392 0 -1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_25_56
timestamp 1751532423
transform 1 0 7616 0 -1 23520
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_25_67
timestamp 1751532440
transform 1 0 8848 0 -1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_25_69
timestamp 1751532423
transform 1 0 9072 0 -1 23520
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_25_72
timestamp 1751532246
transform 1 0 9408 0 -1 23520
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_25_142
timestamp 1751532246
transform 1 0 17248 0 -1 23520
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_25_156
timestamp 1751532440
transform 1 0 18816 0 -1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_25_165
timestamp 1751532440
transform 1 0 19824 0 -1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_25_175
timestamp 1751532312
transform 1 0 20944 0 -1 23520
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_25_219
timestamp 1751532440
transform 1 0 25872 0 -1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_25_223
timestamp 1751532440
transform 1 0 26320 0 -1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_25_252
timestamp 1751532440
transform 1 0 29568 0 -1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_25_256
timestamp 1751532440
transform 1 0 30016 0 -1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_25_258
timestamp 1751532423
transform 1 0 30240 0 -1 23520
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_25_265
timestamp 1751532312
transform 1 0 31024 0 -1 23520
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_25_273
timestamp 1751532246
transform 1 0 31920 0 -1 23520
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_25_277
timestamp 1751532440
transform 1 0 32368 0 -1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_25_279
timestamp 1751532423
transform 1 0 32592 0 -1 23520
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_25_282
timestamp 1751532312
transform 1 0 32928 0 -1 23520
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_25_290
timestamp 1751532246
transform 1 0 33824 0 -1 23520
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_25_294
timestamp 1751532423
transform 1 0 34272 0 -1 23520
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_26_2
timestamp 1751532351
transform 1 0 1568 0 1 23520
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_26_37
timestamp 1751532423
transform 1 0 5488 0 1 23520
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_26_66
timestamp 1751532423
transform 1 0 8736 0 1 23520
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_26_81
timestamp 1751532246
transform 1 0 10416 0 1 23520
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_26_151
timestamp 1751532246
transform 1 0 18256 0 1 23520
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_26_177
timestamp 1751532312
transform 1 0 21168 0 1 23520
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_26_185
timestamp 1751532246
transform 1 0 22064 0 1 23520
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_26_189
timestamp 1751532423
transform 1 0 22512 0 1 23520
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_26_196
timestamp 1751532440
transform 1 0 23296 0 1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_26_225
timestamp 1751532440
transform 1 0 26544 0 1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_26_253
timestamp 1751532351
transform 1 0 29680 0 1 23520
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_26_269
timestamp 1751532351
transform 1 0 31472 0 1 23520
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_26_285
timestamp 1751532312
transform 1 0 33264 0 1 23520
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_26_293
timestamp 1751532440
transform 1 0 34160 0 1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_27_2
timestamp 1751532312
transform 1 0 1568 0 -1 25088
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_27_16
timestamp 1751532246
transform 1 0 3136 0 -1 25088
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_27_20
timestamp 1751532440
transform 1 0 3584 0 -1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_27_22
timestamp 1751532423
transform 1 0 3808 0 -1 25088
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_27_37
timestamp 1751532312
transform 1 0 5488 0 -1 25088
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_27_45
timestamp 1751532440
transform 1 0 6384 0 -1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_27_64
timestamp 1751532246
transform 1 0 8512 0 -1 25088
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_27_68
timestamp 1751532440
transform 1 0 8960 0 -1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_27_104
timestamp 1751532423
transform 1 0 12992 0 -1 25088
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_27_137
timestamp 1751532440
transform 1 0 16688 0 -1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_27_139
timestamp 1751532423
transform 1 0 16912 0 -1 25088
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_27_148
timestamp 1751532246
transform 1 0 17920 0 -1 25088
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_27_190
timestamp 1751532423
transform 1 0 22624 0 -1 25088
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_27_209
timestamp 1751532423
transform 1 0 24752 0 -1 25088
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_27_218
timestamp 1751532312
transform 1 0 25760 0 -1 25088
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_27_228
timestamp 1751532440
transform 1 0 26880 0 -1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_27_256
timestamp 1751532351
transform 1 0 30016 0 -1 25088
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_27_272
timestamp 1751532312
transform 1 0 31808 0 -1 25088
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_27_282
timestamp 1751532312
transform 1 0 32928 0 -1 25088
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_27_290
timestamp 1751532246
transform 1 0 33824 0 -1 25088
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_27_294
timestamp 1751532423
transform 1 0 34272 0 -1 25088
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_28_37
timestamp 1751532440
transform 1 0 5488 0 1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_28_41
timestamp 1751532423
transform 1 0 5936 0 1 25088
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_28_73
timestamp 1751532440
transform 1 0 9520 0 1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_28_77
timestamp 1751532423
transform 1 0 9968 0 1 25088
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_28_111
timestamp 1751532423
transform 1 0 13776 0 1 25088
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_28_147
timestamp 1751532312
transform 1 0 17808 0 1 25088
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_28_162
timestamp 1751532423
transform 1 0 19488 0 1 25088
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_28_173
timestamp 1751532440
transform 1 0 20720 0 1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_28_177
timestamp 1751532351
transform 1 0 21168 0 1 25088
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_28_193
timestamp 1751532440
transform 1 0 22960 0 1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_28_195
timestamp 1751532423
transform 1 0 23184 0 1 25088
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_28_212
timestamp 1751532351
transform 1 0 25088 0 1 25088
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_28_228
timestamp 1751532423
transform 1 0 26880 0 1 25088
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_28_243
timestamp 1751532440
transform 1 0 28560 0 1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_28_274
timestamp 1751532440
transform 1 0 32032 0 1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_28_278
timestamp 1751532351
transform 1 0 32480 0 1 25088
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_28_294
timestamp 1751532423
transform 1 0 34272 0 1 25088
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_29_2
timestamp 1751532246
transform 1 0 1568 0 -1 26656
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_29_6
timestamp 1751532440
transform 1 0 2016 0 -1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_29_69
timestamp 1751532423
transform 1 0 9072 0 -1 26656
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_29_79
timestamp 1751532440
transform 1 0 10192 0 -1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_29_83
timestamp 1751532440
transform 1 0 10640 0 -1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_29_85
timestamp 1751532423
transform 1 0 10864 0 -1 26656
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_29_92
timestamp 1751532440
transform 1 0 11648 0 -1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_29_103
timestamp 1751532440
transform 1 0 12880 0 -1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_29_107
timestamp 1751532351
transform 1 0 13328 0 -1 26656
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_29_123
timestamp 1751532246
transform 1 0 15120 0 -1 26656
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_29_127
timestamp 1751532440
transform 1 0 15568 0 -1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_29_129
timestamp 1751532423
transform 1 0 15792 0 -1 26656
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_29_132
timestamp 1751532440
transform 1 0 16128 0 -1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_29_136
timestamp 1751532246
transform 1 0 16576 0 -1 26656
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_29_169
timestamp 1751532246
transform 1 0 20272 0 -1 26656
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_29_180
timestamp 1751532312
transform 1 0 21504 0 -1 26656
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_29_188
timestamp 1751532246
transform 1 0 22400 0 -1 26656
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_29_198
timestamp 1751532423
transform 1 0 23520 0 -1 26656
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_29_206
timestamp 1751532246
transform 1 0 24416 0 -1 26656
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_29_212
timestamp 1751532312
transform 1 0 25088 0 -1 26656
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_29_220
timestamp 1751532440
transform 1 0 25984 0 -1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_29_222
timestamp 1751532423
transform 1 0 26208 0 -1 26656
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_29_229
timestamp 1751532440
transform 1 0 26992 0 -1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_29_231
timestamp 1751532423
transform 1 0 27216 0 -1 26656
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_29_239
timestamp 1751532440
transform 1 0 28112 0 -1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_29_255
timestamp 1751532351
transform 1 0 29904 0 -1 26656
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_29_271
timestamp 1751532312
transform 1 0 31696 0 -1 26656
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_29_279
timestamp 1751532423
transform 1 0 32592 0 -1 26656
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_29_282
timestamp 1751532312
transform 1 0 32928 0 -1 26656
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_29_290
timestamp 1751532246
transform 1 0 33824 0 -1 26656
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_29_294
timestamp 1751532423
transform 1 0 34272 0 -1 26656
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_30_2
timestamp 1751532351
transform 1 0 1568 0 1 26656
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_30_18
timestamp 1751532351
transform 1 0 3360 0 1 26656
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_30_34
timestamp 1751532423
transform 1 0 5152 0 1 26656
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_30_37
timestamp 1751532440
transform 1 0 5488 0 1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_30_41
timestamp 1751532246
transform 1 0 5936 0 1 26656
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_30_45
timestamp 1751532440
transform 1 0 6384 0 1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_30_47
timestamp 1751532423
transform 1 0 6608 0 1 26656
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_30_54
timestamp 1751532423
transform 1 0 7392 0 1 26656
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_30_82
timestamp 1751532440
transform 1 0 10528 0 1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_30_86
timestamp 1751532351
transform 1 0 10976 0 1 26656
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_30_102
timestamp 1751532440
transform 1 0 12768 0 1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_30_104
timestamp 1751532423
transform 1 0 12992 0 1 26656
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_30_107
timestamp 1751532246
transform 1 0 13328 0 1 26656
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_30_111
timestamp 1751532423
transform 1 0 13776 0 1 26656
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_30_126
timestamp 1751532246
transform 1 0 15456 0 1 26656
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_30_130
timestamp 1751532440
transform 1 0 15904 0 1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_30_132
timestamp 1751532423
transform 1 0 16128 0 1 26656
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_30_147
timestamp 1751532351
transform 1 0 17808 0 1 26656
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_30_163
timestamp 1751532246
transform 1 0 19600 0 1 26656
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_30_167
timestamp 1751532423
transform 1 0 20048 0 1 26656
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_30_204
timestamp 1751532312
transform 1 0 24192 0 1 26656
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_30_239
timestamp 1751532246
transform 1 0 28112 0 1 26656
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_30_243
timestamp 1751532440
transform 1 0 28560 0 1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_30_247
timestamp 1751532351
transform 1 0 29008 0 1 26656
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_30_263
timestamp 1751532351
transform 1 0 30800 0 1 26656
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_30_279
timestamp 1751532351
transform 1 0 32592 0 1 26656
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_31_2
timestamp 1751532351
transform 1 0 1568 0 -1 28224
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_31_18
timestamp 1751532351
transform 1 0 3360 0 -1 28224
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_31_34
timestamp 1751532351
transform 1 0 5152 0 -1 28224
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_31_50
timestamp 1751532312
transform 1 0 6944 0 -1 28224
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_31_58
timestamp 1751532440
transform 1 0 7840 0 -1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_31_66
timestamp 1751532246
transform 1 0 8736 0 -1 28224
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_31_72
timestamp 1751532312
transform 1 0 9408 0 -1 28224
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_31_80
timestamp 1751532246
transform 1 0 10304 0 -1 28224
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_31_84
timestamp 1751532423
transform 1 0 10752 0 -1 28224
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_31_91
timestamp 1751532246
transform 1 0 11536 0 -1 28224
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_31_95
timestamp 1751532423
transform 1 0 11984 0 -1 28224
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_31_107
timestamp 1751532246
transform 1 0 13328 0 -1 28224
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_31_111
timestamp 1751532440
transform 1 0 13776 0 -1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_31_142
timestamp 1751532351
transform 1 0 17248 0 -1 28224
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_31_158
timestamp 1751532351
transform 1 0 19040 0 -1 28224
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_31_174
timestamp 1751532440
transform 1 0 20832 0 -1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_31_176
timestamp 1751532423
transform 1 0 21056 0 -1 28224
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_31_183
timestamp 1751532312
transform 1 0 21840 0 -1 28224
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_31_191
timestamp 1751532246
transform 1 0 22736 0 -1 28224
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_31_195
timestamp 1751532423
transform 1 0 23184 0 -1 28224
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_31_203
timestamp 1751532246
transform 1 0 24080 0 -1 28224
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_31_207
timestamp 1751532440
transform 1 0 24528 0 -1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_31_209
timestamp 1751532423
transform 1 0 24752 0 -1 28224
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_31_219
timestamp 1751532246
transform 1 0 25872 0 -1 28224
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_31_223
timestamp 1751532440
transform 1 0 26320 0 -1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_31_225
timestamp 1751532423
transform 1 0 26544 0 -1 28224
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_31_251
timestamp 1751532351
transform 1 0 29456 0 -1 28224
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_31_267
timestamp 1751532312
transform 1 0 31248 0 -1 28224
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_31_275
timestamp 1751532246
transform 1 0 32144 0 -1 28224
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_31_279
timestamp 1751532423
transform 1 0 32592 0 -1 28224
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_31_282
timestamp 1751532312
transform 1 0 32928 0 -1 28224
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_31_290
timestamp 1751532246
transform 1 0 33824 0 -1 28224
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_31_294
timestamp 1751532423
transform 1 0 34272 0 -1 28224
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_32_2
timestamp 1751532351
transform 1 0 1568 0 1 28224
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_32_18
timestamp 1751532351
transform 1 0 3360 0 1 28224
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_32_34
timestamp 1751532423
transform 1 0 5152 0 1 28224
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_32_37
timestamp 1751532351
transform 1 0 5488 0 1 28224
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_32_53
timestamp 1751532351
transform 1 0 7280 0 1 28224
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_32_69
timestamp 1751532246
transform 1 0 9072 0 1 28224
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_32_73
timestamp 1751532423
transform 1 0 9520 0 1 28224
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_32_101
timestamp 1751532440
transform 1 0 12656 0 1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_32_131
timestamp 1751532312
transform 1 0 16016 0 1 28224
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_32_139
timestamp 1751532440
transform 1 0 16912 0 1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_32_177
timestamp 1751532312
transform 1 0 21168 0 1 28224
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_32_185
timestamp 1751532246
transform 1 0 22064 0 1 28224
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_32_189
timestamp 1751532440
transform 1 0 22512 0 1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_32_197
timestamp 1751532440
transform 1 0 23408 0 1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_32_220
timestamp 1751532246
transform 1 0 25984 0 1 28224
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_32_224
timestamp 1751532423
transform 1 0 26432 0 1 28224
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_32_239
timestamp 1751532246
transform 1 0 28112 0 1 28224
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_32_243
timestamp 1751532440
transform 1 0 28560 0 1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_32_247
timestamp 1751532351
transform 1 0 29008 0 1 28224
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_32_263
timestamp 1751532351
transform 1 0 30800 0 1 28224
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_32_279
timestamp 1751532351
transform 1 0 32592 0 1 28224
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_33_2
timestamp 1751532351
transform 1 0 1568 0 -1 29792
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_33_18
timestamp 1751532351
transform 1 0 3360 0 -1 29792
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_33_34
timestamp 1751532351
transform 1 0 5152 0 -1 29792
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_33_50
timestamp 1751532351
transform 1 0 6944 0 -1 29792
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_33_66
timestamp 1751532246
transform 1 0 8736 0 -1 29792
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_33_72
timestamp 1751532351
transform 1 0 9408 0 -1 29792
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_33_88
timestamp 1751532440
transform 1 0 11200 0 -1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_33_90
timestamp 1751532423
transform 1 0 11424 0 -1 29792
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_33_98
timestamp 1751532423
transform 1 0 12320 0 -1 29792
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_33_113
timestamp 1751532423
transform 1 0 14000 0 -1 29792
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_33_121
timestamp 1751532246
transform 1 0 14896 0 -1 29792
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_33_125
timestamp 1751532440
transform 1 0 15344 0 -1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_33_127
timestamp 1751532423
transform 1 0 15568 0 -1 29792
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_33_135
timestamp 1751532246
transform 1 0 16464 0 -1 29792
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_33_139
timestamp 1751532423
transform 1 0 16912 0 -1 29792
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_33_142
timestamp 1751532246
transform 1 0 17248 0 -1 29792
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_33_146
timestamp 1751532440
transform 1 0 17696 0 -1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_33_179
timestamp 1751532312
transform 1 0 21392 0 -1 29792
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_33_187
timestamp 1751532423
transform 1 0 22288 0 -1 29792
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_33_206
timestamp 1751532246
transform 1 0 24416 0 -1 29792
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_33_223
timestamp 1751532246
transform 1 0 26320 0 -1 29792
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_33_238
timestamp 1751532351
transform 1 0 28000 0 -1 29792
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_33_254
timestamp 1751532351
transform 1 0 29792 0 -1 29792
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_33_270
timestamp 1751532312
transform 1 0 31584 0 -1 29792
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_33_278
timestamp 1751532440
transform 1 0 32480 0 -1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_33_282
timestamp 1751532312
transform 1 0 32928 0 -1 29792
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_33_290
timestamp 1751532246
transform 1 0 33824 0 -1 29792
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_33_294
timestamp 1751532423
transform 1 0 34272 0 -1 29792
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_34_2
timestamp 1751532351
transform 1 0 1568 0 1 29792
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_34_18
timestamp 1751532351
transform 1 0 3360 0 1 29792
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_34_34
timestamp 1751532423
transform 1 0 5152 0 1 29792
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_34_37
timestamp 1751532351
transform 1 0 5488 0 1 29792
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_34_53
timestamp 1751532351
transform 1 0 7280 0 1 29792
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_34_69
timestamp 1751532246
transform 1 0 9072 0 1 29792
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_34_73
timestamp 1751532423
transform 1 0 9520 0 1 29792
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_34_101
timestamp 1751532440
transform 1 0 12656 0 1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_34_121
timestamp 1751532246
transform 1 0 14896 0 1 29792
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_34_125
timestamp 1751532440
transform 1 0 15344 0 1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_34_152
timestamp 1751532440
transform 1 0 18368 0 1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_34_154
timestamp 1751532423
transform 1 0 18592 0 1 29792
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_34_177
timestamp 1751532246
transform 1 0 21168 0 1 29792
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_34_215
timestamp 1751532440
transform 1 0 25424 0 1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_34_217
timestamp 1751532423
transform 1 0 25648 0 1 29792
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_34_247
timestamp 1751532440
transform 1 0 29008 0 1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_34_251
timestamp 1751532351
transform 1 0 29456 0 1 29792
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_34_267
timestamp 1751532351
transform 1 0 31248 0 1 29792
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_34_283
timestamp 1751532312
transform 1 0 33040 0 1 29792
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_34_291
timestamp 1751532246
transform 1 0 33936 0 1 29792
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_35_2
timestamp 1751532351
transform 1 0 1568 0 -1 31360
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_35_18
timestamp 1751532351
transform 1 0 3360 0 -1 31360
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_35_34
timestamp 1751532351
transform 1 0 5152 0 -1 31360
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_35_50
timestamp 1751532351
transform 1 0 6944 0 -1 31360
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_35_66
timestamp 1751532246
transform 1 0 8736 0 -1 31360
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_35_72
timestamp 1751532312
transform 1 0 9408 0 -1 31360
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_35_80
timestamp 1751532246
transform 1 0 10304 0 -1 31360
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_35_84
timestamp 1751532440
transform 1 0 10752 0 -1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_35_142
timestamp 1751532312
transform 1 0 17248 0 -1 31360
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_35_150
timestamp 1751532440
transform 1 0 18144 0 -1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_35_179
timestamp 1751532246
transform 1 0 21392 0 -1 31360
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_35_218
timestamp 1751532312
transform 1 0 25760 0 -1 31360
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_35_226
timestamp 1751532246
transform 1 0 26656 0 -1 31360
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_35_230
timestamp 1751532423
transform 1 0 27104 0 -1 31360
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_35_237
timestamp 1751532351
transform 1 0 27888 0 -1 31360
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_35_253
timestamp 1751532351
transform 1 0 29680 0 -1 31360
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_35_269
timestamp 1751532312
transform 1 0 31472 0 -1 31360
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_35_277
timestamp 1751532440
transform 1 0 32368 0 -1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_35_279
timestamp 1751532423
transform 1 0 32592 0 -1 31360
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_8  FILLER_0_35_282
timestamp 1751532312
transform 1 0 32928 0 -1 31360
box -86 -86 982 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_35_290
timestamp 1751532246
transform 1 0 33824 0 -1 31360
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_35_294
timestamp 1751532423
transform 1 0 34272 0 -1 31360
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_36_2
timestamp 1751532351
transform 1 0 1568 0 1 31360
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_36_18
timestamp 1751532351
transform 1 0 3360 0 1 31360
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_36_36
timestamp 1751532351
transform 1 0 5376 0 1 31360
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_36_52
timestamp 1751532351
transform 1 0 7168 0 1 31360
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_36_70
timestamp 1751532351
transform 1 0 9184 0 1 31360
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_36_86
timestamp 1751532351
transform 1 0 10976 0 1 31360
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_36_111
timestamp 1751532351
transform 1 0 13776 0 1 31360
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__fill_2  FILLER_0_36_133
timestamp 1751532440
transform 1 0 16240 0 1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_36_135
timestamp 1751532423
transform 1 0 16464 0 1 31360
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_36_138
timestamp 1751532351
transform 1 0 16800 0 1 31360
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_36_154
timestamp 1751532246
transform 1 0 18592 0 1 31360
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_36_165
timestamp 1751532246
transform 1 0 19824 0 1 31360
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_36_169
timestamp 1751532423
transform 1 0 20272 0 1 31360
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_36_172
timestamp 1751532351
transform 1 0 20608 0 1 31360
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_36_188
timestamp 1751532351
transform 1 0 22400 0 1 31360
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_36_206
timestamp 1751532351
transform 1 0 24416 0 1 31360
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_36_222
timestamp 1751532351
transform 1 0 26208 0 1 31360
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_36_240
timestamp 1751532351
transform 1 0 28224 0 1 31360
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_36_256
timestamp 1751532351
transform 1 0 30016 0 1 31360
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_16  FILLER_0_36_274
timestamp 1751532351
transform 1 0 32032 0 1 31360
box -86 -86 1878 870
use gf180mcu_as_sc_mcu7t3v3__decap_4  FILLER_0_36_290
timestamp 1751532246
transform 1 0 33824 0 1 31360
box -86 -86 534 870
use gf180mcu_as_sc_mcu7t3v3__fill_1  FILLER_0_36_294
timestamp 1751532423
transform 1 0 34272 0 1 31360
box -86 -86 198 870
use gf180mcu_as_sc_mcu7t3v3__buff_2  input1
timestamp 1751534193
transform 1 0 10864 0 1 3136
box -86 -86 758 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  output2
timestamp 1751661108
transform -1 0 20384 0 1 3136
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  output3
timestamp 1751661108
transform 1 0 25200 0 1 3136
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__clkbuff_12  output4
timestamp 1751661108
transform -1 0 32704 0 -1 4704
box -86 -86 2886 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_0_Left_37 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_as_sc_mcu7t3v3/mag
timestamp 1751532504
transform 1 0 1344 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_0_Right_0
timestamp 1751532504
transform -1 0 34608 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_1_Left_38
timestamp 1751532504
transform 1 0 1344 0 -1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_1_Right_1
timestamp 1751532504
transform -1 0 34608 0 -1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_2_Left_39
timestamp 1751532504
transform 1 0 1344 0 1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_2_Right_2
timestamp 1751532504
transform -1 0 34608 0 1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_3_Left_40
timestamp 1751532504
transform 1 0 1344 0 -1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_3_Right_3
timestamp 1751532504
transform -1 0 34608 0 -1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_4_Left_41
timestamp 1751532504
transform 1 0 1344 0 1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_4_Right_4
timestamp 1751532504
transform -1 0 34608 0 1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_5_Left_42
timestamp 1751532504
transform 1 0 1344 0 -1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_5_Right_5
timestamp 1751532504
transform -1 0 34608 0 -1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_6_Left_43
timestamp 1751532504
transform 1 0 1344 0 1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_6_Right_6
timestamp 1751532504
transform -1 0 34608 0 1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_7_Left_44
timestamp 1751532504
transform 1 0 1344 0 -1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_7_Right_7
timestamp 1751532504
transform -1 0 34608 0 -1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_8_Left_45
timestamp 1751532504
transform 1 0 1344 0 1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_8_Right_8
timestamp 1751532504
transform -1 0 34608 0 1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_9_Left_46
timestamp 1751532504
transform 1 0 1344 0 -1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_9_Right_9
timestamp 1751532504
transform -1 0 34608 0 -1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_10_Left_47
timestamp 1751532504
transform 1 0 1344 0 1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_10_Right_10
timestamp 1751532504
transform -1 0 34608 0 1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_11_Left_48
timestamp 1751532504
transform 1 0 1344 0 -1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_11_Right_11
timestamp 1751532504
transform -1 0 34608 0 -1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_12_Left_49
timestamp 1751532504
transform 1 0 1344 0 1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_12_Right_12
timestamp 1751532504
transform -1 0 34608 0 1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_13_Left_50
timestamp 1751532504
transform 1 0 1344 0 -1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_13_Right_13
timestamp 1751532504
transform -1 0 34608 0 -1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_14_Left_51
timestamp 1751532504
transform 1 0 1344 0 1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_14_Right_14
timestamp 1751532504
transform -1 0 34608 0 1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_15_Left_52
timestamp 1751532504
transform 1 0 1344 0 -1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_15_Right_15
timestamp 1751532504
transform -1 0 34608 0 -1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_16_Left_53
timestamp 1751532504
transform 1 0 1344 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_16_Right_16
timestamp 1751532504
transform -1 0 34608 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_17_Left_54
timestamp 1751532504
transform 1 0 1344 0 -1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_17_Right_17
timestamp 1751532504
transform -1 0 34608 0 -1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_18_Left_55
timestamp 1751532504
transform 1 0 1344 0 1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_18_Right_18
timestamp 1751532504
transform -1 0 34608 0 1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_19_Left_56
timestamp 1751532504
transform 1 0 1344 0 -1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_19_Right_19
timestamp 1751532504
transform -1 0 34608 0 -1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_20_Left_57
timestamp 1751532504
transform 1 0 1344 0 1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_20_Right_20
timestamp 1751532504
transform -1 0 34608 0 1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_21_Left_58
timestamp 1751532504
transform 1 0 1344 0 -1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_21_Right_21
timestamp 1751532504
transform -1 0 34608 0 -1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_22_Left_59
timestamp 1751532504
transform 1 0 1344 0 1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_22_Right_22
timestamp 1751532504
transform -1 0 34608 0 1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_23_Left_60
timestamp 1751532504
transform 1 0 1344 0 -1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_23_Right_23
timestamp 1751532504
transform -1 0 34608 0 -1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_24_Left_61
timestamp 1751532504
transform 1 0 1344 0 1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_24_Right_24
timestamp 1751532504
transform -1 0 34608 0 1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_25_Left_62
timestamp 1751532504
transform 1 0 1344 0 -1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_25_Right_25
timestamp 1751532504
transform -1 0 34608 0 -1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_26_Left_63
timestamp 1751532504
transform 1 0 1344 0 1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_26_Right_26
timestamp 1751532504
transform -1 0 34608 0 1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_27_Left_64
timestamp 1751532504
transform 1 0 1344 0 -1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_27_Right_27
timestamp 1751532504
transform -1 0 34608 0 -1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_28_Left_65
timestamp 1751532504
transform 1 0 1344 0 1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_28_Right_28
timestamp 1751532504
transform -1 0 34608 0 1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_29_Left_66
timestamp 1751532504
transform 1 0 1344 0 -1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_29_Right_29
timestamp 1751532504
transform -1 0 34608 0 -1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_30_Left_67
timestamp 1751532504
transform 1 0 1344 0 1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_30_Right_30
timestamp 1751532504
transform -1 0 34608 0 1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_31_Left_68
timestamp 1751532504
transform 1 0 1344 0 -1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_31_Right_31
timestamp 1751532504
transform -1 0 34608 0 -1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_32_Left_69
timestamp 1751532504
transform 1 0 1344 0 1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_32_Right_32
timestamp 1751532504
transform -1 0 34608 0 1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_33_Left_70
timestamp 1751532504
transform 1 0 1344 0 -1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_33_Right_33
timestamp 1751532504
transform -1 0 34608 0 -1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_34_Left_71
timestamp 1751532504
transform 1 0 1344 0 1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_34_Right_34
timestamp 1751532504
transform -1 0 34608 0 1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_35_Left_72
timestamp 1751532504
transform 1 0 1344 0 -1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_35_Right_35
timestamp 1751532504
transform -1 0 34608 0 -1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_36_Left_73
timestamp 1751532504
transform 1 0 1344 0 1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  PHY_EDGE_ROW_36_Right_36
timestamp 1751532504
transform -1 0 34608 0 1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_0_74
timestamp 1751532504
transform 1 0 5152 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_0_75
timestamp 1751532504
transform 1 0 8960 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_0_76
timestamp 1751532504
transform 1 0 12768 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_0_77
timestamp 1751532504
transform 1 0 16576 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_0_78
timestamp 1751532504
transform 1 0 20384 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_0_79
timestamp 1751532504
transform 1 0 24192 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_0_80
timestamp 1751532504
transform 1 0 28000 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_0_81
timestamp 1751532504
transform 1 0 31808 0 1 3136
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_1_82
timestamp 1751532504
transform 1 0 9184 0 -1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_1_83
timestamp 1751532504
transform 1 0 17024 0 -1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_1_84
timestamp 1751532504
transform 1 0 24864 0 -1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_1_85
timestamp 1751532504
transform 1 0 32704 0 -1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_2_86
timestamp 1751532504
transform 1 0 5264 0 1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_2_87
timestamp 1751532504
transform 1 0 13104 0 1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_2_88
timestamp 1751532504
transform 1 0 20944 0 1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_2_89
timestamp 1751532504
transform 1 0 28784 0 1 4704
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_3_90
timestamp 1751532504
transform 1 0 9184 0 -1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_3_91
timestamp 1751532504
transform 1 0 17024 0 -1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_3_92
timestamp 1751532504
transform 1 0 24864 0 -1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_3_93
timestamp 1751532504
transform 1 0 32704 0 -1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_4_94
timestamp 1751532504
transform 1 0 5264 0 1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_4_95
timestamp 1751532504
transform 1 0 13104 0 1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_4_96
timestamp 1751532504
transform 1 0 20944 0 1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_4_97
timestamp 1751532504
transform 1 0 28784 0 1 6272
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_5_98
timestamp 1751532504
transform 1 0 9184 0 -1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_5_99
timestamp 1751532504
transform 1 0 17024 0 -1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_5_100
timestamp 1751532504
transform 1 0 24864 0 -1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_5_101
timestamp 1751532504
transform 1 0 32704 0 -1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_6_102
timestamp 1751532504
transform 1 0 5264 0 1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_6_103
timestamp 1751532504
transform 1 0 13104 0 1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_6_104
timestamp 1751532504
transform 1 0 20944 0 1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_6_105
timestamp 1751532504
transform 1 0 28784 0 1 7840
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_7_106
timestamp 1751532504
transform 1 0 9184 0 -1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_7_107
timestamp 1751532504
transform 1 0 17024 0 -1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_7_108
timestamp 1751532504
transform 1 0 24864 0 -1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_7_109
timestamp 1751532504
transform 1 0 32704 0 -1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_8_110
timestamp 1751532504
transform 1 0 5264 0 1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_8_111
timestamp 1751532504
transform 1 0 13104 0 1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_8_112
timestamp 1751532504
transform 1 0 20944 0 1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_8_113
timestamp 1751532504
transform 1 0 28784 0 1 9408
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_9_114
timestamp 1751532504
transform 1 0 9184 0 -1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_9_115
timestamp 1751532504
transform 1 0 17024 0 -1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_9_116
timestamp 1751532504
transform 1 0 24864 0 -1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_9_117
timestamp 1751532504
transform 1 0 32704 0 -1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_10_118
timestamp 1751532504
transform 1 0 5264 0 1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_10_119
timestamp 1751532504
transform 1 0 13104 0 1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_10_120
timestamp 1751532504
transform 1 0 20944 0 1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_10_121
timestamp 1751532504
transform 1 0 28784 0 1 10976
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_11_122
timestamp 1751532504
transform 1 0 9184 0 -1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_11_123
timestamp 1751532504
transform 1 0 17024 0 -1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_11_124
timestamp 1751532504
transform 1 0 24864 0 -1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_11_125
timestamp 1751532504
transform 1 0 32704 0 -1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_12_126
timestamp 1751532504
transform 1 0 5264 0 1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_12_127
timestamp 1751532504
transform 1 0 13104 0 1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_12_128
timestamp 1751532504
transform 1 0 20944 0 1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_12_129
timestamp 1751532504
transform 1 0 28784 0 1 12544
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_13_130
timestamp 1751532504
transform 1 0 9184 0 -1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_13_131
timestamp 1751532504
transform 1 0 17024 0 -1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_13_132
timestamp 1751532504
transform 1 0 24864 0 -1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_13_133
timestamp 1751532504
transform 1 0 32704 0 -1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_14_134
timestamp 1751532504
transform 1 0 5264 0 1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_14_135
timestamp 1751532504
transform 1 0 13104 0 1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_14_136
timestamp 1751532504
transform 1 0 20944 0 1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_14_137
timestamp 1751532504
transform 1 0 28784 0 1 14112
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_15_138
timestamp 1751532504
transform 1 0 9184 0 -1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_15_139
timestamp 1751532504
transform 1 0 17024 0 -1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_15_140
timestamp 1751532504
transform 1 0 24864 0 -1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_15_141
timestamp 1751532504
transform 1 0 32704 0 -1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_16_142
timestamp 1751532504
transform 1 0 5264 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_16_143
timestamp 1751532504
transform 1 0 13104 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_16_144
timestamp 1751532504
transform 1 0 20944 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_16_145
timestamp 1751532504
transform 1 0 28784 0 1 15680
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_17_146
timestamp 1751532504
transform 1 0 9184 0 -1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_17_147
timestamp 1751532504
transform 1 0 17024 0 -1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_17_148
timestamp 1751532504
transform 1 0 24864 0 -1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_17_149
timestamp 1751532504
transform 1 0 32704 0 -1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_18_150
timestamp 1751532504
transform 1 0 5264 0 1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_18_151
timestamp 1751532504
transform 1 0 13104 0 1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_18_152
timestamp 1751532504
transform 1 0 20944 0 1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_18_153
timestamp 1751532504
transform 1 0 28784 0 1 17248
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_19_154
timestamp 1751532504
transform 1 0 9184 0 -1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_19_155
timestamp 1751532504
transform 1 0 17024 0 -1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_19_156
timestamp 1751532504
transform 1 0 24864 0 -1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_19_157
timestamp 1751532504
transform 1 0 32704 0 -1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_20_158
timestamp 1751532504
transform 1 0 5264 0 1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_20_159
timestamp 1751532504
transform 1 0 13104 0 1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_20_160
timestamp 1751532504
transform 1 0 20944 0 1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_20_161
timestamp 1751532504
transform 1 0 28784 0 1 18816
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_21_162
timestamp 1751532504
transform 1 0 9184 0 -1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_21_163
timestamp 1751532504
transform 1 0 17024 0 -1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_21_164
timestamp 1751532504
transform 1 0 24864 0 -1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_21_165
timestamp 1751532504
transform 1 0 32704 0 -1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_22_166
timestamp 1751532504
transform 1 0 5264 0 1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_22_167
timestamp 1751532504
transform 1 0 13104 0 1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_22_168
timestamp 1751532504
transform 1 0 20944 0 1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_22_169
timestamp 1751532504
transform 1 0 28784 0 1 20384
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_23_170
timestamp 1751532504
transform 1 0 9184 0 -1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_23_171
timestamp 1751532504
transform 1 0 17024 0 -1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_23_172
timestamp 1751532504
transform 1 0 24864 0 -1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_23_173
timestamp 1751532504
transform 1 0 32704 0 -1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_24_174
timestamp 1751532504
transform 1 0 5264 0 1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_24_175
timestamp 1751532504
transform 1 0 13104 0 1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_24_176
timestamp 1751532504
transform 1 0 20944 0 1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_24_177
timestamp 1751532504
transform 1 0 28784 0 1 21952
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_25_178
timestamp 1751532504
transform 1 0 9184 0 -1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_25_179
timestamp 1751532504
transform 1 0 17024 0 -1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_25_180
timestamp 1751532504
transform 1 0 24864 0 -1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_25_181
timestamp 1751532504
transform 1 0 32704 0 -1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_26_182
timestamp 1751532504
transform 1 0 5264 0 1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_26_183
timestamp 1751532504
transform 1 0 13104 0 1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_26_184
timestamp 1751532504
transform 1 0 20944 0 1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_26_185
timestamp 1751532504
transform 1 0 28784 0 1 23520
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_27_186
timestamp 1751532504
transform 1 0 9184 0 -1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_27_187
timestamp 1751532504
transform 1 0 17024 0 -1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_27_188
timestamp 1751532504
transform 1 0 24864 0 -1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_27_189
timestamp 1751532504
transform 1 0 32704 0 -1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_28_190
timestamp 1751532504
transform 1 0 5264 0 1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_28_191
timestamp 1751532504
transform 1 0 13104 0 1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_28_192
timestamp 1751532504
transform 1 0 20944 0 1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_28_193
timestamp 1751532504
transform 1 0 28784 0 1 25088
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_29_194
timestamp 1751532504
transform 1 0 9184 0 -1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_29_195
timestamp 1751532504
transform 1 0 17024 0 -1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_29_196
timestamp 1751532504
transform 1 0 24864 0 -1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_29_197
timestamp 1751532504
transform 1 0 32704 0 -1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_30_198
timestamp 1751532504
transform 1 0 5264 0 1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_30_199
timestamp 1751532504
transform 1 0 13104 0 1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_30_200
timestamp 1751532504
transform 1 0 20944 0 1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_30_201
timestamp 1751532504
transform 1 0 28784 0 1 26656
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_31_202
timestamp 1751532504
transform 1 0 9184 0 -1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_31_203
timestamp 1751532504
transform 1 0 17024 0 -1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_31_204
timestamp 1751532504
transform 1 0 24864 0 -1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_31_205
timestamp 1751532504
transform 1 0 32704 0 -1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_32_206
timestamp 1751532504
transform 1 0 5264 0 1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_32_207
timestamp 1751532504
transform 1 0 13104 0 1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_32_208
timestamp 1751532504
transform 1 0 20944 0 1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_32_209
timestamp 1751532504
transform 1 0 28784 0 1 28224
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_33_210
timestamp 1751532504
transform 1 0 9184 0 -1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_33_211
timestamp 1751532504
transform 1 0 17024 0 -1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_33_212
timestamp 1751532504
transform 1 0 24864 0 -1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_33_213
timestamp 1751532504
transform 1 0 32704 0 -1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_34_214
timestamp 1751532504
transform 1 0 5264 0 1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_34_215
timestamp 1751532504
transform 1 0 13104 0 1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_34_216
timestamp 1751532504
transform 1 0 20944 0 1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_34_217
timestamp 1751532504
transform 1 0 28784 0 1 29792
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_35_218
timestamp 1751532504
transform 1 0 9184 0 -1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_35_219
timestamp 1751532504
transform 1 0 17024 0 -1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_35_220
timestamp 1751532504
transform 1 0 24864 0 -1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_35_221
timestamp 1751532504
transform 1 0 32704 0 -1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_36_222
timestamp 1751532504
transform 1 0 5152 0 1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_36_223
timestamp 1751532504
transform 1 0 8960 0 1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_36_224
timestamp 1751532504
transform 1 0 12768 0 1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_36_225
timestamp 1751532504
transform 1 0 16576 0 1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_36_226
timestamp 1751532504
transform 1 0 20384 0 1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_36_227
timestamp 1751532504
transform 1 0 24192 0 1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_36_228
timestamp 1751532504
transform 1 0 28000 0 1 31360
box -86 -86 310 870
use gf180mcu_as_sc_mcu7t3v3__tap_2  TAP_TAPCELL_ROW_36_229
timestamp 1751532504
transform 1 0 31808 0 1 31360
box -86 -86 310 870
<< labels >>
flabel metal2 s 17920 0 18032 800 0 FreeSans 448 90 0 0 io_out[0]
port 0 nsew signal output
flabel metal2 s 25088 0 25200 800 0 FreeSans 448 90 0 0 io_out[1]
port 1 nsew signal output
flabel metal2 s 32256 0 32368 800 0 FreeSans 448 90 0 0 io_out[2]
port 2 nsew signal output
flabel metal2 s 10752 0 10864 800 0 FreeSans 448 90 0 0 rst_n
port 3 nsew signal input
flabel metal4 s 5342 3076 5662 32204 0 FreeSans 1280 90 0 0 vdd
port 4 nsew power bidirectional
flabel metal4 s 13658 3076 13978 32204 0 FreeSans 1280 90 0 0 vdd
port 4 nsew power bidirectional
flabel metal4 s 21974 3076 22294 32204 0 FreeSans 1280 90 0 0 vdd
port 4 nsew power bidirectional
flabel metal4 s 30290 3076 30610 32204 0 FreeSans 1280 90 0 0 vdd
port 4 nsew power bidirectional
flabel metal4 s 9500 3076 9820 32204 0 FreeSans 1280 90 0 0 vss
port 5 nsew ground bidirectional
flabel metal4 s 17816 3076 18136 32204 0 FreeSans 1280 90 0 0 vss
port 5 nsew ground bidirectional
flabel metal4 s 26132 3076 26452 32204 0 FreeSans 1280 90 0 0 vss
port 5 nsew ground bidirectional
flabel metal4 s 34448 3076 34768 32204 0 FreeSans 1280 90 0 0 vss
port 5 nsew ground bidirectional
flabel metal2 s 3584 0 3696 800 0 FreeSans 448 90 0 0 wb_clk_i
port 6 nsew signal input
rlabel metal1 17976 32144 17976 32144 0 vdd
rlabel via1 18056 31360 18056 31360 0 vss
rlabel metal2 4256 23240 4256 23240 0 LFSR\[0\]
rlabel metal2 4760 23352 4760 23352 0 LFSR\[1\]
rlabel metal3 5824 24696 5824 24696 0 LFSR\[2\]
rlabel metal2 10248 23968 10248 23968 0 LFSR\[3\]
rlabel metal2 8568 23800 8568 23800 0 LFSR\[4\]
rlabel metal2 8008 26096 8008 26096 0 LFSR\[5\]
rlabel metal2 12712 25592 12712 25592 0 LFSR\[6\]
rlabel metal2 32424 4760 32424 4760 0 OP
rlabel metal2 25816 22008 25816 22008 0 OP_reg
rlabel metal2 19096 12656 19096 12656 0 PC\[0\]
rlabel metal3 14812 13608 14812 13608 0 PC\[1\]
rlabel metal2 11368 13104 11368 13104 0 PC\[2\]
rlabel metal2 16800 4424 16800 4424 0 PC\[3\]
rlabel metal3 17528 5096 17528 5096 0 PC\[4\]
rlabel metal2 4704 4312 4704 4312 0 PC\[5\]
rlabel metal3 16520 8232 16520 8232 0 _0000_
rlabel metal2 8512 8232 8512 8232 0 _0001_
rlabel metal3 7784 14728 7784 14728 0 _0002_
rlabel metal2 3640 13272 3640 13272 0 _0003_
rlabel metal2 3080 14784 3080 14784 0 _0004_
rlabel metal3 6496 14728 6496 14728 0 _0005_
rlabel metal2 21336 8064 21336 8064 0 _0006_
rlabel metal2 20328 9688 20328 9688 0 _0007_
rlabel metal3 24864 11480 24864 11480 0 _0008_
rlabel metal2 24248 7532 24248 7532 0 _0009_
rlabel metal2 23800 5432 23800 5432 0 _0010_
rlabel metal2 21112 3808 21112 3808 0 _0011_
rlabel metal3 26656 4200 26656 4200 0 _0012_
rlabel metal2 33208 3920 33208 3920 0 _0013_
rlabel metal3 32760 6776 32760 6776 0 _0014_
rlabel metal2 26992 5880 26992 5880 0 _0015_
rlabel metal3 29960 8904 29960 8904 0 _0016_
rlabel metal2 26712 10864 26712 10864 0 _0017_
rlabel metal2 33320 9296 33320 9296 0 _0018_
rlabel metal3 30576 12936 30576 12936 0 _0019_
rlabel metal2 33320 14224 33320 14224 0 _0020_
rlabel metal2 32312 16912 32312 16912 0 _0021_
rlabel metal2 33544 19544 33544 19544 0 _0022_
rlabel metal2 28168 20356 28168 20356 0 _0023_
rlabel metal2 27664 13160 27664 13160 0 _0024_
rlabel metal2 23912 13160 23912 13160 0 _0025_
rlabel metal2 27328 16184 27328 16184 0 _0026_
rlabel metal2 25928 19544 25928 19544 0 _0027_
rlabel metal3 31304 21448 31304 21448 0 _0028_
rlabel metal2 5880 10668 5880 10668 0 _0029_
rlabel metal3 4536 12264 4536 12264 0 _0030_
rlabel metal2 5768 9520 5768 9520 0 _0031_
rlabel metal2 7896 6440 7896 6440 0 _0032_
rlabel metal2 3976 6524 3976 6524 0 _0033_
rlabel metal2 2800 5488 2800 5488 0 _0034_
rlabel metal2 23912 20272 23912 20272 0 _0035_
rlabel metal2 23352 21784 23352 21784 0 _0036_
rlabel metal2 2688 22568 2688 22568 0 _0037_
rlabel metal2 2688 24920 2688 24920 0 _0038_
rlabel metal2 4872 25928 4872 25928 0 _0039_
rlabel metal2 11872 21784 11872 21784 0 _0040_
rlabel metal2 8344 27384 8344 27384 0 _0041_
rlabel metal3 6552 26936 6552 26936 0 _0042_
rlabel metal2 10976 25592 10976 25592 0 _0043_
rlabel metal2 17528 25928 17528 25928 0 _0044_
rlabel metal3 24920 24024 24920 24024 0 _0045_
rlabel metal2 28728 23408 28728 23408 0 _0046_
rlabel metal2 29736 25200 29736 25200 0 _0047_
rlabel metal2 26264 26488 26264 26488 0 _0048_
rlabel metal2 27944 30520 27944 30520 0 _0049_
rlabel metal3 24024 30856 24024 30856 0 _0050_
rlabel metal2 22736 28840 22736 28840 0 _0051_
rlabel metal3 21784 27160 21784 27160 0 _0052_
rlabel metal2 21000 25144 21000 25144 0 _0053_
rlabel metal2 10696 19488 10696 19488 0 _0054_
rlabel metal2 10248 17136 10248 17136 0 _0055_
rlabel metal2 14952 20888 14952 20888 0 _0056_
rlabel metal2 16184 16408 16184 16408 0 _0057_
rlabel metal2 22344 16240 22344 16240 0 _0058_
rlabel metal2 19824 15288 19824 15288 0 _0059_
rlabel metal2 19768 20356 19768 20356 0 _0060_
rlabel metal2 22232 18816 22232 18816 0 _0061_
rlabel metal2 14896 23128 14896 23128 0 _0062_
rlabel metal2 21896 12376 21896 12376 0 _0063_
rlabel metal2 11704 29736 11704 29736 0 _0064_
rlabel metal2 11144 28112 11144 28112 0 _0065_
rlabel metal2 13160 31416 13160 31416 0 _0066_
rlabel metal2 14840 27440 14840 27440 0 _0067_
rlabel metal2 14840 31248 14840 31248 0 _0068_
rlabel metal2 21112 28952 21112 28952 0 _0069_
rlabel metal2 20552 31416 20552 31416 0 _0070_
rlabel metal2 21336 16912 21336 16912 0 _0071_
rlabel metal2 22792 17584 22792 17584 0 _0072_
rlabel metal2 21392 19124 21392 19124 0 _0073_
rlabel metal2 19656 18340 19656 18340 0 _0074_
rlabel metal3 18340 17864 18340 17864 0 _0075_
rlabel metal3 18368 15512 18368 15512 0 _0076_
rlabel metal2 17640 29288 17640 29288 0 _0077_
rlabel metal2 17192 27776 17192 27776 0 _0078_
rlabel metal2 12712 27459 12712 27459 0 _0079_
rlabel metal2 15456 29120 15456 29120 0 _0080_
rlabel metal3 15624 27048 15624 27048 0 _0081_
rlabel metal2 16352 24696 16352 24696 0 _0082_
rlabel metal2 19656 24276 19656 24276 0 _0083_
rlabel metal2 24080 26264 24080 26264 0 _0084_
rlabel metal3 26096 25480 26096 25480 0 _0085_
rlabel metal2 23744 24024 23744 24024 0 _0086_
rlabel metal2 18200 22736 18200 22736 0 _0087_
rlabel metal2 22120 24864 22120 24864 0 _0088_
rlabel metal2 19208 22988 19208 22988 0 _0089_
rlabel metal2 17808 22988 17808 22988 0 _0090_
rlabel metal2 17640 22492 17640 22492 0 _0091_
rlabel metal2 16268 20552 16268 20552 0 _0092_
rlabel metal2 16632 19264 16632 19264 0 _0093_
rlabel metal3 17612 19208 17612 19208 0 _0094_
rlabel metal3 18172 21784 18172 21784 0 _0095_
rlabel metal2 17304 21168 17304 21168 0 _0096_
rlabel metal3 16520 15176 16520 15176 0 _0097_
rlabel metal2 17752 13608 17752 13608 0 _0098_
rlabel metal2 16408 10640 16408 10640 0 _0099_
rlabel metal2 15960 10256 15960 10256 0 _0100_
rlabel metal2 11256 6048 11256 6048 0 _0101_
rlabel metal2 11592 5292 11592 5292 0 _0102_
rlabel metal3 11424 5880 11424 5880 0 _0103_
rlabel metal3 12264 6104 12264 6104 0 _0104_
rlabel metal2 17920 12852 17920 12852 0 _0105_
rlabel metal2 16924 11573 16924 11573 0 _0106_
rlabel metal2 18984 12208 18984 12208 0 _0107_
rlabel metal2 16156 11368 16156 11368 0 _0108_
rlabel metal2 14840 11088 14840 11088 0 _0109_
rlabel metal2 12824 7336 12824 7336 0 _0110_
rlabel metal2 5096 12880 5096 12880 0 _0111_
rlabel metal2 24584 25536 24584 25536 0 _0112_
rlabel metal3 18312 21336 18312 21336 0 _0113_
rlabel metal2 18088 13048 18088 13048 0 _0114_
rlabel metal3 18424 12152 18424 12152 0 _0115_
rlabel metal2 17248 5880 17248 5880 0 _0116_
rlabel metal2 16464 6048 16464 6048 0 _0117_
rlabel metal2 18088 4956 18088 4956 0 _0118_
rlabel metal2 19656 5768 19656 5768 0 _0119_
rlabel metal2 17976 16856 17976 16856 0 _0120_
rlabel metal2 17640 6552 17640 6552 0 _0121_
rlabel metal2 15064 6272 15064 6272 0 _0122_
rlabel metal2 11592 6272 11592 6272 0 _0123_
rlabel metal2 6834 5152 6834 5152 0 _0124_
rlabel metal2 8120 5320 8120 5320 0 _0125_
rlabel metal2 18200 12880 18200 12880 0 _0126_
rlabel metal3 18032 12936 18032 12936 0 _0127_
rlabel metal2 14504 11312 14504 11312 0 _0128_
rlabel metal2 12824 10662 12824 10662 0 _0129_
rlabel metal3 4872 6048 4872 6048 0 _0130_
rlabel metal2 12936 10584 12936 10584 0 _0131_
rlabel metal2 7000 4984 7000 4984 0 _0132_
rlabel metal2 11014 4984 11014 4984 0 _0133_
rlabel metal2 18940 5955 18940 5955 0 _0134_
rlabel metal2 18200 5824 18200 5824 0 _0135_
rlabel metal2 17080 6328 17080 6328 0 _0136_
rlabel metal2 11928 5768 11928 5768 0 _0137_
rlabel metal2 12376 5040 12376 5040 0 _0138_
rlabel metal2 13328 6216 13328 6216 0 _0139_
rlabel metal2 5636 4452 5636 4452 0 _0140_
rlabel metal3 5208 3528 5208 3528 0 _0141_
rlabel metal2 3640 4872 3640 4872 0 _0142_
rlabel metal3 4900 6664 4900 6664 0 _0143_
rlabel metal2 6274 5768 6274 5768 0 _0144_
rlabel metal3 4648 5880 4648 5880 0 _0145_
rlabel metal2 16072 8680 16072 8680 0 _0146_
rlabel metal2 13608 9464 13608 9464 0 _0147_
rlabel metal2 4984 7317 4984 7317 0 _0148_
rlabel metal2 7896 7280 7896 7280 0 _0149_
rlabel metal2 14616 6944 14616 6944 0 _0150_
rlabel metal2 14896 6496 14896 6496 0 _0151_
rlabel metal3 12992 11592 12992 11592 0 _0152_
rlabel metal3 11452 12152 11452 12152 0 _0153_
rlabel metal2 5768 12984 5768 12984 0 _0154_
rlabel metal3 9940 9800 9940 9800 0 _0155_
rlabel metal3 12880 7784 12880 7784 0 _0156_
rlabel metal3 13412 6664 13412 6664 0 _0157_
rlabel metal3 14140 6888 14140 6888 0 _0158_
rlabel metal2 7896 8064 7896 8064 0 _0159_
rlabel metal2 3808 5096 3808 5096 0 _0160_
rlabel metal3 12432 8232 12432 8232 0 _0161_
rlabel metal3 11452 6888 11452 6888 0 _0162_
rlabel metal2 10360 13048 10360 13048 0 _0163_
rlabel via2 8008 12170 8008 12170 0 _0164_
rlabel metal2 11480 7924 11480 7924 0 _0165_
rlabel metal2 11592 7812 11592 7812 0 _0166_
rlabel metal2 13944 8120 13944 8120 0 _0167_
rlabel metal2 14896 7728 14896 7728 0 _0168_
rlabel metal4 8120 6272 8120 6272 0 _0169_
rlabel metal2 7784 5544 7784 5544 0 _0170_
rlabel metal2 4816 5096 4816 5096 0 _0171_
rlabel metal3 6272 5992 6272 5992 0 _0172_
rlabel metal2 8288 6580 8288 6580 0 _0173_
rlabel via1 8017 5992 8017 5992 0 _0174_
rlabel metal2 7336 9632 7336 9632 0 _0175_
rlabel metal2 5768 9996 5768 9996 0 _0176_
rlabel metal3 5040 12936 5040 12936 0 _0177_
rlabel metal3 6944 9016 6944 9016 0 _0178_
rlabel metal2 7840 8904 7840 8904 0 _0179_
rlabel metal2 10136 10976 10136 10976 0 _0180_
rlabel metal2 4032 7448 4032 7448 0 _0181_
rlabel metal3 9576 7336 9576 7336 0 _0182_
rlabel metal2 8680 9352 8680 9352 0 _0183_
rlabel metal2 7336 4928 7336 4928 0 _0184_
rlabel metal2 8120 7056 8120 7056 0 _0185_
rlabel metal2 8344 8820 8344 8820 0 _0186_
rlabel metal2 8344 9408 8344 9408 0 _0187_
rlabel metal2 8064 10080 8064 10080 0 _0188_
rlabel metal2 7000 11630 7000 11630 0 _0189_
rlabel metal2 3920 8316 3920 8316 0 _0190_
rlabel metal2 4760 10108 4760 10108 0 _0191_
rlabel metal2 7112 11284 7112 11284 0 _0192_
rlabel metal2 3304 12110 3304 12110 0 _0193_
rlabel via1 7336 11354 7336 11354 0 _0194_
rlabel metal2 7364 7560 7364 7560 0 _0195_
rlabel metal2 8344 10920 8344 10920 0 _0196_
rlabel metal2 7644 10696 7644 10696 0 _0197_
rlabel via1 3584 9782 3584 9782 0 _0198_
rlabel metal2 4088 9128 4088 9128 0 _0199_
rlabel metal2 3136 10192 3136 10192 0 _0200_
rlabel metal2 4312 10360 4312 10360 0 _0201_
rlabel metal2 3080 13440 3080 13440 0 _0202_
rlabel metal2 3080 8750 3080 8750 0 _0203_
rlabel metal2 2408 13216 2408 13216 0 _0204_
rlabel metal2 2632 13104 2632 13104 0 _0205_
rlabel metal2 2744 13020 2744 13020 0 _0206_
rlabel metal2 4032 12292 4032 12292 0 _0207_
rlabel metal2 3864 11592 3864 11592 0 _0208_
rlabel metal2 3668 11592 3668 11592 0 _0209_
rlabel metal2 4778 12096 4778 12096 0 _0210_
rlabel metal2 5208 13403 5208 13403 0 _0211_
rlabel metal2 4312 13104 4312 13104 0 _0212_
rlabel metal2 3864 6076 3864 6076 0 _0213_
rlabel metal2 3304 7448 3304 7448 0 _0214_
rlabel metal2 3640 5964 3640 5964 0 _0215_
rlabel metal2 3136 6216 3136 6216 0 _0216_
rlabel metal2 6440 5152 6440 5152 0 _0217_
rlabel metal2 10136 5572 10136 5572 0 _0218_
rlabel metal2 5880 5992 5880 5992 0 _0219_
rlabel metal2 3360 8680 3360 8680 0 _0220_
rlabel metal2 3416 6986 3416 6986 0 _0221_
rlabel metal3 3276 6664 3276 6664 0 _0222_
rlabel metal2 4984 5292 4984 5292 0 _0223_
rlabel metal3 16632 11368 16632 11368 0 _0224_
rlabel metal2 7784 13048 7784 13048 0 _0225_
rlabel via2 7000 12922 7000 12922 0 _0226_
rlabel metal2 7000 12376 7000 12376 0 _0227_
rlabel metal2 6468 13160 6468 13160 0 _0228_
rlabel metal2 27132 20664 27132 20664 0 _0229_
rlabel metal2 21840 8232 21840 8232 0 _0230_
rlabel metal2 20328 23240 20328 23240 0 _0231_
rlabel metal2 23240 6048 23240 6048 0 _0232_
rlabel metal2 29792 16940 29792 16940 0 _0233_
rlabel metal2 31752 17556 31752 17556 0 _0234_
rlabel metal2 28616 17276 28616 17276 0 _0235_
rlabel metal3 30520 16856 30520 16856 0 _0236_
rlabel metal2 29736 13496 29736 13496 0 _0237_
rlabel metal2 25704 9128 25704 9128 0 _0238_
rlabel metal2 27272 15120 27272 15120 0 _0239_
rlabel via2 23128 9786 23128 9786 0 _0240_
rlabel metal2 29848 6104 29848 6104 0 _0241_
rlabel metal2 25704 10248 25704 10248 0 _0242_
rlabel metal3 28616 9016 28616 9016 0 _0243_
rlabel metal2 29624 10528 29624 10528 0 _0244_
rlabel metal3 28448 5096 28448 5096 0 _0245_
rlabel metal2 29204 5320 29204 5320 0 _0246_
rlabel metal2 29960 10528 29960 10528 0 _0247_
rlabel metal3 24864 10472 24864 10472 0 _0248_
rlabel metal2 23576 13272 23576 13272 0 _0249_
rlabel metal2 28728 13328 28728 13328 0 _0250_
rlabel metal3 28616 8232 28616 8232 0 _0251_
rlabel metal2 27832 5152 27832 5152 0 _0252_
rlabel metal2 22736 23912 22736 23912 0 _0253_
rlabel metal2 23016 22680 23016 22680 0 _0254_
rlabel metal2 22792 10192 22792 10192 0 _0255_
rlabel metal2 21336 10304 21336 10304 0 _0256_
rlabel metal2 30520 15904 30520 15904 0 _0257_
rlabel metal2 24360 7840 24360 7840 0 _0258_
rlabel metal3 24192 10360 24192 10360 0 _0259_
rlabel metal2 24472 7896 24472 7896 0 _0260_
rlabel metal3 23884 7448 23884 7448 0 _0261_
rlabel metal2 24136 7986 24136 7986 0 _0262_
rlabel metal2 23464 6020 23464 6020 0 _0263_
rlabel metal2 23352 5180 23352 5180 0 _0264_
rlabel metal2 23520 4032 23520 4032 0 _0265_
rlabel metal2 23464 5124 23464 5124 0 _0266_
rlabel metal2 28168 6586 28168 6586 0 _0267_
rlabel metal2 22456 5432 22456 5432 0 _0268_
rlabel metal3 21672 3528 21672 3528 0 _0269_
rlabel metal2 28056 5922 28056 5922 0 _0270_
rlabel metal2 28672 3808 28672 3808 0 _0271_
rlabel metal2 28392 4620 28392 4620 0 _0272_
rlabel metal2 28560 8344 28560 8344 0 _0273_
rlabel metal2 30632 4956 30632 4956 0 _0274_
rlabel metal2 30968 5152 30968 5152 0 _0275_
rlabel metal2 31080 4396 31080 4396 0 _0276_
rlabel metal2 31864 6636 31864 6636 0 _0277_
rlabel via1 30398 6664 30398 6664 0 _0278_
rlabel metal2 32312 6524 32312 6524 0 _0279_
rlabel metal2 30632 6384 30632 6384 0 _0280_
rlabel metal3 29960 6720 29960 6720 0 _0281_
rlabel metal2 28392 9072 28392 9072 0 _0282_
rlabel metal2 29568 8708 29568 8708 0 _0283_
rlabel metal2 29624 9836 29624 9836 0 _0284_
rlabel metal2 28000 9772 28000 9772 0 _0285_
rlabel metal2 29400 9744 29400 9744 0 _0286_
rlabel metal2 27496 11060 27496 11060 0 _0287_
rlabel metal2 32760 10920 32760 10920 0 _0288_
rlabel via2 33656 12928 33656 12928 0 _0289_
rlabel metal2 31976 9996 31976 9996 0 _0290_
rlabel metal2 29176 18424 29176 18424 0 _0291_
rlabel metal2 31640 12460 31640 12460 0 _0292_
rlabel metal3 31640 12152 31640 12152 0 _0293_
rlabel metal2 30296 12880 30296 12880 0 _0294_
rlabel metal2 31864 16450 31864 16450 0 _0295_
rlabel metal2 31080 14174 31080 14174 0 _0296_
rlabel metal2 31752 14952 31752 14952 0 _0297_
rlabel metal2 32984 14000 32984 14000 0 _0298_
rlabel metal2 30940 16632 30940 16632 0 _0299_
rlabel metal2 31080 18424 31080 18424 0 _0300_
rlabel metal2 32480 16212 32480 16212 0 _0301_
rlabel metal2 31864 19180 31864 19180 0 _0302_
rlabel metal2 29512 17584 29512 17584 0 _0303_
rlabel metal2 32200 19068 32200 19068 0 _0304_
rlabel metal2 28840 18885 28840 18885 0 _0305_
rlabel metal2 29232 15288 29232 15288 0 _0306_
rlabel via2 27608 17621 27608 17621 0 _0307_
rlabel metal2 28504 20496 28504 20496 0 _0308_
rlabel metal2 28056 14826 28056 14826 0 _0309_
rlabel metal3 28644 14504 28644 14504 0 _0310_
rlabel metal2 28056 13160 28056 13160 0 _0311_
rlabel metal2 25368 14078 25368 14078 0 _0312_
rlabel metal2 26936 16282 26936 16282 0 _0313_
rlabel metal2 27552 15988 27552 15988 0 _0314_
rlabel metal2 27832 17864 27832 17864 0 _0315_
rlabel metal2 28336 16856 28336 16856 0 _0316_
rlabel metal3 29848 19880 29848 19880 0 _0317_
rlabel metal2 26936 19824 26936 19824 0 _0318_
rlabel metal2 31864 20888 31864 20888 0 _0319_
rlabel metal2 30856 20440 30856 20440 0 _0320_
rlabel metal2 30968 22456 30968 22456 0 _0321_
rlabel metal2 20216 26208 20216 26208 0 _0322_
rlabel metal3 22176 21784 22176 21784 0 _0323_
rlabel metal2 17528 19096 17528 19096 0 _0324_
rlabel metal2 20328 18760 20328 18760 0 _0325_
rlabel metal2 20328 17696 20328 17696 0 _0326_
rlabel metal2 22904 20888 22904 20888 0 _0327_
rlabel metal2 20440 20468 20440 20468 0 _0328_
rlabel metal2 22456 20664 22456 20664 0 _0329_
rlabel metal2 23184 20412 23184 20412 0 _0330_
rlabel metal2 16632 23856 16632 23856 0 _0331_
rlabel metal2 8512 23044 8512 23044 0 _0332_
rlabel metal2 11032 24668 11032 24668 0 _0333_
rlabel metal2 8344 23688 8344 23688 0 _0334_
rlabel metal2 8232 23436 8232 23436 0 _0335_
rlabel metal2 9576 22512 9576 22512 0 _0336_
rlabel metal2 23800 21518 23800 21518 0 _0337_
rlabel metal3 24052 22344 24052 22344 0 _0338_
rlabel metal2 22904 22260 22904 22260 0 _0339_
rlabel metal3 4256 21560 4256 21560 0 _0340_
rlabel metal2 2856 19656 2856 19656 0 _0341_
rlabel metal3 5460 20888 5460 20888 0 _0342_
rlabel metal2 4536 18760 4536 18760 0 _0343_
rlabel metal2 5208 18144 5208 18144 0 _0344_
rlabel metal2 7224 19264 7224 19264 0 _0345_
rlabel metal2 3304 18648 3304 18648 0 _0346_
rlabel metal2 4312 18424 4312 18424 0 _0347_
rlabel metal2 3248 19684 3248 19684 0 _0348_
rlabel metal2 3920 21980 3920 21980 0 _0349_
rlabel metal2 4088 22400 4088 22400 0 _0350_
rlabel metal2 16352 24304 16352 24304 0 _0351_
rlabel metal2 16408 25340 16408 25340 0 _0352_
rlabel metal2 15288 25424 15288 25424 0 _0353_
rlabel metal2 16184 25522 16184 25522 0 _0354_
rlabel metal2 3752 22792 3752 22792 0 _0355_
rlabel metal3 3780 22344 3780 22344 0 _0356_
rlabel metal2 5040 21168 5040 21168 0 _0357_
rlabel metal2 2968 19684 2968 19684 0 _0358_
rlabel metal3 4153 19992 4153 19992 0 _0359_
rlabel metal2 4284 21672 4284 21672 0 _0360_
rlabel metal2 6104 23800 6104 23800 0 _0361_
rlabel metal3 5236 23912 5236 23912 0 _0362_
rlabel metal2 5096 24192 5096 24192 0 _0363_
rlabel metal2 3080 24416 3080 24416 0 _0364_
rlabel metal3 6160 19208 6160 19208 0 _0365_
rlabel metal3 8204 19992 8204 19992 0 _0366_
rlabel metal2 7280 17640 7280 17640 0 _0367_
rlabel metal2 7280 18508 7280 18508 0 _0368_
rlabel metal2 7952 19992 7952 19992 0 _0369_
rlabel metal2 7000 21840 7000 21840 0 _0370_
rlabel metal3 8372 23912 8372 23912 0 _0371_
rlabel metal2 7336 24192 7336 24192 0 _0372_
rlabel metal2 6580 24136 6580 24136 0 _0373_
rlabel metal2 21112 20384 21112 20384 0 _0374_
rlabel metal2 12152 25088 12152 25088 0 _0375_
rlabel metal2 15792 18172 15792 18172 0 _0376_
rlabel metal2 22456 24248 22456 24248 0 _0377_
rlabel metal3 18312 24920 18312 24920 0 _0378_
rlabel metal2 6328 18480 6328 18480 0 _0379_
rlabel metal2 8904 21560 8904 21560 0 _0380_
rlabel metal3 12572 22568 12572 22568 0 _0381_
rlabel metal2 13832 22456 13832 22456 0 _0382_
rlabel metal2 12152 21896 12152 21896 0 _0383_
rlabel metal2 5880 19684 5880 19684 0 _0384_
rlabel metal2 4508 20104 4508 20104 0 _0385_
rlabel metal2 8568 18620 8568 18620 0 _0386_
rlabel metal2 9016 22008 9016 22008 0 _0387_
rlabel metal2 5600 19880 5600 19880 0 _0388_
rlabel metal2 6412 21000 6412 21000 0 _0389_
rlabel metal2 8008 24864 8008 24864 0 _0390_
rlabel metal2 7560 24752 7560 24752 0 _0391_
rlabel metal3 8148 24696 8148 24696 0 _0392_
rlabel metal2 6748 18536 6748 18536 0 _0393_
rlabel metal2 7644 19432 7644 19432 0 _0394_
rlabel metal2 7672 22036 7672 22036 0 _0395_
rlabel metal2 8120 25536 8120 25536 0 _0396_
rlabel metal2 8540 25480 8540 25480 0 _0397_
rlabel metal2 7392 27048 7392 27048 0 _0398_
rlabel metal2 7560 22605 7560 22605 0 _0399_
rlabel metal3 8344 22344 8344 22344 0 _0400_
rlabel metal2 9268 22456 9268 22456 0 _0401_
rlabel metal2 21224 17528 21224 17528 0 _0402_
rlabel metal2 12403 23912 12403 23912 0 _0403_
rlabel metal2 11704 24360 11704 24360 0 _0404_
rlabel metal2 12768 24864 12768 24864 0 _0405_
rlabel metal2 17052 25480 17052 25480 0 _0406_
rlabel metal3 23464 24584 23464 24584 0 _0407_
rlabel metal2 24360 24752 24360 24752 0 _0408_
rlabel metal2 24472 24668 24472 24668 0 _0409_
rlabel metal2 27272 23716 27272 23716 0 _0410_
rlabel metal2 28616 26342 28616 26342 0 _0411_
rlabel metal2 28504 23828 28504 23828 0 _0412_
rlabel metal2 28616 25452 28616 25452 0 _0413_
rlabel metal3 29316 26040 29316 26040 0 _0414_
rlabel metal2 29064 24780 29064 24780 0 _0415_
rlabel metal2 23296 29400 23296 29400 0 _0416_
rlabel metal2 27384 26152 27384 26152 0 _0417_
rlabel metal2 27496 28000 27496 28000 0 _0418_
rlabel metal2 26992 26264 26992 26264 0 _0419_
rlabel metal2 27272 29077 27272 29077 0 _0420_
rlabel metal2 28728 28168 28728 28168 0 _0421_
rlabel metal3 28336 29400 28336 29400 0 _0422_
rlabel metal2 27272 30744 27272 30744 0 _0423_
rlabel metal2 25704 28000 25704 28000 0 _0424_
rlabel metal2 24920 30072 24920 30072 0 _0425_
rlabel metal2 25760 30968 25760 30968 0 _0426_
rlabel metal2 23688 29357 23688 29357 0 _0427_
rlabel metal2 24024 29736 24024 29736 0 _0428_
rlabel metal2 23408 28616 23408 28616 0 _0429_
rlabel metal3 21980 27048 21980 27048 0 _0430_
rlabel metal2 20888 26600 20888 26600 0 _0431_
rlabel metal3 21448 26264 21448 26264 0 _0432_
rlabel metal2 21308 26376 21308 26376 0 _0433_
rlabel metal2 20748 24136 20748 24136 0 _0434_
rlabel metal2 16128 18424 16128 18424 0 _0435_
rlabel metal2 12992 19992 12992 19992 0 _0436_
rlabel metal2 11760 19208 11760 19208 0 _0437_
rlabel metal3 12292 17640 12292 17640 0 _0438_
rlabel via1 12161 17864 12161 17864 0 _0439_
rlabel metal2 11592 19544 11592 19544 0 _0440_
rlabel metal2 11172 19208 11172 19208 0 _0441_
rlabel metal2 18368 15428 18368 15428 0 _0442_
rlabel metal2 12712 17192 12712 17192 0 _0443_
rlabel metal2 13328 18228 13328 18228 0 _0444_
rlabel metal2 15624 18480 15624 18480 0 _0445_
rlabel metal2 15288 17920 15288 17920 0 _0446_
rlabel metal2 10920 17584 10920 17584 0 _0447_
rlabel metal2 14448 20608 14448 20608 0 _0448_
rlabel metal2 15512 20468 15512 20468 0 _0449_
rlabel metal2 15176 20446 15176 20446 0 _0450_
rlabel metal3 13272 19208 13272 19208 0 _0451_
rlabel metal2 13776 17780 13776 17780 0 _0452_
rlabel metal2 14504 16408 14504 16408 0 _0453_
rlabel metal2 15232 15624 15232 15624 0 _0454_
rlabel metal2 15260 16856 15260 16856 0 _0455_
rlabel metal2 21728 16968 21728 16968 0 _0456_
rlabel metal2 18536 17080 18536 17080 0 _0457_
rlabel metal2 19292 16856 19292 16856 0 _0458_
rlabel metal3 22232 20776 22232 20776 0 _0459_
rlabel metal3 20748 20776 20748 20776 0 _0460_
rlabel metal2 23072 16968 23072 16968 0 _0461_
rlabel metal2 22064 18368 22064 18368 0 _0462_
rlabel metal2 14616 25424 14616 25424 0 _0463_
rlabel metal3 22008 13160 22008 13160 0 _0464_
rlabel metal2 21756 13720 21756 13720 0 _0465_
rlabel metal2 18984 28896 18984 28896 0 _0466_
rlabel metal3 20412 30072 20412 30072 0 _0467_
rlabel metal3 13524 29176 13524 29176 0 _0468_
rlabel metal3 11928 27832 11928 27832 0 _0469_
rlabel metal2 13496 30184 13496 30184 0 _0470_
rlabel metal2 15960 29478 15960 29478 0 _0471_
rlabel metal2 14952 28784 14952 28784 0 _0472_
rlabel metal2 14952 27488 14952 27488 0 _0473_
rlabel metal2 16072 29848 16072 29848 0 _0474_
rlabel metal2 20216 29512 20216 29512 0 _0475_
rlabel metal2 16240 31752 16240 31752 0 _0476_
rlabel metal2 19208 29357 19208 29357 0 _0477_
rlabel metal2 19544 29456 19544 29456 0 _0478_
rlabel metal2 19656 29484 19656 29484 0 _0479_
rlabel metal2 19992 30520 19992 30520 0 _0480_
rlabel metal3 28476 20776 28476 20776 0 clknet_0_wb_clk_i
rlabel metal2 5740 3640 5740 3640 0 clknet_3_0__leaf_wb_clk_i
rlabel metal2 13832 5208 13832 5208 0 clknet_3_1__leaf_wb_clk_i
rlabel metal2 2296 25760 2296 25760 0 clknet_3_2__leaf_wb_clk_i
rlabel metal2 14168 27832 14168 27832 0 clknet_3_3__leaf_wb_clk_i
rlabel metal3 22932 15176 22932 15176 0 clknet_3_4__leaf_wb_clk_i
rlabel metal2 31024 5712 31024 5712 0 clknet_3_5__leaf_wb_clk_i
rlabel metal2 23464 20720 23464 20720 0 clknet_3_6__leaf_wb_clk_i
rlabel metal2 29036 30184 29036 30184 0 clknet_3_7__leaf_wb_clk_i
rlabel metal2 26264 24472 26264 24472 0 clock_div\[0\]
rlabel metal3 27048 23912 27048 23912 0 clock_div\[1\]
rlabel metal3 28672 25368 28672 25368 0 clock_div\[2\]
rlabel metal2 28504 28000 28504 28000 0 clock_div\[3\]
rlabel metal2 26712 28672 26712 28672 0 clock_div\[4\]
rlabel metal2 24528 28616 24528 28616 0 clock_div\[5\]
rlabel metal2 24136 28994 24136 28994 0 clock_div\[6\]
rlabel metal2 23912 27496 23912 27496 0 clock_div\[7\]
rlabel metal2 18424 24752 18424 24752 0 clock_div\[8\]
rlabel metal3 22456 7560 22456 7560 0 counter\[0\]
rlabel metal2 32088 8316 32088 8316 0 counter\[10\]
rlabel metal2 28616 10136 28616 10136 0 counter\[11\]
rlabel via2 30968 10591 30968 10591 0 counter\[12\]
rlabel metal2 31752 13552 31752 13552 0 counter\[13\]
rlabel metal3 31304 14392 31304 14392 0 counter\[14\]
rlabel metal2 31640 18088 31640 18088 0 counter\[15\]
rlabel metal2 32312 19544 32312 19544 0 counter\[16\]
rlabel metal2 29680 19208 29680 19208 0 counter\[17\]
rlabel metal2 29176 14056 29176 14056 0 counter\[18\]
rlabel metal2 26936 14000 26936 14000 0 counter\[19\]
rlabel metal2 22456 8120 22456 8120 0 counter\[1\]
rlabel metal3 27076 16072 27076 16072 0 counter\[20\]
rlabel metal2 28504 17248 28504 17248 0 counter\[21\]
rlabel metal3 29736 21560 29736 21560 0 counter\[22\]
rlabel metal2 24808 9912 24808 9912 0 counter\[2\]
rlabel metal2 25368 7896 25368 7896 0 counter\[3\]
rlabel metal2 25480 5488 25480 5488 0 counter\[4\]
rlabel metal2 22344 4872 22344 4872 0 counter\[5\]
rlabel metal2 30072 5964 30072 5964 0 counter\[6\]
rlabel metal2 30408 5824 30408 5824 0 counter\[7\]
rlabel metal3 30576 7448 30576 7448 0 counter\[8\]
rlabel metal2 29512 6608 29512 6608 0 counter\[9\]
rlabel metal2 17976 1190 17976 1190 0 io_out[0]
rlabel metal3 25760 3640 25760 3640 0 io_out[1]
rlabel metal2 32312 1414 32312 1414 0 io_out[2]
rlabel metal3 24388 20776 24388 20776 0 just_inc
rlabel metal2 18930 22036 18930 22036 0 just_rst
rlabel metal2 13384 29008 13384 29008 0 master_clk_div\[0\]
rlabel metal2 12712 29071 12712 29071 0 master_clk_div\[1\]
rlabel metal2 14728 30128 14728 30128 0 master_clk_div\[2\]
rlabel metal3 14840 28616 14840 28616 0 master_clk_div\[3\]
rlabel metal2 16856 29792 16856 29792 0 master_clk_div\[4\]
rlabel metal2 18200 29288 18200 29288 0 master_clk_div\[5\]
rlabel metal2 18760 30184 18760 30184 0 master_clk_div\[6\]
rlabel metal2 4872 3472 4872 3472 0 net1
rlabel metal2 20104 4186 20104 4186 0 net2
rlabel metal2 25480 3794 25480 3794 0 net3
rlabel metal2 32536 4437 32536 4437 0 net4
rlabel metal2 25144 6944 25144 6944 0 net5
rlabel metal2 16072 25452 16072 25452 0 prev_clk_div
rlabel metal2 12208 19880 12208 19880 0 rhythm_LFSR\[0\]
rlabel metal2 12152 19292 12152 19292 0 rhythm_LFSR\[1\]
rlabel metal2 16408 20776 16408 20776 0 rhythm_LFSR\[2\]
rlabel metal2 14280 16912 14280 16912 0 rhythm_LFSR\[3\]
rlabel metal2 10780 3416 10780 3416 0 rst_n
rlabel metal2 19992 11984 19992 11984 0 slow_blink
rlabel metal2 22884 16800 22884 16800 0 tempo_LFSR\[0\]
rlabel metal2 21924 16856 21924 16856 0 tempo_LFSR\[1\]
rlabel metal2 21952 20440 21952 20440 0 tempo_LFSR\[2\]
rlabel metal2 21952 19320 21952 19320 0 tempo_LFSR\[3\]
rlabel metal2 18984 9968 18984 9968 0 tune_ROM\[0\]
rlabel metal3 13841 16856 13841 16856 0 tune_ROM\[1\]
rlabel metal3 6048 17640 6048 17640 0 tune_ROM\[2\]
rlabel metal2 4088 17752 4088 17752 0 tune_ROM\[3\]
rlabel metal2 4648 16968 4648 16968 0 tune_ROM\[4\]
rlabel metal2 2632 18816 2632 18816 0 tune_ROM\[5\]
rlabel metal2 3640 2478 3640 2478 0 wb_clk_i
<< properties >>
string FIXED_BBOX 0 0 36000 36000
<< end >>
