module diceroll (io_in,
    rst_n,
    vdd,
    vss,
    wb_clk_i,
    io_out);
 input io_in;
 input rst_n;
 inout vdd;
 inout vss;
 input wb_clk_i;
 output [8:0] io_out;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire _247_;
 wire _248_;
 wire _249_;
 wire _250_;
 wire _251_;
 wire _252_;
 wire _253_;
 wire _254_;
 wire _255_;
 wire _256_;
 wire _257_;
 wire _258_;
 wire _259_;
 wire _260_;
 wire _261_;
 wire _262_;
 wire _263_;
 wire _264_;
 wire _265_;
 wire _266_;
 wire _267_;
 wire _268_;
 wire _269_;
 wire _270_;
 wire _271_;
 wire _272_;
 wire _273_;
 wire _274_;
 wire _275_;
 wire _276_;
 wire _277_;
 wire _278_;
 wire _279_;
 wire _280_;
 wire _281_;
 wire _282_;
 wire _283_;
 wire _284_;
 wire _285_;
 wire _286_;
 wire _287_;
 wire _288_;
 wire _289_;
 wire _290_;
 wire _291_;
 wire _292_;
 wire _293_;
 wire _294_;
 wire _295_;
 wire _296_;
 wire _297_;
 wire _298_;
 wire _299_;
 wire _300_;
 wire _301_;
 wire _302_;
 wire _303_;
 wire _304_;
 wire _305_;
 wire _306_;
 wire _307_;
 wire _308_;
 wire _309_;
 wire _310_;
 wire _311_;
 wire _312_;
 wire _313_;
 wire _314_;
 wire _315_;
 wire _316_;
 wire _317_;
 wire _318_;
 wire _319_;
 wire _320_;
 wire _321_;
 wire _322_;
 wire _323_;
 wire _324_;
 wire _325_;
 wire _326_;
 wire _327_;
 wire _328_;
 wire _329_;
 wire _330_;
 wire _331_;
 wire _332_;
 wire _333_;
 wire _334_;
 wire _335_;
 wire _336_;
 wire _337_;
 wire _338_;
 wire _339_;
 wire _340_;
 wire _341_;
 wire _342_;
 wire _343_;
 wire _344_;
 wire _345_;
 wire _346_;
 wire _347_;
 wire _348_;
 wire _349_;
 wire _350_;
 wire _351_;
 wire _352_;
 wire _353_;
 wire _354_;
 wire _355_;
 wire _356_;
 wire _357_;
 wire _358_;
 wire _359_;
 wire _360_;
 wire _361_;
 wire _362_;
 wire _363_;
 wire _364_;
 wire _365_;
 wire _366_;
 wire \bcd[0] ;
 wire \bcd[1] ;
 wire \bcd[2] ;
 wire \clkdiv[0] ;
 wire \clkdiv[1] ;
 wire \clkdiv[2] ;
 wire \clkdiv[3] ;
 wire \clkdiv[4] ;
 wire \clkdiv[5] ;
 wire \clkdiv[6] ;
 wire \clkdiv[7] ;
 wire clknet_0_wb_clk_i;
 wire clknet_3_0__leaf_wb_clk_i;
 wire clknet_3_1__leaf_wb_clk_i;
 wire clknet_3_2__leaf_wb_clk_i;
 wire clknet_3_3__leaf_wb_clk_i;
 wire clknet_3_4__leaf_wb_clk_i;
 wire clknet_3_5__leaf_wb_clk_i;
 wire clknet_3_6__leaf_wb_clk_i;
 wire clknet_3_7__leaf_wb_clk_i;
 wire \counter[0] ;
 wire \counter[10] ;
 wire \counter[11] ;
 wire \counter[12] ;
 wire \counter[13] ;
 wire \counter[14] ;
 wire \counter[15] ;
 wire \counter[1] ;
 wire \counter[2] ;
 wire \counter[3] ;
 wire \counter[4] ;
 wire \counter[5] ;
 wire \counter[6] ;
 wire \counter[7] ;
 wire \counter[8] ;
 wire \counter[9] ;
 wire dp;
 wire \lfsr[0] ;
 wire \lfsr[10] ;
 wire \lfsr[11] ;
 wire \lfsr[12] ;
 wire \lfsr[13] ;
 wire \lfsr[14] ;
 wire \lfsr[15] ;
 wire \lfsr[1] ;
 wire \lfsr[2] ;
 wire \lfsr[3] ;
 wire \lfsr[4] ;
 wire \lfsr[5] ;
 wire \lfsr[6] ;
 wire \lfsr[7] ;
 wire \lfsr[8] ;
 wire \lfsr[9] ;
 wire \m_clkdiv[0] ;
 wire \m_clkdiv[1] ;
 wire \m_clkdiv[2] ;
 wire \m_clkdiv[3] ;
 wire \m_clkdiv[4] ;
 wire \m_clkdiv[5] ;
 wire \m_clkdiv[6] ;
 wire \m_clkdiv[7] ;
 wire \m_clkdiv[8] ;
 wire \m_clkdiv[9] ;
 wire net1;
 wire net10;
 wire net11;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire \r_counter[0] ;
 wire \r_counter[1] ;
 wire \r_counter[2] ;

 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__367__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(net2));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__385__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(\clkdiv[0] ));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__399__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_091_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__400__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(net1));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__406__B (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(\clkdiv[0] ));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__409__D (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_105_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__429__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_064_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__432__B (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_105_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__434__B (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_129_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__436__B (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_128_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__442__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(net2));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__447__C (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_142_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__452__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_142_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__456__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_146_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__471__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_157_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__472__B (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_158_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__474__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_064_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__476__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_161_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__480__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_158_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__484__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_161_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__494__C (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_175_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__498__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_158_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__502__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_158_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__510__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_161_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__512__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_091_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__514__B (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_190_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__519__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_190_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__521__D (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_157_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__525__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_190_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__526__D (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_146_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__529__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(\lfsr[3] ));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__530__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_142_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__531__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_205_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__536__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(\lfsr[3] ));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__542__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_157_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__546__B (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_217_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__547__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_214_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__564__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_190_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__565__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_129_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__573__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_129_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__577__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_129_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__584__D (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_175_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__588__B (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_128_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__589__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(net1));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__593__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_214_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__598__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_064_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__602__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_258_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__606__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_258_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__608__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_064_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__610__B (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_205_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__611__B (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_267_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__611__D (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_268_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__618__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_258_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__620__B (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_267_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__620__C (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_268_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__625__C (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_258_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__628__B (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_268_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__634__D (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_286_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__635__C (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_286_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__641__B (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_091_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__641__D (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_142_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__642__C (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_293_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__644__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_293_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__660__D (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_293_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__664__B (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_293_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__672__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(\clkdiv[0] ));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__675__B (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_319_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__676__C (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_157_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__682__B (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_128_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__682__D (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_175_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__683__B (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_319_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__684__B (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_128_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__689__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_161_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__692__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_146_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__693__B (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_267_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__699__B (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_319_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__701__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_214_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__706__C (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_205_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__711__B (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_267_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__715__D (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_205_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__716__B (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_319_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__718__B (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_217_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__719__B (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_217_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__720__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_214_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__727__D (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_175_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__729__B (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_105_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__731__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_217_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__731__C (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_146_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__732__C (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(_365_));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__736__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_3_6__leaf_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__737__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_3_6__leaf_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__738__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_3_6__leaf_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__739__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_3_7__leaf_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__741__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_3_1__leaf_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__742__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_3_1__leaf_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__743__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_3_1__leaf_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__744__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_3_1__leaf_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__745__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_3_4__leaf_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__746__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_3_4__leaf_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__747__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_3_4__leaf_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__748__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_3_5__leaf_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__749__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_3_5__leaf_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__750__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_3_4__leaf_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__751__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_3_7__leaf_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__752__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_3_6__leaf_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__753__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_3_6__leaf_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__754__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_3_5__leaf_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__755__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_3_7__leaf_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__756__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_3_5__leaf_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__757__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_3_7__leaf_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__758__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_3_5__leaf_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__759__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_3_5__leaf_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__760__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_3_5__leaf_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__761__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_3_5__leaf_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__762__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_3_5__leaf_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__763__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_3_5__leaf_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__764__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_3_7__leaf_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__765__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_3_7__leaf_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__766__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_3_7__leaf_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__767__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_3_7__leaf_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__768__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_3_7__leaf_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__769__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_3_6__leaf_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__770__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_3_0__leaf_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__771__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_3_0__leaf_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__772__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_3_2__leaf_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__773__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_3_2__leaf_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__774__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_3_2__leaf_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__775__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_3_2__leaf_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__776__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_3_2__leaf_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__777__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_3_2__leaf_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__778__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_3_1__leaf_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__779__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_3_0__leaf_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__780__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_3_0__leaf_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__781__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_3_0__leaf_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__782__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_3_0__leaf_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__783__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_3_0__leaf_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__784__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_3_1__leaf_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__785__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_3_0__leaf_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__786__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_3_4__leaf_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__787__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_3_6__leaf_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__788__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_3_1__leaf_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__789__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_3_2__leaf_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__791__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_3_6__leaf_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__794__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_3_4__leaf_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__795__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_3_4__leaf_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__796__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_3_4__leaf_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__797__CLK (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_3_7__leaf_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA__799__A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(\lfsr[3] ));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA_clkbuf_0_wb_clk_i_A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA_clkbuf_3_0__f_wb_clk_i_A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA_clkbuf_3_1__f_wb_clk_i_A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA_clkbuf_3_2__f_wb_clk_i_A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA_clkbuf_3_3__f_wb_clk_i_A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA_clkbuf_3_4__f_wb_clk_i_A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA_clkbuf_3_5__f_wb_clk_i_A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA_clkbuf_3_6__f_wb_clk_i_A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA_clkbuf_3_7__f_wb_clk_i_A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA_clkload0_A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_3_0__leaf_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA_clkload1_A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_3_1__leaf_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA_clkload2_A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_3_2__leaf_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA_clkload4_A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_3_4__leaf_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA_clkload5_A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(clknet_3_6__leaf_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA_input1_A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(io_in));
 gf180mcu_as_sc_mcu7t3v3__diode_2 ANTENNA_input2_A (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .DIODE(rst_n));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_0_104 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_0_120 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_0_138 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_0_154 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_0_172 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_0_18 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_0_188 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_0_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_0_206 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_0_222 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_0_240 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_0_256 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_0_274 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_0_290 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_0_308 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_0_324 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_0_342 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_0_358 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_0_36 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_0_376 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_0_52 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_0_70 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_0_86 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_10_102 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_10_104 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_10_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_10_123 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_10_139 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_10_155 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_10_170 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_10_174 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_10_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_10_18 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_10_193 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_10_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_10_209 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_10_225 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_10_233 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_10_243 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_10_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_10_25 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_10_263 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_10_279 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_10_295 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_10_311 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_10_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_10_325 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_10_329 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_10_33 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_10_336 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_10_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_10_381 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_10_383 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_10_45 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_10_58 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_10_74 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_10_90 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_10_98 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_11_113 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_11_129 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_11_137 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_11_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_11_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_11_181 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_11_197 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_11_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_11_205 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_11_209 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_11_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_11_228 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_11_244 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_11_260 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_11_276 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_11_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_11_298 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_11_314 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_11_330 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_11_342 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_11_35 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_11_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_11_354 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_11_361 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_11_377 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_11_381 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_11_383 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_11_39 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_11_55 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_11_6 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_11_63 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_11_67 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_11_69 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_11_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_11_88 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_11_96 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_11_98 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_12_111 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_12_115 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_12_131 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_12_139 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_12_143 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_12_173 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_12_18 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_12_188 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_12_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_12_204 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_12_220 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_12_236 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_12_244 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_12_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_12_263 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_12_279 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_12_287 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_12_291 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_12_293 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_12_300 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_12_308 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_12_312 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_12_314 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_12_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_12_325 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_12_327 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_12_335 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_12_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_12_353 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_12_369 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_12_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_12_377 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_12_381 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_12_383 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_12_45 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_12_49 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_12_74 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_12_82 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_12_86 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_13_125 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_13_129 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_13_137 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_13_139 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_13_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_13_158 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_13_18 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_13_183 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_13_199 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_13_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_13_207 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_13_209 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_13_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_13_228 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_13_244 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_13_260 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_13_276 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_13_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_13_286 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_13_315 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_13_319 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_13_335 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_13_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_13_343 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_13_347 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_13_349 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_13_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_13_368 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_13_50 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_13_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_13_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_13_80 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_14_101 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_14_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_14_140 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_14_144 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_14_160 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_14_168 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_14_171 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_14_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_14_18 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_14_193 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_14_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_14_201 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_14_205 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_14_207 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_14_214 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_14_218 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_14_226 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_14_235 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_14_241 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_14_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_14_253 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_14_281 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_14_285 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_14_302 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_14_310 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_14_314 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_14_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_14_325 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_14_329 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_14_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_14_341 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_14_345 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_14_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_14_382 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_14_60 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_14_78 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_15_101 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_15_105 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_15_109 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_15_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_15_146 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_15_162 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_15_178 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_15_18 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_15_194 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_15_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_15_246 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_15_251 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_15_26 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_15_276 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_15_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_15_290 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_15_292 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_15_302 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_15_318 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_15_336 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_15_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_15_368 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_15_55 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_15_59 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_15_67 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_15_69 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_16_101 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_16_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_16_115 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_16_119 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_16_127 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_16_143 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_16_159 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_16_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_16_18 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_16_181 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_16_189 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_16_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_16_201 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_16_209 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_16_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_16_228 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_16_272 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_16_288 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_16_304 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_16_312 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_16_314 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_16_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_16_333 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_16_335 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_16_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_16_342 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_16_358 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_16_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_16_374 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_16_382 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_16_53 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_16_69 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_16_85 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_17_104 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_17_112 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_17_116 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_17_124 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_17_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_17_158 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_17_166 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_17_168 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_17_179 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_17_18 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_17_189 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_17_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_17_205 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_17_209 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_17_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_17_228 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_17_236 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_17_251 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_17_267 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_17_275 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_17_279 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_17_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_17_286 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_17_296 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_17_312 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_17_320 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_17_324 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_17_332 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_17_334 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_17_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_17_345 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_17_349 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_17_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_17_368 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_17_50 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_17_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_17_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_17_88 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_18_102 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_18_104 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_18_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_18_111 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_18_113 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_18_130 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_18_138 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_18_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_18_149 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_18_165 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_18_173 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_18_18 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_18_184 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_18_188 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_18_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_18_204 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_18_220 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_18_228 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_18_234 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_18_242 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_18_244 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_18_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_18_263 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_18_279 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_18_310 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_18_314 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_18_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_18_330 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_18_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_18_346 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_18_350 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_18_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_18_380 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_18_53 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_18_57 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_18_86 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_18_90 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_18_98 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_19_106 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_19_110 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_19_112 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_19_139 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_19_148 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_19_164 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_19_178 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_19_18 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_19_182 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_19_198 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_19_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_19_206 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_19_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_19_220 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_19_241 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_19_243 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_19_253 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_19_255 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_19_270 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_19_278 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_19_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_19_311 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_19_315 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_19_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_19_343 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_19_347 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_19_349 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_19_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_19_358 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_19_374 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_19_382 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_19_50 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_19_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_19_78 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_19_82 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_19_98 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_1_104 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_1_120 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_1_136 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_1_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_1_158 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_1_162 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_1_164 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_1_172 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_1_18 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_1_188 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_1_196 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_1_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_1_200 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_1_207 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_1_209 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_1_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_1_255 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_1_259 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_1_275 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_1_279 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_1_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_1_298 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_1_314 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_1_330 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_1_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_1_346 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_1_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_1_368 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_1_50 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_1_52 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_1_59 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_1_67 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_1_69 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_1_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_1_88 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_20_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_20_123 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_20_139 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_20_143 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_20_145 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_20_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_20_193 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_20_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_20_209 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_20_223 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_20_239 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_20_243 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_20_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_20_263 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_20_279 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_20_295 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_20_309 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_20_31 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_20_313 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_20_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_20_333 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_20_337 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_20_344 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_20_348 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_20_350 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_20_361 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_20_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_20_377 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_20_381 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_20_383 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_20_53 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_20_80 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_20_82 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_20_89 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_21_10 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_21_102 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_21_118 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_21_134 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_21_138 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_21_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_21_158 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_21_174 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_21_190 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_21_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_21_20 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_21_206 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_21_245 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_21_249 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_21_265 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_21_273 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_21_278 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_21_286 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_21_302 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_21_315 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_21_331 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_21_347 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_21_349 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_21_35 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_21_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_21_368 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_21_46 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_21_62 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_21_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_21_80 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_21_98 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_22_114 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_22_130 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_22_146 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_22_162 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_22_170 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_22_174 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_22_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_22_18 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_22_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_22_208 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_22_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_22_228 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_22_244 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_22_254 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_22_270 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_22_286 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_22_302 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_22_310 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_22_314 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_22_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_22_333 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_22_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_22_349 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_22_361 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_22_377 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_22_381 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_22_383 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_22_44 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_22_60 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_22_76 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_22_84 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_22_88 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_22_97 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_23_101 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_23_117 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_23_125 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_23_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_23_158 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_23_160 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_23_170 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_23_18 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_23_186 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_23_194 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_23_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_23_201 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_23_209 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_23_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_23_228 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_23_236 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_23_240 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_23_254 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_23_270 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_23_278 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_23_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_23_290 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_23_324 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_23_328 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_23_336 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_23_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_23_362 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_23_366 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_23_371 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_23_379 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_23_383 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_23_50 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_23_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_23_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_23_97 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_24_102 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_24_104 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_24_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_24_115 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_24_119 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_24_137 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_24_141 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_24_143 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_24_167 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_24_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_24_18 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_24_193 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_24_197 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_24_199 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_24_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_24_207 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_24_223 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_24_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_24_26 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_24_263 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_24_303 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_24_314 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_24_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_24_333 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_24_345 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_24_349 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_24_380 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_24_44 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_24_52 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_24_56 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_24_58 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_24_86 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_24_90 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_24_98 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_25_104 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_25_112 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_25_116 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_25_127 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_25_131 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_25_139 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_25_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_25_146 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_25_148 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_25_156 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_25_172 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_25_176 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_25_18 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_25_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_25_205 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_25_209 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_25_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_25_228 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_25_244 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_25_262 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_25_278 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_25_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_25_298 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_25_31 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_25_314 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_25_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_25_33 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_25_333 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_25_349 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_25_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_25_368 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_25_48 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_25_64 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_25_68 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_25_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_25_88 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_26_10 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_26_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_26_115 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_26_119 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_26_121 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_26_130 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_26_146 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_26_162 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_26_170 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_26_174 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_26_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_26_185 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_26_189 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_26_191 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_26_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_26_20 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_26_211 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_26_215 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_26_231 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_26_239 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_26_243 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_26_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_26_263 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_26_279 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_26_28 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_26_295 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_26_30 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_26_303 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_26_313 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_26_33 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_26_330 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_26_338 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_26_346 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_26_350 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_26_366 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_26_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_26_382 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_26_53 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_26_69 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_26_79 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_26_87 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_26_97 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_27_104 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_27_108 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_27_120 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_27_124 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_27_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_27_158 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_27_170 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_27_186 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_27_190 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_27_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_27_204 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_27_208 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_27_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_27_228 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_27_244 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_27_260 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_27_276 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_27_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_27_290 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_27_292 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_27_299 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_27_315 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_27_32 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_27_331 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_27_347 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_27_349 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_27_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_27_36 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_27_368 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_27_38 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_27_4 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_27_52 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_27_68 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_27_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_27_88 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_28_102 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_28_104 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_28_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_28_109 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_28_124 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_28_140 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_28_148 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_28_157 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_28_169 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_28_173 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_28_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_28_18 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_28_185 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_28_189 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_28_191 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_28_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_28_216 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_28_220 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_28_236 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_28_244 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_28_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_28_251 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_28_266 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_28_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_28_298 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_28_314 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_28_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_28_333 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_28_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_28_349 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_28_365 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_28_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_28_371 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_28_379 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_28_383 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_28_53 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_28_79 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_28_86 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_29_106 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_29_115 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_29_127 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_29_135 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_29_139 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_29_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_29_146 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_29_148 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_29_166 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_29_18 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_29_182 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_29_186 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_29_188 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_29_193 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_29_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_29_201 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_29_203 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_29_206 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_29_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_29_228 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_29_236 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_29_238 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_29_264 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_29_268 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_29_276 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_29_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_29_290 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_29_297 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_29_305 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_29_309 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_29_311 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_29_318 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_29_325 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_29_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_29_341 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_29_345 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_29_347 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_29_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_29_354 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_29_382 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_29_50 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_29_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_29_82 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_29_98 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_2_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_2_138 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_2_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_2_172 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_2_174 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_2_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_2_18 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_2_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_2_220 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_2_224 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_2_232 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_2_236 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_2_243 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_2_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_2_263 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_2_272 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_2_300 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_2_304 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_2_312 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_2_314 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_2_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_2_333 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_2_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_2_349 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_2_365 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_2_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_2_381 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_2_383 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_2_45 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_2_73 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_2_77 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_30_104 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_30_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_30_122 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_30_126 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_30_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_30_150 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_30_154 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_30_158 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_30_174 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_30_18 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_30_183 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_30_187 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_30_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_30_201 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_30_217 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_30_233 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_30_237 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_30_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_30_260 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_30_276 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_30_292 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_30_296 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_30_298 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_30_311 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_30_329 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_30_333 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_30_335 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_30_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_30_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_30_364 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_30_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_30_380 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_30_41 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_30_56 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_30_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_30_88 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_31_103 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_31_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_31_123 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_31_139 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_31_153 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_31_157 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_31_173 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_31_18 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_31_189 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_31_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_31_205 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_31_207 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_31_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_31_214 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_31_229 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_31_259 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_31_275 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_31_279 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_31_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_31_290 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_31_292 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_31_295 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_31_299 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_31_303 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_31_311 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_31_313 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_31_322 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_31_334 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_31_341 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_31_349 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_31_36 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_31_362 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_31_378 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_31_382 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_31_40 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_31_44 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_31_60 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_31_68 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_31_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_31_87 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_32_103 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_32_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_32_123 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_32_139 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_32_155 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_32_164 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_32_168 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_32_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_32_181 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_32_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_32_209 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_32_213 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_32_221 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_32_233 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_32_241 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_32_257 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_32_265 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_32_31 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_32_313 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_32_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_32_333 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_32_349 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_32_365 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_32_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_32_381 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_32_383 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_32_53 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_32_55 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_32_63 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_32_71 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_32_95 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_33_111 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_33_119 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_33_130 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_33_134 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_33_138 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_33_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_33_158 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_33_166 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_33_18 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_33_182 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_33_186 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_33_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_33_202 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_33_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_33_234 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_33_250 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_33_26 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_33_266 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_33_274 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_33_278 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_33_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_33_289 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_33_305 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_33_321 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_33_337 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_33_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_33_347 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_33_349 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_33_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_33_368 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_33_38 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_33_40 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_33_55 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_33_63 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_33_67 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_33_69 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_33_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_33_76 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_33_87 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_33_95 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_34_100 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_34_104 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_34_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_34_115 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_34_119 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_34_131 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_34_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_34_146 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_34_162 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_34_164 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_34_172 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_34_174 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_34_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_34_18 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_34_181 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_34_197 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_34_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_34_213 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_34_221 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_34_223 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_34_235 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_34_243 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_34_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_34_263 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_34_279 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_34_295 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_34_311 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_34_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_34_333 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_34_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_34_365 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_34_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_34_381 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_34_383 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_34_53 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_34_57 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_34_59 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_35_126 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_35_130 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_35_138 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_35_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_35_146 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_35_161 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_35_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_35_18 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_35_193 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_35_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_35_209 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_35_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_35_220 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_35_222 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_35_249 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_35_265 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_35_273 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_35_277 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_35_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_35_333 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_35_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_35_341 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_35_345 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_35_349 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_35_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_35_354 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_35_382 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_35_50 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_35_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_35_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_35_86 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_35_90 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_36_101 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_36_139 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_36_147 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_36_163 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_36_171 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_36_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_36_18 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_36_185 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_36_187 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_36_194 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_36_198 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_36_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_36_214 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_36_222 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_36_230 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_36_234 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_36_237 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_36_272 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_36_280 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_36_284 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_36_321 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_36_337 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_36_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_36_365 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_36_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_36_381 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_36_383 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_36_39 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_36_42 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_36_44 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_36_59 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_36_67 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_36_71 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_36_73 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_37_104 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_37_120 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_37_128 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_37_134 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_37_138 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_37_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_37_158 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_37_174 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_37_18 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_37_182 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_37_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_37_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_37_216 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_37_22 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_37_232 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_37_240 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_37_242 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_37_270 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_37_274 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_37_278 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_37_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_37_298 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_37_306 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_37_310 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_37_327 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_37_343 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_37_347 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_37_349 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_37_362 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_37_378 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_37_38 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_37_382 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_37_50 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_37_54 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_37_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_37_88 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_38_103 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_38_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_38_123 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_38_139 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_38_147 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_38_159 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_38_163 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_38_171 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_38_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_38_187 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_38_191 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_38_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_38_210 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_38_226 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_38_242 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_38_244 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_38_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_38_256 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_38_272 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_38_276 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_38_284 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_38_300 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_38_308 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_38_31 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_38_312 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_38_314 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_38_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_38_333 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_38_349 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_38_365 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_38_381 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_38_383 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_38_51 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_38_59 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_38_67 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_38_83 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_38_99 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_39_10 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_39_104 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_39_108 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_39_121 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_39_125 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_39_129 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_39_14 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_39_166 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_39_170 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_39_174 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_39_176 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_39_185 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_39_191 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_39_195 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_39_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_39_202 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_39_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_39_22 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_39_228 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_39_230 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_39_244 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_39_252 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_39_254 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_39_265 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_39_273 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_39_277 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_39_279 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_39_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_39_298 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_39_302 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_39_313 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_39_329 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_39_345 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_39_349 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_39_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_39_368 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_39_44 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_39_60 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_39_68 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_39_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_39_88 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_3_105 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_3_115 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_3_131 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_3_139 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_3_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_3_158 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_3_18 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_3_183 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_3_194 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_3_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_3_205 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_3_209 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_3_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_3_228 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_3_257 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_3_261 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_3_275 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_3_279 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_3_288 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_3_304 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_3_320 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_3_336 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_3_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_3_344 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_3_348 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_3_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_3_368 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_3_50 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_3_54 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_3_76 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_3_92 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_40_100 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_40_104 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_40_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_40_111 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_40_126 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_40_134 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_40_149 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_40_151 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_40_162 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_40_170 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_40_174 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_40_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_40_18 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_40_193 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_40_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_40_221 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_40_225 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_40_230 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_40_261 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_40_277 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_40_293 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_40_309 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_40_314 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_40_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_40_321 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_40_329 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_40_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_40_340 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_40_351 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_40_363 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_40_371 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_40_379 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_40_383 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_40_48 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_40_52 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_40_68 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_40_84 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_41_104 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_41_122 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_41_138 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_41_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_41_150 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_41_158 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_41_174 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_41_18 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_41_190 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_41_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_41_206 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_41_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_41_228 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_41_236 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_41_240 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_41_242 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_41_260 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_41_276 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_41_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_41_290 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_41_332 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_41_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_41_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_41_354 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_41_382 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_41_42 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_41_50 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_41_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_41_86 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_41_96 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_42_103 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_42_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_42_123 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_42_139 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_42_147 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_42_151 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_42_154 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_42_158 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_42_165 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_42_173 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_42_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_42_18 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_42_193 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_42_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_42_219 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_42_235 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_42_243 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_42_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_42_290 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_42_294 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_42_310 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_42_314 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_42_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_42_321 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_42_337 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_42_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_42_341 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_42_343 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_42_354 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_42_358 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_42_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_42_374 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_42_382 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_42_45 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_42_73 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_42_75 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_43_108 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_43_124 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_43_179 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_43_18 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_43_183 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_43_199 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_43_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_43_20 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_43_207 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_43_209 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_43_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_43_228 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_43_232 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_43_240 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_43_256 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_43_272 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_43_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_43_298 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_43_31 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_43_314 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_43_330 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_43_346 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_43_35 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_43_356 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_43_372 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_43_380 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_43_51 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_43_67 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_43_69 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_43_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_43_76 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_43_92 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_44_101 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_44_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_44_123 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_44_139 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_44_155 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_44_171 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_44_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_44_18 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_44_193 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_44_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_44_20 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_44_205 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_44_221 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_44_237 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_44_260 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_44_276 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_44_292 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_44_308 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_44_31 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_44_312 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_44_314 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_44_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_44_333 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_44_337 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_44_339 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_44_369 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_44_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_44_377 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_44_381 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_44_383 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_44_53 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_44_69 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_44_85 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_45_10 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_45_104 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_45_114 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_45_122 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_45_126 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_45_128 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_45_135 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_45_139 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_45_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_45_158 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_45_174 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_45_190 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_45_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_45_208 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_45_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_45_228 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_45_236 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_45_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_45_263 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_45_279 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_45_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_45_298 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_45_306 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_45_319 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_45_335 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_45_343 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_45_347 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_45_349 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_45_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_45_368 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_45_38 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_45_54 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_45_61 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_45_69 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_45_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_45_88 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_46_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_46_109 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_46_116 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_46_124 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_46_126 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_46_154 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_46_162 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_46_172 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_46_174 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_46_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_46_18 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_46_193 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_46_195 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_46_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_46_209 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_46_225 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_46_241 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_46_254 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_46_26 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_46_261 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_46_277 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_46_284 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_46_300 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_46_308 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_46_312 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_46_314 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_46_323 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_46_339 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_46_347 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_46_357 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_46_365 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_46_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_46_372 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_46_376 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_46_53 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_46_61 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_46_63 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_47_118 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_47_134 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_47_138 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_47_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_47_150 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_47_179 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_47_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_47_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_47_216 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_47_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_47_251 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_47_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_47_284 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_47_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_47_345 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_47_347 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_47_379 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_47_38 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_47_383 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_47_6 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_47_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_47_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_47_88 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_47_90 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_48_101 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_48_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_48_123 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_48_139 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_48_155 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_48_171 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_48_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_48_18 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_48_193 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_48_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_48_209 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_48_225 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_48_241 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_48_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_48_263 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_48_279 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_48_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_48_298 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_48_306 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_48_310 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_48_314 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_48_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_48_333 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_48_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_48_349 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_48_357 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_48_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_48_53 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_48_69 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_48_85 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_49_101 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_49_104 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_49_106 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_49_132 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_49_138 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_49_140 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_49_166 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_49_172 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_49_174 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_49_18 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_49_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_49_200 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_49_206 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_49_208 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_49_234 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_49_240 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_49_242 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_49_26 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_49_268 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_49_274 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_49_276 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_49_30 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_49_302 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_49_308 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_49_310 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_49_336 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_49_342 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_49_344 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_49_36 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_49_370 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_49_376 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_49_38 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_49_45 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_49_61 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_49_65 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_49_70 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_49_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_49_79 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_49_95 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_49_99 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_4_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_4_123 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_4_139 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_4_155 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_4_163 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_4_167 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_4_171 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_4_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_4_18 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_4_193 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_4_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_4_209 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_4_225 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_4_241 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_4_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_4_255 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_4_259 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_4_261 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_4_276 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_4_292 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_4_308 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_4_312 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_4_314 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_4_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_4_333 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_4_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_4_349 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_4_365 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_4_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_4_381 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_4_383 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_4_53 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_4_64 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_4_80 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_4_96 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_4_98 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_5_104 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_5_112 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_5_121 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_5_137 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_5_139 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_5_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_5_146 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_5_153 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_5_161 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_5_165 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_5_174 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_5_178 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_5_18 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_5_180 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_5_188 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_5_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_5_204 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_5_208 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_5_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_5_228 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_5_244 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_5_260 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_5_276 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_5_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_5_298 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_5_314 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_5_330 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_5_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_5_346 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_5_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_5_368 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_5_50 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_5_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_5_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_5_88 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_6_117 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_6_121 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_6_129 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_6_173 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_6_18 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_6_191 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_6_199 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_6_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_6_207 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_6_223 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_6_239 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_6_243 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_6_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_6_263 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_6_279 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_6_295 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_6_311 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_6_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_6_333 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_6_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_6_349 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_6_365 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_6_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_6_381 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_6_383 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_6_53 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_6_69 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_6_77 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_6_81 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_6_89 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_7_114 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_7_130 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_7_138 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_7_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_7_158 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_7_169 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_7_175 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_7_18 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_7_191 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_7_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_7_207 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_7_209 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_7_219 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_7_22 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_7_223 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_7_227 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_7_231 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_7_234 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_7_250 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_7_266 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_7_270 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_7_272 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_7_29 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_7_295 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_7_311 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_7_327 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_7_343 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_7_347 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_7_349 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_7_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_7_368 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_7_45 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_7_49 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_7_62 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_7_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_8_100 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_8_104 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_8_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_8_123 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_8_139 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_8_155 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_8_171 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_8_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_8_193 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_8_197 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_8_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_8_232 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_8_241 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_8_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_8_255 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_8_259 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_8_262 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_8_281 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_8_312 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_8_314 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_8_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_8_321 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_8_337 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_8_353 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_8_369 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_8_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_8_377 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_8_381 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_8_383 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_8_41 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_8_49 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_8_6 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_8_71 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_8_87 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_8_89 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_8_92 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_9_106 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_9_122 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_9_138 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_9_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_9_158 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_9_174 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_9_18 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_9_182 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_9_191 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_9_199 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_9_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_9_203 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_9_205 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_9_222 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_9_226 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_9_230 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_1 FILLER_0_9_232 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_9_274 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_9_278 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_9_289 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_9_305 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_9_313 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_9_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_9_344 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_9_348 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_9_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_9_368 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_16 FILLER_0_9_50 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_9_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_9_78 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_8 FILLER_0_9_82 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__decap_4 FILLER_0_9_90 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__fill_2 FILLER_0_9_94 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_0_Left_50 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_0_Right_0 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_10_Left_60 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_10_Right_10 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_11_Left_61 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_11_Right_11 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_12_Left_62 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_12_Right_12 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_13_Left_63 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_13_Right_13 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_14_Left_64 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_14_Right_14 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_15_Left_65 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_15_Right_15 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_16_Left_66 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_16_Right_16 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_17_Left_67 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_17_Right_17 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_18_Left_68 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_18_Right_18 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_19_Left_69 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_19_Right_19 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_1_Left_51 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_1_Right_1 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_20_Left_70 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_20_Right_20 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_21_Left_71 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_21_Right_21 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_22_Left_72 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_22_Right_22 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_23_Left_73 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_23_Right_23 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_24_Left_74 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_24_Right_24 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_25_Left_75 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_25_Right_25 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_26_Left_76 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_26_Right_26 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_27_Left_77 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_27_Right_27 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_28_Left_78 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_28_Right_28 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_29_Left_79 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_29_Right_29 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_2_Left_52 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_2_Right_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_30_Left_80 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_30_Right_30 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_31_Left_81 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_31_Right_31 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_32_Left_82 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_32_Right_32 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_33_Left_83 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_33_Right_33 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_34_Left_84 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_34_Right_34 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_35_Left_85 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_35_Right_35 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_36_Left_86 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_36_Right_36 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_37_Left_87 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_37_Right_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_38_Left_88 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_38_Right_38 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_39_Left_89 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_39_Right_39 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_3_Left_53 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_3_Right_3 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_40_Left_90 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_40_Right_40 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_41_Left_91 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_41_Right_41 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_42_Left_92 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_42_Right_42 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_43_Left_93 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_43_Right_43 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_44_Left_94 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_44_Right_44 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_45_Left_95 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_45_Right_45 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_46_Left_96 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_46_Right_46 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_47_Left_97 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_47_Right_47 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_48_Left_98 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_48_Right_48 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_49_Left_99 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_49_Right_49 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_4_Left_54 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_4_Right_4 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_5_Left_55 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_5_Right_5 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_6_Left_56 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_6_Right_6 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_7_Left_57 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_7_Right_7 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_8_Left_58 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_8_Right_8 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_9_Left_59 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 PHY_EDGE_ROW_9_Right_9 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_0_100 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_0_101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_0_102 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_0_103 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_0_104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_0_105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_0_106 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_0_107 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_0_108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_0_109 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_0_110 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_10_156 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_10_157 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_10_158 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_10_159 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_10_160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_11_161 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_11_162 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_11_163 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_11_164 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_11_165 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_12_166 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_12_167 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_12_168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_12_169 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_12_170 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_13_171 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_13_172 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_13_173 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_13_174 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_13_175 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_14_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_14_177 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_14_178 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_14_179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_14_180 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_15_181 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_15_182 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_15_183 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_15_184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_15_185 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_16_186 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_16_187 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_16_188 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_16_189 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_16_190 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_17_191 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_17_192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_17_193 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_17_194 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_17_195 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_18_196 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_18_197 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_18_198 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_18_199 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_18_200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_19_201 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_19_202 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_19_203 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_19_204 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_19_205 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_1_111 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_1_112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_1_113 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_1_114 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_1_115 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_20_206 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_20_207 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_20_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_20_209 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_20_210 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_21_211 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_21_212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_21_213 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_21_214 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_21_215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_22_216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_22_217 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_22_218 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_22_219 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_22_220 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_23_221 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_23_222 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_23_223 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_23_224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_23_225 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_24_226 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_24_227 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_24_228 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_24_229 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_24_230 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_25_231 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_25_232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_25_233 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_25_234 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_25_235 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_26_236 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_26_237 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_26_238 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_26_239 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_26_240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_27_241 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_27_242 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_27_243 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_27_244 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_27_245 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_28_246 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_28_247 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_28_248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_28_249 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_28_250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_29_251 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_29_252 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_29_253 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_29_254 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_29_255 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_2_116 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_2_117 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_2_118 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_2_119 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_2_120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_30_256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_30_257 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_30_258 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_30_259 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_30_260 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_31_261 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_31_262 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_31_263 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_31_264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_31_265 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_32_266 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_32_267 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_32_268 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_32_269 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_32_270 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_33_271 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_33_272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_33_273 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_33_274 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_33_275 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_34_276 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_34_277 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_34_278 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_34_279 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_34_280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_35_281 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_35_282 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_35_283 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_35_284 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_35_285 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_36_286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_36_287 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_36_288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_36_289 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_36_290 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_37_291 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_37_292 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_37_293 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_37_294 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_37_295 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_38_296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_38_297 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_38_298 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_38_299 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_38_300 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_39_301 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_39_302 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_39_303 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_39_304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_39_305 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_3_121 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_3_122 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_3_123 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_3_124 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_3_125 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_40_306 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_40_307 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_40_308 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_40_309 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_40_310 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_41_311 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_41_312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_41_313 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_41_314 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_41_315 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_42_316 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_42_317 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_42_318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_42_319 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_42_320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_43_321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_43_322 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_43_323 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_43_324 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_43_325 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_44_326 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_44_327 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_44_328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_44_329 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_44_330 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_45_331 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_45_332 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_45_333 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_45_334 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_45_335 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_46_336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_46_337 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_46_338 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_46_339 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_46_340 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_47_341 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_47_342 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_47_343 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_47_344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_47_345 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_48_346 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_48_347 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_48_348 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_48_349 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_48_350 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_49_351 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_49_352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_49_353 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_49_354 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_49_355 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_49_356 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_49_357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_49_358 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_49_359 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_49_360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_49_361 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_4_126 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_4_127 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_4_128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_4_129 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_4_130 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_5_131 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_5_132 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_5_133 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_5_134 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_5_135 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_6_136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_6_137 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_6_138 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_6_139 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_6_140 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_7_141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_7_142 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_7_143 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_7_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_7_145 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_8_146 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_8_147 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_8_148 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_8_149 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_8_150 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_9_151 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_9_152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_9_153 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_9_154 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__tap_2 TAP_TAPCELL_ROW_9_155 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _367_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(net2),
    .Y(_064_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _368_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_065_),
    .A(\bcd[2] ));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _369_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\clkdiv[2] ),
    .Y(_066_));
 gf180mcu_as_sc_mcu7t3v3__nand2b_2 _370_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_067_),
    .B(_066_),
    .A(\counter[2] ));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _371_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\clkdiv[4] ),
    .Y(_068_));
 gf180mcu_as_sc_mcu7t3v3__nand2b_2 _372_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_069_),
    .B(_068_),
    .A(\counter[4] ));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _373_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(\counter[6] ),
    .A(\clkdiv[6] ),
    .Y(_070_));
 gf180mcu_as_sc_mcu7t3v3__nand3_2 _374_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_067_),
    .B(_069_),
    .C(_070_),
    .Y(_071_));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _375_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(\counter[1] ),
    .A(\clkdiv[1] ),
    .Y(_072_));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _376_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(\counter[5] ),
    .A(\clkdiv[5] ),
    .Y(_073_));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _377_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_074_),
    .B(_073_),
    .A(_072_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _378_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\counter[2] ),
    .Y(_075_));
 gf180mcu_as_sc_mcu7t3v3__nand2b_2 _379_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_076_),
    .B(_075_),
    .A(\clkdiv[2] ));
 gf180mcu_as_sc_mcu7t3v3__nand2b_2 _380_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_077_),
    .B(\counter[4] ),
    .A(\clkdiv[4] ));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _381_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(\counter[7] ),
    .A(\clkdiv[7] ),
    .Y(_078_));
 gf180mcu_as_sc_mcu7t3v3__nand3_2 _382_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_076_),
    .B(_077_),
    .C(_078_),
    .Y(_079_));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _383_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_071_),
    .B(_074_),
    .C(_079_),
    .Y(_080_));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _384_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(\counter[3] ),
    .A(\clkdiv[3] ),
    .Y(_081_));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _385_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(\counter[0] ),
    .A(\clkdiv[0] ),
    .Y(_082_));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _386_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_083_),
    .B(_082_),
    .A(_081_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _387_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_084_),
    .A(\counter[12] ));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _388_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\counter[15] ),
    .B(\counter[14] ),
    .C(\counter[13] ),
    .Y(_085_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _389_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_086_),
    .B(\counter[10] ),
    .A(\counter[11] ));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _390_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_087_),
    .B(\counter[8] ),
    .A(\counter[9] ));
 gf180mcu_as_sc_mcu7t3v3__nand4_2 _391_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_084_),
    .B(_085_),
    .C(_086_),
    .D(_087_),
    .Y(_088_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _392_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_089_),
    .B(_088_),
    .A(_083_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _393_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(\m_clkdiv[6] ),
    .A(\m_clkdiv[7] ),
    .Y(_090_));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _394_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\m_clkdiv[9] ),
    .B(\m_clkdiv[8] ),
    .C(_090_),
    .Y(_091_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _395_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(\m_clkdiv[0] ),
    .A(\m_clkdiv[1] ),
    .Y(_092_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _396_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(\m_clkdiv[5] ),
    .A(\m_clkdiv[2] ),
    .Y(_093_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _397_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(\m_clkdiv[4] ),
    .A(\m_clkdiv[3] ),
    .Y(_094_));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _398_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_092_),
    .B(_093_),
    .C(_094_),
    .Y(_095_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _399_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_095_),
    .A(_091_),
    .Y(_096_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _400_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_097_),
    .A(net1));
 gf180mcu_as_sc_mcu7t3v3__nor2b_2 _401_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_098_),
    .B(\clkdiv[4] ),
    .A(\clkdiv[5] ));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _402_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\clkdiv[3] ),
    .Y(_099_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _403_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_100_),
    .B(\clkdiv[2] ),
    .A(_099_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _404_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\clkdiv[7] ),
    .Y(_101_));
 gf180mcu_as_sc_mcu7t3v3__nor2b_2 _405_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_102_),
    .B(\clkdiv[6] ),
    .A(_101_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _406_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_103_),
    .B(\clkdiv[0] ),
    .A(\clkdiv[1] ));
 gf180mcu_as_sc_mcu7t3v3__nand4_2 _407_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_098_),
    .B(_100_),
    .C(_102_),
    .D(_103_),
    .Y(_104_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _408_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_104_),
    .A(_097_),
    .Y(_105_));
 gf180mcu_as_sc_mcu7t3v3__nand4_2 _409_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_080_),
    .B(_089_),
    .C(_096_),
    .D(_105_),
    .Y(_106_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _410_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_106_),
    .Y(_107_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _411_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\r_counter[1] ),
    .Y(_108_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _412_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_109_),
    .A(\lfsr[1] ));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _413_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_109_),
    .A(_108_),
    .Y(_110_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _414_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(\lfsr[0] ),
    .A(\r_counter[0] ),
    .Y(_111_));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _415_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_111_),
    .A(_110_),
    .Y(_112_));
 gf180mcu_as_sc_mcu7t3v3__maj3_2 _416_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_113_),
    .A(\r_counter[1] ),
    .B(\lfsr[1] ),
    .C(_111_));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _417_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(\lfsr[2] ),
    .A(\r_counter[2] ),
    .Y(_114_));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _418_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_114_),
    .A(_113_),
    .Y(_115_));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _419_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_116_),
    .B(_115_),
    .A(_112_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _420_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_117_),
    .A(\lfsr[2] ));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _421_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_117_),
    .A(\r_counter[2] ),
    .Y(_118_));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _422_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_118_),
    .A(_113_),
    .Y(_119_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _423_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\r_counter[0] ),
    .Y(_120_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _424_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_121_),
    .A(\lfsr[0] ));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _425_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_121_),
    .A(_120_),
    .Y(_122_));
 gf180mcu_as_sc_mcu7t3v3__nand3_2 _426_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_110_),
    .B(_119_),
    .C(_122_),
    .Y(_123_));
 gf180mcu_as_sc_mcu7t3v3__nor2b_2 _427_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_124_),
    .B(_106_),
    .A(_123_));
 gf180mcu_as_sc_mcu7t3v3__aoi22_4 _428_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_125_),
    .A(_065_),
    .B(_107_),
    .C(_116_),
    .D(_124_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _429_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_125_),
    .A(_064_),
    .Y(_126_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _430_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_126_),
    .Y(_019_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _431_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_089_),
    .A(_080_),
    .Y(_127_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _432_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_105_),
    .A(_096_),
    .Y(_128_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _433_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\lfsr[0] ),
    .Y(_129_));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _434_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_129_),
    .A(_120_),
    .Y(_130_));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _435_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_131_),
    .B(_130_),
    .A(_112_));
 gf180mcu_as_sc_mcu7t3v3__nand4_2 _436_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_127_),
    .B(_128_),
    .C(_123_),
    .D(_131_),
    .Y(_132_));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _437_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_133_),
    .B(_107_),
    .A(\bcd[1] ));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _438_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_134_),
    .B(_133_),
    .A(_132_));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _439_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_135_),
    .B(_130_),
    .A(_119_));
 gf180mcu_as_sc_mcu7t3v3__nand3_2 _440_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_110_),
    .B(_115_),
    .C(_122_),
    .Y(_136_));
 gf180mcu_as_sc_mcu7t3v3__ao31_2 _441_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .D(_107_),
    .A(_131_),
    .B(_135_),
    .C(_136_),
    .Y(_137_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _442_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_138_),
    .A(net2));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _443_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_139_),
    .C(_138_),
    .B(_107_),
    .A(\bcd[0] ));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _444_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_140_),
    .B(_139_),
    .A(_137_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _445_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_140_),
    .A(_134_),
    .Y(_141_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _446_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_138_),
    .Y(_142_));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _447_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_143_),
    .A(_132_),
    .B(_133_),
    .C(_142_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _448_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_140_),
    .Y(_017_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _449_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_144_),
    .C(_125_),
    .B(_017_),
    .A(_143_));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _450_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_145_),
    .A(_019_),
    .B(_141_),
    .C(_144_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _451_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_145_),
    .Y(_000_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _452_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_142_),
    .Y(_146_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _453_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_106_),
    .Y(_147_));
 gf180mcu_as_sc_mcu7t3v3__ao22_2 _454_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_065_),
    .B(_147_),
    .C(_116_),
    .D(_124_),
    .Y(_148_));
 gf180mcu_as_sc_mcu7t3v3__aoi22_2 _455_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_149_),
    .A(_132_),
    .B(_133_),
    .C(_137_),
    .D(_139_));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _456_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_146_),
    .B(_148_),
    .C(_149_),
    .Y(_150_));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _457_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_151_),
    .A(_141_),
    .B(_150_),
    .C(_144_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _458_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_151_),
    .Y(_001_));
 gf180mcu_as_sc_mcu7t3v3__aoi31_2 _459_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_125_),
    .B(_132_),
    .C(_133_),
    .Y(_002_),
    .D(_017_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _460_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_152_),
    .B(_017_),
    .A(_134_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _461_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_150_),
    .A(_152_),
    .Y(_153_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _462_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_153_),
    .Y(_003_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _463_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_018_),
    .A(_143_));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _464_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_154_),
    .A(_148_),
    .B(_018_),
    .C(_150_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _465_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_154_),
    .Y(_004_));
 gf180mcu_as_sc_mcu7t3v3__nand4_2 _466_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_148_),
    .B(_018_),
    .C(_137_),
    .D(_139_),
    .Y(_155_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _467_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_155_),
    .Y(_005_));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _468_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_006_),
    .B(_150_),
    .A(_141_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _469_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_138_),
    .Y(_156_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _470_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_156_),
    .Y(_157_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _471_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_157_),
    .Y(_158_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _472_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_007_),
    .B(_158_),
    .A(\m_clkdiv[0] ));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _473_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(\m_clkdiv[0] ),
    .A(\m_clkdiv[1] ),
    .Y(_159_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _474_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_064_),
    .Y(_160_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _475_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_160_),
    .Y(_161_));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _476_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_162_),
    .B(_092_),
    .A(_161_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _477_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_008_),
    .B(_162_),
    .A(_159_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _478_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_163_),
    .B(_159_),
    .A(\m_clkdiv[2] ));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _479_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_159_),
    .A(\m_clkdiv[2] ),
    .Y(_164_));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _480_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_158_),
    .B(_163_),
    .C(_164_),
    .Y(_165_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _481_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_165_),
    .Y(_009_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _482_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_164_),
    .A(\m_clkdiv[3] ),
    .Y(_166_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _483_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_164_),
    .A(\m_clkdiv[3] ),
    .Y(_167_));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _484_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_168_),
    .B(_167_),
    .A(_161_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _485_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_010_),
    .B(_168_),
    .A(_166_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _486_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_166_),
    .A(\m_clkdiv[4] ),
    .Y(_169_));
 gf180mcu_as_sc_mcu7t3v3__nand4_2 _487_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\m_clkdiv[3] ),
    .B(\m_clkdiv[2] ),
    .C(\m_clkdiv[4] ),
    .D(_159_),
    .Y(_170_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _488_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_170_),
    .A(_160_),
    .Y(_171_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _489_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_171_),
    .A(_169_),
    .Y(_172_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _490_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_172_),
    .Y(_011_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _491_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_173_),
    .A(\m_clkdiv[5] ));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _492_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_174_),
    .B(_170_),
    .A(_173_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _493_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_156_),
    .Y(_175_));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _494_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_176_),
    .A(_173_),
    .B(_170_),
    .C(_175_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _495_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_012_),
    .B(_176_),
    .A(_174_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _496_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_177_),
    .B(_174_),
    .A(\m_clkdiv[6] ));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _497_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_174_),
    .A(\m_clkdiv[6] ),
    .Y(_178_));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _498_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_158_),
    .B(_177_),
    .C(_178_),
    .Y(_179_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _499_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_179_),
    .Y(_013_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _500_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_180_),
    .B(_178_),
    .A(\m_clkdiv[7] ));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _501_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_178_),
    .A(\m_clkdiv[7] ),
    .Y(_181_));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _502_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_158_),
    .B(_180_),
    .C(_181_),
    .Y(_182_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _503_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_182_),
    .Y(_014_));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _504_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_183_),
    .B(_181_),
    .A(\m_clkdiv[8] ));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _505_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_181_),
    .A(\m_clkdiv[8] ),
    .Y(_184_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _506_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_184_),
    .A(_160_),
    .Y(_185_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _507_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_185_),
    .A(_183_),
    .Y(_186_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _508_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_186_),
    .Y(_015_));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _509_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_183_),
    .A(\m_clkdiv[9] ),
    .Y(_187_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _510_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_187_),
    .A(_161_),
    .Y(_188_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _511_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_188_),
    .Y(_016_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _512_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_091_),
    .Y(_189_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _513_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_095_),
    .Y(_190_));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _514_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_191_),
    .B(_190_),
    .A(_189_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _515_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_191_),
    .Y(_192_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _516_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_192_),
    .Y(_193_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _517_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_189_),
    .Y(_194_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _518_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_194_),
    .Y(_195_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _519_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_190_),
    .Y(_196_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _520_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_196_),
    .Y(_197_));
 gf180mcu_as_sc_mcu7t3v3__ao31_2 _521_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .D(_157_),
    .A(_109_),
    .B(_195_),
    .C(_197_),
    .Y(_198_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _522_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_020_),
    .C(_198_),
    .B(_193_),
    .A(_121_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _523_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_192_),
    .Y(_199_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _524_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_189_),
    .Y(_200_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _525_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_190_),
    .Y(_201_));
 gf180mcu_as_sc_mcu7t3v3__ao31_2 _526_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .D(_146_),
    .A(\lfsr[2] ),
    .B(_200_),
    .C(_201_),
    .Y(_202_));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _527_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_203_),
    .A(\lfsr[1] ),
    .B(_199_),
    .C(_202_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _528_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_203_),
    .Y(_021_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _529_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_204_),
    .A(\lfsr[3] ));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _530_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_142_),
    .Y(_205_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _531_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_205_),
    .Y(_206_));
 gf180mcu_as_sc_mcu7t3v3__ao31_2 _532_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .D(_206_),
    .A(_204_),
    .B(_195_),
    .C(_197_),
    .Y(_207_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _533_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_022_),
    .C(_207_),
    .B(_193_),
    .A(_117_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _534_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_156_),
    .Y(_208_));
 gf180mcu_as_sc_mcu7t3v3__ao31_2 _535_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .D(_208_),
    .A(\lfsr[4] ),
    .B(_200_),
    .C(_201_),
    .Y(_209_));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _536_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_210_),
    .A(\lfsr[3] ),
    .B(_199_),
    .C(_209_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _537_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_210_),
    .Y(_023_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _538_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_192_),
    .Y(_211_));
 gf180mcu_as_sc_mcu7t3v3__ao31_2 _539_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .D(_208_),
    .A(\lfsr[5] ),
    .B(_194_),
    .C(_196_),
    .Y(_212_));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _540_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_213_),
    .A(\lfsr[4] ),
    .B(_211_),
    .C(_212_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _541_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_213_),
    .Y(_024_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _542_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_157_),
    .Y(_214_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _543_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_215_),
    .B(_211_),
    .A(\lfsr[6] ));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _544_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_096_),
    .Y(_216_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _545_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_216_),
    .Y(_217_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _546_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_218_),
    .B(_217_),
    .A(\lfsr[5] ));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _547_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_214_),
    .B(_215_),
    .C(_218_),
    .Y(_219_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _548_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_219_),
    .Y(_025_));
 gf180mcu_as_sc_mcu7t3v3__ao31_2 _549_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .D(_208_),
    .A(\lfsr[7] ),
    .B(_194_),
    .C(_196_),
    .Y(_220_));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _550_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_221_),
    .A(\lfsr[6] ),
    .B(_211_),
    .C(_220_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _551_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_221_),
    .Y(_026_));
 gf180mcu_as_sc_mcu7t3v3__ao31_2 _552_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .D(_208_),
    .A(\lfsr[8] ),
    .B(_194_),
    .C(_196_),
    .Y(_222_));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _553_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_223_),
    .A(\lfsr[7] ),
    .B(_211_),
    .C(_222_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _554_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_223_),
    .Y(_027_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _555_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_224_),
    .A(\lfsr[8] ));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _556_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_225_),
    .A(\lfsr[9] ));
 gf180mcu_as_sc_mcu7t3v3__ao31_2 _557_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .D(_206_),
    .A(_225_),
    .B(_195_),
    .C(_197_),
    .Y(_226_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _558_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_028_),
    .C(_226_),
    .B(_193_),
    .A(_224_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _559_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_227_),
    .A(\lfsr[10] ));
 gf180mcu_as_sc_mcu7t3v3__ao31_2 _560_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .D(_206_),
    .A(_227_),
    .B(_195_),
    .C(_197_),
    .Y(_228_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _561_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_029_),
    .C(_228_),
    .B(_193_),
    .A(_225_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _562_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_192_),
    .Y(_229_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _563_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_189_),
    .Y(_230_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _564_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_190_),
    .Y(_231_));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _565_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(\lfsr[11] ),
    .A(_129_),
    .Y(_232_));
 gf180mcu_as_sc_mcu7t3v3__ao31_2 _566_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .D(_206_),
    .A(_230_),
    .B(_231_),
    .C(_232_),
    .Y(_233_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _567_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_030_),
    .C(_233_),
    .B(_229_),
    .A(_227_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _568_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_234_),
    .A(\lfsr[11] ));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _569_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_235_),
    .A(\lfsr[12] ));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _570_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_156_),
    .Y(_236_));
 gf180mcu_as_sc_mcu7t3v3__ao31_2 _571_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .D(_236_),
    .A(_235_),
    .B(_230_),
    .C(_231_),
    .Y(_237_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _572_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_031_),
    .C(_237_),
    .B(_229_),
    .A(_234_));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _573_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(\lfsr[13] ),
    .A(_129_),
    .Y(_238_));
 gf180mcu_as_sc_mcu7t3v3__ao31_2 _574_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .D(_236_),
    .A(_200_),
    .B(_201_),
    .C(_238_),
    .Y(_239_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _575_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_032_),
    .C(_239_),
    .B(_229_),
    .A(_235_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _576_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_240_),
    .A(\lfsr[13] ));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _577_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(\lfsr[14] ),
    .A(_129_),
    .Y(_241_));
 gf180mcu_as_sc_mcu7t3v3__ao31_2 _578_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .D(_236_),
    .A(_200_),
    .B(_201_),
    .C(_241_),
    .Y(_242_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _579_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_033_),
    .C(_242_),
    .B(_229_),
    .A(_240_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _580_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_243_),
    .A(\lfsr[14] ));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _581_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_244_),
    .A(\lfsr[15] ));
 gf180mcu_as_sc_mcu7t3v3__ao31_2 _582_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .D(_236_),
    .A(_244_),
    .B(_230_),
    .C(_231_),
    .Y(_245_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _583_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_034_),
    .C(_245_),
    .B(_199_),
    .A(_243_));
 gf180mcu_as_sc_mcu7t3v3__ao31_2 _584_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .D(_175_),
    .A(_121_),
    .B(_230_),
    .C(_231_),
    .Y(_246_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _585_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_035_),
    .C(_246_),
    .B(_199_),
    .A(_244_));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _586_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_247_),
    .B(_089_),
    .A(_080_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _587_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\counter[0] ),
    .Y(_248_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _588_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_249_),
    .C(_248_),
    .B(_128_),
    .A(_247_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _589_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(net1),
    .Y(_250_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _590_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_104_),
    .A(_250_),
    .Y(_251_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _591_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_251_),
    .A(_216_),
    .Y(_252_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _592_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_252_),
    .A(_248_),
    .Y(_253_));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _593_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_214_),
    .B(_249_),
    .C(_253_),
    .Y(_254_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _594_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_254_),
    .Y(_036_));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _595_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_255_),
    .B(_251_),
    .A(_096_));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _596_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_256_),
    .A(_097_),
    .B(_247_),
    .C(_255_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _597_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_256_),
    .Y(_257_));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _598_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_258_),
    .B(_257_),
    .A(_064_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _599_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_259_),
    .B(_253_),
    .A(\counter[1] ));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _600_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_248_),
    .A(\counter[1] ),
    .Y(_260_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _601_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_260_),
    .A(_252_),
    .Y(_261_));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _602_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_258_),
    .B(_259_),
    .C(_261_),
    .Y(_262_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _603_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_262_),
    .Y(_037_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _604_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_261_),
    .A(_075_),
    .Y(_263_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _605_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_264_),
    .B(_261_),
    .A(_075_));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _606_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_258_),
    .B(_263_),
    .C(_264_),
    .Y(_265_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _607_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_265_),
    .Y(_038_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _608_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_256_),
    .A(_064_),
    .Y(_266_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _609_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_266_),
    .Y(_267_));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _610_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_250_),
    .B(_205_),
    .C(_127_),
    .Y(_268_));
 gf180mcu_as_sc_mcu7t3v3__aoi22_2 _611_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_269_),
    .A(\counter[3] ),
    .B(_267_),
    .C(_263_),
    .D(_268_));
 gf180mcu_as_sc_mcu7t3v3__nand4_2 _612_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\counter[3] ),
    .B(_075_),
    .C(\counter[1] ),
    .D(_248_),
    .Y(_270_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _613_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_271_),
    .B(_270_),
    .A(_255_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _614_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_039_),
    .B(_271_),
    .A(_269_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _615_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\counter[4] ),
    .Y(_272_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _616_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_273_),
    .B(_271_),
    .A(_272_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _617_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_271_),
    .A(_272_),
    .Y(_274_));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _618_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_258_),
    .B(_273_),
    .C(_274_),
    .Y(_275_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _619_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_275_),
    .Y(_040_));
 gf180mcu_as_sc_mcu7t3v3__aoi22_2 _620_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_276_),
    .A(\counter[5] ),
    .B(_267_),
    .C(_268_),
    .D(_274_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _621_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_272_),
    .A(\counter[5] ),
    .Y(_277_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _622_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_277_),
    .A(_271_),
    .Y(_278_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _623_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_041_),
    .B(_278_),
    .A(_276_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _624_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\counter[6] ),
    .Y(_279_));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _625_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_280_),
    .A(_279_),
    .B(_278_),
    .C(_258_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _626_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_281_),
    .B(_278_),
    .A(_279_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _627_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_042_),
    .B(_281_),
    .A(_280_));
 gf180mcu_as_sc_mcu7t3v3__nand2b_2 _628_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_282_),
    .B(_268_),
    .A(\counter[7] ));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _629_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_283_),
    .C(\counter[7] ),
    .B(_278_),
    .A(_279_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _630_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_043_),
    .C(_283_),
    .B(_282_),
    .A(_280_));
 gf180mcu_as_sc_mcu7t3v3__nand3_2 _631_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_279_),
    .B(\counter[5] ),
    .C(_272_),
    .Y(_284_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _632_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_285_),
    .B(_284_),
    .A(_270_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _633_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_285_),
    .A(\counter[7] ),
    .Y(_286_));
 gf180mcu_as_sc_mcu7t3v3__nand4_2 _634_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\counter[8] ),
    .B(_216_),
    .C(_251_),
    .D(_286_),
    .Y(_287_));
 gf180mcu_as_sc_mcu7t3v3__ao31_2 _635_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .D(\counter[8] ),
    .A(_216_),
    .B(_251_),
    .C(_286_),
    .Y(_288_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _636_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_288_),
    .A(_266_),
    .Y(_289_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _637_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_289_),
    .A(_287_),
    .Y(_290_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _638_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_290_),
    .Y(_044_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _639_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_291_),
    .A(\counter[9] ));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _640_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_292_),
    .B(_287_),
    .A(_291_));
 gf180mcu_as_sc_mcu7t3v3__ao31_2 _641_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .D(_142_),
    .A(_250_),
    .B(_091_),
    .C(_095_),
    .Y(_293_));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _642_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_294_),
    .A(_291_),
    .B(_287_),
    .C(_293_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _643_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_045_),
    .B(_294_),
    .A(_292_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _644_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_293_),
    .Y(_295_));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _645_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_292_),
    .A(\counter[10] ),
    .Y(_296_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _646_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_046_),
    .B(_296_),
    .A(_295_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _647_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_297_),
    .C(\counter[11] ),
    .B(_292_),
    .A(\counter[10] ));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _648_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_298_),
    .B(\counter[10] ),
    .A(\counter[11] ));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _649_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_291_),
    .B(_287_),
    .C(_298_),
    .Y(_299_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _650_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_299_),
    .Y(_300_));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _651_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_295_),
    .B(_297_),
    .C(_300_),
    .Y(_301_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _652_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_301_),
    .Y(_047_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _653_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\counter[12] ),
    .Y(_302_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _654_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_303_),
    .B(_300_),
    .A(_302_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _655_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_300_),
    .A(_302_),
    .Y(_304_));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _656_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_295_),
    .B(_303_),
    .C(_304_),
    .Y(_305_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _657_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_305_),
    .Y(_048_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _658_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\counter[13] ),
    .Y(_306_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _659_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_307_),
    .B(_304_),
    .A(_306_));
 gf180mcu_as_sc_mcu7t3v3__ao31_2 _660_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .D(_293_),
    .A(_306_),
    .B(_302_),
    .C(_300_),
    .Y(_308_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _661_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_049_),
    .B(_308_),
    .A(_307_));
 gf180mcu_as_sc_mcu7t3v3__nand4_2 _662_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\counter[14] ),
    .B(_306_),
    .C(_302_),
    .D(_299_),
    .Y(_309_));
 gf180mcu_as_sc_mcu7t3v3__ao31_2 _663_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .D(\counter[14] ),
    .A(_306_),
    .B(\counter[12] ),
    .C(_299_),
    .Y(_310_));
 gf180mcu_as_sc_mcu7t3v3__nor2b_2 _664_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_311_),
    .B(_293_),
    .A(_310_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _665_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_311_),
    .A(_309_),
    .Y(_312_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _666_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_312_),
    .Y(_050_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _667_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_313_),
    .A(\counter[15] ));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _668_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_309_),
    .A(_313_),
    .Y(_314_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _669_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_315_),
    .C(_295_),
    .B(_309_),
    .A(_313_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _670_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_315_),
    .A(_314_),
    .Y(_316_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _671_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_316_),
    .Y(_051_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _672_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\clkdiv[0] ),
    .Y(_317_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _673_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_318_),
    .A(_317_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _674_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_257_),
    .Y(_319_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _675_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_319_),
    .A(_318_),
    .Y(_320_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _676_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_321_),
    .C(_157_),
    .B(_147_),
    .A(_318_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _677_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_321_),
    .A(_320_),
    .Y(_322_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _678_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_322_),
    .Y(_052_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _679_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\clkdiv[1] ),
    .Y(_323_));
 gf180mcu_as_sc_mcu7t3v3__inv_2 _680_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_324_),
    .A(_323_));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _681_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_317_),
    .A(_323_),
    .Y(_325_));
 gf180mcu_as_sc_mcu7t3v3__ao31_2 _682_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .D(_175_),
    .A(_127_),
    .B(_128_),
    .C(_325_),
    .Y(_326_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _683_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_053_),
    .C(_326_),
    .B(_319_),
    .A(_324_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _684_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_128_),
    .A(_127_),
    .Y(_327_));
 gf180mcu_as_sc_mcu7t3v3__nand3_2 _685_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_066_),
    .B(_323_),
    .C(_317_),
    .Y(_328_));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _686_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_329_),
    .A(_323_),
    .B(_317_),
    .C(_066_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _687_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_257_),
    .A(_066_),
    .Y(_330_));
 gf180mcu_as_sc_mcu7t3v3__ao31_2 _688_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .D(_330_),
    .A(_327_),
    .B(_328_),
    .C(_329_),
    .Y(_331_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _689_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_331_),
    .A(_161_),
    .Y(_332_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _690_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_332_),
    .Y(_054_));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _691_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_328_),
    .A(_099_),
    .Y(_333_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _692_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_334_),
    .B(_147_),
    .A(_146_));
 gf180mcu_as_sc_mcu7t3v3__ao22_2 _693_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_099_),
    .B(_267_),
    .C(_333_),
    .D(_334_),
    .Y(_335_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _694_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_335_),
    .Y(_055_));
 gf180mcu_as_sc_mcu7t3v3__nor2b_2 _695_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_336_),
    .B(_328_),
    .A(_099_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _696_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_336_),
    .A(_068_),
    .Y(_337_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _697_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_337_),
    .Y(_338_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _698_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_339_),
    .B(_338_),
    .A(_147_));
 gf180mcu_as_sc_mcu7t3v3__aoi21_2 _699_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_340_),
    .C(_339_),
    .B(_319_),
    .A(_068_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _700_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_341_),
    .B(_336_),
    .A(_068_));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _701_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_214_),
    .B(_340_),
    .C(_341_),
    .Y(_342_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _702_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_342_),
    .Y(_056_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _703_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\clkdiv[5] ),
    .Y(_343_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _704_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_338_),
    .A(_343_),
    .Y(_344_));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _705_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_345_),
    .B(_338_),
    .A(_343_));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _706_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_346_),
    .A(_343_),
    .B(_257_),
    .C(_205_));
 gf180mcu_as_sc_mcu7t3v3__ao31_2 _707_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .D(_346_),
    .A(_327_),
    .B(_344_),
    .C(_345_),
    .Y(_347_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _708_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_347_),
    .Y(_057_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _709_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\clkdiv[6] ),
    .Y(_348_));
 gf180mcu_as_sc_mcu7t3v3__xnor2_2 _710_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_345_),
    .A(_348_),
    .Y(_349_));
 gf180mcu_as_sc_mcu7t3v3__ao22_2 _711_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_348_),
    .B(_267_),
    .C(_349_),
    .D(_334_),
    .Y(_350_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _712_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_350_),
    .Y(_058_));
 gf180mcu_as_sc_mcu7t3v3__ao31_2 _713_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .D(_101_),
    .A(_348_),
    .B(\clkdiv[5] ),
    .C(_337_),
    .Y(_351_));
 gf180mcu_as_sc_mcu7t3v3__nand4_2 _714_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_101_),
    .B(_348_),
    .C(_343_),
    .D(_338_),
    .Y(_352_));
 gf180mcu_as_sc_mcu7t3v3__ao31_2 _715_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .D(_205_),
    .A(_327_),
    .B(_351_),
    .C(_352_),
    .Y(_353_));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _716_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_354_),
    .A(_101_),
    .B(_319_),
    .C(_353_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _717_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_354_),
    .Y(_059_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _718_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_355_),
    .B(_217_),
    .A(_120_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _719_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_217_),
    .A(_120_),
    .Y(_356_));
 gf180mcu_as_sc_mcu7t3v3__nor3_2 _720_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_214_),
    .B(_355_),
    .C(_356_),
    .Y(_357_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _721_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_357_),
    .Y(_060_));
 gf180mcu_as_sc_mcu7t3v3__and2_2 _722_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_356_),
    .A(_108_),
    .Y(_358_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _723_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_356_),
    .A(_108_),
    .Y(_359_));
 gf180mcu_as_sc_mcu7t3v3__nand2_2 _724_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_360_),
    .B(_359_),
    .A(_160_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _725_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_061_),
    .B(_360_),
    .A(_358_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _726_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_361_),
    .B(_358_),
    .A(\r_counter[2] ));
 gf180mcu_as_sc_mcu7t3v3__ao31_2 _727_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .D(_175_),
    .A(\r_counter[2] ),
    .B(_108_),
    .C(_356_),
    .Y(_362_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _728_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_062_),
    .B(_362_),
    .A(_361_));
 gf180mcu_as_sc_mcu7t3v3__or2_2 _729_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .B(_105_),
    .A(_191_),
    .Y(_363_));
 gf180mcu_as_sc_mcu7t3v3__nor2_2 _730_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_364_),
    .B(_104_),
    .A(_250_));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _731_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_365_),
    .A(_217_),
    .B(_364_),
    .C(_146_));
 gf180mcu_as_sc_mcu7t3v3__ao21_2 _732_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .Y(_366_),
    .A(dp),
    .B(_363_),
    .C(_365_));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _733_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(_366_),
    .Y(_063_));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _734_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_3_3__leaf_wb_clk_i),
    .D(_005_),
    .Q(net5));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _735_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_3_3__leaf_wb_clk_i),
    .D(_000_),
    .Q(net3));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _736_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_3_6__leaf_wb_clk_i),
    .D(_001_),
    .Q(net6));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _737_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_3_6__leaf_wb_clk_i),
    .D(_002_),
    .Q(net7));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _738_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_3_6__leaf_wb_clk_i),
    .D(_003_),
    .Q(net8));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _739_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_3_7__leaf_wb_clk_i),
    .D(_004_),
    .Q(net9));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _740_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_3_3__leaf_wb_clk_i),
    .D(_006_),
    .Q(net4));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _741_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_3_1__leaf_wb_clk_i),
    .D(_007_),
    .Q(\m_clkdiv[0] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _742_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_3_1__leaf_wb_clk_i),
    .D(_008_),
    .Q(\m_clkdiv[1] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _743_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_3_1__leaf_wb_clk_i),
    .D(_009_),
    .Q(\m_clkdiv[2] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _744_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_3_1__leaf_wb_clk_i),
    .D(_010_),
    .Q(\m_clkdiv[3] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _745_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_3_4__leaf_wb_clk_i),
    .D(_011_),
    .Q(\m_clkdiv[4] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _746_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_3_4__leaf_wb_clk_i),
    .D(_012_),
    .Q(\m_clkdiv[5] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _747_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_3_4__leaf_wb_clk_i),
    .D(_013_),
    .Q(\m_clkdiv[6] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _748_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_3_5__leaf_wb_clk_i),
    .D(_014_),
    .Q(\m_clkdiv[7] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _749_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_3_5__leaf_wb_clk_i),
    .D(_015_),
    .Q(\m_clkdiv[8] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _750_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_3_4__leaf_wb_clk_i),
    .D(_016_),
    .Q(\m_clkdiv[9] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _751_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_3_7__leaf_wb_clk_i),
    .D(_017_),
    .Q(\bcd[0] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _752_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_3_6__leaf_wb_clk_i),
    .D(_018_),
    .Q(\bcd[1] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _753_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_3_6__leaf_wb_clk_i),
    .D(_019_),
    .Q(\bcd[2] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _754_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_3_5__leaf_wb_clk_i),
    .D(_020_),
    .Q(\lfsr[0] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _755_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_3_7__leaf_wb_clk_i),
    .D(_021_),
    .Q(\lfsr[1] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _756_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_3_5__leaf_wb_clk_i),
    .D(_022_),
    .Q(\lfsr[2] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _757_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_3_7__leaf_wb_clk_i),
    .D(_023_),
    .Q(\lfsr[3] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _758_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_3_5__leaf_wb_clk_i),
    .D(_024_),
    .Q(\lfsr[4] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _759_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_3_5__leaf_wb_clk_i),
    .D(_025_),
    .Q(\lfsr[5] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _760_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_3_5__leaf_wb_clk_i),
    .D(_026_),
    .Q(\lfsr[6] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _761_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_3_5__leaf_wb_clk_i),
    .D(_027_),
    .Q(\lfsr[7] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _762_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_3_5__leaf_wb_clk_i),
    .D(_028_),
    .Q(\lfsr[8] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _763_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_3_5__leaf_wb_clk_i),
    .D(_029_),
    .Q(\lfsr[9] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _764_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_3_7__leaf_wb_clk_i),
    .D(_030_),
    .Q(\lfsr[10] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _765_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_3_7__leaf_wb_clk_i),
    .D(_031_),
    .Q(\lfsr[11] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _766_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_3_7__leaf_wb_clk_i),
    .D(_032_),
    .Q(\lfsr[12] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _767_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_3_7__leaf_wb_clk_i),
    .D(_033_),
    .Q(\lfsr[13] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _768_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_3_7__leaf_wb_clk_i),
    .D(_034_),
    .Q(\lfsr[14] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _769_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_3_6__leaf_wb_clk_i),
    .D(_035_),
    .Q(\lfsr[15] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _770_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_3_0__leaf_wb_clk_i),
    .D(_036_),
    .Q(\counter[0] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _771_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_3_0__leaf_wb_clk_i),
    .D(_037_),
    .Q(\counter[1] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _772_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_3_2__leaf_wb_clk_i),
    .D(_038_),
    .Q(\counter[2] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _773_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_3_2__leaf_wb_clk_i),
    .D(_039_),
    .Q(\counter[3] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _774_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_3_2__leaf_wb_clk_i),
    .D(_040_),
    .Q(\counter[4] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _775_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_3_2__leaf_wb_clk_i),
    .D(_041_),
    .Q(\counter[5] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _776_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_3_2__leaf_wb_clk_i),
    .D(_042_),
    .Q(\counter[6] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _777_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_3_2__leaf_wb_clk_i),
    .D(_043_),
    .Q(\counter[7] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _778_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_3_1__leaf_wb_clk_i),
    .D(_044_),
    .Q(\counter[8] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _779_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_3_0__leaf_wb_clk_i),
    .D(_045_),
    .Q(\counter[9] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _780_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_3_0__leaf_wb_clk_i),
    .D(_046_),
    .Q(\counter[10] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _781_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_3_0__leaf_wb_clk_i),
    .D(_047_),
    .Q(\counter[11] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _782_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_3_0__leaf_wb_clk_i),
    .D(_048_),
    .Q(\counter[12] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _783_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_3_0__leaf_wb_clk_i),
    .D(_049_),
    .Q(\counter[13] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _784_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_3_1__leaf_wb_clk_i),
    .D(_050_),
    .Q(\counter[14] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _785_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_3_0__leaf_wb_clk_i),
    .D(_051_),
    .Q(\counter[15] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _786_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_3_4__leaf_wb_clk_i),
    .D(_052_),
    .Q(\clkdiv[0] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _787_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_3_6__leaf_wb_clk_i),
    .D(_053_),
    .Q(\clkdiv[1] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _788_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_3_1__leaf_wb_clk_i),
    .D(_054_),
    .Q(\clkdiv[2] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _789_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_3_2__leaf_wb_clk_i),
    .D(_055_),
    .Q(\clkdiv[3] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _790_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_3_3__leaf_wb_clk_i),
    .D(_056_),
    .Q(\clkdiv[4] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _791_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_3_6__leaf_wb_clk_i),
    .D(_057_),
    .Q(\clkdiv[5] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _792_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_3_3__leaf_wb_clk_i),
    .D(_058_),
    .Q(\clkdiv[6] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _793_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_3_3__leaf_wb_clk_i),
    .D(_059_),
    .Q(\clkdiv[7] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _794_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_3_4__leaf_wb_clk_i),
    .D(_060_),
    .Q(\r_counter[0] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _795_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_3_4__leaf_wb_clk_i),
    .D(_061_),
    .Q(\r_counter[1] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _796_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_3_4__leaf_wb_clk_i),
    .D(_062_),
    .Q(\r_counter[2] ));
 gf180mcu_as_sc_mcu7t3v3__dfxtp_2 _797_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .CLK(clknet_3_7__leaf_wb_clk_i),
    .D(_063_),
    .Q(dp));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _798_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(dp),
    .Y(net10));
 gf180mcu_as_sc_mcu7t3v3__buff_2 _799_ (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(\lfsr[3] ),
    .Y(net11));
 gf180mcu_as_sc_mcu7t3v3__clkbuff_12 clkbuf_0_wb_clk_i (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(wb_clk_i),
    .Y(clknet_0_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__clkbuff_12 clkbuf_3_0__f_wb_clk_i (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(clknet_0_wb_clk_i),
    .Y(clknet_3_0__leaf_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__clkbuff_12 clkbuf_3_1__f_wb_clk_i (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(clknet_0_wb_clk_i),
    .Y(clknet_3_1__leaf_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__clkbuff_12 clkbuf_3_2__f_wb_clk_i (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(clknet_0_wb_clk_i),
    .Y(clknet_3_2__leaf_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__clkbuff_12 clkbuf_3_3__f_wb_clk_i (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(clknet_0_wb_clk_i),
    .Y(clknet_3_3__leaf_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__clkbuff_12 clkbuf_3_4__f_wb_clk_i (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(clknet_0_wb_clk_i),
    .Y(clknet_3_4__leaf_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__clkbuff_12 clkbuf_3_5__f_wb_clk_i (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(clknet_0_wb_clk_i),
    .Y(clknet_3_5__leaf_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__clkbuff_12 clkbuf_3_6__f_wb_clk_i (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(clknet_0_wb_clk_i),
    .Y(clknet_3_6__leaf_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__clkbuff_12 clkbuf_3_7__f_wb_clk_i (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(clknet_0_wb_clk_i),
    .Y(clknet_3_7__leaf_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__inv_2 clkload0 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(clknet_3_0__leaf_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__inv_4 clkload1 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(clknet_3_1__leaf_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__inv_4 clkload2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(clknet_3_2__leaf_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__clkbuff_12 clkload3 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(clknet_3_3__leaf_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__inv_2 clkload4 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(clknet_3_4__leaf_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__inv_2 clkload5 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(clknet_3_6__leaf_wb_clk_i));
 gf180mcu_as_sc_mcu7t3v3__buff_2 input1 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(io_in),
    .Y(net1));
 gf180mcu_as_sc_mcu7t3v3__buff_2 input2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(rst_n),
    .Y(net2));
 gf180mcu_as_sc_mcu7t3v3__clkbuff_12 output10 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(net10),
    .Y(io_out[7]));
 gf180mcu_as_sc_mcu7t3v3__clkbuff_12 output11 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(net11),
    .Y(io_out[8]));
 gf180mcu_as_sc_mcu7t3v3__clkbuff_12 output3 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(net3),
    .Y(io_out[0]));
 gf180mcu_as_sc_mcu7t3v3__clkbuff_12 output4 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(net4),
    .Y(io_out[1]));
 gf180mcu_as_sc_mcu7t3v3__clkbuff_12 output5 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(net5),
    .Y(io_out[2]));
 gf180mcu_as_sc_mcu7t3v3__clkbuff_12 output6 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(net6),
    .Y(io_out[3]));
 gf180mcu_as_sc_mcu7t3v3__clkbuff_12 output7 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(net7),
    .Y(io_out[4]));
 gf180mcu_as_sc_mcu7t3v3__clkbuff_12 output8 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(net8),
    .Y(io_out[5]));
 gf180mcu_as_sc_mcu7t3v3__clkbuff_12 output9 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss),
    .A(net9),
    .Y(io_out[6]));
endmodule
