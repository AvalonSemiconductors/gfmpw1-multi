magic
tech gf180mcuD
timestamp 1638034600
<< fillblock >>
rect 0 -3522 3000 0
<< metal4 >>
rect 0 -2250 6 -2244
rect 0 -2256 6 -2250
rect 0 -2262 6 -2256
rect 0 -2268 6 -2262
rect 0 -2274 6 -2268
rect 0 -2280 6 -2274
rect 0 -2286 6 -2280
rect 0 -2292 6 -2286
rect 0 -2298 6 -2292
rect 0 -2304 6 -2298
rect 0 -2310 6 -2304
rect 0 -2316 6 -2310
rect 0 -2322 6 -2316
rect 0 -2328 6 -2322
rect 0 -2334 6 -2328
rect 0 -2340 6 -2334
rect 0 -2346 6 -2340
rect 0 -2352 6 -2346
rect 0 -2358 6 -2352
rect 0 -2364 6 -2358
rect 0 -2370 6 -2364
rect 0 -2376 6 -2370
rect 6 -2178 12 -2172
rect 6 -2184 12 -2178
rect 6 -2190 12 -2184
rect 6 -2196 12 -2190
rect 6 -2202 12 -2196
rect 6 -2208 12 -2202
rect 6 -2214 12 -2208
rect 6 -2220 12 -2214
rect 6 -2226 12 -2220
rect 6 -2232 12 -2226
rect 6 -2238 12 -2232
rect 6 -2244 12 -2238
rect 6 -2250 12 -2244
rect 6 -2256 12 -2250
rect 6 -2262 12 -2256
rect 6 -2268 12 -2262
rect 6 -2274 12 -2268
rect 6 -2280 12 -2274
rect 6 -2286 12 -2280
rect 6 -2292 12 -2286
rect 6 -2298 12 -2292
rect 6 -2304 12 -2298
rect 6 -2310 12 -2304
rect 6 -2316 12 -2310
rect 6 -2322 12 -2316
rect 6 -2328 12 -2322
rect 6 -2334 12 -2328
rect 6 -2340 12 -2334
rect 6 -2346 12 -2340
rect 6 -2352 12 -2346
rect 6 -2358 12 -2352
rect 6 -2364 12 -2358
rect 6 -2370 12 -2364
rect 6 -2376 12 -2370
rect 6 -2382 12 -2376
rect 6 -2388 12 -2382
rect 6 -2394 12 -2388
rect 6 -2400 12 -2394
rect 6 -2406 12 -2400
rect 6 -2412 12 -2406
rect 6 -2418 12 -2412
rect 6 -2424 12 -2418
rect 6 -2430 12 -2424
rect 6 -2436 12 -2430
rect 6 -2442 12 -2436
rect 6 -2448 12 -2442
rect 12 -2136 18 -2130
rect 12 -2142 18 -2136
rect 12 -2148 18 -2142
rect 12 -2154 18 -2148
rect 12 -2160 18 -2154
rect 12 -2166 18 -2160
rect 12 -2172 18 -2166
rect 12 -2178 18 -2172
rect 12 -2184 18 -2178
rect 12 -2190 18 -2184
rect 12 -2196 18 -2190
rect 12 -2202 18 -2196
rect 12 -2208 18 -2202
rect 12 -2214 18 -2208
rect 12 -2220 18 -2214
rect 12 -2226 18 -2220
rect 12 -2232 18 -2226
rect 12 -2238 18 -2232
rect 12 -2244 18 -2238
rect 12 -2250 18 -2244
rect 12 -2256 18 -2250
rect 12 -2262 18 -2256
rect 12 -2268 18 -2262
rect 12 -2274 18 -2268
rect 12 -2280 18 -2274
rect 12 -2286 18 -2280
rect 12 -2292 18 -2286
rect 12 -2298 18 -2292
rect 12 -2304 18 -2298
rect 12 -2310 18 -2304
rect 12 -2316 18 -2310
rect 12 -2322 18 -2316
rect 12 -2328 18 -2322
rect 12 -2334 18 -2328
rect 12 -2340 18 -2334
rect 12 -2346 18 -2340
rect 12 -2352 18 -2346
rect 12 -2358 18 -2352
rect 12 -2364 18 -2358
rect 12 -2370 18 -2364
rect 12 -2376 18 -2370
rect 12 -2382 18 -2376
rect 12 -2388 18 -2382
rect 12 -2394 18 -2388
rect 12 -2400 18 -2394
rect 12 -2406 18 -2400
rect 12 -2412 18 -2406
rect 12 -2418 18 -2412
rect 12 -2424 18 -2418
rect 12 -2430 18 -2424
rect 12 -2436 18 -2430
rect 12 -2442 18 -2436
rect 12 -2448 18 -2442
rect 12 -2454 18 -2448
rect 12 -2460 18 -2454
rect 12 -2466 18 -2460
rect 12 -2472 18 -2466
rect 12 -2478 18 -2472
rect 12 -2484 18 -2478
rect 12 -2490 18 -2484
rect 18 -2100 24 -2094
rect 18 -2106 24 -2100
rect 18 -2112 24 -2106
rect 18 -2118 24 -2112
rect 18 -2124 24 -2118
rect 18 -2130 24 -2124
rect 18 -2136 24 -2130
rect 18 -2142 24 -2136
rect 18 -2148 24 -2142
rect 18 -2154 24 -2148
rect 18 -2160 24 -2154
rect 18 -2166 24 -2160
rect 18 -2172 24 -2166
rect 18 -2178 24 -2172
rect 18 -2184 24 -2178
rect 18 -2190 24 -2184
rect 18 -2196 24 -2190
rect 18 -2202 24 -2196
rect 18 -2208 24 -2202
rect 18 -2214 24 -2208
rect 18 -2220 24 -2214
rect 18 -2226 24 -2220
rect 18 -2232 24 -2226
rect 18 -2238 24 -2232
rect 18 -2244 24 -2238
rect 18 -2250 24 -2244
rect 18 -2256 24 -2250
rect 18 -2262 24 -2256
rect 18 -2268 24 -2262
rect 18 -2274 24 -2268
rect 18 -2280 24 -2274
rect 18 -2286 24 -2280
rect 18 -2292 24 -2286
rect 18 -2298 24 -2292
rect 18 -2304 24 -2298
rect 18 -2310 24 -2304
rect 18 -2316 24 -2310
rect 18 -2322 24 -2316
rect 18 -2328 24 -2322
rect 18 -2334 24 -2328
rect 18 -2340 24 -2334
rect 18 -2346 24 -2340
rect 18 -2352 24 -2346
rect 18 -2358 24 -2352
rect 18 -2364 24 -2358
rect 18 -2370 24 -2364
rect 18 -2376 24 -2370
rect 18 -2382 24 -2376
rect 18 -2388 24 -2382
rect 18 -2394 24 -2388
rect 18 -2400 24 -2394
rect 18 -2406 24 -2400
rect 18 -2412 24 -2406
rect 18 -2418 24 -2412
rect 18 -2424 24 -2418
rect 18 -2430 24 -2424
rect 18 -2436 24 -2430
rect 18 -2442 24 -2436
rect 18 -2448 24 -2442
rect 18 -2454 24 -2448
rect 18 -2460 24 -2454
rect 18 -2466 24 -2460
rect 18 -2472 24 -2466
rect 18 -2478 24 -2472
rect 18 -2484 24 -2478
rect 18 -2490 24 -2484
rect 18 -2496 24 -2490
rect 18 -2502 24 -2496
rect 18 -2508 24 -2502
rect 18 -2514 24 -2508
rect 18 -2520 24 -2514
rect 18 -2526 24 -2520
rect 24 -2070 30 -2064
rect 24 -2076 30 -2070
rect 24 -2082 30 -2076
rect 24 -2088 30 -2082
rect 24 -2094 30 -2088
rect 24 -2100 30 -2094
rect 24 -2106 30 -2100
rect 24 -2112 30 -2106
rect 24 -2118 30 -2112
rect 24 -2124 30 -2118
rect 24 -2130 30 -2124
rect 24 -2136 30 -2130
rect 24 -2142 30 -2136
rect 24 -2148 30 -2142
rect 24 -2154 30 -2148
rect 24 -2160 30 -2154
rect 24 -2166 30 -2160
rect 24 -2172 30 -2166
rect 24 -2178 30 -2172
rect 24 -2184 30 -2178
rect 24 -2190 30 -2184
rect 24 -2196 30 -2190
rect 24 -2202 30 -2196
rect 24 -2208 30 -2202
rect 24 -2214 30 -2208
rect 24 -2220 30 -2214
rect 24 -2226 30 -2220
rect 24 -2232 30 -2226
rect 24 -2238 30 -2232
rect 24 -2244 30 -2238
rect 24 -2250 30 -2244
rect 24 -2256 30 -2250
rect 24 -2262 30 -2256
rect 24 -2268 30 -2262
rect 24 -2274 30 -2268
rect 24 -2280 30 -2274
rect 24 -2286 30 -2280
rect 24 -2292 30 -2286
rect 24 -2298 30 -2292
rect 24 -2304 30 -2298
rect 24 -2310 30 -2304
rect 24 -2316 30 -2310
rect 24 -2322 30 -2316
rect 24 -2328 30 -2322
rect 24 -2334 30 -2328
rect 24 -2340 30 -2334
rect 24 -2346 30 -2340
rect 24 -2352 30 -2346
rect 24 -2358 30 -2352
rect 24 -2364 30 -2358
rect 24 -2370 30 -2364
rect 24 -2376 30 -2370
rect 24 -2382 30 -2376
rect 24 -2388 30 -2382
rect 24 -2394 30 -2388
rect 24 -2400 30 -2394
rect 24 -2406 30 -2400
rect 24 -2412 30 -2406
rect 24 -2418 30 -2412
rect 24 -2424 30 -2418
rect 24 -2430 30 -2424
rect 24 -2436 30 -2430
rect 24 -2442 30 -2436
rect 24 -2448 30 -2442
rect 24 -2454 30 -2448
rect 24 -2460 30 -2454
rect 24 -2466 30 -2460
rect 24 -2472 30 -2466
rect 24 -2478 30 -2472
rect 24 -2484 30 -2478
rect 24 -2490 30 -2484
rect 24 -2496 30 -2490
rect 24 -2502 30 -2496
rect 24 -2508 30 -2502
rect 24 -2514 30 -2508
rect 24 -2520 30 -2514
rect 24 -2526 30 -2520
rect 24 -2532 30 -2526
rect 24 -2538 30 -2532
rect 24 -2544 30 -2538
rect 24 -2550 30 -2544
rect 24 -2556 30 -2550
rect 24 -2562 30 -2556
rect 30 -2040 36 -2034
rect 30 -2046 36 -2040
rect 30 -2052 36 -2046
rect 30 -2058 36 -2052
rect 30 -2064 36 -2058
rect 30 -2070 36 -2064
rect 30 -2076 36 -2070
rect 30 -2082 36 -2076
rect 30 -2088 36 -2082
rect 30 -2094 36 -2088
rect 30 -2100 36 -2094
rect 30 -2106 36 -2100
rect 30 -2112 36 -2106
rect 30 -2118 36 -2112
rect 30 -2124 36 -2118
rect 30 -2130 36 -2124
rect 30 -2136 36 -2130
rect 30 -2142 36 -2136
rect 30 -2148 36 -2142
rect 30 -2154 36 -2148
rect 30 -2160 36 -2154
rect 30 -2166 36 -2160
rect 30 -2172 36 -2166
rect 30 -2178 36 -2172
rect 30 -2184 36 -2178
rect 30 -2190 36 -2184
rect 30 -2196 36 -2190
rect 30 -2202 36 -2196
rect 30 -2208 36 -2202
rect 30 -2214 36 -2208
rect 30 -2220 36 -2214
rect 30 -2226 36 -2220
rect 30 -2232 36 -2226
rect 30 -2238 36 -2232
rect 30 -2244 36 -2238
rect 30 -2250 36 -2244
rect 30 -2256 36 -2250
rect 30 -2262 36 -2256
rect 30 -2268 36 -2262
rect 30 -2274 36 -2268
rect 30 -2280 36 -2274
rect 30 -2286 36 -2280
rect 30 -2292 36 -2286
rect 30 -2298 36 -2292
rect 30 -2304 36 -2298
rect 30 -2310 36 -2304
rect 30 -2316 36 -2310
rect 30 -2322 36 -2316
rect 30 -2328 36 -2322
rect 30 -2334 36 -2328
rect 30 -2340 36 -2334
rect 30 -2346 36 -2340
rect 30 -2352 36 -2346
rect 30 -2358 36 -2352
rect 30 -2364 36 -2358
rect 30 -2370 36 -2364
rect 30 -2376 36 -2370
rect 30 -2382 36 -2376
rect 30 -2388 36 -2382
rect 30 -2394 36 -2388
rect 30 -2400 36 -2394
rect 30 -2406 36 -2400
rect 30 -2412 36 -2406
rect 30 -2418 36 -2412
rect 30 -2424 36 -2418
rect 30 -2430 36 -2424
rect 30 -2436 36 -2430
rect 30 -2442 36 -2436
rect 30 -2448 36 -2442
rect 30 -2454 36 -2448
rect 30 -2460 36 -2454
rect 30 -2466 36 -2460
rect 30 -2472 36 -2466
rect 30 -2478 36 -2472
rect 30 -2484 36 -2478
rect 30 -2490 36 -2484
rect 30 -2496 36 -2490
rect 30 -2502 36 -2496
rect 30 -2508 36 -2502
rect 30 -2514 36 -2508
rect 30 -2520 36 -2514
rect 30 -2526 36 -2520
rect 30 -2532 36 -2526
rect 30 -2538 36 -2532
rect 30 -2544 36 -2538
rect 30 -2550 36 -2544
rect 30 -2556 36 -2550
rect 30 -2562 36 -2556
rect 30 -2568 36 -2562
rect 30 -2574 36 -2568
rect 30 -2580 36 -2574
rect 30 -2586 36 -2580
rect 36 -2016 42 -2010
rect 36 -2022 42 -2016
rect 36 -2028 42 -2022
rect 36 -2034 42 -2028
rect 36 -2040 42 -2034
rect 36 -2046 42 -2040
rect 36 -2052 42 -2046
rect 36 -2058 42 -2052
rect 36 -2064 42 -2058
rect 36 -2070 42 -2064
rect 36 -2076 42 -2070
rect 36 -2082 42 -2076
rect 36 -2088 42 -2082
rect 36 -2094 42 -2088
rect 36 -2100 42 -2094
rect 36 -2106 42 -2100
rect 36 -2112 42 -2106
rect 36 -2118 42 -2112
rect 36 -2124 42 -2118
rect 36 -2130 42 -2124
rect 36 -2136 42 -2130
rect 36 -2142 42 -2136
rect 36 -2148 42 -2142
rect 36 -2154 42 -2148
rect 36 -2160 42 -2154
rect 36 -2166 42 -2160
rect 36 -2172 42 -2166
rect 36 -2178 42 -2172
rect 36 -2184 42 -2178
rect 36 -2190 42 -2184
rect 36 -2196 42 -2190
rect 36 -2202 42 -2196
rect 36 -2208 42 -2202
rect 36 -2214 42 -2208
rect 36 -2220 42 -2214
rect 36 -2226 42 -2220
rect 36 -2232 42 -2226
rect 36 -2238 42 -2232
rect 36 -2244 42 -2238
rect 36 -2250 42 -2244
rect 36 -2256 42 -2250
rect 36 -2262 42 -2256
rect 36 -2268 42 -2262
rect 36 -2274 42 -2268
rect 36 -2280 42 -2274
rect 36 -2286 42 -2280
rect 36 -2292 42 -2286
rect 36 -2298 42 -2292
rect 36 -2304 42 -2298
rect 36 -2310 42 -2304
rect 36 -2316 42 -2310
rect 36 -2322 42 -2316
rect 36 -2328 42 -2322
rect 36 -2334 42 -2328
rect 36 -2340 42 -2334
rect 36 -2346 42 -2340
rect 36 -2352 42 -2346
rect 36 -2358 42 -2352
rect 36 -2364 42 -2358
rect 36 -2370 42 -2364
rect 36 -2376 42 -2370
rect 36 -2382 42 -2376
rect 36 -2388 42 -2382
rect 36 -2394 42 -2388
rect 36 -2400 42 -2394
rect 36 -2406 42 -2400
rect 36 -2412 42 -2406
rect 36 -2418 42 -2412
rect 36 -2424 42 -2418
rect 36 -2430 42 -2424
rect 36 -2436 42 -2430
rect 36 -2442 42 -2436
rect 36 -2448 42 -2442
rect 36 -2454 42 -2448
rect 36 -2460 42 -2454
rect 36 -2466 42 -2460
rect 36 -2472 42 -2466
rect 36 -2478 42 -2472
rect 36 -2484 42 -2478
rect 36 -2490 42 -2484
rect 36 -2496 42 -2490
rect 36 -2502 42 -2496
rect 36 -2508 42 -2502
rect 36 -2514 42 -2508
rect 36 -2520 42 -2514
rect 36 -2526 42 -2520
rect 36 -2532 42 -2526
rect 36 -2538 42 -2532
rect 36 -2544 42 -2538
rect 36 -2550 42 -2544
rect 36 -2556 42 -2550
rect 36 -2562 42 -2556
rect 36 -2568 42 -2562
rect 36 -2574 42 -2568
rect 36 -2580 42 -2574
rect 36 -2586 42 -2580
rect 36 -2592 42 -2586
rect 36 -2598 42 -2592
rect 36 -2604 42 -2598
rect 36 -2610 42 -2604
rect 42 -1992 48 -1986
rect 42 -1998 48 -1992
rect 42 -2004 48 -1998
rect 42 -2010 48 -2004
rect 42 -2016 48 -2010
rect 42 -2022 48 -2016
rect 42 -2028 48 -2022
rect 42 -2034 48 -2028
rect 42 -2040 48 -2034
rect 42 -2046 48 -2040
rect 42 -2052 48 -2046
rect 42 -2058 48 -2052
rect 42 -2064 48 -2058
rect 42 -2070 48 -2064
rect 42 -2076 48 -2070
rect 42 -2082 48 -2076
rect 42 -2088 48 -2082
rect 42 -2094 48 -2088
rect 42 -2100 48 -2094
rect 42 -2106 48 -2100
rect 42 -2112 48 -2106
rect 42 -2118 48 -2112
rect 42 -2124 48 -2118
rect 42 -2130 48 -2124
rect 42 -2136 48 -2130
rect 42 -2142 48 -2136
rect 42 -2148 48 -2142
rect 42 -2154 48 -2148
rect 42 -2160 48 -2154
rect 42 -2166 48 -2160
rect 42 -2172 48 -2166
rect 42 -2178 48 -2172
rect 42 -2184 48 -2178
rect 42 -2190 48 -2184
rect 42 -2196 48 -2190
rect 42 -2202 48 -2196
rect 42 -2208 48 -2202
rect 42 -2214 48 -2208
rect 42 -2220 48 -2214
rect 42 -2226 48 -2220
rect 42 -2232 48 -2226
rect 42 -2238 48 -2232
rect 42 -2244 48 -2238
rect 42 -2250 48 -2244
rect 42 -2256 48 -2250
rect 42 -2262 48 -2256
rect 42 -2268 48 -2262
rect 42 -2274 48 -2268
rect 42 -2280 48 -2274
rect 42 -2286 48 -2280
rect 42 -2292 48 -2286
rect 42 -2298 48 -2292
rect 42 -2304 48 -2298
rect 42 -2310 48 -2304
rect 42 -2316 48 -2310
rect 42 -2322 48 -2316
rect 42 -2328 48 -2322
rect 42 -2334 48 -2328
rect 42 -2340 48 -2334
rect 42 -2346 48 -2340
rect 42 -2352 48 -2346
rect 42 -2358 48 -2352
rect 42 -2364 48 -2358
rect 42 -2370 48 -2364
rect 42 -2376 48 -2370
rect 42 -2382 48 -2376
rect 42 -2388 48 -2382
rect 42 -2394 48 -2388
rect 42 -2400 48 -2394
rect 42 -2406 48 -2400
rect 42 -2412 48 -2406
rect 42 -2418 48 -2412
rect 42 -2424 48 -2418
rect 42 -2430 48 -2424
rect 42 -2436 48 -2430
rect 42 -2442 48 -2436
rect 42 -2448 48 -2442
rect 42 -2454 48 -2448
rect 42 -2460 48 -2454
rect 42 -2466 48 -2460
rect 42 -2472 48 -2466
rect 42 -2478 48 -2472
rect 42 -2484 48 -2478
rect 42 -2490 48 -2484
rect 42 -2496 48 -2490
rect 42 -2502 48 -2496
rect 42 -2508 48 -2502
rect 42 -2514 48 -2508
rect 42 -2520 48 -2514
rect 42 -2526 48 -2520
rect 42 -2532 48 -2526
rect 42 -2538 48 -2532
rect 42 -2544 48 -2538
rect 42 -2550 48 -2544
rect 42 -2556 48 -2550
rect 42 -2562 48 -2556
rect 42 -2568 48 -2562
rect 42 -2574 48 -2568
rect 42 -2580 48 -2574
rect 42 -2586 48 -2580
rect 42 -2592 48 -2586
rect 42 -2598 48 -2592
rect 42 -2604 48 -2598
rect 42 -2610 48 -2604
rect 42 -2616 48 -2610
rect 42 -2622 48 -2616
rect 42 -2628 48 -2622
rect 42 -2634 48 -2628
rect 48 -1974 54 -1968
rect 48 -1980 54 -1974
rect 48 -1986 54 -1980
rect 48 -1992 54 -1986
rect 48 -1998 54 -1992
rect 48 -2004 54 -1998
rect 48 -2010 54 -2004
rect 48 -2016 54 -2010
rect 48 -2022 54 -2016
rect 48 -2028 54 -2022
rect 48 -2034 54 -2028
rect 48 -2040 54 -2034
rect 48 -2046 54 -2040
rect 48 -2052 54 -2046
rect 48 -2058 54 -2052
rect 48 -2064 54 -2058
rect 48 -2070 54 -2064
rect 48 -2076 54 -2070
rect 48 -2082 54 -2076
rect 48 -2088 54 -2082
rect 48 -2094 54 -2088
rect 48 -2100 54 -2094
rect 48 -2106 54 -2100
rect 48 -2112 54 -2106
rect 48 -2118 54 -2112
rect 48 -2124 54 -2118
rect 48 -2130 54 -2124
rect 48 -2136 54 -2130
rect 48 -2142 54 -2136
rect 48 -2148 54 -2142
rect 48 -2154 54 -2148
rect 48 -2160 54 -2154
rect 48 -2166 54 -2160
rect 48 -2172 54 -2166
rect 48 -2178 54 -2172
rect 48 -2184 54 -2178
rect 48 -2190 54 -2184
rect 48 -2196 54 -2190
rect 48 -2202 54 -2196
rect 48 -2208 54 -2202
rect 48 -2214 54 -2208
rect 48 -2220 54 -2214
rect 48 -2226 54 -2220
rect 48 -2232 54 -2226
rect 48 -2238 54 -2232
rect 48 -2244 54 -2238
rect 48 -2250 54 -2244
rect 48 -2256 54 -2250
rect 48 -2262 54 -2256
rect 48 -2268 54 -2262
rect 48 -2274 54 -2268
rect 48 -2280 54 -2274
rect 48 -2286 54 -2280
rect 48 -2292 54 -2286
rect 48 -2298 54 -2292
rect 48 -2304 54 -2298
rect 48 -2310 54 -2304
rect 48 -2316 54 -2310
rect 48 -2322 54 -2316
rect 48 -2328 54 -2322
rect 48 -2334 54 -2328
rect 48 -2340 54 -2334
rect 48 -2346 54 -2340
rect 48 -2352 54 -2346
rect 48 -2358 54 -2352
rect 48 -2364 54 -2358
rect 48 -2370 54 -2364
rect 48 -2376 54 -2370
rect 48 -2382 54 -2376
rect 48 -2388 54 -2382
rect 48 -2394 54 -2388
rect 48 -2400 54 -2394
rect 48 -2406 54 -2400
rect 48 -2412 54 -2406
rect 48 -2418 54 -2412
rect 48 -2424 54 -2418
rect 48 -2430 54 -2424
rect 48 -2436 54 -2430
rect 48 -2442 54 -2436
rect 48 -2448 54 -2442
rect 48 -2454 54 -2448
rect 48 -2460 54 -2454
rect 48 -2466 54 -2460
rect 48 -2472 54 -2466
rect 48 -2478 54 -2472
rect 48 -2484 54 -2478
rect 48 -2490 54 -2484
rect 48 -2496 54 -2490
rect 48 -2502 54 -2496
rect 48 -2508 54 -2502
rect 48 -2514 54 -2508
rect 48 -2520 54 -2514
rect 48 -2526 54 -2520
rect 48 -2532 54 -2526
rect 48 -2538 54 -2532
rect 48 -2544 54 -2538
rect 48 -2550 54 -2544
rect 48 -2556 54 -2550
rect 48 -2562 54 -2556
rect 48 -2568 54 -2562
rect 48 -2574 54 -2568
rect 48 -2580 54 -2574
rect 48 -2586 54 -2580
rect 48 -2592 54 -2586
rect 48 -2598 54 -2592
rect 48 -2604 54 -2598
rect 48 -2610 54 -2604
rect 48 -2616 54 -2610
rect 48 -2622 54 -2616
rect 48 -2628 54 -2622
rect 48 -2634 54 -2628
rect 48 -2640 54 -2634
rect 48 -2646 54 -2640
rect 48 -2652 54 -2646
rect 54 -1950 60 -1944
rect 54 -1956 60 -1950
rect 54 -1962 60 -1956
rect 54 -1968 60 -1962
rect 54 -1974 60 -1968
rect 54 -1980 60 -1974
rect 54 -1986 60 -1980
rect 54 -1992 60 -1986
rect 54 -1998 60 -1992
rect 54 -2004 60 -1998
rect 54 -2010 60 -2004
rect 54 -2016 60 -2010
rect 54 -2022 60 -2016
rect 54 -2028 60 -2022
rect 54 -2034 60 -2028
rect 54 -2040 60 -2034
rect 54 -2046 60 -2040
rect 54 -2052 60 -2046
rect 54 -2058 60 -2052
rect 54 -2064 60 -2058
rect 54 -2070 60 -2064
rect 54 -2076 60 -2070
rect 54 -2082 60 -2076
rect 54 -2088 60 -2082
rect 54 -2094 60 -2088
rect 54 -2100 60 -2094
rect 54 -2106 60 -2100
rect 54 -2112 60 -2106
rect 54 -2118 60 -2112
rect 54 -2124 60 -2118
rect 54 -2130 60 -2124
rect 54 -2136 60 -2130
rect 54 -2142 60 -2136
rect 54 -2148 60 -2142
rect 54 -2154 60 -2148
rect 54 -2160 60 -2154
rect 54 -2166 60 -2160
rect 54 -2172 60 -2166
rect 54 -2178 60 -2172
rect 54 -2184 60 -2178
rect 54 -2190 60 -2184
rect 54 -2196 60 -2190
rect 54 -2202 60 -2196
rect 54 -2208 60 -2202
rect 54 -2214 60 -2208
rect 54 -2220 60 -2214
rect 54 -2226 60 -2220
rect 54 -2232 60 -2226
rect 54 -2238 60 -2232
rect 54 -2244 60 -2238
rect 54 -2250 60 -2244
rect 54 -2256 60 -2250
rect 54 -2262 60 -2256
rect 54 -2268 60 -2262
rect 54 -2274 60 -2268
rect 54 -2280 60 -2274
rect 54 -2286 60 -2280
rect 54 -2292 60 -2286
rect 54 -2298 60 -2292
rect 54 -2304 60 -2298
rect 54 -2310 60 -2304
rect 54 -2316 60 -2310
rect 54 -2322 60 -2316
rect 54 -2328 60 -2322
rect 54 -2334 60 -2328
rect 54 -2340 60 -2334
rect 54 -2346 60 -2340
rect 54 -2352 60 -2346
rect 54 -2358 60 -2352
rect 54 -2364 60 -2358
rect 54 -2370 60 -2364
rect 54 -2376 60 -2370
rect 54 -2382 60 -2376
rect 54 -2388 60 -2382
rect 54 -2394 60 -2388
rect 54 -2400 60 -2394
rect 54 -2406 60 -2400
rect 54 -2412 60 -2406
rect 54 -2418 60 -2412
rect 54 -2424 60 -2418
rect 54 -2430 60 -2424
rect 54 -2436 60 -2430
rect 54 -2442 60 -2436
rect 54 -2448 60 -2442
rect 54 -2454 60 -2448
rect 54 -2460 60 -2454
rect 54 -2466 60 -2460
rect 54 -2472 60 -2466
rect 54 -2478 60 -2472
rect 54 -2484 60 -2478
rect 54 -2490 60 -2484
rect 54 -2496 60 -2490
rect 54 -2502 60 -2496
rect 54 -2508 60 -2502
rect 54 -2514 60 -2508
rect 54 -2520 60 -2514
rect 54 -2526 60 -2520
rect 54 -2532 60 -2526
rect 54 -2538 60 -2532
rect 54 -2544 60 -2538
rect 54 -2550 60 -2544
rect 54 -2556 60 -2550
rect 54 -2562 60 -2556
rect 54 -2568 60 -2562
rect 54 -2574 60 -2568
rect 54 -2580 60 -2574
rect 54 -2586 60 -2580
rect 54 -2592 60 -2586
rect 54 -2598 60 -2592
rect 54 -2604 60 -2598
rect 54 -2610 60 -2604
rect 54 -2616 60 -2610
rect 54 -2622 60 -2616
rect 54 -2628 60 -2622
rect 54 -2634 60 -2628
rect 54 -2640 60 -2634
rect 54 -2646 60 -2640
rect 54 -2652 60 -2646
rect 54 -2658 60 -2652
rect 54 -2664 60 -2658
rect 54 -2670 60 -2664
rect 54 -2676 60 -2670
rect 60 -1932 66 -1926
rect 60 -1938 66 -1932
rect 60 -1944 66 -1938
rect 60 -1950 66 -1944
rect 60 -1956 66 -1950
rect 60 -1962 66 -1956
rect 60 -1968 66 -1962
rect 60 -1974 66 -1968
rect 60 -1980 66 -1974
rect 60 -1986 66 -1980
rect 60 -1992 66 -1986
rect 60 -1998 66 -1992
rect 60 -2004 66 -1998
rect 60 -2010 66 -2004
rect 60 -2016 66 -2010
rect 60 -2022 66 -2016
rect 60 -2028 66 -2022
rect 60 -2034 66 -2028
rect 60 -2040 66 -2034
rect 60 -2046 66 -2040
rect 60 -2052 66 -2046
rect 60 -2058 66 -2052
rect 60 -2064 66 -2058
rect 60 -2070 66 -2064
rect 60 -2076 66 -2070
rect 60 -2082 66 -2076
rect 60 -2088 66 -2082
rect 60 -2094 66 -2088
rect 60 -2100 66 -2094
rect 60 -2106 66 -2100
rect 60 -2112 66 -2106
rect 60 -2118 66 -2112
rect 60 -2124 66 -2118
rect 60 -2130 66 -2124
rect 60 -2136 66 -2130
rect 60 -2142 66 -2136
rect 60 -2148 66 -2142
rect 60 -2154 66 -2148
rect 60 -2160 66 -2154
rect 60 -2166 66 -2160
rect 60 -2172 66 -2166
rect 60 -2178 66 -2172
rect 60 -2184 66 -2178
rect 60 -2190 66 -2184
rect 60 -2196 66 -2190
rect 60 -2202 66 -2196
rect 60 -2208 66 -2202
rect 60 -2214 66 -2208
rect 60 -2220 66 -2214
rect 60 -2226 66 -2220
rect 60 -2232 66 -2226
rect 60 -2238 66 -2232
rect 60 -2244 66 -2238
rect 60 -2250 66 -2244
rect 60 -2256 66 -2250
rect 60 -2262 66 -2256
rect 60 -2268 66 -2262
rect 60 -2274 66 -2268
rect 60 -2280 66 -2274
rect 60 -2286 66 -2280
rect 60 -2292 66 -2286
rect 60 -2298 66 -2292
rect 60 -2304 66 -2298
rect 60 -2310 66 -2304
rect 60 -2316 66 -2310
rect 60 -2322 66 -2316
rect 60 -2328 66 -2322
rect 60 -2334 66 -2328
rect 60 -2340 66 -2334
rect 60 -2346 66 -2340
rect 60 -2352 66 -2346
rect 60 -2358 66 -2352
rect 60 -2364 66 -2358
rect 60 -2370 66 -2364
rect 60 -2376 66 -2370
rect 60 -2382 66 -2376
rect 60 -2388 66 -2382
rect 60 -2394 66 -2388
rect 60 -2400 66 -2394
rect 60 -2406 66 -2400
rect 60 -2412 66 -2406
rect 60 -2418 66 -2412
rect 60 -2424 66 -2418
rect 60 -2430 66 -2424
rect 60 -2436 66 -2430
rect 60 -2442 66 -2436
rect 60 -2448 66 -2442
rect 60 -2454 66 -2448
rect 60 -2460 66 -2454
rect 60 -2466 66 -2460
rect 60 -2472 66 -2466
rect 60 -2478 66 -2472
rect 60 -2484 66 -2478
rect 60 -2490 66 -2484
rect 60 -2496 66 -2490
rect 60 -2502 66 -2496
rect 60 -2508 66 -2502
rect 60 -2514 66 -2508
rect 60 -2520 66 -2514
rect 60 -2526 66 -2520
rect 60 -2532 66 -2526
rect 60 -2538 66 -2532
rect 60 -2544 66 -2538
rect 60 -2550 66 -2544
rect 60 -2556 66 -2550
rect 60 -2562 66 -2556
rect 60 -2568 66 -2562
rect 60 -2574 66 -2568
rect 60 -2580 66 -2574
rect 60 -2586 66 -2580
rect 60 -2592 66 -2586
rect 60 -2598 66 -2592
rect 60 -2604 66 -2598
rect 60 -2610 66 -2604
rect 60 -2616 66 -2610
rect 60 -2622 66 -2616
rect 60 -2628 66 -2622
rect 60 -2634 66 -2628
rect 60 -2640 66 -2634
rect 60 -2646 66 -2640
rect 60 -2652 66 -2646
rect 60 -2658 66 -2652
rect 60 -2664 66 -2658
rect 60 -2670 66 -2664
rect 60 -2676 66 -2670
rect 60 -2682 66 -2676
rect 60 -2688 66 -2682
rect 60 -2694 66 -2688
rect 66 -1914 72 -1908
rect 66 -1920 72 -1914
rect 66 -1926 72 -1920
rect 66 -1932 72 -1926
rect 66 -1938 72 -1932
rect 66 -1944 72 -1938
rect 66 -1950 72 -1944
rect 66 -1956 72 -1950
rect 66 -1962 72 -1956
rect 66 -1968 72 -1962
rect 66 -1974 72 -1968
rect 66 -1980 72 -1974
rect 66 -1986 72 -1980
rect 66 -1992 72 -1986
rect 66 -1998 72 -1992
rect 66 -2004 72 -1998
rect 66 -2010 72 -2004
rect 66 -2016 72 -2010
rect 66 -2022 72 -2016
rect 66 -2028 72 -2022
rect 66 -2034 72 -2028
rect 66 -2040 72 -2034
rect 66 -2046 72 -2040
rect 66 -2052 72 -2046
rect 66 -2058 72 -2052
rect 66 -2064 72 -2058
rect 66 -2070 72 -2064
rect 66 -2076 72 -2070
rect 66 -2082 72 -2076
rect 66 -2088 72 -2082
rect 66 -2094 72 -2088
rect 66 -2100 72 -2094
rect 66 -2106 72 -2100
rect 66 -2112 72 -2106
rect 66 -2118 72 -2112
rect 66 -2124 72 -2118
rect 66 -2130 72 -2124
rect 66 -2136 72 -2130
rect 66 -2142 72 -2136
rect 66 -2148 72 -2142
rect 66 -2154 72 -2148
rect 66 -2160 72 -2154
rect 66 -2166 72 -2160
rect 66 -2172 72 -2166
rect 66 -2178 72 -2172
rect 66 -2184 72 -2178
rect 66 -2190 72 -2184
rect 66 -2196 72 -2190
rect 66 -2202 72 -2196
rect 66 -2208 72 -2202
rect 66 -2214 72 -2208
rect 66 -2220 72 -2214
rect 66 -2226 72 -2220
rect 66 -2232 72 -2226
rect 66 -2238 72 -2232
rect 66 -2244 72 -2238
rect 66 -2250 72 -2244
rect 66 -2256 72 -2250
rect 66 -2262 72 -2256
rect 66 -2268 72 -2262
rect 66 -2274 72 -2268
rect 66 -2280 72 -2274
rect 66 -2286 72 -2280
rect 66 -2292 72 -2286
rect 66 -2298 72 -2292
rect 66 -2304 72 -2298
rect 66 -2310 72 -2304
rect 66 -2316 72 -2310
rect 66 -2322 72 -2316
rect 66 -2328 72 -2322
rect 66 -2334 72 -2328
rect 66 -2340 72 -2334
rect 66 -2346 72 -2340
rect 66 -2352 72 -2346
rect 66 -2358 72 -2352
rect 66 -2364 72 -2358
rect 66 -2370 72 -2364
rect 66 -2376 72 -2370
rect 66 -2382 72 -2376
rect 66 -2388 72 -2382
rect 66 -2394 72 -2388
rect 66 -2400 72 -2394
rect 66 -2406 72 -2400
rect 66 -2412 72 -2406
rect 66 -2418 72 -2412
rect 66 -2424 72 -2418
rect 66 -2430 72 -2424
rect 66 -2436 72 -2430
rect 66 -2442 72 -2436
rect 66 -2448 72 -2442
rect 66 -2454 72 -2448
rect 66 -2460 72 -2454
rect 66 -2466 72 -2460
rect 66 -2472 72 -2466
rect 66 -2478 72 -2472
rect 66 -2484 72 -2478
rect 66 -2490 72 -2484
rect 66 -2496 72 -2490
rect 66 -2502 72 -2496
rect 66 -2508 72 -2502
rect 66 -2514 72 -2508
rect 66 -2520 72 -2514
rect 66 -2526 72 -2520
rect 66 -2532 72 -2526
rect 66 -2538 72 -2532
rect 66 -2544 72 -2538
rect 66 -2550 72 -2544
rect 66 -2556 72 -2550
rect 66 -2562 72 -2556
rect 66 -2568 72 -2562
rect 66 -2574 72 -2568
rect 66 -2580 72 -2574
rect 66 -2586 72 -2580
rect 66 -2592 72 -2586
rect 66 -2598 72 -2592
rect 66 -2604 72 -2598
rect 66 -2610 72 -2604
rect 66 -2616 72 -2610
rect 66 -2622 72 -2616
rect 66 -2628 72 -2622
rect 66 -2634 72 -2628
rect 66 -2640 72 -2634
rect 66 -2646 72 -2640
rect 66 -2652 72 -2646
rect 66 -2658 72 -2652
rect 66 -2664 72 -2658
rect 66 -2670 72 -2664
rect 66 -2676 72 -2670
rect 66 -2682 72 -2676
rect 66 -2688 72 -2682
rect 66 -2694 72 -2688
rect 66 -2700 72 -2694
rect 66 -2706 72 -2700
rect 66 -2712 72 -2706
rect 72 -1902 78 -1896
rect 72 -1908 78 -1902
rect 72 -1914 78 -1908
rect 72 -1920 78 -1914
rect 72 -1926 78 -1920
rect 72 -1932 78 -1926
rect 72 -1938 78 -1932
rect 72 -1944 78 -1938
rect 72 -1950 78 -1944
rect 72 -1956 78 -1950
rect 72 -1962 78 -1956
rect 72 -1968 78 -1962
rect 72 -1974 78 -1968
rect 72 -1980 78 -1974
rect 72 -1986 78 -1980
rect 72 -1992 78 -1986
rect 72 -1998 78 -1992
rect 72 -2004 78 -1998
rect 72 -2010 78 -2004
rect 72 -2016 78 -2010
rect 72 -2022 78 -2016
rect 72 -2028 78 -2022
rect 72 -2034 78 -2028
rect 72 -2040 78 -2034
rect 72 -2046 78 -2040
rect 72 -2052 78 -2046
rect 72 -2058 78 -2052
rect 72 -2064 78 -2058
rect 72 -2070 78 -2064
rect 72 -2076 78 -2070
rect 72 -2082 78 -2076
rect 72 -2088 78 -2082
rect 72 -2094 78 -2088
rect 72 -2100 78 -2094
rect 72 -2106 78 -2100
rect 72 -2112 78 -2106
rect 72 -2118 78 -2112
rect 72 -2124 78 -2118
rect 72 -2130 78 -2124
rect 72 -2136 78 -2130
rect 72 -2142 78 -2136
rect 72 -2148 78 -2142
rect 72 -2154 78 -2148
rect 72 -2160 78 -2154
rect 72 -2166 78 -2160
rect 72 -2172 78 -2166
rect 72 -2178 78 -2172
rect 72 -2184 78 -2178
rect 72 -2190 78 -2184
rect 72 -2196 78 -2190
rect 72 -2202 78 -2196
rect 72 -2208 78 -2202
rect 72 -2214 78 -2208
rect 72 -2220 78 -2214
rect 72 -2226 78 -2220
rect 72 -2232 78 -2226
rect 72 -2238 78 -2232
rect 72 -2244 78 -2238
rect 72 -2250 78 -2244
rect 72 -2256 78 -2250
rect 72 -2262 78 -2256
rect 72 -2268 78 -2262
rect 72 -2274 78 -2268
rect 72 -2280 78 -2274
rect 72 -2286 78 -2280
rect 72 -2292 78 -2286
rect 72 -2298 78 -2292
rect 72 -2304 78 -2298
rect 72 -2310 78 -2304
rect 72 -2316 78 -2310
rect 72 -2322 78 -2316
rect 72 -2328 78 -2322
rect 72 -2334 78 -2328
rect 72 -2340 78 -2334
rect 72 -2346 78 -2340
rect 72 -2352 78 -2346
rect 72 -2358 78 -2352
rect 72 -2364 78 -2358
rect 72 -2370 78 -2364
rect 72 -2376 78 -2370
rect 72 -2382 78 -2376
rect 72 -2388 78 -2382
rect 72 -2394 78 -2388
rect 72 -2400 78 -2394
rect 72 -2406 78 -2400
rect 72 -2412 78 -2406
rect 72 -2418 78 -2412
rect 72 -2424 78 -2418
rect 72 -2430 78 -2424
rect 72 -2436 78 -2430
rect 72 -2442 78 -2436
rect 72 -2448 78 -2442
rect 72 -2454 78 -2448
rect 72 -2460 78 -2454
rect 72 -2466 78 -2460
rect 72 -2472 78 -2466
rect 72 -2478 78 -2472
rect 72 -2484 78 -2478
rect 72 -2490 78 -2484
rect 72 -2496 78 -2490
rect 72 -2502 78 -2496
rect 72 -2508 78 -2502
rect 72 -2514 78 -2508
rect 72 -2520 78 -2514
rect 72 -2526 78 -2520
rect 72 -2532 78 -2526
rect 72 -2538 78 -2532
rect 72 -2544 78 -2538
rect 72 -2550 78 -2544
rect 72 -2556 78 -2550
rect 72 -2562 78 -2556
rect 72 -2568 78 -2562
rect 72 -2574 78 -2568
rect 72 -2580 78 -2574
rect 72 -2586 78 -2580
rect 72 -2592 78 -2586
rect 72 -2598 78 -2592
rect 72 -2604 78 -2598
rect 72 -2610 78 -2604
rect 72 -2616 78 -2610
rect 72 -2622 78 -2616
rect 72 -2628 78 -2622
rect 72 -2634 78 -2628
rect 72 -2640 78 -2634
rect 72 -2646 78 -2640
rect 72 -2652 78 -2646
rect 72 -2658 78 -2652
rect 72 -2664 78 -2658
rect 72 -2670 78 -2664
rect 72 -2676 78 -2670
rect 72 -2682 78 -2676
rect 72 -2688 78 -2682
rect 72 -2694 78 -2688
rect 72 -2700 78 -2694
rect 72 -2706 78 -2700
rect 72 -2712 78 -2706
rect 72 -2718 78 -2712
rect 72 -2724 78 -2718
rect 78 -1884 84 -1878
rect 78 -1890 84 -1884
rect 78 -1896 84 -1890
rect 78 -1902 84 -1896
rect 78 -1908 84 -1902
rect 78 -1914 84 -1908
rect 78 -1920 84 -1914
rect 78 -1926 84 -1920
rect 78 -1932 84 -1926
rect 78 -1938 84 -1932
rect 78 -1944 84 -1938
rect 78 -1950 84 -1944
rect 78 -1956 84 -1950
rect 78 -1962 84 -1956
rect 78 -1968 84 -1962
rect 78 -1974 84 -1968
rect 78 -1980 84 -1974
rect 78 -1986 84 -1980
rect 78 -1992 84 -1986
rect 78 -1998 84 -1992
rect 78 -2004 84 -1998
rect 78 -2010 84 -2004
rect 78 -2016 84 -2010
rect 78 -2022 84 -2016
rect 78 -2028 84 -2022
rect 78 -2034 84 -2028
rect 78 -2040 84 -2034
rect 78 -2046 84 -2040
rect 78 -2052 84 -2046
rect 78 -2058 84 -2052
rect 78 -2064 84 -2058
rect 78 -2070 84 -2064
rect 78 -2076 84 -2070
rect 78 -2082 84 -2076
rect 78 -2088 84 -2082
rect 78 -2094 84 -2088
rect 78 -2100 84 -2094
rect 78 -2106 84 -2100
rect 78 -2112 84 -2106
rect 78 -2118 84 -2112
rect 78 -2124 84 -2118
rect 78 -2130 84 -2124
rect 78 -2136 84 -2130
rect 78 -2142 84 -2136
rect 78 -2148 84 -2142
rect 78 -2154 84 -2148
rect 78 -2160 84 -2154
rect 78 -2166 84 -2160
rect 78 -2172 84 -2166
rect 78 -2178 84 -2172
rect 78 -2184 84 -2178
rect 78 -2190 84 -2184
rect 78 -2196 84 -2190
rect 78 -2202 84 -2196
rect 78 -2208 84 -2202
rect 78 -2214 84 -2208
rect 78 -2220 84 -2214
rect 78 -2226 84 -2220
rect 78 -2232 84 -2226
rect 78 -2238 84 -2232
rect 78 -2244 84 -2238
rect 78 -2250 84 -2244
rect 78 -2256 84 -2250
rect 78 -2262 84 -2256
rect 78 -2268 84 -2262
rect 78 -2274 84 -2268
rect 78 -2280 84 -2274
rect 78 -2286 84 -2280
rect 78 -2292 84 -2286
rect 78 -2298 84 -2292
rect 78 -2304 84 -2298
rect 78 -2310 84 -2304
rect 78 -2316 84 -2310
rect 78 -2322 84 -2316
rect 78 -2328 84 -2322
rect 78 -2334 84 -2328
rect 78 -2340 84 -2334
rect 78 -2346 84 -2340
rect 78 -2352 84 -2346
rect 78 -2358 84 -2352
rect 78 -2364 84 -2358
rect 78 -2370 84 -2364
rect 78 -2376 84 -2370
rect 78 -2382 84 -2376
rect 78 -2388 84 -2382
rect 78 -2394 84 -2388
rect 78 -2400 84 -2394
rect 78 -2406 84 -2400
rect 78 -2412 84 -2406
rect 78 -2418 84 -2412
rect 78 -2424 84 -2418
rect 78 -2430 84 -2424
rect 78 -2436 84 -2430
rect 78 -2442 84 -2436
rect 78 -2448 84 -2442
rect 78 -2454 84 -2448
rect 78 -2460 84 -2454
rect 78 -2466 84 -2460
rect 78 -2472 84 -2466
rect 78 -2478 84 -2472
rect 78 -2484 84 -2478
rect 78 -2490 84 -2484
rect 78 -2496 84 -2490
rect 78 -2502 84 -2496
rect 78 -2508 84 -2502
rect 78 -2514 84 -2508
rect 78 -2520 84 -2514
rect 78 -2526 84 -2520
rect 78 -2532 84 -2526
rect 78 -2538 84 -2532
rect 78 -2544 84 -2538
rect 78 -2550 84 -2544
rect 78 -2556 84 -2550
rect 78 -2562 84 -2556
rect 78 -2568 84 -2562
rect 78 -2574 84 -2568
rect 78 -2580 84 -2574
rect 78 -2586 84 -2580
rect 78 -2592 84 -2586
rect 78 -2598 84 -2592
rect 78 -2604 84 -2598
rect 78 -2610 84 -2604
rect 78 -2616 84 -2610
rect 78 -2622 84 -2616
rect 78 -2628 84 -2622
rect 78 -2634 84 -2628
rect 78 -2640 84 -2634
rect 78 -2646 84 -2640
rect 78 -2652 84 -2646
rect 78 -2658 84 -2652
rect 78 -2664 84 -2658
rect 78 -2670 84 -2664
rect 78 -2676 84 -2670
rect 78 -2682 84 -2676
rect 78 -2688 84 -2682
rect 78 -2694 84 -2688
rect 78 -2700 84 -2694
rect 78 -2706 84 -2700
rect 78 -2712 84 -2706
rect 78 -2718 84 -2712
rect 78 -2724 84 -2718
rect 78 -2730 84 -2724
rect 78 -2736 84 -2730
rect 78 -2742 84 -2736
rect 84 -1866 90 -1860
rect 84 -1872 90 -1866
rect 84 -1878 90 -1872
rect 84 -1884 90 -1878
rect 84 -1890 90 -1884
rect 84 -1896 90 -1890
rect 84 -1902 90 -1896
rect 84 -1908 90 -1902
rect 84 -1914 90 -1908
rect 84 -1920 90 -1914
rect 84 -1926 90 -1920
rect 84 -1932 90 -1926
rect 84 -1938 90 -1932
rect 84 -1944 90 -1938
rect 84 -1950 90 -1944
rect 84 -1956 90 -1950
rect 84 -1962 90 -1956
rect 84 -1968 90 -1962
rect 84 -1974 90 -1968
rect 84 -1980 90 -1974
rect 84 -1986 90 -1980
rect 84 -1992 90 -1986
rect 84 -1998 90 -1992
rect 84 -2004 90 -1998
rect 84 -2010 90 -2004
rect 84 -2016 90 -2010
rect 84 -2022 90 -2016
rect 84 -2028 90 -2022
rect 84 -2034 90 -2028
rect 84 -2040 90 -2034
rect 84 -2046 90 -2040
rect 84 -2052 90 -2046
rect 84 -2058 90 -2052
rect 84 -2064 90 -2058
rect 84 -2070 90 -2064
rect 84 -2076 90 -2070
rect 84 -2082 90 -2076
rect 84 -2088 90 -2082
rect 84 -2094 90 -2088
rect 84 -2100 90 -2094
rect 84 -2106 90 -2100
rect 84 -2112 90 -2106
rect 84 -2118 90 -2112
rect 84 -2124 90 -2118
rect 84 -2130 90 -2124
rect 84 -2136 90 -2130
rect 84 -2142 90 -2136
rect 84 -2148 90 -2142
rect 84 -2154 90 -2148
rect 84 -2160 90 -2154
rect 84 -2166 90 -2160
rect 84 -2172 90 -2166
rect 84 -2178 90 -2172
rect 84 -2184 90 -2178
rect 84 -2190 90 -2184
rect 84 -2196 90 -2190
rect 84 -2202 90 -2196
rect 84 -2208 90 -2202
rect 84 -2214 90 -2208
rect 84 -2220 90 -2214
rect 84 -2226 90 -2220
rect 84 -2232 90 -2226
rect 84 -2238 90 -2232
rect 84 -2244 90 -2238
rect 84 -2250 90 -2244
rect 84 -2256 90 -2250
rect 84 -2262 90 -2256
rect 84 -2268 90 -2262
rect 84 -2274 90 -2268
rect 84 -2280 90 -2274
rect 84 -2286 90 -2280
rect 84 -2292 90 -2286
rect 84 -2298 90 -2292
rect 84 -2304 90 -2298
rect 84 -2310 90 -2304
rect 84 -2316 90 -2310
rect 84 -2322 90 -2316
rect 84 -2328 90 -2322
rect 84 -2334 90 -2328
rect 84 -2340 90 -2334
rect 84 -2346 90 -2340
rect 84 -2352 90 -2346
rect 84 -2358 90 -2352
rect 84 -2364 90 -2358
rect 84 -2370 90 -2364
rect 84 -2376 90 -2370
rect 84 -2382 90 -2376
rect 84 -2388 90 -2382
rect 84 -2394 90 -2388
rect 84 -2400 90 -2394
rect 84 -2406 90 -2400
rect 84 -2412 90 -2406
rect 84 -2418 90 -2412
rect 84 -2424 90 -2418
rect 84 -2430 90 -2424
rect 84 -2436 90 -2430
rect 84 -2442 90 -2436
rect 84 -2448 90 -2442
rect 84 -2454 90 -2448
rect 84 -2460 90 -2454
rect 84 -2466 90 -2460
rect 84 -2472 90 -2466
rect 84 -2478 90 -2472
rect 84 -2484 90 -2478
rect 84 -2490 90 -2484
rect 84 -2496 90 -2490
rect 84 -2502 90 -2496
rect 84 -2508 90 -2502
rect 84 -2514 90 -2508
rect 84 -2520 90 -2514
rect 84 -2526 90 -2520
rect 84 -2532 90 -2526
rect 84 -2538 90 -2532
rect 84 -2544 90 -2538
rect 84 -2550 90 -2544
rect 84 -2556 90 -2550
rect 84 -2562 90 -2556
rect 84 -2568 90 -2562
rect 84 -2574 90 -2568
rect 84 -2580 90 -2574
rect 84 -2586 90 -2580
rect 84 -2592 90 -2586
rect 84 -2598 90 -2592
rect 84 -2604 90 -2598
rect 84 -2610 90 -2604
rect 84 -2616 90 -2610
rect 84 -2622 90 -2616
rect 84 -2628 90 -2622
rect 84 -2634 90 -2628
rect 84 -2640 90 -2634
rect 84 -2646 90 -2640
rect 84 -2652 90 -2646
rect 84 -2658 90 -2652
rect 84 -2664 90 -2658
rect 84 -2670 90 -2664
rect 84 -2676 90 -2670
rect 84 -2682 90 -2676
rect 84 -2688 90 -2682
rect 84 -2694 90 -2688
rect 84 -2700 90 -2694
rect 84 -2706 90 -2700
rect 84 -2712 90 -2706
rect 84 -2718 90 -2712
rect 84 -2724 90 -2718
rect 84 -2730 90 -2724
rect 84 -2736 90 -2730
rect 84 -2742 90 -2736
rect 84 -2748 90 -2742
rect 84 -2754 90 -2748
rect 84 -2760 90 -2754
rect 90 -1854 96 -1848
rect 90 -1860 96 -1854
rect 90 -1866 96 -1860
rect 90 -1872 96 -1866
rect 90 -1878 96 -1872
rect 90 -1884 96 -1878
rect 90 -1890 96 -1884
rect 90 -1896 96 -1890
rect 90 -1902 96 -1896
rect 90 -1908 96 -1902
rect 90 -1914 96 -1908
rect 90 -1920 96 -1914
rect 90 -1926 96 -1920
rect 90 -1932 96 -1926
rect 90 -1938 96 -1932
rect 90 -1944 96 -1938
rect 90 -1950 96 -1944
rect 90 -1956 96 -1950
rect 90 -1962 96 -1956
rect 90 -1968 96 -1962
rect 90 -1974 96 -1968
rect 90 -1980 96 -1974
rect 90 -1986 96 -1980
rect 90 -1992 96 -1986
rect 90 -1998 96 -1992
rect 90 -2004 96 -1998
rect 90 -2010 96 -2004
rect 90 -2016 96 -2010
rect 90 -2022 96 -2016
rect 90 -2028 96 -2022
rect 90 -2034 96 -2028
rect 90 -2040 96 -2034
rect 90 -2046 96 -2040
rect 90 -2052 96 -2046
rect 90 -2058 96 -2052
rect 90 -2064 96 -2058
rect 90 -2070 96 -2064
rect 90 -2076 96 -2070
rect 90 -2082 96 -2076
rect 90 -2088 96 -2082
rect 90 -2094 96 -2088
rect 90 -2100 96 -2094
rect 90 -2106 96 -2100
rect 90 -2112 96 -2106
rect 90 -2118 96 -2112
rect 90 -2124 96 -2118
rect 90 -2130 96 -2124
rect 90 -2136 96 -2130
rect 90 -2142 96 -2136
rect 90 -2148 96 -2142
rect 90 -2154 96 -2148
rect 90 -2160 96 -2154
rect 90 -2166 96 -2160
rect 90 -2172 96 -2166
rect 90 -2178 96 -2172
rect 90 -2184 96 -2178
rect 90 -2190 96 -2184
rect 90 -2196 96 -2190
rect 90 -2202 96 -2196
rect 90 -2208 96 -2202
rect 90 -2214 96 -2208
rect 90 -2220 96 -2214
rect 90 -2226 96 -2220
rect 90 -2232 96 -2226
rect 90 -2238 96 -2232
rect 90 -2244 96 -2238
rect 90 -2250 96 -2244
rect 90 -2256 96 -2250
rect 90 -2262 96 -2256
rect 90 -2268 96 -2262
rect 90 -2274 96 -2268
rect 90 -2280 96 -2274
rect 90 -2286 96 -2280
rect 90 -2292 96 -2286
rect 90 -2298 96 -2292
rect 90 -2304 96 -2298
rect 90 -2310 96 -2304
rect 90 -2316 96 -2310
rect 90 -2322 96 -2316
rect 90 -2328 96 -2322
rect 90 -2334 96 -2328
rect 90 -2340 96 -2334
rect 90 -2346 96 -2340
rect 90 -2352 96 -2346
rect 90 -2358 96 -2352
rect 90 -2364 96 -2358
rect 90 -2370 96 -2364
rect 90 -2376 96 -2370
rect 90 -2382 96 -2376
rect 90 -2388 96 -2382
rect 90 -2394 96 -2388
rect 90 -2400 96 -2394
rect 90 -2406 96 -2400
rect 90 -2412 96 -2406
rect 90 -2418 96 -2412
rect 90 -2424 96 -2418
rect 90 -2430 96 -2424
rect 90 -2436 96 -2430
rect 90 -2442 96 -2436
rect 90 -2448 96 -2442
rect 90 -2454 96 -2448
rect 90 -2460 96 -2454
rect 90 -2466 96 -2460
rect 90 -2472 96 -2466
rect 90 -2478 96 -2472
rect 90 -2484 96 -2478
rect 90 -2490 96 -2484
rect 90 -2496 96 -2490
rect 90 -2502 96 -2496
rect 90 -2508 96 -2502
rect 90 -2514 96 -2508
rect 90 -2520 96 -2514
rect 90 -2526 96 -2520
rect 90 -2532 96 -2526
rect 90 -2538 96 -2532
rect 90 -2544 96 -2538
rect 90 -2550 96 -2544
rect 90 -2556 96 -2550
rect 90 -2562 96 -2556
rect 90 -2568 96 -2562
rect 90 -2574 96 -2568
rect 90 -2580 96 -2574
rect 90 -2586 96 -2580
rect 90 -2592 96 -2586
rect 90 -2598 96 -2592
rect 90 -2604 96 -2598
rect 90 -2610 96 -2604
rect 90 -2616 96 -2610
rect 90 -2622 96 -2616
rect 90 -2628 96 -2622
rect 90 -2634 96 -2628
rect 90 -2640 96 -2634
rect 90 -2646 96 -2640
rect 90 -2652 96 -2646
rect 90 -2658 96 -2652
rect 90 -2664 96 -2658
rect 90 -2670 96 -2664
rect 90 -2676 96 -2670
rect 90 -2682 96 -2676
rect 90 -2688 96 -2682
rect 90 -2694 96 -2688
rect 90 -2700 96 -2694
rect 90 -2706 96 -2700
rect 90 -2712 96 -2706
rect 90 -2718 96 -2712
rect 90 -2724 96 -2718
rect 90 -2730 96 -2724
rect 90 -2736 96 -2730
rect 90 -2742 96 -2736
rect 90 -2748 96 -2742
rect 90 -2754 96 -2748
rect 90 -2760 96 -2754
rect 90 -2766 96 -2760
rect 90 -2772 96 -2766
rect 96 -1842 102 -1836
rect 96 -1848 102 -1842
rect 96 -1854 102 -1848
rect 96 -1860 102 -1854
rect 96 -1866 102 -1860
rect 96 -1872 102 -1866
rect 96 -1878 102 -1872
rect 96 -1884 102 -1878
rect 96 -1890 102 -1884
rect 96 -1896 102 -1890
rect 96 -1902 102 -1896
rect 96 -1908 102 -1902
rect 96 -1914 102 -1908
rect 96 -1920 102 -1914
rect 96 -1926 102 -1920
rect 96 -1932 102 -1926
rect 96 -1938 102 -1932
rect 96 -1944 102 -1938
rect 96 -1950 102 -1944
rect 96 -1956 102 -1950
rect 96 -1962 102 -1956
rect 96 -1968 102 -1962
rect 96 -1974 102 -1968
rect 96 -1980 102 -1974
rect 96 -1986 102 -1980
rect 96 -1992 102 -1986
rect 96 -1998 102 -1992
rect 96 -2004 102 -1998
rect 96 -2010 102 -2004
rect 96 -2016 102 -2010
rect 96 -2022 102 -2016
rect 96 -2028 102 -2022
rect 96 -2034 102 -2028
rect 96 -2040 102 -2034
rect 96 -2046 102 -2040
rect 96 -2052 102 -2046
rect 96 -2058 102 -2052
rect 96 -2064 102 -2058
rect 96 -2070 102 -2064
rect 96 -2076 102 -2070
rect 96 -2082 102 -2076
rect 96 -2088 102 -2082
rect 96 -2094 102 -2088
rect 96 -2100 102 -2094
rect 96 -2106 102 -2100
rect 96 -2112 102 -2106
rect 96 -2118 102 -2112
rect 96 -2124 102 -2118
rect 96 -2130 102 -2124
rect 96 -2136 102 -2130
rect 96 -2142 102 -2136
rect 96 -2148 102 -2142
rect 96 -2154 102 -2148
rect 96 -2160 102 -2154
rect 96 -2166 102 -2160
rect 96 -2172 102 -2166
rect 96 -2178 102 -2172
rect 96 -2184 102 -2178
rect 96 -2190 102 -2184
rect 96 -2196 102 -2190
rect 96 -2202 102 -2196
rect 96 -2208 102 -2202
rect 96 -2214 102 -2208
rect 96 -2220 102 -2214
rect 96 -2226 102 -2220
rect 96 -2232 102 -2226
rect 96 -2238 102 -2232
rect 96 -2244 102 -2238
rect 96 -2250 102 -2244
rect 96 -2256 102 -2250
rect 96 -2262 102 -2256
rect 96 -2268 102 -2262
rect 96 -2274 102 -2268
rect 96 -2280 102 -2274
rect 96 -2286 102 -2280
rect 96 -2292 102 -2286
rect 96 -2298 102 -2292
rect 96 -2304 102 -2298
rect 96 -2310 102 -2304
rect 96 -2316 102 -2310
rect 96 -2322 102 -2316
rect 96 -2328 102 -2322
rect 96 -2334 102 -2328
rect 96 -2340 102 -2334
rect 96 -2346 102 -2340
rect 96 -2352 102 -2346
rect 96 -2358 102 -2352
rect 96 -2364 102 -2358
rect 96 -2370 102 -2364
rect 96 -2376 102 -2370
rect 96 -2382 102 -2376
rect 96 -2388 102 -2382
rect 96 -2394 102 -2388
rect 96 -2400 102 -2394
rect 96 -2406 102 -2400
rect 96 -2412 102 -2406
rect 96 -2418 102 -2412
rect 96 -2424 102 -2418
rect 96 -2430 102 -2424
rect 96 -2436 102 -2430
rect 96 -2442 102 -2436
rect 96 -2448 102 -2442
rect 96 -2454 102 -2448
rect 96 -2460 102 -2454
rect 96 -2466 102 -2460
rect 96 -2472 102 -2466
rect 96 -2478 102 -2472
rect 96 -2484 102 -2478
rect 96 -2490 102 -2484
rect 96 -2496 102 -2490
rect 96 -2502 102 -2496
rect 96 -2508 102 -2502
rect 96 -2514 102 -2508
rect 96 -2520 102 -2514
rect 96 -2526 102 -2520
rect 96 -2532 102 -2526
rect 96 -2538 102 -2532
rect 96 -2544 102 -2538
rect 96 -2550 102 -2544
rect 96 -2556 102 -2550
rect 96 -2562 102 -2556
rect 96 -2568 102 -2562
rect 96 -2574 102 -2568
rect 96 -2580 102 -2574
rect 96 -2586 102 -2580
rect 96 -2592 102 -2586
rect 96 -2598 102 -2592
rect 96 -2604 102 -2598
rect 96 -2610 102 -2604
rect 96 -2616 102 -2610
rect 96 -2622 102 -2616
rect 96 -2628 102 -2622
rect 96 -2634 102 -2628
rect 96 -2640 102 -2634
rect 96 -2646 102 -2640
rect 96 -2652 102 -2646
rect 96 -2658 102 -2652
rect 96 -2664 102 -2658
rect 96 -2670 102 -2664
rect 96 -2676 102 -2670
rect 96 -2682 102 -2676
rect 96 -2688 102 -2682
rect 96 -2694 102 -2688
rect 96 -2700 102 -2694
rect 96 -2706 102 -2700
rect 96 -2712 102 -2706
rect 96 -2718 102 -2712
rect 96 -2724 102 -2718
rect 96 -2730 102 -2724
rect 96 -2736 102 -2730
rect 96 -2742 102 -2736
rect 96 -2748 102 -2742
rect 96 -2754 102 -2748
rect 96 -2760 102 -2754
rect 96 -2766 102 -2760
rect 96 -2772 102 -2766
rect 96 -2778 102 -2772
rect 96 -2784 102 -2778
rect 96 -2790 102 -2784
rect 102 -1824 108 -1818
rect 102 -1830 108 -1824
rect 102 -1836 108 -1830
rect 102 -1842 108 -1836
rect 102 -1848 108 -1842
rect 102 -1854 108 -1848
rect 102 -1860 108 -1854
rect 102 -1866 108 -1860
rect 102 -1872 108 -1866
rect 102 -1878 108 -1872
rect 102 -1884 108 -1878
rect 102 -1890 108 -1884
rect 102 -1896 108 -1890
rect 102 -1902 108 -1896
rect 102 -1908 108 -1902
rect 102 -1914 108 -1908
rect 102 -1920 108 -1914
rect 102 -1926 108 -1920
rect 102 -1932 108 -1926
rect 102 -1938 108 -1932
rect 102 -1944 108 -1938
rect 102 -1950 108 -1944
rect 102 -1956 108 -1950
rect 102 -1962 108 -1956
rect 102 -1968 108 -1962
rect 102 -1974 108 -1968
rect 102 -1980 108 -1974
rect 102 -1986 108 -1980
rect 102 -1992 108 -1986
rect 102 -1998 108 -1992
rect 102 -2004 108 -1998
rect 102 -2010 108 -2004
rect 102 -2016 108 -2010
rect 102 -2022 108 -2016
rect 102 -2028 108 -2022
rect 102 -2034 108 -2028
rect 102 -2040 108 -2034
rect 102 -2046 108 -2040
rect 102 -2052 108 -2046
rect 102 -2058 108 -2052
rect 102 -2064 108 -2058
rect 102 -2070 108 -2064
rect 102 -2076 108 -2070
rect 102 -2082 108 -2076
rect 102 -2088 108 -2082
rect 102 -2094 108 -2088
rect 102 -2100 108 -2094
rect 102 -2106 108 -2100
rect 102 -2112 108 -2106
rect 102 -2118 108 -2112
rect 102 -2124 108 -2118
rect 102 -2130 108 -2124
rect 102 -2136 108 -2130
rect 102 -2142 108 -2136
rect 102 -2148 108 -2142
rect 102 -2154 108 -2148
rect 102 -2160 108 -2154
rect 102 -2166 108 -2160
rect 102 -2172 108 -2166
rect 102 -2178 108 -2172
rect 102 -2184 108 -2178
rect 102 -2190 108 -2184
rect 102 -2196 108 -2190
rect 102 -2202 108 -2196
rect 102 -2208 108 -2202
rect 102 -2214 108 -2208
rect 102 -2220 108 -2214
rect 102 -2226 108 -2220
rect 102 -2232 108 -2226
rect 102 -2238 108 -2232
rect 102 -2244 108 -2238
rect 102 -2250 108 -2244
rect 102 -2256 108 -2250
rect 102 -2262 108 -2256
rect 102 -2268 108 -2262
rect 102 -2274 108 -2268
rect 102 -2280 108 -2274
rect 102 -2286 108 -2280
rect 102 -2292 108 -2286
rect 102 -2298 108 -2292
rect 102 -2304 108 -2298
rect 102 -2310 108 -2304
rect 102 -2316 108 -2310
rect 102 -2322 108 -2316
rect 102 -2328 108 -2322
rect 102 -2334 108 -2328
rect 102 -2340 108 -2334
rect 102 -2346 108 -2340
rect 102 -2352 108 -2346
rect 102 -2358 108 -2352
rect 102 -2364 108 -2358
rect 102 -2370 108 -2364
rect 102 -2376 108 -2370
rect 102 -2382 108 -2376
rect 102 -2388 108 -2382
rect 102 -2394 108 -2388
rect 102 -2400 108 -2394
rect 102 -2406 108 -2400
rect 102 -2412 108 -2406
rect 102 -2418 108 -2412
rect 102 -2424 108 -2418
rect 102 -2430 108 -2424
rect 102 -2436 108 -2430
rect 102 -2442 108 -2436
rect 102 -2448 108 -2442
rect 102 -2454 108 -2448
rect 102 -2460 108 -2454
rect 102 -2466 108 -2460
rect 102 -2472 108 -2466
rect 102 -2478 108 -2472
rect 102 -2484 108 -2478
rect 102 -2490 108 -2484
rect 102 -2496 108 -2490
rect 102 -2502 108 -2496
rect 102 -2508 108 -2502
rect 102 -2514 108 -2508
rect 102 -2520 108 -2514
rect 102 -2526 108 -2520
rect 102 -2532 108 -2526
rect 102 -2538 108 -2532
rect 102 -2544 108 -2538
rect 102 -2550 108 -2544
rect 102 -2556 108 -2550
rect 102 -2562 108 -2556
rect 102 -2568 108 -2562
rect 102 -2574 108 -2568
rect 102 -2580 108 -2574
rect 102 -2586 108 -2580
rect 102 -2592 108 -2586
rect 102 -2598 108 -2592
rect 102 -2604 108 -2598
rect 102 -2610 108 -2604
rect 102 -2616 108 -2610
rect 102 -2622 108 -2616
rect 102 -2628 108 -2622
rect 102 -2634 108 -2628
rect 102 -2640 108 -2634
rect 102 -2646 108 -2640
rect 102 -2652 108 -2646
rect 102 -2658 108 -2652
rect 102 -2664 108 -2658
rect 102 -2670 108 -2664
rect 102 -2676 108 -2670
rect 102 -2682 108 -2676
rect 102 -2688 108 -2682
rect 102 -2694 108 -2688
rect 102 -2700 108 -2694
rect 102 -2706 108 -2700
rect 102 -2712 108 -2706
rect 102 -2718 108 -2712
rect 102 -2724 108 -2718
rect 102 -2730 108 -2724
rect 102 -2736 108 -2730
rect 102 -2742 108 -2736
rect 102 -2748 108 -2742
rect 102 -2754 108 -2748
rect 102 -2760 108 -2754
rect 102 -2766 108 -2760
rect 102 -2772 108 -2766
rect 102 -2778 108 -2772
rect 102 -2784 108 -2778
rect 102 -2790 108 -2784
rect 102 -2796 108 -2790
rect 102 -2802 108 -2796
rect 108 -1812 114 -1806
rect 108 -1818 114 -1812
rect 108 -1824 114 -1818
rect 108 -1830 114 -1824
rect 108 -1836 114 -1830
rect 108 -1842 114 -1836
rect 108 -1848 114 -1842
rect 108 -1854 114 -1848
rect 108 -1860 114 -1854
rect 108 -1866 114 -1860
rect 108 -1872 114 -1866
rect 108 -1878 114 -1872
rect 108 -1884 114 -1878
rect 108 -1890 114 -1884
rect 108 -1896 114 -1890
rect 108 -1902 114 -1896
rect 108 -1908 114 -1902
rect 108 -1914 114 -1908
rect 108 -1920 114 -1914
rect 108 -1926 114 -1920
rect 108 -1932 114 -1926
rect 108 -1938 114 -1932
rect 108 -1944 114 -1938
rect 108 -1950 114 -1944
rect 108 -1956 114 -1950
rect 108 -1962 114 -1956
rect 108 -1968 114 -1962
rect 108 -1974 114 -1968
rect 108 -1980 114 -1974
rect 108 -1986 114 -1980
rect 108 -1992 114 -1986
rect 108 -1998 114 -1992
rect 108 -2004 114 -1998
rect 108 -2010 114 -2004
rect 108 -2016 114 -2010
rect 108 -2022 114 -2016
rect 108 -2028 114 -2022
rect 108 -2034 114 -2028
rect 108 -2040 114 -2034
rect 108 -2046 114 -2040
rect 108 -2052 114 -2046
rect 108 -2058 114 -2052
rect 108 -2064 114 -2058
rect 108 -2070 114 -2064
rect 108 -2076 114 -2070
rect 108 -2082 114 -2076
rect 108 -2088 114 -2082
rect 108 -2094 114 -2088
rect 108 -2100 114 -2094
rect 108 -2106 114 -2100
rect 108 -2112 114 -2106
rect 108 -2118 114 -2112
rect 108 -2124 114 -2118
rect 108 -2130 114 -2124
rect 108 -2136 114 -2130
rect 108 -2142 114 -2136
rect 108 -2148 114 -2142
rect 108 -2154 114 -2148
rect 108 -2160 114 -2154
rect 108 -2166 114 -2160
rect 108 -2172 114 -2166
rect 108 -2178 114 -2172
rect 108 -2184 114 -2178
rect 108 -2190 114 -2184
rect 108 -2196 114 -2190
rect 108 -2202 114 -2196
rect 108 -2208 114 -2202
rect 108 -2214 114 -2208
rect 108 -2220 114 -2214
rect 108 -2226 114 -2220
rect 108 -2232 114 -2226
rect 108 -2238 114 -2232
rect 108 -2244 114 -2238
rect 108 -2250 114 -2244
rect 108 -2256 114 -2250
rect 108 -2262 114 -2256
rect 108 -2268 114 -2262
rect 108 -2274 114 -2268
rect 108 -2280 114 -2274
rect 108 -2286 114 -2280
rect 108 -2292 114 -2286
rect 108 -2298 114 -2292
rect 108 -2304 114 -2298
rect 108 -2310 114 -2304
rect 108 -2316 114 -2310
rect 108 -2322 114 -2316
rect 108 -2328 114 -2322
rect 108 -2334 114 -2328
rect 108 -2340 114 -2334
rect 108 -2346 114 -2340
rect 108 -2352 114 -2346
rect 108 -2358 114 -2352
rect 108 -2364 114 -2358
rect 108 -2370 114 -2364
rect 108 -2376 114 -2370
rect 108 -2382 114 -2376
rect 108 -2388 114 -2382
rect 108 -2394 114 -2388
rect 108 -2400 114 -2394
rect 108 -2406 114 -2400
rect 108 -2412 114 -2406
rect 108 -2418 114 -2412
rect 108 -2424 114 -2418
rect 108 -2430 114 -2424
rect 108 -2436 114 -2430
rect 108 -2442 114 -2436
rect 108 -2448 114 -2442
rect 108 -2454 114 -2448
rect 108 -2460 114 -2454
rect 108 -2466 114 -2460
rect 108 -2472 114 -2466
rect 108 -2478 114 -2472
rect 108 -2484 114 -2478
rect 108 -2490 114 -2484
rect 108 -2496 114 -2490
rect 108 -2502 114 -2496
rect 108 -2508 114 -2502
rect 108 -2514 114 -2508
rect 108 -2520 114 -2514
rect 108 -2526 114 -2520
rect 108 -2532 114 -2526
rect 108 -2538 114 -2532
rect 108 -2544 114 -2538
rect 108 -2550 114 -2544
rect 108 -2556 114 -2550
rect 108 -2562 114 -2556
rect 108 -2568 114 -2562
rect 108 -2574 114 -2568
rect 108 -2580 114 -2574
rect 108 -2586 114 -2580
rect 108 -2592 114 -2586
rect 108 -2598 114 -2592
rect 108 -2604 114 -2598
rect 108 -2610 114 -2604
rect 108 -2616 114 -2610
rect 108 -2622 114 -2616
rect 108 -2628 114 -2622
rect 108 -2634 114 -2628
rect 108 -2640 114 -2634
rect 108 -2646 114 -2640
rect 108 -2652 114 -2646
rect 108 -2658 114 -2652
rect 108 -2664 114 -2658
rect 108 -2670 114 -2664
rect 108 -2676 114 -2670
rect 108 -2682 114 -2676
rect 108 -2688 114 -2682
rect 108 -2694 114 -2688
rect 108 -2700 114 -2694
rect 108 -2706 114 -2700
rect 108 -2712 114 -2706
rect 108 -2718 114 -2712
rect 108 -2724 114 -2718
rect 108 -2730 114 -2724
rect 108 -2736 114 -2730
rect 108 -2742 114 -2736
rect 108 -2748 114 -2742
rect 108 -2754 114 -2748
rect 108 -2760 114 -2754
rect 108 -2766 114 -2760
rect 108 -2772 114 -2766
rect 108 -2778 114 -2772
rect 108 -2784 114 -2778
rect 108 -2790 114 -2784
rect 108 -2796 114 -2790
rect 108 -2802 114 -2796
rect 108 -2808 114 -2802
rect 108 -2814 114 -2808
rect 114 -1800 120 -1794
rect 114 -1806 120 -1800
rect 114 -1812 120 -1806
rect 114 -1818 120 -1812
rect 114 -1824 120 -1818
rect 114 -1830 120 -1824
rect 114 -1836 120 -1830
rect 114 -1842 120 -1836
rect 114 -1848 120 -1842
rect 114 -1854 120 -1848
rect 114 -1860 120 -1854
rect 114 -1866 120 -1860
rect 114 -1872 120 -1866
rect 114 -1878 120 -1872
rect 114 -1884 120 -1878
rect 114 -1890 120 -1884
rect 114 -1896 120 -1890
rect 114 -1902 120 -1896
rect 114 -1908 120 -1902
rect 114 -1914 120 -1908
rect 114 -1920 120 -1914
rect 114 -1926 120 -1920
rect 114 -1932 120 -1926
rect 114 -1938 120 -1932
rect 114 -1944 120 -1938
rect 114 -1950 120 -1944
rect 114 -1956 120 -1950
rect 114 -1962 120 -1956
rect 114 -1968 120 -1962
rect 114 -1974 120 -1968
rect 114 -1980 120 -1974
rect 114 -1986 120 -1980
rect 114 -1992 120 -1986
rect 114 -1998 120 -1992
rect 114 -2004 120 -1998
rect 114 -2010 120 -2004
rect 114 -2016 120 -2010
rect 114 -2022 120 -2016
rect 114 -2028 120 -2022
rect 114 -2034 120 -2028
rect 114 -2040 120 -2034
rect 114 -2046 120 -2040
rect 114 -2052 120 -2046
rect 114 -2058 120 -2052
rect 114 -2064 120 -2058
rect 114 -2070 120 -2064
rect 114 -2076 120 -2070
rect 114 -2082 120 -2076
rect 114 -2088 120 -2082
rect 114 -2094 120 -2088
rect 114 -2100 120 -2094
rect 114 -2106 120 -2100
rect 114 -2112 120 -2106
rect 114 -2118 120 -2112
rect 114 -2124 120 -2118
rect 114 -2130 120 -2124
rect 114 -2136 120 -2130
rect 114 -2142 120 -2136
rect 114 -2148 120 -2142
rect 114 -2154 120 -2148
rect 114 -2160 120 -2154
rect 114 -2166 120 -2160
rect 114 -2172 120 -2166
rect 114 -2178 120 -2172
rect 114 -2184 120 -2178
rect 114 -2190 120 -2184
rect 114 -2196 120 -2190
rect 114 -2202 120 -2196
rect 114 -2208 120 -2202
rect 114 -2214 120 -2208
rect 114 -2220 120 -2214
rect 114 -2226 120 -2220
rect 114 -2232 120 -2226
rect 114 -2238 120 -2232
rect 114 -2244 120 -2238
rect 114 -2250 120 -2244
rect 114 -2256 120 -2250
rect 114 -2262 120 -2256
rect 114 -2268 120 -2262
rect 114 -2274 120 -2268
rect 114 -2280 120 -2274
rect 114 -2286 120 -2280
rect 114 -2292 120 -2286
rect 114 -2298 120 -2292
rect 114 -2304 120 -2298
rect 114 -2310 120 -2304
rect 114 -2316 120 -2310
rect 114 -2322 120 -2316
rect 114 -2328 120 -2322
rect 114 -2334 120 -2328
rect 114 -2340 120 -2334
rect 114 -2346 120 -2340
rect 114 -2352 120 -2346
rect 114 -2358 120 -2352
rect 114 -2364 120 -2358
rect 114 -2370 120 -2364
rect 114 -2376 120 -2370
rect 114 -2382 120 -2376
rect 114 -2388 120 -2382
rect 114 -2394 120 -2388
rect 114 -2400 120 -2394
rect 114 -2406 120 -2400
rect 114 -2412 120 -2406
rect 114 -2418 120 -2412
rect 114 -2424 120 -2418
rect 114 -2430 120 -2424
rect 114 -2436 120 -2430
rect 114 -2442 120 -2436
rect 114 -2448 120 -2442
rect 114 -2454 120 -2448
rect 114 -2460 120 -2454
rect 114 -2466 120 -2460
rect 114 -2472 120 -2466
rect 114 -2478 120 -2472
rect 114 -2484 120 -2478
rect 114 -2490 120 -2484
rect 114 -2496 120 -2490
rect 114 -2502 120 -2496
rect 114 -2508 120 -2502
rect 114 -2514 120 -2508
rect 114 -2520 120 -2514
rect 114 -2526 120 -2520
rect 114 -2532 120 -2526
rect 114 -2538 120 -2532
rect 114 -2544 120 -2538
rect 114 -2550 120 -2544
rect 114 -2556 120 -2550
rect 114 -2562 120 -2556
rect 114 -2568 120 -2562
rect 114 -2574 120 -2568
rect 114 -2580 120 -2574
rect 114 -2586 120 -2580
rect 114 -2592 120 -2586
rect 114 -2598 120 -2592
rect 114 -2604 120 -2598
rect 114 -2610 120 -2604
rect 114 -2616 120 -2610
rect 114 -2622 120 -2616
rect 114 -2628 120 -2622
rect 114 -2634 120 -2628
rect 114 -2640 120 -2634
rect 114 -2646 120 -2640
rect 114 -2652 120 -2646
rect 114 -2658 120 -2652
rect 114 -2664 120 -2658
rect 114 -2670 120 -2664
rect 114 -2676 120 -2670
rect 114 -2682 120 -2676
rect 114 -2688 120 -2682
rect 114 -2694 120 -2688
rect 114 -2700 120 -2694
rect 114 -2706 120 -2700
rect 114 -2712 120 -2706
rect 114 -2718 120 -2712
rect 114 -2724 120 -2718
rect 114 -2730 120 -2724
rect 114 -2736 120 -2730
rect 114 -2742 120 -2736
rect 114 -2748 120 -2742
rect 114 -2754 120 -2748
rect 114 -2760 120 -2754
rect 114 -2766 120 -2760
rect 114 -2772 120 -2766
rect 114 -2778 120 -2772
rect 114 -2784 120 -2778
rect 114 -2790 120 -2784
rect 114 -2796 120 -2790
rect 114 -2802 120 -2796
rect 114 -2808 120 -2802
rect 114 -2814 120 -2808
rect 114 -2820 120 -2814
rect 114 -2826 120 -2820
rect 120 -1788 126 -1782
rect 120 -1794 126 -1788
rect 120 -1800 126 -1794
rect 120 -1806 126 -1800
rect 120 -1812 126 -1806
rect 120 -1818 126 -1812
rect 120 -1824 126 -1818
rect 120 -1830 126 -1824
rect 120 -1836 126 -1830
rect 120 -1842 126 -1836
rect 120 -1848 126 -1842
rect 120 -1854 126 -1848
rect 120 -1860 126 -1854
rect 120 -1866 126 -1860
rect 120 -1872 126 -1866
rect 120 -1878 126 -1872
rect 120 -1884 126 -1878
rect 120 -1890 126 -1884
rect 120 -1896 126 -1890
rect 120 -1902 126 -1896
rect 120 -1908 126 -1902
rect 120 -1914 126 -1908
rect 120 -1920 126 -1914
rect 120 -1926 126 -1920
rect 120 -1932 126 -1926
rect 120 -1938 126 -1932
rect 120 -1944 126 -1938
rect 120 -1950 126 -1944
rect 120 -1956 126 -1950
rect 120 -1962 126 -1956
rect 120 -1968 126 -1962
rect 120 -1974 126 -1968
rect 120 -1980 126 -1974
rect 120 -1986 126 -1980
rect 120 -1992 126 -1986
rect 120 -1998 126 -1992
rect 120 -2004 126 -1998
rect 120 -2010 126 -2004
rect 120 -2016 126 -2010
rect 120 -2022 126 -2016
rect 120 -2028 126 -2022
rect 120 -2034 126 -2028
rect 120 -2040 126 -2034
rect 120 -2046 126 -2040
rect 120 -2052 126 -2046
rect 120 -2058 126 -2052
rect 120 -2064 126 -2058
rect 120 -2070 126 -2064
rect 120 -2076 126 -2070
rect 120 -2082 126 -2076
rect 120 -2088 126 -2082
rect 120 -2094 126 -2088
rect 120 -2100 126 -2094
rect 120 -2106 126 -2100
rect 120 -2112 126 -2106
rect 120 -2118 126 -2112
rect 120 -2124 126 -2118
rect 120 -2130 126 -2124
rect 120 -2136 126 -2130
rect 120 -2142 126 -2136
rect 120 -2148 126 -2142
rect 120 -2154 126 -2148
rect 120 -2160 126 -2154
rect 120 -2166 126 -2160
rect 120 -2172 126 -2166
rect 120 -2178 126 -2172
rect 120 -2184 126 -2178
rect 120 -2190 126 -2184
rect 120 -2196 126 -2190
rect 120 -2202 126 -2196
rect 120 -2208 126 -2202
rect 120 -2214 126 -2208
rect 120 -2220 126 -2214
rect 120 -2226 126 -2220
rect 120 -2232 126 -2226
rect 120 -2238 126 -2232
rect 120 -2244 126 -2238
rect 120 -2250 126 -2244
rect 120 -2256 126 -2250
rect 120 -2262 126 -2256
rect 120 -2268 126 -2262
rect 120 -2274 126 -2268
rect 120 -2280 126 -2274
rect 120 -2286 126 -2280
rect 120 -2292 126 -2286
rect 120 -2298 126 -2292
rect 120 -2304 126 -2298
rect 120 -2310 126 -2304
rect 120 -2316 126 -2310
rect 120 -2322 126 -2316
rect 120 -2328 126 -2322
rect 120 -2334 126 -2328
rect 120 -2340 126 -2334
rect 120 -2346 126 -2340
rect 120 -2352 126 -2346
rect 120 -2358 126 -2352
rect 120 -2364 126 -2358
rect 120 -2370 126 -2364
rect 120 -2376 126 -2370
rect 120 -2382 126 -2376
rect 120 -2388 126 -2382
rect 120 -2394 126 -2388
rect 120 -2400 126 -2394
rect 120 -2406 126 -2400
rect 120 -2412 126 -2406
rect 120 -2418 126 -2412
rect 120 -2424 126 -2418
rect 120 -2430 126 -2424
rect 120 -2436 126 -2430
rect 120 -2442 126 -2436
rect 120 -2448 126 -2442
rect 120 -2454 126 -2448
rect 120 -2460 126 -2454
rect 120 -2466 126 -2460
rect 120 -2472 126 -2466
rect 120 -2478 126 -2472
rect 120 -2484 126 -2478
rect 120 -2490 126 -2484
rect 120 -2496 126 -2490
rect 120 -2502 126 -2496
rect 120 -2508 126 -2502
rect 120 -2514 126 -2508
rect 120 -2520 126 -2514
rect 120 -2526 126 -2520
rect 120 -2532 126 -2526
rect 120 -2538 126 -2532
rect 120 -2544 126 -2538
rect 120 -2550 126 -2544
rect 120 -2556 126 -2550
rect 120 -2562 126 -2556
rect 120 -2568 126 -2562
rect 120 -2574 126 -2568
rect 120 -2580 126 -2574
rect 120 -2586 126 -2580
rect 120 -2592 126 -2586
rect 120 -2598 126 -2592
rect 120 -2604 126 -2598
rect 120 -2610 126 -2604
rect 120 -2616 126 -2610
rect 120 -2622 126 -2616
rect 120 -2628 126 -2622
rect 120 -2634 126 -2628
rect 120 -2640 126 -2634
rect 120 -2646 126 -2640
rect 120 -2652 126 -2646
rect 120 -2658 126 -2652
rect 120 -2664 126 -2658
rect 120 -2670 126 -2664
rect 120 -2676 126 -2670
rect 120 -2682 126 -2676
rect 120 -2688 126 -2682
rect 120 -2694 126 -2688
rect 120 -2700 126 -2694
rect 120 -2706 126 -2700
rect 120 -2712 126 -2706
rect 120 -2718 126 -2712
rect 120 -2724 126 -2718
rect 120 -2730 126 -2724
rect 120 -2736 126 -2730
rect 120 -2742 126 -2736
rect 120 -2748 126 -2742
rect 120 -2754 126 -2748
rect 120 -2760 126 -2754
rect 120 -2766 126 -2760
rect 120 -2772 126 -2766
rect 120 -2778 126 -2772
rect 120 -2784 126 -2778
rect 120 -2790 126 -2784
rect 120 -2796 126 -2790
rect 120 -2802 126 -2796
rect 120 -2808 126 -2802
rect 120 -2814 126 -2808
rect 120 -2820 126 -2814
rect 120 -2826 126 -2820
rect 120 -2832 126 -2826
rect 120 -2838 126 -2832
rect 126 -1776 132 -1770
rect 126 -1782 132 -1776
rect 126 -1788 132 -1782
rect 126 -1794 132 -1788
rect 126 -1800 132 -1794
rect 126 -1806 132 -1800
rect 126 -1812 132 -1806
rect 126 -1818 132 -1812
rect 126 -1824 132 -1818
rect 126 -1830 132 -1824
rect 126 -1836 132 -1830
rect 126 -1842 132 -1836
rect 126 -1848 132 -1842
rect 126 -1854 132 -1848
rect 126 -1860 132 -1854
rect 126 -1866 132 -1860
rect 126 -1872 132 -1866
rect 126 -1878 132 -1872
rect 126 -1884 132 -1878
rect 126 -1890 132 -1884
rect 126 -1896 132 -1890
rect 126 -1902 132 -1896
rect 126 -1908 132 -1902
rect 126 -1914 132 -1908
rect 126 -1920 132 -1914
rect 126 -1926 132 -1920
rect 126 -1932 132 -1926
rect 126 -1938 132 -1932
rect 126 -1944 132 -1938
rect 126 -1950 132 -1944
rect 126 -1956 132 -1950
rect 126 -1962 132 -1956
rect 126 -1968 132 -1962
rect 126 -1974 132 -1968
rect 126 -1980 132 -1974
rect 126 -1986 132 -1980
rect 126 -1992 132 -1986
rect 126 -1998 132 -1992
rect 126 -2004 132 -1998
rect 126 -2010 132 -2004
rect 126 -2016 132 -2010
rect 126 -2022 132 -2016
rect 126 -2028 132 -2022
rect 126 -2034 132 -2028
rect 126 -2040 132 -2034
rect 126 -2046 132 -2040
rect 126 -2052 132 -2046
rect 126 -2058 132 -2052
rect 126 -2064 132 -2058
rect 126 -2070 132 -2064
rect 126 -2076 132 -2070
rect 126 -2082 132 -2076
rect 126 -2088 132 -2082
rect 126 -2094 132 -2088
rect 126 -2100 132 -2094
rect 126 -2106 132 -2100
rect 126 -2112 132 -2106
rect 126 -2118 132 -2112
rect 126 -2124 132 -2118
rect 126 -2130 132 -2124
rect 126 -2136 132 -2130
rect 126 -2142 132 -2136
rect 126 -2148 132 -2142
rect 126 -2154 132 -2148
rect 126 -2160 132 -2154
rect 126 -2166 132 -2160
rect 126 -2172 132 -2166
rect 126 -2178 132 -2172
rect 126 -2184 132 -2178
rect 126 -2190 132 -2184
rect 126 -2196 132 -2190
rect 126 -2202 132 -2196
rect 126 -2208 132 -2202
rect 126 -2214 132 -2208
rect 126 -2220 132 -2214
rect 126 -2226 132 -2220
rect 126 -2232 132 -2226
rect 126 -2238 132 -2232
rect 126 -2244 132 -2238
rect 126 -2250 132 -2244
rect 126 -2256 132 -2250
rect 126 -2262 132 -2256
rect 126 -2268 132 -2262
rect 126 -2274 132 -2268
rect 126 -2280 132 -2274
rect 126 -2286 132 -2280
rect 126 -2292 132 -2286
rect 126 -2298 132 -2292
rect 126 -2304 132 -2298
rect 126 -2310 132 -2304
rect 126 -2316 132 -2310
rect 126 -2322 132 -2316
rect 126 -2328 132 -2322
rect 126 -2334 132 -2328
rect 126 -2340 132 -2334
rect 126 -2346 132 -2340
rect 126 -2352 132 -2346
rect 126 -2358 132 -2352
rect 126 -2364 132 -2358
rect 126 -2370 132 -2364
rect 126 -2376 132 -2370
rect 126 -2382 132 -2376
rect 126 -2388 132 -2382
rect 126 -2394 132 -2388
rect 126 -2400 132 -2394
rect 126 -2406 132 -2400
rect 126 -2412 132 -2406
rect 126 -2418 132 -2412
rect 126 -2424 132 -2418
rect 126 -2430 132 -2424
rect 126 -2436 132 -2430
rect 126 -2442 132 -2436
rect 126 -2448 132 -2442
rect 126 -2454 132 -2448
rect 126 -2460 132 -2454
rect 126 -2466 132 -2460
rect 126 -2472 132 -2466
rect 126 -2478 132 -2472
rect 126 -2484 132 -2478
rect 126 -2490 132 -2484
rect 126 -2496 132 -2490
rect 126 -2502 132 -2496
rect 126 -2508 132 -2502
rect 126 -2514 132 -2508
rect 126 -2520 132 -2514
rect 126 -2526 132 -2520
rect 126 -2532 132 -2526
rect 126 -2538 132 -2532
rect 126 -2544 132 -2538
rect 126 -2550 132 -2544
rect 126 -2556 132 -2550
rect 126 -2562 132 -2556
rect 126 -2568 132 -2562
rect 126 -2574 132 -2568
rect 126 -2580 132 -2574
rect 126 -2586 132 -2580
rect 126 -2592 132 -2586
rect 126 -2598 132 -2592
rect 126 -2604 132 -2598
rect 126 -2610 132 -2604
rect 126 -2616 132 -2610
rect 126 -2622 132 -2616
rect 126 -2628 132 -2622
rect 126 -2634 132 -2628
rect 126 -2640 132 -2634
rect 126 -2646 132 -2640
rect 126 -2652 132 -2646
rect 126 -2658 132 -2652
rect 126 -2664 132 -2658
rect 126 -2670 132 -2664
rect 126 -2676 132 -2670
rect 126 -2682 132 -2676
rect 126 -2688 132 -2682
rect 126 -2694 132 -2688
rect 126 -2700 132 -2694
rect 126 -2706 132 -2700
rect 126 -2712 132 -2706
rect 126 -2718 132 -2712
rect 126 -2724 132 -2718
rect 126 -2730 132 -2724
rect 126 -2736 132 -2730
rect 126 -2742 132 -2736
rect 126 -2748 132 -2742
rect 126 -2754 132 -2748
rect 126 -2760 132 -2754
rect 126 -2766 132 -2760
rect 126 -2772 132 -2766
rect 126 -2778 132 -2772
rect 126 -2784 132 -2778
rect 126 -2790 132 -2784
rect 126 -2796 132 -2790
rect 126 -2802 132 -2796
rect 126 -2808 132 -2802
rect 126 -2814 132 -2808
rect 126 -2820 132 -2814
rect 126 -2826 132 -2820
rect 126 -2832 132 -2826
rect 126 -2838 132 -2832
rect 126 -2844 132 -2838
rect 126 -2850 132 -2844
rect 132 -1764 138 -1758
rect 132 -1770 138 -1764
rect 132 -1776 138 -1770
rect 132 -1782 138 -1776
rect 132 -1788 138 -1782
rect 132 -1794 138 -1788
rect 132 -1800 138 -1794
rect 132 -1806 138 -1800
rect 132 -1812 138 -1806
rect 132 -1818 138 -1812
rect 132 -1824 138 -1818
rect 132 -1830 138 -1824
rect 132 -1836 138 -1830
rect 132 -1842 138 -1836
rect 132 -1848 138 -1842
rect 132 -1854 138 -1848
rect 132 -1860 138 -1854
rect 132 -1866 138 -1860
rect 132 -1872 138 -1866
rect 132 -1878 138 -1872
rect 132 -1884 138 -1878
rect 132 -1890 138 -1884
rect 132 -1896 138 -1890
rect 132 -1902 138 -1896
rect 132 -1908 138 -1902
rect 132 -1914 138 -1908
rect 132 -1920 138 -1914
rect 132 -1926 138 -1920
rect 132 -1932 138 -1926
rect 132 -1938 138 -1932
rect 132 -1944 138 -1938
rect 132 -1950 138 -1944
rect 132 -1956 138 -1950
rect 132 -1962 138 -1956
rect 132 -1968 138 -1962
rect 132 -1974 138 -1968
rect 132 -1980 138 -1974
rect 132 -1986 138 -1980
rect 132 -1992 138 -1986
rect 132 -1998 138 -1992
rect 132 -2004 138 -1998
rect 132 -2010 138 -2004
rect 132 -2016 138 -2010
rect 132 -2022 138 -2016
rect 132 -2028 138 -2022
rect 132 -2034 138 -2028
rect 132 -2040 138 -2034
rect 132 -2046 138 -2040
rect 132 -2052 138 -2046
rect 132 -2058 138 -2052
rect 132 -2064 138 -2058
rect 132 -2070 138 -2064
rect 132 -2076 138 -2070
rect 132 -2082 138 -2076
rect 132 -2088 138 -2082
rect 132 -2094 138 -2088
rect 132 -2100 138 -2094
rect 132 -2106 138 -2100
rect 132 -2112 138 -2106
rect 132 -2118 138 -2112
rect 132 -2124 138 -2118
rect 132 -2130 138 -2124
rect 132 -2136 138 -2130
rect 132 -2142 138 -2136
rect 132 -2148 138 -2142
rect 132 -2154 138 -2148
rect 132 -2160 138 -2154
rect 132 -2166 138 -2160
rect 132 -2172 138 -2166
rect 132 -2178 138 -2172
rect 132 -2184 138 -2178
rect 132 -2190 138 -2184
rect 132 -2196 138 -2190
rect 132 -2202 138 -2196
rect 132 -2208 138 -2202
rect 132 -2214 138 -2208
rect 132 -2220 138 -2214
rect 132 -2226 138 -2220
rect 132 -2232 138 -2226
rect 132 -2238 138 -2232
rect 132 -2244 138 -2238
rect 132 -2250 138 -2244
rect 132 -2256 138 -2250
rect 132 -2262 138 -2256
rect 132 -2268 138 -2262
rect 132 -2274 138 -2268
rect 132 -2280 138 -2274
rect 132 -2286 138 -2280
rect 132 -2292 138 -2286
rect 132 -2298 138 -2292
rect 132 -2304 138 -2298
rect 132 -2310 138 -2304
rect 132 -2316 138 -2310
rect 132 -2322 138 -2316
rect 132 -2328 138 -2322
rect 132 -2334 138 -2328
rect 132 -2340 138 -2334
rect 132 -2346 138 -2340
rect 132 -2352 138 -2346
rect 132 -2358 138 -2352
rect 132 -2364 138 -2358
rect 132 -2370 138 -2364
rect 132 -2376 138 -2370
rect 132 -2382 138 -2376
rect 132 -2388 138 -2382
rect 132 -2394 138 -2388
rect 132 -2400 138 -2394
rect 132 -2406 138 -2400
rect 132 -2412 138 -2406
rect 132 -2418 138 -2412
rect 132 -2424 138 -2418
rect 132 -2430 138 -2424
rect 132 -2436 138 -2430
rect 132 -2442 138 -2436
rect 132 -2448 138 -2442
rect 132 -2454 138 -2448
rect 132 -2460 138 -2454
rect 132 -2466 138 -2460
rect 132 -2472 138 -2466
rect 132 -2478 138 -2472
rect 132 -2484 138 -2478
rect 132 -2490 138 -2484
rect 132 -2496 138 -2490
rect 132 -2502 138 -2496
rect 132 -2508 138 -2502
rect 132 -2514 138 -2508
rect 132 -2520 138 -2514
rect 132 -2526 138 -2520
rect 132 -2532 138 -2526
rect 132 -2538 138 -2532
rect 132 -2544 138 -2538
rect 132 -2550 138 -2544
rect 132 -2556 138 -2550
rect 132 -2562 138 -2556
rect 132 -2568 138 -2562
rect 132 -2574 138 -2568
rect 132 -2580 138 -2574
rect 132 -2586 138 -2580
rect 132 -2592 138 -2586
rect 132 -2598 138 -2592
rect 132 -2604 138 -2598
rect 132 -2610 138 -2604
rect 132 -2616 138 -2610
rect 132 -2622 138 -2616
rect 132 -2628 138 -2622
rect 132 -2634 138 -2628
rect 132 -2640 138 -2634
rect 132 -2646 138 -2640
rect 132 -2652 138 -2646
rect 132 -2658 138 -2652
rect 132 -2664 138 -2658
rect 132 -2670 138 -2664
rect 132 -2676 138 -2670
rect 132 -2682 138 -2676
rect 132 -2688 138 -2682
rect 132 -2694 138 -2688
rect 132 -2700 138 -2694
rect 132 -2706 138 -2700
rect 132 -2712 138 -2706
rect 132 -2718 138 -2712
rect 132 -2724 138 -2718
rect 132 -2730 138 -2724
rect 132 -2736 138 -2730
rect 132 -2742 138 -2736
rect 132 -2748 138 -2742
rect 132 -2754 138 -2748
rect 132 -2760 138 -2754
rect 132 -2766 138 -2760
rect 132 -2772 138 -2766
rect 132 -2778 138 -2772
rect 132 -2784 138 -2778
rect 132 -2790 138 -2784
rect 132 -2796 138 -2790
rect 132 -2802 138 -2796
rect 132 -2808 138 -2802
rect 132 -2814 138 -2808
rect 132 -2820 138 -2814
rect 132 -2826 138 -2820
rect 132 -2832 138 -2826
rect 132 -2838 138 -2832
rect 132 -2844 138 -2838
rect 132 -2850 138 -2844
rect 132 -2856 138 -2850
rect 132 -2862 138 -2856
rect 138 -1752 144 -1746
rect 138 -1758 144 -1752
rect 138 -1764 144 -1758
rect 138 -1770 144 -1764
rect 138 -1776 144 -1770
rect 138 -1782 144 -1776
rect 138 -1788 144 -1782
rect 138 -1794 144 -1788
rect 138 -1800 144 -1794
rect 138 -1806 144 -1800
rect 138 -1812 144 -1806
rect 138 -1818 144 -1812
rect 138 -1824 144 -1818
rect 138 -1830 144 -1824
rect 138 -1836 144 -1830
rect 138 -1842 144 -1836
rect 138 -1848 144 -1842
rect 138 -1854 144 -1848
rect 138 -1860 144 -1854
rect 138 -1866 144 -1860
rect 138 -1872 144 -1866
rect 138 -1878 144 -1872
rect 138 -1884 144 -1878
rect 138 -1890 144 -1884
rect 138 -1896 144 -1890
rect 138 -1902 144 -1896
rect 138 -1908 144 -1902
rect 138 -1914 144 -1908
rect 138 -1920 144 -1914
rect 138 -1926 144 -1920
rect 138 -1932 144 -1926
rect 138 -1938 144 -1932
rect 138 -1944 144 -1938
rect 138 -1950 144 -1944
rect 138 -1956 144 -1950
rect 138 -1962 144 -1956
rect 138 -1968 144 -1962
rect 138 -1974 144 -1968
rect 138 -1980 144 -1974
rect 138 -1986 144 -1980
rect 138 -1992 144 -1986
rect 138 -1998 144 -1992
rect 138 -2004 144 -1998
rect 138 -2010 144 -2004
rect 138 -2016 144 -2010
rect 138 -2022 144 -2016
rect 138 -2028 144 -2022
rect 138 -2034 144 -2028
rect 138 -2040 144 -2034
rect 138 -2046 144 -2040
rect 138 -2052 144 -2046
rect 138 -2058 144 -2052
rect 138 -2064 144 -2058
rect 138 -2070 144 -2064
rect 138 -2076 144 -2070
rect 138 -2082 144 -2076
rect 138 -2088 144 -2082
rect 138 -2094 144 -2088
rect 138 -2100 144 -2094
rect 138 -2106 144 -2100
rect 138 -2112 144 -2106
rect 138 -2118 144 -2112
rect 138 -2124 144 -2118
rect 138 -2130 144 -2124
rect 138 -2136 144 -2130
rect 138 -2142 144 -2136
rect 138 -2148 144 -2142
rect 138 -2154 144 -2148
rect 138 -2160 144 -2154
rect 138 -2166 144 -2160
rect 138 -2172 144 -2166
rect 138 -2178 144 -2172
rect 138 -2184 144 -2178
rect 138 -2190 144 -2184
rect 138 -2196 144 -2190
rect 138 -2202 144 -2196
rect 138 -2208 144 -2202
rect 138 -2214 144 -2208
rect 138 -2220 144 -2214
rect 138 -2226 144 -2220
rect 138 -2232 144 -2226
rect 138 -2238 144 -2232
rect 138 -2244 144 -2238
rect 138 -2250 144 -2244
rect 138 -2256 144 -2250
rect 138 -2262 144 -2256
rect 138 -2268 144 -2262
rect 138 -2274 144 -2268
rect 138 -2280 144 -2274
rect 138 -2286 144 -2280
rect 138 -2292 144 -2286
rect 138 -2298 144 -2292
rect 138 -2304 144 -2298
rect 138 -2310 144 -2304
rect 138 -2316 144 -2310
rect 138 -2322 144 -2316
rect 138 -2328 144 -2322
rect 138 -2334 144 -2328
rect 138 -2340 144 -2334
rect 138 -2346 144 -2340
rect 138 -2352 144 -2346
rect 138 -2358 144 -2352
rect 138 -2364 144 -2358
rect 138 -2370 144 -2364
rect 138 -2376 144 -2370
rect 138 -2382 144 -2376
rect 138 -2388 144 -2382
rect 138 -2394 144 -2388
rect 138 -2400 144 -2394
rect 138 -2406 144 -2400
rect 138 -2412 144 -2406
rect 138 -2418 144 -2412
rect 138 -2424 144 -2418
rect 138 -2430 144 -2424
rect 138 -2436 144 -2430
rect 138 -2442 144 -2436
rect 138 -2448 144 -2442
rect 138 -2454 144 -2448
rect 138 -2460 144 -2454
rect 138 -2466 144 -2460
rect 138 -2472 144 -2466
rect 138 -2478 144 -2472
rect 138 -2484 144 -2478
rect 138 -2490 144 -2484
rect 138 -2496 144 -2490
rect 138 -2502 144 -2496
rect 138 -2508 144 -2502
rect 138 -2514 144 -2508
rect 138 -2520 144 -2514
rect 138 -2526 144 -2520
rect 138 -2532 144 -2526
rect 138 -2538 144 -2532
rect 138 -2544 144 -2538
rect 138 -2550 144 -2544
rect 138 -2556 144 -2550
rect 138 -2562 144 -2556
rect 138 -2568 144 -2562
rect 138 -2574 144 -2568
rect 138 -2580 144 -2574
rect 138 -2586 144 -2580
rect 138 -2592 144 -2586
rect 138 -2598 144 -2592
rect 138 -2604 144 -2598
rect 138 -2610 144 -2604
rect 138 -2616 144 -2610
rect 138 -2622 144 -2616
rect 138 -2628 144 -2622
rect 138 -2634 144 -2628
rect 138 -2640 144 -2634
rect 138 -2646 144 -2640
rect 138 -2652 144 -2646
rect 138 -2658 144 -2652
rect 138 -2664 144 -2658
rect 138 -2670 144 -2664
rect 138 -2676 144 -2670
rect 138 -2682 144 -2676
rect 138 -2688 144 -2682
rect 138 -2694 144 -2688
rect 138 -2700 144 -2694
rect 138 -2706 144 -2700
rect 138 -2712 144 -2706
rect 138 -2718 144 -2712
rect 138 -2724 144 -2718
rect 138 -2730 144 -2724
rect 138 -2736 144 -2730
rect 138 -2742 144 -2736
rect 138 -2748 144 -2742
rect 138 -2754 144 -2748
rect 138 -2760 144 -2754
rect 138 -2766 144 -2760
rect 138 -2772 144 -2766
rect 138 -2778 144 -2772
rect 138 -2784 144 -2778
rect 138 -2790 144 -2784
rect 138 -2796 144 -2790
rect 138 -2802 144 -2796
rect 138 -2808 144 -2802
rect 138 -2814 144 -2808
rect 138 -2820 144 -2814
rect 138 -2826 144 -2820
rect 138 -2832 144 -2826
rect 138 -2838 144 -2832
rect 138 -2844 144 -2838
rect 138 -2850 144 -2844
rect 138 -2856 144 -2850
rect 138 -2862 144 -2856
rect 138 -2868 144 -2862
rect 138 -2874 144 -2868
rect 144 -1740 150 -1734
rect 144 -1746 150 -1740
rect 144 -1752 150 -1746
rect 144 -1758 150 -1752
rect 144 -1764 150 -1758
rect 144 -1770 150 -1764
rect 144 -1776 150 -1770
rect 144 -1782 150 -1776
rect 144 -1788 150 -1782
rect 144 -1794 150 -1788
rect 144 -1800 150 -1794
rect 144 -1806 150 -1800
rect 144 -1812 150 -1806
rect 144 -1818 150 -1812
rect 144 -1824 150 -1818
rect 144 -1830 150 -1824
rect 144 -1836 150 -1830
rect 144 -1842 150 -1836
rect 144 -1848 150 -1842
rect 144 -1854 150 -1848
rect 144 -1860 150 -1854
rect 144 -1866 150 -1860
rect 144 -1872 150 -1866
rect 144 -1878 150 -1872
rect 144 -1884 150 -1878
rect 144 -1890 150 -1884
rect 144 -1896 150 -1890
rect 144 -1902 150 -1896
rect 144 -1908 150 -1902
rect 144 -1914 150 -1908
rect 144 -1920 150 -1914
rect 144 -1926 150 -1920
rect 144 -1932 150 -1926
rect 144 -1938 150 -1932
rect 144 -1944 150 -1938
rect 144 -1950 150 -1944
rect 144 -1956 150 -1950
rect 144 -1962 150 -1956
rect 144 -1968 150 -1962
rect 144 -1974 150 -1968
rect 144 -1980 150 -1974
rect 144 -1986 150 -1980
rect 144 -1992 150 -1986
rect 144 -1998 150 -1992
rect 144 -2004 150 -1998
rect 144 -2010 150 -2004
rect 144 -2016 150 -2010
rect 144 -2022 150 -2016
rect 144 -2028 150 -2022
rect 144 -2034 150 -2028
rect 144 -2040 150 -2034
rect 144 -2046 150 -2040
rect 144 -2052 150 -2046
rect 144 -2058 150 -2052
rect 144 -2064 150 -2058
rect 144 -2070 150 -2064
rect 144 -2076 150 -2070
rect 144 -2082 150 -2076
rect 144 -2088 150 -2082
rect 144 -2094 150 -2088
rect 144 -2100 150 -2094
rect 144 -2106 150 -2100
rect 144 -2112 150 -2106
rect 144 -2118 150 -2112
rect 144 -2124 150 -2118
rect 144 -2130 150 -2124
rect 144 -2136 150 -2130
rect 144 -2142 150 -2136
rect 144 -2148 150 -2142
rect 144 -2154 150 -2148
rect 144 -2160 150 -2154
rect 144 -2166 150 -2160
rect 144 -2172 150 -2166
rect 144 -2178 150 -2172
rect 144 -2184 150 -2178
rect 144 -2190 150 -2184
rect 144 -2196 150 -2190
rect 144 -2202 150 -2196
rect 144 -2208 150 -2202
rect 144 -2214 150 -2208
rect 144 -2220 150 -2214
rect 144 -2226 150 -2220
rect 144 -2232 150 -2226
rect 144 -2238 150 -2232
rect 144 -2244 150 -2238
rect 144 -2250 150 -2244
rect 144 -2256 150 -2250
rect 144 -2262 150 -2256
rect 144 -2268 150 -2262
rect 144 -2274 150 -2268
rect 144 -2280 150 -2274
rect 144 -2286 150 -2280
rect 144 -2292 150 -2286
rect 144 -2298 150 -2292
rect 144 -2304 150 -2298
rect 144 -2310 150 -2304
rect 144 -2316 150 -2310
rect 144 -2322 150 -2316
rect 144 -2328 150 -2322
rect 144 -2334 150 -2328
rect 144 -2340 150 -2334
rect 144 -2346 150 -2340
rect 144 -2352 150 -2346
rect 144 -2358 150 -2352
rect 144 -2364 150 -2358
rect 144 -2370 150 -2364
rect 144 -2376 150 -2370
rect 144 -2382 150 -2376
rect 144 -2388 150 -2382
rect 144 -2394 150 -2388
rect 144 -2400 150 -2394
rect 144 -2406 150 -2400
rect 144 -2412 150 -2406
rect 144 -2418 150 -2412
rect 144 -2424 150 -2418
rect 144 -2430 150 -2424
rect 144 -2436 150 -2430
rect 144 -2442 150 -2436
rect 144 -2448 150 -2442
rect 144 -2454 150 -2448
rect 144 -2460 150 -2454
rect 144 -2466 150 -2460
rect 144 -2472 150 -2466
rect 144 -2478 150 -2472
rect 144 -2484 150 -2478
rect 144 -2490 150 -2484
rect 144 -2496 150 -2490
rect 144 -2502 150 -2496
rect 144 -2508 150 -2502
rect 144 -2514 150 -2508
rect 144 -2520 150 -2514
rect 144 -2526 150 -2520
rect 144 -2532 150 -2526
rect 144 -2538 150 -2532
rect 144 -2544 150 -2538
rect 144 -2550 150 -2544
rect 144 -2556 150 -2550
rect 144 -2562 150 -2556
rect 144 -2568 150 -2562
rect 144 -2574 150 -2568
rect 144 -2580 150 -2574
rect 144 -2586 150 -2580
rect 144 -2592 150 -2586
rect 144 -2598 150 -2592
rect 144 -2604 150 -2598
rect 144 -2610 150 -2604
rect 144 -2616 150 -2610
rect 144 -2622 150 -2616
rect 144 -2628 150 -2622
rect 144 -2634 150 -2628
rect 144 -2640 150 -2634
rect 144 -2646 150 -2640
rect 144 -2652 150 -2646
rect 144 -2658 150 -2652
rect 144 -2664 150 -2658
rect 144 -2670 150 -2664
rect 144 -2676 150 -2670
rect 144 -2682 150 -2676
rect 144 -2688 150 -2682
rect 144 -2694 150 -2688
rect 144 -2700 150 -2694
rect 144 -2706 150 -2700
rect 144 -2712 150 -2706
rect 144 -2718 150 -2712
rect 144 -2724 150 -2718
rect 144 -2730 150 -2724
rect 144 -2736 150 -2730
rect 144 -2742 150 -2736
rect 144 -2748 150 -2742
rect 144 -2754 150 -2748
rect 144 -2760 150 -2754
rect 144 -2766 150 -2760
rect 144 -2772 150 -2766
rect 144 -2778 150 -2772
rect 144 -2784 150 -2778
rect 144 -2790 150 -2784
rect 144 -2796 150 -2790
rect 144 -2802 150 -2796
rect 144 -2808 150 -2802
rect 144 -2814 150 -2808
rect 144 -2820 150 -2814
rect 144 -2826 150 -2820
rect 144 -2832 150 -2826
rect 144 -2838 150 -2832
rect 144 -2844 150 -2838
rect 144 -2850 150 -2844
rect 144 -2856 150 -2850
rect 144 -2862 150 -2856
rect 144 -2868 150 -2862
rect 144 -2874 150 -2868
rect 144 -2880 150 -2874
rect 144 -2886 150 -2880
rect 150 -1728 156 -1722
rect 150 -1734 156 -1728
rect 150 -1740 156 -1734
rect 150 -1746 156 -1740
rect 150 -1752 156 -1746
rect 150 -1758 156 -1752
rect 150 -1764 156 -1758
rect 150 -1770 156 -1764
rect 150 -1776 156 -1770
rect 150 -1782 156 -1776
rect 150 -1788 156 -1782
rect 150 -1794 156 -1788
rect 150 -1800 156 -1794
rect 150 -1806 156 -1800
rect 150 -1812 156 -1806
rect 150 -1818 156 -1812
rect 150 -1824 156 -1818
rect 150 -1830 156 -1824
rect 150 -1836 156 -1830
rect 150 -1842 156 -1836
rect 150 -1848 156 -1842
rect 150 -1854 156 -1848
rect 150 -1860 156 -1854
rect 150 -1866 156 -1860
rect 150 -1872 156 -1866
rect 150 -1878 156 -1872
rect 150 -1884 156 -1878
rect 150 -1890 156 -1884
rect 150 -1896 156 -1890
rect 150 -1902 156 -1896
rect 150 -1908 156 -1902
rect 150 -1914 156 -1908
rect 150 -1920 156 -1914
rect 150 -1926 156 -1920
rect 150 -1932 156 -1926
rect 150 -1938 156 -1932
rect 150 -1944 156 -1938
rect 150 -1950 156 -1944
rect 150 -1956 156 -1950
rect 150 -1962 156 -1956
rect 150 -1968 156 -1962
rect 150 -1974 156 -1968
rect 150 -1980 156 -1974
rect 150 -1986 156 -1980
rect 150 -1992 156 -1986
rect 150 -1998 156 -1992
rect 150 -2004 156 -1998
rect 150 -2010 156 -2004
rect 150 -2016 156 -2010
rect 150 -2022 156 -2016
rect 150 -2028 156 -2022
rect 150 -2034 156 -2028
rect 150 -2040 156 -2034
rect 150 -2046 156 -2040
rect 150 -2052 156 -2046
rect 150 -2058 156 -2052
rect 150 -2064 156 -2058
rect 150 -2070 156 -2064
rect 150 -2076 156 -2070
rect 150 -2082 156 -2076
rect 150 -2088 156 -2082
rect 150 -2094 156 -2088
rect 150 -2100 156 -2094
rect 150 -2106 156 -2100
rect 150 -2112 156 -2106
rect 150 -2118 156 -2112
rect 150 -2124 156 -2118
rect 150 -2130 156 -2124
rect 150 -2136 156 -2130
rect 150 -2142 156 -2136
rect 150 -2148 156 -2142
rect 150 -2154 156 -2148
rect 150 -2160 156 -2154
rect 150 -2166 156 -2160
rect 150 -2172 156 -2166
rect 150 -2178 156 -2172
rect 150 -2184 156 -2178
rect 150 -2190 156 -2184
rect 150 -2196 156 -2190
rect 150 -2202 156 -2196
rect 150 -2208 156 -2202
rect 150 -2214 156 -2208
rect 150 -2220 156 -2214
rect 150 -2226 156 -2220
rect 150 -2232 156 -2226
rect 150 -2238 156 -2232
rect 150 -2244 156 -2238
rect 150 -2250 156 -2244
rect 150 -2256 156 -2250
rect 150 -2262 156 -2256
rect 150 -2268 156 -2262
rect 150 -2274 156 -2268
rect 150 -2280 156 -2274
rect 150 -2286 156 -2280
rect 150 -2292 156 -2286
rect 150 -2298 156 -2292
rect 150 -2304 156 -2298
rect 150 -2310 156 -2304
rect 150 -2316 156 -2310
rect 150 -2322 156 -2316
rect 150 -2328 156 -2322
rect 150 -2334 156 -2328
rect 150 -2340 156 -2334
rect 150 -2346 156 -2340
rect 150 -2352 156 -2346
rect 150 -2358 156 -2352
rect 150 -2364 156 -2358
rect 150 -2370 156 -2364
rect 150 -2376 156 -2370
rect 150 -2382 156 -2376
rect 150 -2388 156 -2382
rect 150 -2394 156 -2388
rect 150 -2400 156 -2394
rect 150 -2406 156 -2400
rect 150 -2412 156 -2406
rect 150 -2418 156 -2412
rect 150 -2424 156 -2418
rect 150 -2430 156 -2424
rect 150 -2436 156 -2430
rect 150 -2442 156 -2436
rect 150 -2448 156 -2442
rect 150 -2454 156 -2448
rect 150 -2460 156 -2454
rect 150 -2466 156 -2460
rect 150 -2472 156 -2466
rect 150 -2478 156 -2472
rect 150 -2484 156 -2478
rect 150 -2490 156 -2484
rect 150 -2496 156 -2490
rect 150 -2502 156 -2496
rect 150 -2508 156 -2502
rect 150 -2514 156 -2508
rect 150 -2520 156 -2514
rect 150 -2526 156 -2520
rect 150 -2532 156 -2526
rect 150 -2538 156 -2532
rect 150 -2544 156 -2538
rect 150 -2550 156 -2544
rect 150 -2556 156 -2550
rect 150 -2562 156 -2556
rect 150 -2568 156 -2562
rect 150 -2574 156 -2568
rect 150 -2580 156 -2574
rect 150 -2586 156 -2580
rect 150 -2592 156 -2586
rect 150 -2598 156 -2592
rect 150 -2604 156 -2598
rect 150 -2610 156 -2604
rect 150 -2616 156 -2610
rect 150 -2622 156 -2616
rect 150 -2628 156 -2622
rect 150 -2634 156 -2628
rect 150 -2640 156 -2634
rect 150 -2646 156 -2640
rect 150 -2652 156 -2646
rect 150 -2658 156 -2652
rect 150 -2664 156 -2658
rect 150 -2670 156 -2664
rect 150 -2676 156 -2670
rect 150 -2682 156 -2676
rect 150 -2688 156 -2682
rect 150 -2694 156 -2688
rect 150 -2700 156 -2694
rect 150 -2706 156 -2700
rect 150 -2712 156 -2706
rect 150 -2718 156 -2712
rect 150 -2724 156 -2718
rect 150 -2730 156 -2724
rect 150 -2736 156 -2730
rect 150 -2742 156 -2736
rect 150 -2748 156 -2742
rect 150 -2754 156 -2748
rect 150 -2760 156 -2754
rect 150 -2766 156 -2760
rect 150 -2772 156 -2766
rect 150 -2778 156 -2772
rect 150 -2784 156 -2778
rect 150 -2790 156 -2784
rect 150 -2796 156 -2790
rect 150 -2802 156 -2796
rect 150 -2808 156 -2802
rect 150 -2814 156 -2808
rect 150 -2820 156 -2814
rect 150 -2826 156 -2820
rect 150 -2832 156 -2826
rect 150 -2838 156 -2832
rect 150 -2844 156 -2838
rect 150 -2850 156 -2844
rect 150 -2856 156 -2850
rect 150 -2862 156 -2856
rect 150 -2868 156 -2862
rect 150 -2874 156 -2868
rect 150 -2880 156 -2874
rect 150 -2886 156 -2880
rect 150 -2892 156 -2886
rect 150 -2898 156 -2892
rect 156 -1716 162 -1710
rect 156 -1722 162 -1716
rect 156 -1728 162 -1722
rect 156 -1734 162 -1728
rect 156 -1740 162 -1734
rect 156 -1746 162 -1740
rect 156 -1752 162 -1746
rect 156 -1758 162 -1752
rect 156 -1764 162 -1758
rect 156 -1770 162 -1764
rect 156 -1776 162 -1770
rect 156 -1782 162 -1776
rect 156 -1788 162 -1782
rect 156 -1794 162 -1788
rect 156 -1800 162 -1794
rect 156 -1806 162 -1800
rect 156 -1812 162 -1806
rect 156 -1818 162 -1812
rect 156 -1824 162 -1818
rect 156 -1830 162 -1824
rect 156 -1836 162 -1830
rect 156 -1842 162 -1836
rect 156 -1848 162 -1842
rect 156 -1854 162 -1848
rect 156 -1860 162 -1854
rect 156 -1866 162 -1860
rect 156 -1872 162 -1866
rect 156 -1878 162 -1872
rect 156 -1884 162 -1878
rect 156 -1890 162 -1884
rect 156 -1896 162 -1890
rect 156 -1902 162 -1896
rect 156 -1908 162 -1902
rect 156 -1914 162 -1908
rect 156 -1920 162 -1914
rect 156 -1926 162 -1920
rect 156 -1932 162 -1926
rect 156 -1938 162 -1932
rect 156 -1944 162 -1938
rect 156 -1950 162 -1944
rect 156 -1956 162 -1950
rect 156 -1962 162 -1956
rect 156 -1968 162 -1962
rect 156 -1974 162 -1968
rect 156 -1980 162 -1974
rect 156 -1986 162 -1980
rect 156 -1992 162 -1986
rect 156 -1998 162 -1992
rect 156 -2004 162 -1998
rect 156 -2010 162 -2004
rect 156 -2016 162 -2010
rect 156 -2022 162 -2016
rect 156 -2028 162 -2022
rect 156 -2034 162 -2028
rect 156 -2040 162 -2034
rect 156 -2046 162 -2040
rect 156 -2052 162 -2046
rect 156 -2058 162 -2052
rect 156 -2064 162 -2058
rect 156 -2070 162 -2064
rect 156 -2076 162 -2070
rect 156 -2082 162 -2076
rect 156 -2088 162 -2082
rect 156 -2094 162 -2088
rect 156 -2100 162 -2094
rect 156 -2106 162 -2100
rect 156 -2112 162 -2106
rect 156 -2118 162 -2112
rect 156 -2124 162 -2118
rect 156 -2130 162 -2124
rect 156 -2136 162 -2130
rect 156 -2142 162 -2136
rect 156 -2148 162 -2142
rect 156 -2154 162 -2148
rect 156 -2160 162 -2154
rect 156 -2166 162 -2160
rect 156 -2172 162 -2166
rect 156 -2178 162 -2172
rect 156 -2184 162 -2178
rect 156 -2190 162 -2184
rect 156 -2196 162 -2190
rect 156 -2202 162 -2196
rect 156 -2208 162 -2202
rect 156 -2214 162 -2208
rect 156 -2220 162 -2214
rect 156 -2226 162 -2220
rect 156 -2232 162 -2226
rect 156 -2238 162 -2232
rect 156 -2244 162 -2238
rect 156 -2250 162 -2244
rect 156 -2256 162 -2250
rect 156 -2262 162 -2256
rect 156 -2268 162 -2262
rect 156 -2274 162 -2268
rect 156 -2280 162 -2274
rect 156 -2286 162 -2280
rect 156 -2292 162 -2286
rect 156 -2298 162 -2292
rect 156 -2304 162 -2298
rect 156 -2310 162 -2304
rect 156 -2316 162 -2310
rect 156 -2322 162 -2316
rect 156 -2328 162 -2322
rect 156 -2334 162 -2328
rect 156 -2340 162 -2334
rect 156 -2346 162 -2340
rect 156 -2352 162 -2346
rect 156 -2358 162 -2352
rect 156 -2364 162 -2358
rect 156 -2370 162 -2364
rect 156 -2376 162 -2370
rect 156 -2382 162 -2376
rect 156 -2388 162 -2382
rect 156 -2394 162 -2388
rect 156 -2400 162 -2394
rect 156 -2406 162 -2400
rect 156 -2412 162 -2406
rect 156 -2418 162 -2412
rect 156 -2424 162 -2418
rect 156 -2430 162 -2424
rect 156 -2436 162 -2430
rect 156 -2442 162 -2436
rect 156 -2448 162 -2442
rect 156 -2454 162 -2448
rect 156 -2460 162 -2454
rect 156 -2466 162 -2460
rect 156 -2472 162 -2466
rect 156 -2478 162 -2472
rect 156 -2484 162 -2478
rect 156 -2490 162 -2484
rect 156 -2496 162 -2490
rect 156 -2502 162 -2496
rect 156 -2508 162 -2502
rect 156 -2514 162 -2508
rect 156 -2520 162 -2514
rect 156 -2526 162 -2520
rect 156 -2532 162 -2526
rect 156 -2538 162 -2532
rect 156 -2544 162 -2538
rect 156 -2550 162 -2544
rect 156 -2556 162 -2550
rect 156 -2562 162 -2556
rect 156 -2568 162 -2562
rect 156 -2574 162 -2568
rect 156 -2580 162 -2574
rect 156 -2586 162 -2580
rect 156 -2592 162 -2586
rect 156 -2598 162 -2592
rect 156 -2604 162 -2598
rect 156 -2610 162 -2604
rect 156 -2616 162 -2610
rect 156 -2622 162 -2616
rect 156 -2628 162 -2622
rect 156 -2634 162 -2628
rect 156 -2640 162 -2634
rect 156 -2646 162 -2640
rect 156 -2652 162 -2646
rect 156 -2658 162 -2652
rect 156 -2664 162 -2658
rect 156 -2670 162 -2664
rect 156 -2676 162 -2670
rect 156 -2682 162 -2676
rect 156 -2688 162 -2682
rect 156 -2694 162 -2688
rect 156 -2700 162 -2694
rect 156 -2706 162 -2700
rect 156 -2712 162 -2706
rect 156 -2718 162 -2712
rect 156 -2724 162 -2718
rect 156 -2730 162 -2724
rect 156 -2736 162 -2730
rect 156 -2742 162 -2736
rect 156 -2748 162 -2742
rect 156 -2754 162 -2748
rect 156 -2760 162 -2754
rect 156 -2766 162 -2760
rect 156 -2772 162 -2766
rect 156 -2778 162 -2772
rect 156 -2784 162 -2778
rect 156 -2790 162 -2784
rect 156 -2796 162 -2790
rect 156 -2802 162 -2796
rect 156 -2808 162 -2802
rect 156 -2814 162 -2808
rect 156 -2820 162 -2814
rect 156 -2826 162 -2820
rect 156 -2832 162 -2826
rect 156 -2838 162 -2832
rect 156 -2844 162 -2838
rect 156 -2850 162 -2844
rect 156 -2856 162 -2850
rect 156 -2862 162 -2856
rect 156 -2868 162 -2862
rect 156 -2874 162 -2868
rect 156 -2880 162 -2874
rect 156 -2886 162 -2880
rect 156 -2892 162 -2886
rect 156 -2898 162 -2892
rect 156 -2904 162 -2898
rect 156 -2910 162 -2904
rect 162 -1710 168 -1704
rect 162 -1716 168 -1710
rect 162 -1722 168 -1716
rect 162 -1728 168 -1722
rect 162 -1734 168 -1728
rect 162 -1740 168 -1734
rect 162 -1746 168 -1740
rect 162 -1752 168 -1746
rect 162 -1758 168 -1752
rect 162 -1764 168 -1758
rect 162 -1770 168 -1764
rect 162 -1776 168 -1770
rect 162 -1782 168 -1776
rect 162 -1788 168 -1782
rect 162 -1794 168 -1788
rect 162 -1800 168 -1794
rect 162 -1806 168 -1800
rect 162 -1812 168 -1806
rect 162 -1818 168 -1812
rect 162 -1824 168 -1818
rect 162 -1830 168 -1824
rect 162 -1836 168 -1830
rect 162 -1842 168 -1836
rect 162 -1848 168 -1842
rect 162 -1854 168 -1848
rect 162 -1860 168 -1854
rect 162 -1866 168 -1860
rect 162 -1872 168 -1866
rect 162 -1878 168 -1872
rect 162 -1884 168 -1878
rect 162 -1890 168 -1884
rect 162 -1896 168 -1890
rect 162 -1902 168 -1896
rect 162 -1908 168 -1902
rect 162 -1914 168 -1908
rect 162 -1920 168 -1914
rect 162 -1926 168 -1920
rect 162 -1932 168 -1926
rect 162 -1938 168 -1932
rect 162 -1944 168 -1938
rect 162 -1950 168 -1944
rect 162 -1956 168 -1950
rect 162 -1962 168 -1956
rect 162 -1968 168 -1962
rect 162 -1974 168 -1968
rect 162 -1980 168 -1974
rect 162 -1986 168 -1980
rect 162 -1992 168 -1986
rect 162 -1998 168 -1992
rect 162 -2004 168 -1998
rect 162 -2010 168 -2004
rect 162 -2016 168 -2010
rect 162 -2022 168 -2016
rect 162 -2028 168 -2022
rect 162 -2034 168 -2028
rect 162 -2040 168 -2034
rect 162 -2046 168 -2040
rect 162 -2052 168 -2046
rect 162 -2058 168 -2052
rect 162 -2064 168 -2058
rect 162 -2070 168 -2064
rect 162 -2076 168 -2070
rect 162 -2082 168 -2076
rect 162 -2088 168 -2082
rect 162 -2094 168 -2088
rect 162 -2100 168 -2094
rect 162 -2106 168 -2100
rect 162 -2112 168 -2106
rect 162 -2118 168 -2112
rect 162 -2124 168 -2118
rect 162 -2130 168 -2124
rect 162 -2136 168 -2130
rect 162 -2142 168 -2136
rect 162 -2148 168 -2142
rect 162 -2154 168 -2148
rect 162 -2160 168 -2154
rect 162 -2166 168 -2160
rect 162 -2172 168 -2166
rect 162 -2178 168 -2172
rect 162 -2184 168 -2178
rect 162 -2190 168 -2184
rect 162 -2196 168 -2190
rect 162 -2202 168 -2196
rect 162 -2208 168 -2202
rect 162 -2214 168 -2208
rect 162 -2220 168 -2214
rect 162 -2226 168 -2220
rect 162 -2232 168 -2226
rect 162 -2238 168 -2232
rect 162 -2244 168 -2238
rect 162 -2250 168 -2244
rect 162 -2256 168 -2250
rect 162 -2262 168 -2256
rect 162 -2268 168 -2262
rect 162 -2274 168 -2268
rect 162 -2280 168 -2274
rect 162 -2286 168 -2280
rect 162 -2292 168 -2286
rect 162 -2298 168 -2292
rect 162 -2304 168 -2298
rect 162 -2310 168 -2304
rect 162 -2316 168 -2310
rect 162 -2322 168 -2316
rect 162 -2328 168 -2322
rect 162 -2334 168 -2328
rect 162 -2340 168 -2334
rect 162 -2346 168 -2340
rect 162 -2352 168 -2346
rect 162 -2358 168 -2352
rect 162 -2364 168 -2358
rect 162 -2370 168 -2364
rect 162 -2376 168 -2370
rect 162 -2382 168 -2376
rect 162 -2388 168 -2382
rect 162 -2394 168 -2388
rect 162 -2400 168 -2394
rect 162 -2406 168 -2400
rect 162 -2412 168 -2406
rect 162 -2418 168 -2412
rect 162 -2424 168 -2418
rect 162 -2430 168 -2424
rect 162 -2436 168 -2430
rect 162 -2442 168 -2436
rect 162 -2448 168 -2442
rect 162 -2454 168 -2448
rect 162 -2460 168 -2454
rect 162 -2466 168 -2460
rect 162 -2472 168 -2466
rect 162 -2478 168 -2472
rect 162 -2484 168 -2478
rect 162 -2490 168 -2484
rect 162 -2496 168 -2490
rect 162 -2502 168 -2496
rect 162 -2508 168 -2502
rect 162 -2514 168 -2508
rect 162 -2520 168 -2514
rect 162 -2526 168 -2520
rect 162 -2532 168 -2526
rect 162 -2538 168 -2532
rect 162 -2544 168 -2538
rect 162 -2550 168 -2544
rect 162 -2556 168 -2550
rect 162 -2562 168 -2556
rect 162 -2568 168 -2562
rect 162 -2574 168 -2568
rect 162 -2580 168 -2574
rect 162 -2586 168 -2580
rect 162 -2592 168 -2586
rect 162 -2598 168 -2592
rect 162 -2604 168 -2598
rect 162 -2610 168 -2604
rect 162 -2616 168 -2610
rect 162 -2622 168 -2616
rect 162 -2628 168 -2622
rect 162 -2634 168 -2628
rect 162 -2640 168 -2634
rect 162 -2646 168 -2640
rect 162 -2652 168 -2646
rect 162 -2658 168 -2652
rect 162 -2664 168 -2658
rect 162 -2670 168 -2664
rect 162 -2676 168 -2670
rect 162 -2682 168 -2676
rect 162 -2688 168 -2682
rect 162 -2694 168 -2688
rect 162 -2700 168 -2694
rect 162 -2706 168 -2700
rect 162 -2712 168 -2706
rect 162 -2718 168 -2712
rect 162 -2724 168 -2718
rect 162 -2730 168 -2724
rect 162 -2736 168 -2730
rect 162 -2742 168 -2736
rect 162 -2748 168 -2742
rect 162 -2754 168 -2748
rect 162 -2760 168 -2754
rect 162 -2766 168 -2760
rect 162 -2772 168 -2766
rect 162 -2778 168 -2772
rect 162 -2784 168 -2778
rect 162 -2790 168 -2784
rect 162 -2796 168 -2790
rect 162 -2802 168 -2796
rect 162 -2808 168 -2802
rect 162 -2814 168 -2808
rect 162 -2820 168 -2814
rect 162 -2826 168 -2820
rect 162 -2832 168 -2826
rect 162 -2838 168 -2832
rect 162 -2844 168 -2838
rect 162 -2850 168 -2844
rect 162 -2856 168 -2850
rect 162 -2862 168 -2856
rect 162 -2868 168 -2862
rect 162 -2874 168 -2868
rect 162 -2880 168 -2874
rect 162 -2886 168 -2880
rect 162 -2892 168 -2886
rect 162 -2898 168 -2892
rect 162 -2904 168 -2898
rect 162 -2910 168 -2904
rect 162 -2916 168 -2910
rect 168 -1698 174 -1692
rect 168 -1704 174 -1698
rect 168 -1710 174 -1704
rect 168 -1716 174 -1710
rect 168 -1722 174 -1716
rect 168 -1728 174 -1722
rect 168 -1734 174 -1728
rect 168 -1740 174 -1734
rect 168 -1746 174 -1740
rect 168 -1752 174 -1746
rect 168 -1758 174 -1752
rect 168 -1764 174 -1758
rect 168 -1770 174 -1764
rect 168 -1776 174 -1770
rect 168 -1782 174 -1776
rect 168 -1788 174 -1782
rect 168 -1794 174 -1788
rect 168 -1800 174 -1794
rect 168 -1806 174 -1800
rect 168 -1812 174 -1806
rect 168 -1818 174 -1812
rect 168 -1824 174 -1818
rect 168 -1830 174 -1824
rect 168 -1836 174 -1830
rect 168 -1842 174 -1836
rect 168 -1848 174 -1842
rect 168 -1854 174 -1848
rect 168 -1860 174 -1854
rect 168 -1866 174 -1860
rect 168 -1872 174 -1866
rect 168 -1878 174 -1872
rect 168 -1884 174 -1878
rect 168 -1890 174 -1884
rect 168 -1896 174 -1890
rect 168 -1902 174 -1896
rect 168 -1908 174 -1902
rect 168 -1914 174 -1908
rect 168 -1920 174 -1914
rect 168 -1926 174 -1920
rect 168 -1932 174 -1926
rect 168 -1938 174 -1932
rect 168 -1944 174 -1938
rect 168 -1950 174 -1944
rect 168 -1956 174 -1950
rect 168 -1962 174 -1956
rect 168 -1968 174 -1962
rect 168 -1974 174 -1968
rect 168 -1980 174 -1974
rect 168 -1986 174 -1980
rect 168 -1992 174 -1986
rect 168 -1998 174 -1992
rect 168 -2004 174 -1998
rect 168 -2010 174 -2004
rect 168 -2016 174 -2010
rect 168 -2022 174 -2016
rect 168 -2028 174 -2022
rect 168 -2034 174 -2028
rect 168 -2040 174 -2034
rect 168 -2046 174 -2040
rect 168 -2052 174 -2046
rect 168 -2058 174 -2052
rect 168 -2064 174 -2058
rect 168 -2070 174 -2064
rect 168 -2076 174 -2070
rect 168 -2082 174 -2076
rect 168 -2088 174 -2082
rect 168 -2094 174 -2088
rect 168 -2100 174 -2094
rect 168 -2106 174 -2100
rect 168 -2112 174 -2106
rect 168 -2118 174 -2112
rect 168 -2124 174 -2118
rect 168 -2130 174 -2124
rect 168 -2136 174 -2130
rect 168 -2142 174 -2136
rect 168 -2148 174 -2142
rect 168 -2154 174 -2148
rect 168 -2160 174 -2154
rect 168 -2166 174 -2160
rect 168 -2172 174 -2166
rect 168 -2178 174 -2172
rect 168 -2184 174 -2178
rect 168 -2190 174 -2184
rect 168 -2196 174 -2190
rect 168 -2202 174 -2196
rect 168 -2208 174 -2202
rect 168 -2214 174 -2208
rect 168 -2220 174 -2214
rect 168 -2226 174 -2220
rect 168 -2232 174 -2226
rect 168 -2238 174 -2232
rect 168 -2244 174 -2238
rect 168 -2250 174 -2244
rect 168 -2256 174 -2250
rect 168 -2262 174 -2256
rect 168 -2268 174 -2262
rect 168 -2274 174 -2268
rect 168 -2280 174 -2274
rect 168 -2286 174 -2280
rect 168 -2292 174 -2286
rect 168 -2298 174 -2292
rect 168 -2304 174 -2298
rect 168 -2310 174 -2304
rect 168 -2316 174 -2310
rect 168 -2322 174 -2316
rect 168 -2328 174 -2322
rect 168 -2334 174 -2328
rect 168 -2340 174 -2334
rect 168 -2346 174 -2340
rect 168 -2352 174 -2346
rect 168 -2358 174 -2352
rect 168 -2364 174 -2358
rect 168 -2370 174 -2364
rect 168 -2376 174 -2370
rect 168 -2382 174 -2376
rect 168 -2388 174 -2382
rect 168 -2394 174 -2388
rect 168 -2400 174 -2394
rect 168 -2406 174 -2400
rect 168 -2412 174 -2406
rect 168 -2418 174 -2412
rect 168 -2424 174 -2418
rect 168 -2430 174 -2424
rect 168 -2436 174 -2430
rect 168 -2442 174 -2436
rect 168 -2448 174 -2442
rect 168 -2454 174 -2448
rect 168 -2460 174 -2454
rect 168 -2466 174 -2460
rect 168 -2472 174 -2466
rect 168 -2478 174 -2472
rect 168 -2484 174 -2478
rect 168 -2490 174 -2484
rect 168 -2496 174 -2490
rect 168 -2502 174 -2496
rect 168 -2508 174 -2502
rect 168 -2514 174 -2508
rect 168 -2520 174 -2514
rect 168 -2526 174 -2520
rect 168 -2532 174 -2526
rect 168 -2538 174 -2532
rect 168 -2544 174 -2538
rect 168 -2550 174 -2544
rect 168 -2556 174 -2550
rect 168 -2562 174 -2556
rect 168 -2568 174 -2562
rect 168 -2574 174 -2568
rect 168 -2580 174 -2574
rect 168 -2586 174 -2580
rect 168 -2592 174 -2586
rect 168 -2598 174 -2592
rect 168 -2604 174 -2598
rect 168 -2610 174 -2604
rect 168 -2616 174 -2610
rect 168 -2622 174 -2616
rect 168 -2628 174 -2622
rect 168 -2634 174 -2628
rect 168 -2640 174 -2634
rect 168 -2646 174 -2640
rect 168 -2652 174 -2646
rect 168 -2658 174 -2652
rect 168 -2664 174 -2658
rect 168 -2670 174 -2664
rect 168 -2676 174 -2670
rect 168 -2682 174 -2676
rect 168 -2688 174 -2682
rect 168 -2694 174 -2688
rect 168 -2700 174 -2694
rect 168 -2706 174 -2700
rect 168 -2712 174 -2706
rect 168 -2718 174 -2712
rect 168 -2724 174 -2718
rect 168 -2730 174 -2724
rect 168 -2736 174 -2730
rect 168 -2742 174 -2736
rect 168 -2748 174 -2742
rect 168 -2754 174 -2748
rect 168 -2760 174 -2754
rect 168 -2766 174 -2760
rect 168 -2772 174 -2766
rect 168 -2778 174 -2772
rect 168 -2784 174 -2778
rect 168 -2790 174 -2784
rect 168 -2796 174 -2790
rect 168 -2802 174 -2796
rect 168 -2808 174 -2802
rect 168 -2814 174 -2808
rect 168 -2820 174 -2814
rect 168 -2826 174 -2820
rect 168 -2832 174 -2826
rect 168 -2838 174 -2832
rect 168 -2844 174 -2838
rect 168 -2850 174 -2844
rect 168 -2856 174 -2850
rect 168 -2862 174 -2856
rect 168 -2868 174 -2862
rect 168 -2874 174 -2868
rect 168 -2880 174 -2874
rect 168 -2886 174 -2880
rect 168 -2892 174 -2886
rect 168 -2898 174 -2892
rect 168 -2904 174 -2898
rect 168 -2910 174 -2904
rect 168 -2916 174 -2910
rect 168 -2922 174 -2916
rect 168 -2928 174 -2922
rect 174 -1686 180 -1680
rect 174 -1692 180 -1686
rect 174 -1698 180 -1692
rect 174 -1704 180 -1698
rect 174 -1710 180 -1704
rect 174 -1716 180 -1710
rect 174 -1722 180 -1716
rect 174 -1728 180 -1722
rect 174 -1734 180 -1728
rect 174 -1740 180 -1734
rect 174 -1746 180 -1740
rect 174 -1752 180 -1746
rect 174 -1758 180 -1752
rect 174 -1764 180 -1758
rect 174 -1770 180 -1764
rect 174 -1776 180 -1770
rect 174 -1782 180 -1776
rect 174 -1788 180 -1782
rect 174 -1794 180 -1788
rect 174 -1800 180 -1794
rect 174 -1806 180 -1800
rect 174 -1812 180 -1806
rect 174 -1818 180 -1812
rect 174 -1824 180 -1818
rect 174 -1830 180 -1824
rect 174 -1836 180 -1830
rect 174 -1842 180 -1836
rect 174 -1848 180 -1842
rect 174 -1854 180 -1848
rect 174 -1860 180 -1854
rect 174 -1866 180 -1860
rect 174 -1872 180 -1866
rect 174 -1878 180 -1872
rect 174 -1884 180 -1878
rect 174 -1890 180 -1884
rect 174 -1896 180 -1890
rect 174 -1902 180 -1896
rect 174 -1908 180 -1902
rect 174 -1914 180 -1908
rect 174 -1920 180 -1914
rect 174 -1926 180 -1920
rect 174 -1932 180 -1926
rect 174 -1938 180 -1932
rect 174 -1944 180 -1938
rect 174 -1950 180 -1944
rect 174 -1956 180 -1950
rect 174 -1962 180 -1956
rect 174 -1968 180 -1962
rect 174 -1974 180 -1968
rect 174 -1980 180 -1974
rect 174 -1986 180 -1980
rect 174 -1992 180 -1986
rect 174 -1998 180 -1992
rect 174 -2004 180 -1998
rect 174 -2010 180 -2004
rect 174 -2016 180 -2010
rect 174 -2022 180 -2016
rect 174 -2028 180 -2022
rect 174 -2034 180 -2028
rect 174 -2040 180 -2034
rect 174 -2046 180 -2040
rect 174 -2052 180 -2046
rect 174 -2058 180 -2052
rect 174 -2064 180 -2058
rect 174 -2070 180 -2064
rect 174 -2076 180 -2070
rect 174 -2082 180 -2076
rect 174 -2088 180 -2082
rect 174 -2094 180 -2088
rect 174 -2100 180 -2094
rect 174 -2106 180 -2100
rect 174 -2112 180 -2106
rect 174 -2118 180 -2112
rect 174 -2124 180 -2118
rect 174 -2130 180 -2124
rect 174 -2136 180 -2130
rect 174 -2142 180 -2136
rect 174 -2148 180 -2142
rect 174 -2154 180 -2148
rect 174 -2160 180 -2154
rect 174 -2166 180 -2160
rect 174 -2172 180 -2166
rect 174 -2178 180 -2172
rect 174 -2184 180 -2178
rect 174 -2190 180 -2184
rect 174 -2196 180 -2190
rect 174 -2202 180 -2196
rect 174 -2208 180 -2202
rect 174 -2214 180 -2208
rect 174 -2220 180 -2214
rect 174 -2226 180 -2220
rect 174 -2232 180 -2226
rect 174 -2238 180 -2232
rect 174 -2244 180 -2238
rect 174 -2250 180 -2244
rect 174 -2256 180 -2250
rect 174 -2262 180 -2256
rect 174 -2268 180 -2262
rect 174 -2274 180 -2268
rect 174 -2280 180 -2274
rect 174 -2286 180 -2280
rect 174 -2292 180 -2286
rect 174 -2298 180 -2292
rect 174 -2304 180 -2298
rect 174 -2310 180 -2304
rect 174 -2316 180 -2310
rect 174 -2322 180 -2316
rect 174 -2328 180 -2322
rect 174 -2334 180 -2328
rect 174 -2340 180 -2334
rect 174 -2346 180 -2340
rect 174 -2352 180 -2346
rect 174 -2358 180 -2352
rect 174 -2364 180 -2358
rect 174 -2370 180 -2364
rect 174 -2376 180 -2370
rect 174 -2382 180 -2376
rect 174 -2388 180 -2382
rect 174 -2394 180 -2388
rect 174 -2400 180 -2394
rect 174 -2406 180 -2400
rect 174 -2412 180 -2406
rect 174 -2418 180 -2412
rect 174 -2424 180 -2418
rect 174 -2430 180 -2424
rect 174 -2436 180 -2430
rect 174 -2442 180 -2436
rect 174 -2448 180 -2442
rect 174 -2454 180 -2448
rect 174 -2460 180 -2454
rect 174 -2466 180 -2460
rect 174 -2472 180 -2466
rect 174 -2478 180 -2472
rect 174 -2484 180 -2478
rect 174 -2490 180 -2484
rect 174 -2496 180 -2490
rect 174 -2502 180 -2496
rect 174 -2508 180 -2502
rect 174 -2514 180 -2508
rect 174 -2520 180 -2514
rect 174 -2526 180 -2520
rect 174 -2532 180 -2526
rect 174 -2538 180 -2532
rect 174 -2544 180 -2538
rect 174 -2550 180 -2544
rect 174 -2556 180 -2550
rect 174 -2562 180 -2556
rect 174 -2568 180 -2562
rect 174 -2574 180 -2568
rect 174 -2580 180 -2574
rect 174 -2586 180 -2580
rect 174 -2592 180 -2586
rect 174 -2598 180 -2592
rect 174 -2604 180 -2598
rect 174 -2610 180 -2604
rect 174 -2616 180 -2610
rect 174 -2622 180 -2616
rect 174 -2628 180 -2622
rect 174 -2634 180 -2628
rect 174 -2640 180 -2634
rect 174 -2646 180 -2640
rect 174 -2652 180 -2646
rect 174 -2658 180 -2652
rect 174 -2664 180 -2658
rect 174 -2670 180 -2664
rect 174 -2676 180 -2670
rect 174 -2682 180 -2676
rect 174 -2688 180 -2682
rect 174 -2694 180 -2688
rect 174 -2700 180 -2694
rect 174 -2706 180 -2700
rect 174 -2712 180 -2706
rect 174 -2718 180 -2712
rect 174 -2724 180 -2718
rect 174 -2730 180 -2724
rect 174 -2736 180 -2730
rect 174 -2742 180 -2736
rect 174 -2748 180 -2742
rect 174 -2754 180 -2748
rect 174 -2760 180 -2754
rect 174 -2766 180 -2760
rect 174 -2772 180 -2766
rect 174 -2778 180 -2772
rect 174 -2784 180 -2778
rect 174 -2790 180 -2784
rect 174 -2796 180 -2790
rect 174 -2802 180 -2796
rect 174 -2808 180 -2802
rect 174 -2814 180 -2808
rect 174 -2820 180 -2814
rect 174 -2826 180 -2820
rect 174 -2832 180 -2826
rect 174 -2838 180 -2832
rect 174 -2844 180 -2838
rect 174 -2850 180 -2844
rect 174 -2856 180 -2850
rect 174 -2862 180 -2856
rect 174 -2868 180 -2862
rect 174 -2874 180 -2868
rect 174 -2880 180 -2874
rect 174 -2886 180 -2880
rect 174 -2892 180 -2886
rect 174 -2898 180 -2892
rect 174 -2904 180 -2898
rect 174 -2910 180 -2904
rect 174 -2916 180 -2910
rect 174 -2922 180 -2916
rect 174 -2928 180 -2922
rect 174 -2934 180 -2928
rect 174 -2940 180 -2934
rect 180 -1680 186 -1674
rect 180 -1686 186 -1680
rect 180 -1692 186 -1686
rect 180 -1698 186 -1692
rect 180 -1704 186 -1698
rect 180 -1710 186 -1704
rect 180 -1716 186 -1710
rect 180 -1722 186 -1716
rect 180 -1728 186 -1722
rect 180 -1734 186 -1728
rect 180 -1740 186 -1734
rect 180 -1746 186 -1740
rect 180 -1752 186 -1746
rect 180 -1758 186 -1752
rect 180 -1764 186 -1758
rect 180 -1770 186 -1764
rect 180 -1776 186 -1770
rect 180 -1782 186 -1776
rect 180 -1788 186 -1782
rect 180 -1794 186 -1788
rect 180 -1800 186 -1794
rect 180 -1806 186 -1800
rect 180 -1812 186 -1806
rect 180 -1818 186 -1812
rect 180 -1824 186 -1818
rect 180 -1830 186 -1824
rect 180 -1836 186 -1830
rect 180 -1842 186 -1836
rect 180 -1848 186 -1842
rect 180 -1854 186 -1848
rect 180 -1860 186 -1854
rect 180 -1866 186 -1860
rect 180 -1872 186 -1866
rect 180 -1878 186 -1872
rect 180 -1884 186 -1878
rect 180 -1890 186 -1884
rect 180 -1896 186 -1890
rect 180 -1902 186 -1896
rect 180 -1908 186 -1902
rect 180 -1914 186 -1908
rect 180 -1920 186 -1914
rect 180 -1926 186 -1920
rect 180 -1932 186 -1926
rect 180 -1938 186 -1932
rect 180 -1944 186 -1938
rect 180 -1950 186 -1944
rect 180 -1956 186 -1950
rect 180 -1962 186 -1956
rect 180 -1968 186 -1962
rect 180 -1974 186 -1968
rect 180 -1980 186 -1974
rect 180 -1986 186 -1980
rect 180 -1992 186 -1986
rect 180 -1998 186 -1992
rect 180 -2004 186 -1998
rect 180 -2010 186 -2004
rect 180 -2016 186 -2010
rect 180 -2022 186 -2016
rect 180 -2028 186 -2022
rect 180 -2034 186 -2028
rect 180 -2040 186 -2034
rect 180 -2046 186 -2040
rect 180 -2052 186 -2046
rect 180 -2058 186 -2052
rect 180 -2064 186 -2058
rect 180 -2070 186 -2064
rect 180 -2076 186 -2070
rect 180 -2082 186 -2076
rect 180 -2088 186 -2082
rect 180 -2094 186 -2088
rect 180 -2100 186 -2094
rect 180 -2106 186 -2100
rect 180 -2112 186 -2106
rect 180 -2118 186 -2112
rect 180 -2124 186 -2118
rect 180 -2130 186 -2124
rect 180 -2136 186 -2130
rect 180 -2142 186 -2136
rect 180 -2148 186 -2142
rect 180 -2154 186 -2148
rect 180 -2160 186 -2154
rect 180 -2166 186 -2160
rect 180 -2172 186 -2166
rect 180 -2178 186 -2172
rect 180 -2184 186 -2178
rect 180 -2190 186 -2184
rect 180 -2196 186 -2190
rect 180 -2202 186 -2196
rect 180 -2208 186 -2202
rect 180 -2214 186 -2208
rect 180 -2220 186 -2214
rect 180 -2226 186 -2220
rect 180 -2232 186 -2226
rect 180 -2238 186 -2232
rect 180 -2244 186 -2238
rect 180 -2250 186 -2244
rect 180 -2256 186 -2250
rect 180 -2262 186 -2256
rect 180 -2268 186 -2262
rect 180 -2274 186 -2268
rect 180 -2280 186 -2274
rect 180 -2286 186 -2280
rect 180 -2292 186 -2286
rect 180 -2298 186 -2292
rect 180 -2304 186 -2298
rect 180 -2310 186 -2304
rect 180 -2316 186 -2310
rect 180 -2322 186 -2316
rect 180 -2328 186 -2322
rect 180 -2334 186 -2328
rect 180 -2340 186 -2334
rect 180 -2346 186 -2340
rect 180 -2352 186 -2346
rect 180 -2358 186 -2352
rect 180 -2364 186 -2358
rect 180 -2370 186 -2364
rect 180 -2376 186 -2370
rect 180 -2382 186 -2376
rect 180 -2388 186 -2382
rect 180 -2394 186 -2388
rect 180 -2400 186 -2394
rect 180 -2406 186 -2400
rect 180 -2412 186 -2406
rect 180 -2418 186 -2412
rect 180 -2424 186 -2418
rect 180 -2430 186 -2424
rect 180 -2436 186 -2430
rect 180 -2442 186 -2436
rect 180 -2448 186 -2442
rect 180 -2454 186 -2448
rect 180 -2460 186 -2454
rect 180 -2466 186 -2460
rect 180 -2472 186 -2466
rect 180 -2478 186 -2472
rect 180 -2484 186 -2478
rect 180 -2490 186 -2484
rect 180 -2496 186 -2490
rect 180 -2502 186 -2496
rect 180 -2508 186 -2502
rect 180 -2514 186 -2508
rect 180 -2520 186 -2514
rect 180 -2526 186 -2520
rect 180 -2532 186 -2526
rect 180 -2538 186 -2532
rect 180 -2544 186 -2538
rect 180 -2550 186 -2544
rect 180 -2556 186 -2550
rect 180 -2562 186 -2556
rect 180 -2568 186 -2562
rect 180 -2574 186 -2568
rect 180 -2580 186 -2574
rect 180 -2586 186 -2580
rect 180 -2592 186 -2586
rect 180 -2598 186 -2592
rect 180 -2604 186 -2598
rect 180 -2610 186 -2604
rect 180 -2616 186 -2610
rect 180 -2622 186 -2616
rect 180 -2628 186 -2622
rect 180 -2634 186 -2628
rect 180 -2640 186 -2634
rect 180 -2646 186 -2640
rect 180 -2652 186 -2646
rect 180 -2658 186 -2652
rect 180 -2664 186 -2658
rect 180 -2670 186 -2664
rect 180 -2676 186 -2670
rect 180 -2682 186 -2676
rect 180 -2688 186 -2682
rect 180 -2694 186 -2688
rect 180 -2700 186 -2694
rect 180 -2706 186 -2700
rect 180 -2712 186 -2706
rect 180 -2718 186 -2712
rect 180 -2724 186 -2718
rect 180 -2730 186 -2724
rect 180 -2736 186 -2730
rect 180 -2742 186 -2736
rect 180 -2748 186 -2742
rect 180 -2754 186 -2748
rect 180 -2760 186 -2754
rect 180 -2766 186 -2760
rect 180 -2772 186 -2766
rect 180 -2778 186 -2772
rect 180 -2784 186 -2778
rect 180 -2790 186 -2784
rect 180 -2796 186 -2790
rect 180 -2802 186 -2796
rect 180 -2808 186 -2802
rect 180 -2814 186 -2808
rect 180 -2820 186 -2814
rect 180 -2826 186 -2820
rect 180 -2832 186 -2826
rect 180 -2838 186 -2832
rect 180 -2844 186 -2838
rect 180 -2850 186 -2844
rect 180 -2856 186 -2850
rect 180 -2862 186 -2856
rect 180 -2868 186 -2862
rect 180 -2874 186 -2868
rect 180 -2880 186 -2874
rect 180 -2886 186 -2880
rect 180 -2892 186 -2886
rect 180 -2898 186 -2892
rect 180 -2904 186 -2898
rect 180 -2910 186 -2904
rect 180 -2916 186 -2910
rect 180 -2922 186 -2916
rect 180 -2928 186 -2922
rect 180 -2934 186 -2928
rect 180 -2940 186 -2934
rect 180 -2946 186 -2940
rect 186 -1668 192 -1662
rect 186 -1674 192 -1668
rect 186 -1680 192 -1674
rect 186 -1686 192 -1680
rect 186 -1692 192 -1686
rect 186 -1698 192 -1692
rect 186 -1704 192 -1698
rect 186 -1710 192 -1704
rect 186 -1716 192 -1710
rect 186 -1722 192 -1716
rect 186 -1728 192 -1722
rect 186 -1734 192 -1728
rect 186 -1740 192 -1734
rect 186 -1746 192 -1740
rect 186 -1752 192 -1746
rect 186 -1758 192 -1752
rect 186 -1764 192 -1758
rect 186 -1770 192 -1764
rect 186 -1776 192 -1770
rect 186 -1782 192 -1776
rect 186 -1788 192 -1782
rect 186 -1794 192 -1788
rect 186 -1800 192 -1794
rect 186 -1806 192 -1800
rect 186 -1812 192 -1806
rect 186 -1818 192 -1812
rect 186 -1824 192 -1818
rect 186 -1830 192 -1824
rect 186 -1836 192 -1830
rect 186 -1842 192 -1836
rect 186 -1848 192 -1842
rect 186 -1854 192 -1848
rect 186 -1860 192 -1854
rect 186 -1866 192 -1860
rect 186 -1872 192 -1866
rect 186 -1878 192 -1872
rect 186 -1884 192 -1878
rect 186 -1890 192 -1884
rect 186 -1896 192 -1890
rect 186 -1902 192 -1896
rect 186 -1908 192 -1902
rect 186 -1914 192 -1908
rect 186 -1920 192 -1914
rect 186 -1926 192 -1920
rect 186 -1932 192 -1926
rect 186 -1938 192 -1932
rect 186 -1944 192 -1938
rect 186 -1950 192 -1944
rect 186 -1956 192 -1950
rect 186 -1962 192 -1956
rect 186 -1968 192 -1962
rect 186 -1974 192 -1968
rect 186 -1980 192 -1974
rect 186 -1986 192 -1980
rect 186 -1992 192 -1986
rect 186 -1998 192 -1992
rect 186 -2004 192 -1998
rect 186 -2010 192 -2004
rect 186 -2016 192 -2010
rect 186 -2022 192 -2016
rect 186 -2028 192 -2022
rect 186 -2034 192 -2028
rect 186 -2040 192 -2034
rect 186 -2046 192 -2040
rect 186 -2052 192 -2046
rect 186 -2058 192 -2052
rect 186 -2064 192 -2058
rect 186 -2070 192 -2064
rect 186 -2076 192 -2070
rect 186 -2082 192 -2076
rect 186 -2088 192 -2082
rect 186 -2094 192 -2088
rect 186 -2100 192 -2094
rect 186 -2106 192 -2100
rect 186 -2112 192 -2106
rect 186 -2118 192 -2112
rect 186 -2124 192 -2118
rect 186 -2130 192 -2124
rect 186 -2136 192 -2130
rect 186 -2142 192 -2136
rect 186 -2148 192 -2142
rect 186 -2154 192 -2148
rect 186 -2160 192 -2154
rect 186 -2166 192 -2160
rect 186 -2172 192 -2166
rect 186 -2178 192 -2172
rect 186 -2184 192 -2178
rect 186 -2190 192 -2184
rect 186 -2196 192 -2190
rect 186 -2202 192 -2196
rect 186 -2208 192 -2202
rect 186 -2214 192 -2208
rect 186 -2220 192 -2214
rect 186 -2226 192 -2220
rect 186 -2232 192 -2226
rect 186 -2238 192 -2232
rect 186 -2244 192 -2238
rect 186 -2250 192 -2244
rect 186 -2256 192 -2250
rect 186 -2262 192 -2256
rect 186 -2268 192 -2262
rect 186 -2274 192 -2268
rect 186 -2280 192 -2274
rect 186 -2286 192 -2280
rect 186 -2292 192 -2286
rect 186 -2298 192 -2292
rect 186 -2304 192 -2298
rect 186 -2310 192 -2304
rect 186 -2316 192 -2310
rect 186 -2322 192 -2316
rect 186 -2328 192 -2322
rect 186 -2334 192 -2328
rect 186 -2340 192 -2334
rect 186 -2346 192 -2340
rect 186 -2352 192 -2346
rect 186 -2358 192 -2352
rect 186 -2364 192 -2358
rect 186 -2370 192 -2364
rect 186 -2376 192 -2370
rect 186 -2382 192 -2376
rect 186 -2388 192 -2382
rect 186 -2394 192 -2388
rect 186 -2400 192 -2394
rect 186 -2406 192 -2400
rect 186 -2412 192 -2406
rect 186 -2418 192 -2412
rect 186 -2424 192 -2418
rect 186 -2430 192 -2424
rect 186 -2436 192 -2430
rect 186 -2442 192 -2436
rect 186 -2448 192 -2442
rect 186 -2454 192 -2448
rect 186 -2460 192 -2454
rect 186 -2466 192 -2460
rect 186 -2472 192 -2466
rect 186 -2478 192 -2472
rect 186 -2484 192 -2478
rect 186 -2490 192 -2484
rect 186 -2496 192 -2490
rect 186 -2502 192 -2496
rect 186 -2508 192 -2502
rect 186 -2514 192 -2508
rect 186 -2520 192 -2514
rect 186 -2526 192 -2520
rect 186 -2532 192 -2526
rect 186 -2538 192 -2532
rect 186 -2544 192 -2538
rect 186 -2550 192 -2544
rect 186 -2556 192 -2550
rect 186 -2562 192 -2556
rect 186 -2568 192 -2562
rect 186 -2574 192 -2568
rect 186 -2580 192 -2574
rect 186 -2586 192 -2580
rect 186 -2592 192 -2586
rect 186 -2598 192 -2592
rect 186 -2604 192 -2598
rect 186 -2610 192 -2604
rect 186 -2616 192 -2610
rect 186 -2622 192 -2616
rect 186 -2628 192 -2622
rect 186 -2634 192 -2628
rect 186 -2640 192 -2634
rect 186 -2646 192 -2640
rect 186 -2652 192 -2646
rect 186 -2658 192 -2652
rect 186 -2664 192 -2658
rect 186 -2670 192 -2664
rect 186 -2676 192 -2670
rect 186 -2682 192 -2676
rect 186 -2688 192 -2682
rect 186 -2694 192 -2688
rect 186 -2700 192 -2694
rect 186 -2706 192 -2700
rect 186 -2712 192 -2706
rect 186 -2718 192 -2712
rect 186 -2724 192 -2718
rect 186 -2730 192 -2724
rect 186 -2736 192 -2730
rect 186 -2742 192 -2736
rect 186 -2748 192 -2742
rect 186 -2754 192 -2748
rect 186 -2760 192 -2754
rect 186 -2766 192 -2760
rect 186 -2772 192 -2766
rect 186 -2778 192 -2772
rect 186 -2784 192 -2778
rect 186 -2790 192 -2784
rect 186 -2796 192 -2790
rect 186 -2802 192 -2796
rect 186 -2808 192 -2802
rect 186 -2814 192 -2808
rect 186 -2820 192 -2814
rect 186 -2826 192 -2820
rect 186 -2832 192 -2826
rect 186 -2838 192 -2832
rect 186 -2844 192 -2838
rect 186 -2850 192 -2844
rect 186 -2856 192 -2850
rect 186 -2862 192 -2856
rect 186 -2868 192 -2862
rect 186 -2874 192 -2868
rect 186 -2880 192 -2874
rect 186 -2886 192 -2880
rect 186 -2892 192 -2886
rect 186 -2898 192 -2892
rect 186 -2904 192 -2898
rect 186 -2910 192 -2904
rect 186 -2916 192 -2910
rect 186 -2922 192 -2916
rect 186 -2928 192 -2922
rect 186 -2934 192 -2928
rect 186 -2940 192 -2934
rect 186 -2946 192 -2940
rect 186 -2952 192 -2946
rect 186 -2958 192 -2952
rect 192 -1662 198 -1656
rect 192 -1668 198 -1662
rect 192 -1674 198 -1668
rect 192 -1680 198 -1674
rect 192 -1686 198 -1680
rect 192 -1692 198 -1686
rect 192 -1698 198 -1692
rect 192 -1704 198 -1698
rect 192 -1710 198 -1704
rect 192 -1716 198 -1710
rect 192 -1722 198 -1716
rect 192 -1728 198 -1722
rect 192 -1734 198 -1728
rect 192 -1740 198 -1734
rect 192 -1746 198 -1740
rect 192 -1752 198 -1746
rect 192 -1758 198 -1752
rect 192 -1764 198 -1758
rect 192 -1770 198 -1764
rect 192 -1776 198 -1770
rect 192 -1782 198 -1776
rect 192 -1788 198 -1782
rect 192 -1794 198 -1788
rect 192 -1800 198 -1794
rect 192 -1806 198 -1800
rect 192 -1812 198 -1806
rect 192 -1818 198 -1812
rect 192 -1824 198 -1818
rect 192 -1830 198 -1824
rect 192 -1836 198 -1830
rect 192 -1842 198 -1836
rect 192 -1848 198 -1842
rect 192 -1854 198 -1848
rect 192 -1860 198 -1854
rect 192 -1866 198 -1860
rect 192 -1872 198 -1866
rect 192 -1878 198 -1872
rect 192 -1884 198 -1878
rect 192 -1890 198 -1884
rect 192 -1896 198 -1890
rect 192 -1902 198 -1896
rect 192 -1908 198 -1902
rect 192 -1914 198 -1908
rect 192 -1920 198 -1914
rect 192 -1926 198 -1920
rect 192 -1932 198 -1926
rect 192 -1938 198 -1932
rect 192 -1944 198 -1938
rect 192 -1950 198 -1944
rect 192 -1956 198 -1950
rect 192 -1962 198 -1956
rect 192 -1968 198 -1962
rect 192 -1974 198 -1968
rect 192 -1980 198 -1974
rect 192 -1986 198 -1980
rect 192 -1992 198 -1986
rect 192 -1998 198 -1992
rect 192 -2004 198 -1998
rect 192 -2010 198 -2004
rect 192 -2016 198 -2010
rect 192 -2022 198 -2016
rect 192 -2028 198 -2022
rect 192 -2034 198 -2028
rect 192 -2040 198 -2034
rect 192 -2046 198 -2040
rect 192 -2052 198 -2046
rect 192 -2058 198 -2052
rect 192 -2064 198 -2058
rect 192 -2070 198 -2064
rect 192 -2076 198 -2070
rect 192 -2082 198 -2076
rect 192 -2088 198 -2082
rect 192 -2094 198 -2088
rect 192 -2100 198 -2094
rect 192 -2106 198 -2100
rect 192 -2112 198 -2106
rect 192 -2118 198 -2112
rect 192 -2124 198 -2118
rect 192 -2130 198 -2124
rect 192 -2136 198 -2130
rect 192 -2142 198 -2136
rect 192 -2148 198 -2142
rect 192 -2154 198 -2148
rect 192 -2160 198 -2154
rect 192 -2166 198 -2160
rect 192 -2172 198 -2166
rect 192 -2178 198 -2172
rect 192 -2184 198 -2178
rect 192 -2190 198 -2184
rect 192 -2196 198 -2190
rect 192 -2202 198 -2196
rect 192 -2208 198 -2202
rect 192 -2214 198 -2208
rect 192 -2220 198 -2214
rect 192 -2226 198 -2220
rect 192 -2232 198 -2226
rect 192 -2238 198 -2232
rect 192 -2244 198 -2238
rect 192 -2250 198 -2244
rect 192 -2256 198 -2250
rect 192 -2262 198 -2256
rect 192 -2268 198 -2262
rect 192 -2274 198 -2268
rect 192 -2280 198 -2274
rect 192 -2286 198 -2280
rect 192 -2292 198 -2286
rect 192 -2298 198 -2292
rect 192 -2304 198 -2298
rect 192 -2310 198 -2304
rect 192 -2316 198 -2310
rect 192 -2322 198 -2316
rect 192 -2328 198 -2322
rect 192 -2334 198 -2328
rect 192 -2340 198 -2334
rect 192 -2346 198 -2340
rect 192 -2352 198 -2346
rect 192 -2358 198 -2352
rect 192 -2364 198 -2358
rect 192 -2370 198 -2364
rect 192 -2376 198 -2370
rect 192 -2382 198 -2376
rect 192 -2388 198 -2382
rect 192 -2394 198 -2388
rect 192 -2400 198 -2394
rect 192 -2406 198 -2400
rect 192 -2412 198 -2406
rect 192 -2418 198 -2412
rect 192 -2424 198 -2418
rect 192 -2430 198 -2424
rect 192 -2436 198 -2430
rect 192 -2442 198 -2436
rect 192 -2448 198 -2442
rect 192 -2454 198 -2448
rect 192 -2460 198 -2454
rect 192 -2466 198 -2460
rect 192 -2472 198 -2466
rect 192 -2478 198 -2472
rect 192 -2484 198 -2478
rect 192 -2490 198 -2484
rect 192 -2496 198 -2490
rect 192 -2502 198 -2496
rect 192 -2508 198 -2502
rect 192 -2514 198 -2508
rect 192 -2520 198 -2514
rect 192 -2526 198 -2520
rect 192 -2532 198 -2526
rect 192 -2538 198 -2532
rect 192 -2544 198 -2538
rect 192 -2550 198 -2544
rect 192 -2556 198 -2550
rect 192 -2562 198 -2556
rect 192 -2568 198 -2562
rect 192 -2574 198 -2568
rect 192 -2580 198 -2574
rect 192 -2586 198 -2580
rect 192 -2592 198 -2586
rect 192 -2598 198 -2592
rect 192 -2604 198 -2598
rect 192 -2610 198 -2604
rect 192 -2616 198 -2610
rect 192 -2622 198 -2616
rect 192 -2628 198 -2622
rect 192 -2634 198 -2628
rect 192 -2640 198 -2634
rect 192 -2646 198 -2640
rect 192 -2652 198 -2646
rect 192 -2658 198 -2652
rect 192 -2664 198 -2658
rect 192 -2670 198 -2664
rect 192 -2676 198 -2670
rect 192 -2682 198 -2676
rect 192 -2688 198 -2682
rect 192 -2694 198 -2688
rect 192 -2700 198 -2694
rect 192 -2706 198 -2700
rect 192 -2712 198 -2706
rect 192 -2718 198 -2712
rect 192 -2724 198 -2718
rect 192 -2730 198 -2724
rect 192 -2736 198 -2730
rect 192 -2742 198 -2736
rect 192 -2748 198 -2742
rect 192 -2754 198 -2748
rect 192 -2760 198 -2754
rect 192 -2766 198 -2760
rect 192 -2772 198 -2766
rect 192 -2778 198 -2772
rect 192 -2784 198 -2778
rect 192 -2790 198 -2784
rect 192 -2796 198 -2790
rect 192 -2802 198 -2796
rect 192 -2808 198 -2802
rect 192 -2814 198 -2808
rect 192 -2820 198 -2814
rect 192 -2826 198 -2820
rect 192 -2832 198 -2826
rect 192 -2838 198 -2832
rect 192 -2844 198 -2838
rect 192 -2850 198 -2844
rect 192 -2856 198 -2850
rect 192 -2862 198 -2856
rect 192 -2868 198 -2862
rect 192 -2874 198 -2868
rect 192 -2880 198 -2874
rect 192 -2886 198 -2880
rect 192 -2892 198 -2886
rect 192 -2898 198 -2892
rect 192 -2904 198 -2898
rect 192 -2910 198 -2904
rect 192 -2916 198 -2910
rect 192 -2922 198 -2916
rect 192 -2928 198 -2922
rect 192 -2934 198 -2928
rect 192 -2940 198 -2934
rect 192 -2946 198 -2940
rect 192 -2952 198 -2946
rect 192 -2958 198 -2952
rect 192 -2964 198 -2958
rect 192 -2970 198 -2964
rect 198 -1650 204 -1644
rect 198 -1656 204 -1650
rect 198 -1662 204 -1656
rect 198 -1668 204 -1662
rect 198 -1674 204 -1668
rect 198 -1680 204 -1674
rect 198 -1686 204 -1680
rect 198 -1692 204 -1686
rect 198 -1698 204 -1692
rect 198 -1704 204 -1698
rect 198 -1710 204 -1704
rect 198 -1716 204 -1710
rect 198 -1722 204 -1716
rect 198 -1728 204 -1722
rect 198 -1734 204 -1728
rect 198 -1740 204 -1734
rect 198 -1746 204 -1740
rect 198 -1752 204 -1746
rect 198 -1758 204 -1752
rect 198 -1764 204 -1758
rect 198 -1770 204 -1764
rect 198 -1776 204 -1770
rect 198 -1782 204 -1776
rect 198 -1788 204 -1782
rect 198 -1794 204 -1788
rect 198 -1800 204 -1794
rect 198 -1806 204 -1800
rect 198 -1812 204 -1806
rect 198 -1818 204 -1812
rect 198 -1824 204 -1818
rect 198 -1830 204 -1824
rect 198 -1836 204 -1830
rect 198 -1842 204 -1836
rect 198 -1848 204 -1842
rect 198 -1854 204 -1848
rect 198 -1860 204 -1854
rect 198 -1866 204 -1860
rect 198 -1872 204 -1866
rect 198 -1878 204 -1872
rect 198 -1884 204 -1878
rect 198 -1890 204 -1884
rect 198 -1896 204 -1890
rect 198 -1902 204 -1896
rect 198 -1908 204 -1902
rect 198 -1914 204 -1908
rect 198 -1920 204 -1914
rect 198 -1926 204 -1920
rect 198 -1932 204 -1926
rect 198 -1938 204 -1932
rect 198 -1944 204 -1938
rect 198 -1950 204 -1944
rect 198 -1956 204 -1950
rect 198 -1962 204 -1956
rect 198 -1968 204 -1962
rect 198 -1974 204 -1968
rect 198 -1980 204 -1974
rect 198 -1986 204 -1980
rect 198 -1992 204 -1986
rect 198 -1998 204 -1992
rect 198 -2004 204 -1998
rect 198 -2010 204 -2004
rect 198 -2016 204 -2010
rect 198 -2022 204 -2016
rect 198 -2028 204 -2022
rect 198 -2034 204 -2028
rect 198 -2040 204 -2034
rect 198 -2046 204 -2040
rect 198 -2052 204 -2046
rect 198 -2058 204 -2052
rect 198 -2064 204 -2058
rect 198 -2070 204 -2064
rect 198 -2076 204 -2070
rect 198 -2082 204 -2076
rect 198 -2088 204 -2082
rect 198 -2094 204 -2088
rect 198 -2100 204 -2094
rect 198 -2106 204 -2100
rect 198 -2112 204 -2106
rect 198 -2118 204 -2112
rect 198 -2124 204 -2118
rect 198 -2130 204 -2124
rect 198 -2136 204 -2130
rect 198 -2142 204 -2136
rect 198 -2148 204 -2142
rect 198 -2154 204 -2148
rect 198 -2160 204 -2154
rect 198 -2166 204 -2160
rect 198 -2172 204 -2166
rect 198 -2178 204 -2172
rect 198 -2184 204 -2178
rect 198 -2190 204 -2184
rect 198 -2196 204 -2190
rect 198 -2202 204 -2196
rect 198 -2208 204 -2202
rect 198 -2214 204 -2208
rect 198 -2220 204 -2214
rect 198 -2226 204 -2220
rect 198 -2232 204 -2226
rect 198 -2238 204 -2232
rect 198 -2244 204 -2238
rect 198 -2250 204 -2244
rect 198 -2256 204 -2250
rect 198 -2262 204 -2256
rect 198 -2268 204 -2262
rect 198 -2274 204 -2268
rect 198 -2280 204 -2274
rect 198 -2286 204 -2280
rect 198 -2292 204 -2286
rect 198 -2298 204 -2292
rect 198 -2304 204 -2298
rect 198 -2310 204 -2304
rect 198 -2316 204 -2310
rect 198 -2322 204 -2316
rect 198 -2328 204 -2322
rect 198 -2334 204 -2328
rect 198 -2340 204 -2334
rect 198 -2346 204 -2340
rect 198 -2352 204 -2346
rect 198 -2358 204 -2352
rect 198 -2364 204 -2358
rect 198 -2370 204 -2364
rect 198 -2376 204 -2370
rect 198 -2382 204 -2376
rect 198 -2388 204 -2382
rect 198 -2394 204 -2388
rect 198 -2400 204 -2394
rect 198 -2406 204 -2400
rect 198 -2412 204 -2406
rect 198 -2418 204 -2412
rect 198 -2424 204 -2418
rect 198 -2430 204 -2424
rect 198 -2436 204 -2430
rect 198 -2442 204 -2436
rect 198 -2448 204 -2442
rect 198 -2454 204 -2448
rect 198 -2460 204 -2454
rect 198 -2466 204 -2460
rect 198 -2472 204 -2466
rect 198 -2478 204 -2472
rect 198 -2484 204 -2478
rect 198 -2490 204 -2484
rect 198 -2496 204 -2490
rect 198 -2502 204 -2496
rect 198 -2508 204 -2502
rect 198 -2514 204 -2508
rect 198 -2520 204 -2514
rect 198 -2526 204 -2520
rect 198 -2532 204 -2526
rect 198 -2538 204 -2532
rect 198 -2544 204 -2538
rect 198 -2550 204 -2544
rect 198 -2556 204 -2550
rect 198 -2562 204 -2556
rect 198 -2568 204 -2562
rect 198 -2574 204 -2568
rect 198 -2580 204 -2574
rect 198 -2586 204 -2580
rect 198 -2592 204 -2586
rect 198 -2598 204 -2592
rect 198 -2604 204 -2598
rect 198 -2610 204 -2604
rect 198 -2616 204 -2610
rect 198 -2622 204 -2616
rect 198 -2628 204 -2622
rect 198 -2634 204 -2628
rect 198 -2640 204 -2634
rect 198 -2646 204 -2640
rect 198 -2652 204 -2646
rect 198 -2658 204 -2652
rect 198 -2664 204 -2658
rect 198 -2670 204 -2664
rect 198 -2676 204 -2670
rect 198 -2682 204 -2676
rect 198 -2688 204 -2682
rect 198 -2694 204 -2688
rect 198 -2700 204 -2694
rect 198 -2706 204 -2700
rect 198 -2712 204 -2706
rect 198 -2718 204 -2712
rect 198 -2724 204 -2718
rect 198 -2730 204 -2724
rect 198 -2736 204 -2730
rect 198 -2742 204 -2736
rect 198 -2748 204 -2742
rect 198 -2754 204 -2748
rect 198 -2760 204 -2754
rect 198 -2766 204 -2760
rect 198 -2772 204 -2766
rect 198 -2778 204 -2772
rect 198 -2784 204 -2778
rect 198 -2790 204 -2784
rect 198 -2796 204 -2790
rect 198 -2802 204 -2796
rect 198 -2808 204 -2802
rect 198 -2814 204 -2808
rect 198 -2820 204 -2814
rect 198 -2826 204 -2820
rect 198 -2832 204 -2826
rect 198 -2838 204 -2832
rect 198 -2844 204 -2838
rect 198 -2850 204 -2844
rect 198 -2856 204 -2850
rect 198 -2862 204 -2856
rect 198 -2868 204 -2862
rect 198 -2874 204 -2868
rect 198 -2880 204 -2874
rect 198 -2886 204 -2880
rect 198 -2892 204 -2886
rect 198 -2898 204 -2892
rect 198 -2904 204 -2898
rect 198 -2910 204 -2904
rect 198 -2916 204 -2910
rect 198 -2922 204 -2916
rect 198 -2928 204 -2922
rect 198 -2934 204 -2928
rect 198 -2940 204 -2934
rect 198 -2946 204 -2940
rect 198 -2952 204 -2946
rect 198 -2958 204 -2952
rect 198 -2964 204 -2958
rect 198 -2970 204 -2964
rect 198 -2976 204 -2970
rect 204 -1638 210 -1632
rect 204 -1644 210 -1638
rect 204 -1650 210 -1644
rect 204 -1656 210 -1650
rect 204 -1662 210 -1656
rect 204 -1668 210 -1662
rect 204 -1674 210 -1668
rect 204 -1680 210 -1674
rect 204 -1686 210 -1680
rect 204 -1692 210 -1686
rect 204 -1698 210 -1692
rect 204 -1704 210 -1698
rect 204 -1710 210 -1704
rect 204 -1716 210 -1710
rect 204 -1722 210 -1716
rect 204 -1728 210 -1722
rect 204 -1734 210 -1728
rect 204 -1740 210 -1734
rect 204 -1746 210 -1740
rect 204 -1752 210 -1746
rect 204 -1758 210 -1752
rect 204 -1764 210 -1758
rect 204 -1770 210 -1764
rect 204 -1776 210 -1770
rect 204 -1782 210 -1776
rect 204 -1788 210 -1782
rect 204 -1794 210 -1788
rect 204 -1800 210 -1794
rect 204 -1806 210 -1800
rect 204 -1812 210 -1806
rect 204 -1818 210 -1812
rect 204 -1824 210 -1818
rect 204 -1830 210 -1824
rect 204 -1836 210 -1830
rect 204 -1842 210 -1836
rect 204 -1848 210 -1842
rect 204 -1854 210 -1848
rect 204 -1860 210 -1854
rect 204 -1866 210 -1860
rect 204 -1872 210 -1866
rect 204 -1878 210 -1872
rect 204 -1884 210 -1878
rect 204 -1890 210 -1884
rect 204 -1896 210 -1890
rect 204 -1902 210 -1896
rect 204 -1908 210 -1902
rect 204 -1914 210 -1908
rect 204 -1920 210 -1914
rect 204 -1926 210 -1920
rect 204 -1932 210 -1926
rect 204 -1938 210 -1932
rect 204 -1944 210 -1938
rect 204 -1950 210 -1944
rect 204 -1956 210 -1950
rect 204 -1962 210 -1956
rect 204 -1968 210 -1962
rect 204 -1974 210 -1968
rect 204 -1980 210 -1974
rect 204 -1986 210 -1980
rect 204 -1992 210 -1986
rect 204 -1998 210 -1992
rect 204 -2004 210 -1998
rect 204 -2010 210 -2004
rect 204 -2016 210 -2010
rect 204 -2022 210 -2016
rect 204 -2028 210 -2022
rect 204 -2034 210 -2028
rect 204 -2040 210 -2034
rect 204 -2046 210 -2040
rect 204 -2052 210 -2046
rect 204 -2058 210 -2052
rect 204 -2064 210 -2058
rect 204 -2070 210 -2064
rect 204 -2076 210 -2070
rect 204 -2082 210 -2076
rect 204 -2088 210 -2082
rect 204 -2094 210 -2088
rect 204 -2100 210 -2094
rect 204 -2106 210 -2100
rect 204 -2112 210 -2106
rect 204 -2118 210 -2112
rect 204 -2124 210 -2118
rect 204 -2130 210 -2124
rect 204 -2136 210 -2130
rect 204 -2142 210 -2136
rect 204 -2148 210 -2142
rect 204 -2154 210 -2148
rect 204 -2160 210 -2154
rect 204 -2166 210 -2160
rect 204 -2172 210 -2166
rect 204 -2178 210 -2172
rect 204 -2184 210 -2178
rect 204 -2190 210 -2184
rect 204 -2196 210 -2190
rect 204 -2202 210 -2196
rect 204 -2208 210 -2202
rect 204 -2214 210 -2208
rect 204 -2220 210 -2214
rect 204 -2226 210 -2220
rect 204 -2232 210 -2226
rect 204 -2238 210 -2232
rect 204 -2244 210 -2238
rect 204 -2250 210 -2244
rect 204 -2256 210 -2250
rect 204 -2262 210 -2256
rect 204 -2268 210 -2262
rect 204 -2274 210 -2268
rect 204 -2280 210 -2274
rect 204 -2286 210 -2280
rect 204 -2292 210 -2286
rect 204 -2298 210 -2292
rect 204 -2304 210 -2298
rect 204 -2310 210 -2304
rect 204 -2316 210 -2310
rect 204 -2322 210 -2316
rect 204 -2328 210 -2322
rect 204 -2334 210 -2328
rect 204 -2340 210 -2334
rect 204 -2346 210 -2340
rect 204 -2352 210 -2346
rect 204 -2358 210 -2352
rect 204 -2364 210 -2358
rect 204 -2370 210 -2364
rect 204 -2376 210 -2370
rect 204 -2382 210 -2376
rect 204 -2388 210 -2382
rect 204 -2394 210 -2388
rect 204 -2400 210 -2394
rect 204 -2406 210 -2400
rect 204 -2412 210 -2406
rect 204 -2418 210 -2412
rect 204 -2424 210 -2418
rect 204 -2430 210 -2424
rect 204 -2436 210 -2430
rect 204 -2442 210 -2436
rect 204 -2448 210 -2442
rect 204 -2454 210 -2448
rect 204 -2460 210 -2454
rect 204 -2466 210 -2460
rect 204 -2472 210 -2466
rect 204 -2478 210 -2472
rect 204 -2484 210 -2478
rect 204 -2490 210 -2484
rect 204 -2496 210 -2490
rect 204 -2502 210 -2496
rect 204 -2508 210 -2502
rect 204 -2514 210 -2508
rect 204 -2520 210 -2514
rect 204 -2526 210 -2520
rect 204 -2532 210 -2526
rect 204 -2538 210 -2532
rect 204 -2544 210 -2538
rect 204 -2550 210 -2544
rect 204 -2556 210 -2550
rect 204 -2562 210 -2556
rect 204 -2568 210 -2562
rect 204 -2574 210 -2568
rect 204 -2580 210 -2574
rect 204 -2586 210 -2580
rect 204 -2592 210 -2586
rect 204 -2598 210 -2592
rect 204 -2604 210 -2598
rect 204 -2610 210 -2604
rect 204 -2616 210 -2610
rect 204 -2622 210 -2616
rect 204 -2628 210 -2622
rect 204 -2634 210 -2628
rect 204 -2640 210 -2634
rect 204 -2646 210 -2640
rect 204 -2652 210 -2646
rect 204 -2658 210 -2652
rect 204 -2664 210 -2658
rect 204 -2670 210 -2664
rect 204 -2676 210 -2670
rect 204 -2682 210 -2676
rect 204 -2688 210 -2682
rect 204 -2694 210 -2688
rect 204 -2700 210 -2694
rect 204 -2706 210 -2700
rect 204 -2712 210 -2706
rect 204 -2718 210 -2712
rect 204 -2724 210 -2718
rect 204 -2730 210 -2724
rect 204 -2736 210 -2730
rect 204 -2742 210 -2736
rect 204 -2748 210 -2742
rect 204 -2754 210 -2748
rect 204 -2760 210 -2754
rect 204 -2766 210 -2760
rect 204 -2772 210 -2766
rect 204 -2778 210 -2772
rect 204 -2784 210 -2778
rect 204 -2790 210 -2784
rect 204 -2796 210 -2790
rect 204 -2802 210 -2796
rect 204 -2808 210 -2802
rect 204 -2814 210 -2808
rect 204 -2820 210 -2814
rect 204 -2826 210 -2820
rect 204 -2832 210 -2826
rect 204 -2838 210 -2832
rect 204 -2844 210 -2838
rect 204 -2850 210 -2844
rect 204 -2856 210 -2850
rect 204 -2862 210 -2856
rect 204 -2868 210 -2862
rect 204 -2874 210 -2868
rect 204 -2880 210 -2874
rect 204 -2886 210 -2880
rect 204 -2892 210 -2886
rect 204 -2898 210 -2892
rect 204 -2904 210 -2898
rect 204 -2910 210 -2904
rect 204 -2916 210 -2910
rect 204 -2922 210 -2916
rect 204 -2928 210 -2922
rect 204 -2934 210 -2928
rect 204 -2940 210 -2934
rect 204 -2946 210 -2940
rect 204 -2952 210 -2946
rect 204 -2958 210 -2952
rect 204 -2964 210 -2958
rect 204 -2970 210 -2964
rect 204 -2976 210 -2970
rect 204 -2982 210 -2976
rect 204 -2988 210 -2982
rect 210 -1632 216 -1626
rect 210 -1638 216 -1632
rect 210 -1644 216 -1638
rect 210 -1650 216 -1644
rect 210 -1656 216 -1650
rect 210 -1662 216 -1656
rect 210 -1668 216 -1662
rect 210 -1674 216 -1668
rect 210 -1680 216 -1674
rect 210 -1686 216 -1680
rect 210 -1692 216 -1686
rect 210 -1698 216 -1692
rect 210 -1704 216 -1698
rect 210 -1710 216 -1704
rect 210 -1716 216 -1710
rect 210 -1722 216 -1716
rect 210 -1728 216 -1722
rect 210 -1734 216 -1728
rect 210 -1740 216 -1734
rect 210 -1746 216 -1740
rect 210 -1752 216 -1746
rect 210 -1758 216 -1752
rect 210 -1764 216 -1758
rect 210 -1770 216 -1764
rect 210 -1776 216 -1770
rect 210 -1782 216 -1776
rect 210 -1788 216 -1782
rect 210 -1794 216 -1788
rect 210 -1800 216 -1794
rect 210 -1806 216 -1800
rect 210 -1812 216 -1806
rect 210 -1818 216 -1812
rect 210 -1824 216 -1818
rect 210 -1830 216 -1824
rect 210 -1836 216 -1830
rect 210 -1842 216 -1836
rect 210 -1848 216 -1842
rect 210 -1854 216 -1848
rect 210 -1860 216 -1854
rect 210 -1866 216 -1860
rect 210 -1872 216 -1866
rect 210 -1878 216 -1872
rect 210 -1884 216 -1878
rect 210 -1890 216 -1884
rect 210 -1896 216 -1890
rect 210 -1902 216 -1896
rect 210 -1908 216 -1902
rect 210 -1914 216 -1908
rect 210 -1920 216 -1914
rect 210 -1926 216 -1920
rect 210 -1932 216 -1926
rect 210 -1938 216 -1932
rect 210 -1944 216 -1938
rect 210 -1950 216 -1944
rect 210 -1956 216 -1950
rect 210 -1962 216 -1956
rect 210 -1968 216 -1962
rect 210 -1974 216 -1968
rect 210 -1980 216 -1974
rect 210 -1986 216 -1980
rect 210 -1992 216 -1986
rect 210 -1998 216 -1992
rect 210 -2004 216 -1998
rect 210 -2010 216 -2004
rect 210 -2016 216 -2010
rect 210 -2022 216 -2016
rect 210 -2028 216 -2022
rect 210 -2034 216 -2028
rect 210 -2040 216 -2034
rect 210 -2046 216 -2040
rect 210 -2052 216 -2046
rect 210 -2058 216 -2052
rect 210 -2064 216 -2058
rect 210 -2070 216 -2064
rect 210 -2076 216 -2070
rect 210 -2082 216 -2076
rect 210 -2088 216 -2082
rect 210 -2094 216 -2088
rect 210 -2100 216 -2094
rect 210 -2106 216 -2100
rect 210 -2112 216 -2106
rect 210 -2118 216 -2112
rect 210 -2124 216 -2118
rect 210 -2130 216 -2124
rect 210 -2136 216 -2130
rect 210 -2142 216 -2136
rect 210 -2148 216 -2142
rect 210 -2154 216 -2148
rect 210 -2160 216 -2154
rect 210 -2166 216 -2160
rect 210 -2172 216 -2166
rect 210 -2178 216 -2172
rect 210 -2184 216 -2178
rect 210 -2190 216 -2184
rect 210 -2196 216 -2190
rect 210 -2202 216 -2196
rect 210 -2208 216 -2202
rect 210 -2214 216 -2208
rect 210 -2220 216 -2214
rect 210 -2226 216 -2220
rect 210 -2232 216 -2226
rect 210 -2394 216 -2388
rect 210 -2400 216 -2394
rect 210 -2406 216 -2400
rect 210 -2412 216 -2406
rect 210 -2418 216 -2412
rect 210 -2424 216 -2418
rect 210 -2430 216 -2424
rect 210 -2436 216 -2430
rect 210 -2442 216 -2436
rect 210 -2448 216 -2442
rect 210 -2454 216 -2448
rect 210 -2460 216 -2454
rect 210 -2466 216 -2460
rect 210 -2472 216 -2466
rect 210 -2478 216 -2472
rect 210 -2484 216 -2478
rect 210 -2490 216 -2484
rect 210 -2496 216 -2490
rect 210 -2502 216 -2496
rect 210 -2508 216 -2502
rect 210 -2514 216 -2508
rect 210 -2520 216 -2514
rect 210 -2526 216 -2520
rect 210 -2532 216 -2526
rect 210 -2538 216 -2532
rect 210 -2544 216 -2538
rect 210 -2550 216 -2544
rect 210 -2556 216 -2550
rect 210 -2562 216 -2556
rect 210 -2568 216 -2562
rect 210 -2574 216 -2568
rect 210 -2580 216 -2574
rect 210 -2586 216 -2580
rect 210 -2592 216 -2586
rect 210 -2598 216 -2592
rect 210 -2604 216 -2598
rect 210 -2610 216 -2604
rect 210 -2616 216 -2610
rect 210 -2622 216 -2616
rect 210 -2628 216 -2622
rect 210 -2634 216 -2628
rect 210 -2640 216 -2634
rect 210 -2646 216 -2640
rect 210 -2652 216 -2646
rect 210 -2658 216 -2652
rect 210 -2664 216 -2658
rect 210 -2670 216 -2664
rect 210 -2676 216 -2670
rect 210 -2682 216 -2676
rect 210 -2688 216 -2682
rect 210 -2694 216 -2688
rect 210 -2700 216 -2694
rect 210 -2706 216 -2700
rect 210 -2712 216 -2706
rect 210 -2718 216 -2712
rect 210 -2724 216 -2718
rect 210 -2730 216 -2724
rect 210 -2736 216 -2730
rect 210 -2742 216 -2736
rect 210 -2748 216 -2742
rect 210 -2754 216 -2748
rect 210 -2760 216 -2754
rect 210 -2766 216 -2760
rect 210 -2772 216 -2766
rect 210 -2778 216 -2772
rect 210 -2784 216 -2778
rect 210 -2790 216 -2784
rect 210 -2796 216 -2790
rect 210 -2802 216 -2796
rect 210 -2808 216 -2802
rect 210 -2814 216 -2808
rect 210 -2820 216 -2814
rect 210 -2826 216 -2820
rect 210 -2832 216 -2826
rect 210 -2838 216 -2832
rect 210 -2844 216 -2838
rect 210 -2850 216 -2844
rect 210 -2856 216 -2850
rect 210 -2862 216 -2856
rect 210 -2868 216 -2862
rect 210 -2874 216 -2868
rect 210 -2880 216 -2874
rect 210 -2886 216 -2880
rect 210 -2892 216 -2886
rect 210 -2898 216 -2892
rect 210 -2904 216 -2898
rect 210 -2910 216 -2904
rect 210 -2916 216 -2910
rect 210 -2922 216 -2916
rect 210 -2928 216 -2922
rect 210 -2934 216 -2928
rect 210 -2940 216 -2934
rect 210 -2946 216 -2940
rect 210 -2952 216 -2946
rect 210 -2958 216 -2952
rect 210 -2964 216 -2958
rect 210 -2970 216 -2964
rect 210 -2976 216 -2970
rect 210 -2982 216 -2976
rect 210 -2988 216 -2982
rect 210 -2994 216 -2988
rect 216 -1626 222 -1620
rect 216 -1632 222 -1626
rect 216 -1638 222 -1632
rect 216 -1644 222 -1638
rect 216 -1650 222 -1644
rect 216 -1656 222 -1650
rect 216 -1662 222 -1656
rect 216 -1668 222 -1662
rect 216 -1674 222 -1668
rect 216 -1680 222 -1674
rect 216 -1686 222 -1680
rect 216 -1692 222 -1686
rect 216 -1698 222 -1692
rect 216 -1704 222 -1698
rect 216 -1710 222 -1704
rect 216 -1716 222 -1710
rect 216 -1722 222 -1716
rect 216 -1728 222 -1722
rect 216 -1734 222 -1728
rect 216 -1740 222 -1734
rect 216 -1746 222 -1740
rect 216 -1752 222 -1746
rect 216 -1758 222 -1752
rect 216 -1764 222 -1758
rect 216 -1770 222 -1764
rect 216 -1776 222 -1770
rect 216 -1782 222 -1776
rect 216 -1788 222 -1782
rect 216 -1794 222 -1788
rect 216 -1800 222 -1794
rect 216 -1806 222 -1800
rect 216 -1812 222 -1806
rect 216 -1818 222 -1812
rect 216 -1824 222 -1818
rect 216 -1830 222 -1824
rect 216 -1836 222 -1830
rect 216 -1842 222 -1836
rect 216 -1848 222 -1842
rect 216 -1854 222 -1848
rect 216 -1860 222 -1854
rect 216 -1866 222 -1860
rect 216 -1872 222 -1866
rect 216 -1878 222 -1872
rect 216 -1884 222 -1878
rect 216 -1890 222 -1884
rect 216 -1896 222 -1890
rect 216 -1902 222 -1896
rect 216 -1908 222 -1902
rect 216 -1914 222 -1908
rect 216 -1920 222 -1914
rect 216 -1926 222 -1920
rect 216 -1932 222 -1926
rect 216 -1938 222 -1932
rect 216 -1944 222 -1938
rect 216 -1950 222 -1944
rect 216 -1956 222 -1950
rect 216 -1962 222 -1956
rect 216 -1968 222 -1962
rect 216 -1974 222 -1968
rect 216 -1980 222 -1974
rect 216 -1986 222 -1980
rect 216 -1992 222 -1986
rect 216 -1998 222 -1992
rect 216 -2004 222 -1998
rect 216 -2010 222 -2004
rect 216 -2016 222 -2010
rect 216 -2022 222 -2016
rect 216 -2028 222 -2022
rect 216 -2034 222 -2028
rect 216 -2040 222 -2034
rect 216 -2046 222 -2040
rect 216 -2052 222 -2046
rect 216 -2058 222 -2052
rect 216 -2064 222 -2058
rect 216 -2070 222 -2064
rect 216 -2076 222 -2070
rect 216 -2082 222 -2076
rect 216 -2088 222 -2082
rect 216 -2094 222 -2088
rect 216 -2100 222 -2094
rect 216 -2106 222 -2100
rect 216 -2112 222 -2106
rect 216 -2118 222 -2112
rect 216 -2124 222 -2118
rect 216 -2130 222 -2124
rect 216 -2136 222 -2130
rect 216 -2142 222 -2136
rect 216 -2148 222 -2142
rect 216 -2154 222 -2148
rect 216 -2160 222 -2154
rect 216 -2166 222 -2160
rect 216 -2172 222 -2166
rect 216 -2178 222 -2172
rect 216 -2454 222 -2448
rect 216 -2460 222 -2454
rect 216 -2466 222 -2460
rect 216 -2472 222 -2466
rect 216 -2478 222 -2472
rect 216 -2484 222 -2478
rect 216 -2490 222 -2484
rect 216 -2496 222 -2490
rect 216 -2502 222 -2496
rect 216 -2508 222 -2502
rect 216 -2514 222 -2508
rect 216 -2520 222 -2514
rect 216 -2526 222 -2520
rect 216 -2532 222 -2526
rect 216 -2538 222 -2532
rect 216 -2544 222 -2538
rect 216 -2550 222 -2544
rect 216 -2556 222 -2550
rect 216 -2562 222 -2556
rect 216 -2568 222 -2562
rect 216 -2574 222 -2568
rect 216 -2580 222 -2574
rect 216 -2586 222 -2580
rect 216 -2592 222 -2586
rect 216 -2598 222 -2592
rect 216 -2604 222 -2598
rect 216 -2610 222 -2604
rect 216 -2616 222 -2610
rect 216 -2622 222 -2616
rect 216 -2628 222 -2622
rect 216 -2634 222 -2628
rect 216 -2640 222 -2634
rect 216 -2646 222 -2640
rect 216 -2652 222 -2646
rect 216 -2658 222 -2652
rect 216 -2664 222 -2658
rect 216 -2670 222 -2664
rect 216 -2676 222 -2670
rect 216 -2682 222 -2676
rect 216 -2688 222 -2682
rect 216 -2694 222 -2688
rect 216 -2700 222 -2694
rect 216 -2706 222 -2700
rect 216 -2712 222 -2706
rect 216 -2718 222 -2712
rect 216 -2724 222 -2718
rect 216 -2730 222 -2724
rect 216 -2736 222 -2730
rect 216 -2742 222 -2736
rect 216 -2748 222 -2742
rect 216 -2754 222 -2748
rect 216 -2760 222 -2754
rect 216 -2766 222 -2760
rect 216 -2772 222 -2766
rect 216 -2778 222 -2772
rect 216 -2784 222 -2778
rect 216 -2790 222 -2784
rect 216 -2796 222 -2790
rect 216 -2802 222 -2796
rect 216 -2808 222 -2802
rect 216 -2814 222 -2808
rect 216 -2820 222 -2814
rect 216 -2826 222 -2820
rect 216 -2832 222 -2826
rect 216 -2838 222 -2832
rect 216 -2844 222 -2838
rect 216 -2850 222 -2844
rect 216 -2856 222 -2850
rect 216 -2862 222 -2856
rect 216 -2868 222 -2862
rect 216 -2874 222 -2868
rect 216 -2880 222 -2874
rect 216 -2886 222 -2880
rect 216 -2892 222 -2886
rect 216 -2898 222 -2892
rect 216 -2904 222 -2898
rect 216 -2910 222 -2904
rect 216 -2916 222 -2910
rect 216 -2922 222 -2916
rect 216 -2928 222 -2922
rect 216 -2934 222 -2928
rect 216 -2940 222 -2934
rect 216 -2946 222 -2940
rect 216 -2952 222 -2946
rect 216 -2958 222 -2952
rect 216 -2964 222 -2958
rect 216 -2970 222 -2964
rect 216 -2976 222 -2970
rect 216 -2982 222 -2976
rect 216 -2988 222 -2982
rect 216 -2994 222 -2988
rect 216 -3000 222 -2994
rect 216 -3006 222 -3000
rect 222 -1614 228 -1608
rect 222 -1620 228 -1614
rect 222 -1626 228 -1620
rect 222 -1632 228 -1626
rect 222 -1638 228 -1632
rect 222 -1644 228 -1638
rect 222 -1650 228 -1644
rect 222 -1656 228 -1650
rect 222 -1662 228 -1656
rect 222 -1668 228 -1662
rect 222 -1674 228 -1668
rect 222 -1680 228 -1674
rect 222 -1686 228 -1680
rect 222 -1692 228 -1686
rect 222 -1698 228 -1692
rect 222 -1704 228 -1698
rect 222 -1710 228 -1704
rect 222 -1716 228 -1710
rect 222 -1722 228 -1716
rect 222 -1728 228 -1722
rect 222 -1734 228 -1728
rect 222 -1740 228 -1734
rect 222 -1746 228 -1740
rect 222 -1752 228 -1746
rect 222 -1758 228 -1752
rect 222 -1764 228 -1758
rect 222 -1770 228 -1764
rect 222 -1776 228 -1770
rect 222 -1782 228 -1776
rect 222 -1788 228 -1782
rect 222 -1794 228 -1788
rect 222 -1800 228 -1794
rect 222 -1806 228 -1800
rect 222 -1812 228 -1806
rect 222 -1818 228 -1812
rect 222 -1824 228 -1818
rect 222 -1830 228 -1824
rect 222 -1836 228 -1830
rect 222 -1842 228 -1836
rect 222 -1848 228 -1842
rect 222 -1854 228 -1848
rect 222 -1860 228 -1854
rect 222 -1866 228 -1860
rect 222 -1872 228 -1866
rect 222 -1878 228 -1872
rect 222 -1884 228 -1878
rect 222 -1890 228 -1884
rect 222 -1896 228 -1890
rect 222 -1902 228 -1896
rect 222 -1908 228 -1902
rect 222 -1914 228 -1908
rect 222 -1920 228 -1914
rect 222 -1926 228 -1920
rect 222 -1932 228 -1926
rect 222 -1938 228 -1932
rect 222 -1944 228 -1938
rect 222 -1950 228 -1944
rect 222 -1956 228 -1950
rect 222 -1962 228 -1956
rect 222 -1968 228 -1962
rect 222 -1974 228 -1968
rect 222 -1980 228 -1974
rect 222 -1986 228 -1980
rect 222 -1992 228 -1986
rect 222 -1998 228 -1992
rect 222 -2004 228 -1998
rect 222 -2010 228 -2004
rect 222 -2016 228 -2010
rect 222 -2022 228 -2016
rect 222 -2028 228 -2022
rect 222 -2034 228 -2028
rect 222 -2040 228 -2034
rect 222 -2046 228 -2040
rect 222 -2052 228 -2046
rect 222 -2058 228 -2052
rect 222 -2064 228 -2058
rect 222 -2070 228 -2064
rect 222 -2076 228 -2070
rect 222 -2082 228 -2076
rect 222 -2088 228 -2082
rect 222 -2094 228 -2088
rect 222 -2100 228 -2094
rect 222 -2106 228 -2100
rect 222 -2112 228 -2106
rect 222 -2118 228 -2112
rect 222 -2124 228 -2118
rect 222 -2130 228 -2124
rect 222 -2136 228 -2130
rect 222 -2490 228 -2484
rect 222 -2496 228 -2490
rect 222 -2502 228 -2496
rect 222 -2508 228 -2502
rect 222 -2514 228 -2508
rect 222 -2520 228 -2514
rect 222 -2526 228 -2520
rect 222 -2532 228 -2526
rect 222 -2538 228 -2532
rect 222 -2544 228 -2538
rect 222 -2550 228 -2544
rect 222 -2556 228 -2550
rect 222 -2562 228 -2556
rect 222 -2568 228 -2562
rect 222 -2574 228 -2568
rect 222 -2580 228 -2574
rect 222 -2586 228 -2580
rect 222 -2592 228 -2586
rect 222 -2598 228 -2592
rect 222 -2604 228 -2598
rect 222 -2610 228 -2604
rect 222 -2616 228 -2610
rect 222 -2622 228 -2616
rect 222 -2628 228 -2622
rect 222 -2634 228 -2628
rect 222 -2640 228 -2634
rect 222 -2646 228 -2640
rect 222 -2652 228 -2646
rect 222 -2658 228 -2652
rect 222 -2664 228 -2658
rect 222 -2670 228 -2664
rect 222 -2676 228 -2670
rect 222 -2682 228 -2676
rect 222 -2688 228 -2682
rect 222 -2694 228 -2688
rect 222 -2700 228 -2694
rect 222 -2706 228 -2700
rect 222 -2712 228 -2706
rect 222 -2718 228 -2712
rect 222 -2724 228 -2718
rect 222 -2730 228 -2724
rect 222 -2736 228 -2730
rect 222 -2742 228 -2736
rect 222 -2748 228 -2742
rect 222 -2754 228 -2748
rect 222 -2760 228 -2754
rect 222 -2766 228 -2760
rect 222 -2772 228 -2766
rect 222 -2778 228 -2772
rect 222 -2784 228 -2778
rect 222 -2790 228 -2784
rect 222 -2796 228 -2790
rect 222 -2802 228 -2796
rect 222 -2808 228 -2802
rect 222 -2814 228 -2808
rect 222 -2820 228 -2814
rect 222 -2826 228 -2820
rect 222 -2832 228 -2826
rect 222 -2838 228 -2832
rect 222 -2844 228 -2838
rect 222 -2850 228 -2844
rect 222 -2856 228 -2850
rect 222 -2862 228 -2856
rect 222 -2868 228 -2862
rect 222 -2874 228 -2868
rect 222 -2880 228 -2874
rect 222 -2886 228 -2880
rect 222 -2892 228 -2886
rect 222 -2898 228 -2892
rect 222 -2904 228 -2898
rect 222 -2910 228 -2904
rect 222 -2916 228 -2910
rect 222 -2922 228 -2916
rect 222 -2928 228 -2922
rect 222 -2934 228 -2928
rect 222 -2940 228 -2934
rect 222 -2946 228 -2940
rect 222 -2952 228 -2946
rect 222 -2958 228 -2952
rect 222 -2964 228 -2958
rect 222 -2970 228 -2964
rect 222 -2976 228 -2970
rect 222 -2982 228 -2976
rect 222 -2988 228 -2982
rect 222 -2994 228 -2988
rect 222 -3000 228 -2994
rect 222 -3006 228 -3000
rect 222 -3012 228 -3006
rect 228 -1608 234 -1602
rect 228 -1614 234 -1608
rect 228 -1620 234 -1614
rect 228 -1626 234 -1620
rect 228 -1632 234 -1626
rect 228 -1638 234 -1632
rect 228 -1644 234 -1638
rect 228 -1650 234 -1644
rect 228 -1656 234 -1650
rect 228 -1662 234 -1656
rect 228 -1668 234 -1662
rect 228 -1674 234 -1668
rect 228 -1680 234 -1674
rect 228 -1686 234 -1680
rect 228 -1692 234 -1686
rect 228 -1698 234 -1692
rect 228 -1704 234 -1698
rect 228 -1710 234 -1704
rect 228 -1716 234 -1710
rect 228 -1722 234 -1716
rect 228 -1728 234 -1722
rect 228 -1734 234 -1728
rect 228 -1740 234 -1734
rect 228 -1746 234 -1740
rect 228 -1752 234 -1746
rect 228 -1758 234 -1752
rect 228 -1764 234 -1758
rect 228 -1770 234 -1764
rect 228 -1776 234 -1770
rect 228 -1782 234 -1776
rect 228 -1788 234 -1782
rect 228 -1794 234 -1788
rect 228 -1800 234 -1794
rect 228 -1806 234 -1800
rect 228 -1812 234 -1806
rect 228 -1818 234 -1812
rect 228 -1824 234 -1818
rect 228 -1830 234 -1824
rect 228 -1836 234 -1830
rect 228 -1842 234 -1836
rect 228 -1848 234 -1842
rect 228 -1854 234 -1848
rect 228 -1860 234 -1854
rect 228 -1866 234 -1860
rect 228 -1872 234 -1866
rect 228 -1878 234 -1872
rect 228 -1884 234 -1878
rect 228 -1890 234 -1884
rect 228 -1896 234 -1890
rect 228 -1902 234 -1896
rect 228 -1908 234 -1902
rect 228 -1914 234 -1908
rect 228 -1920 234 -1914
rect 228 -1926 234 -1920
rect 228 -1932 234 -1926
rect 228 -1938 234 -1932
rect 228 -1944 234 -1938
rect 228 -1950 234 -1944
rect 228 -1956 234 -1950
rect 228 -1962 234 -1956
rect 228 -1968 234 -1962
rect 228 -1974 234 -1968
rect 228 -1980 234 -1974
rect 228 -1986 234 -1980
rect 228 -1992 234 -1986
rect 228 -1998 234 -1992
rect 228 -2004 234 -1998
rect 228 -2010 234 -2004
rect 228 -2016 234 -2010
rect 228 -2022 234 -2016
rect 228 -2028 234 -2022
rect 228 -2034 234 -2028
rect 228 -2040 234 -2034
rect 228 -2046 234 -2040
rect 228 -2052 234 -2046
rect 228 -2058 234 -2052
rect 228 -2064 234 -2058
rect 228 -2070 234 -2064
rect 228 -2076 234 -2070
rect 228 -2082 234 -2076
rect 228 -2088 234 -2082
rect 228 -2094 234 -2088
rect 228 -2100 234 -2094
rect 228 -2106 234 -2100
rect 228 -2520 234 -2514
rect 228 -2526 234 -2520
rect 228 -2532 234 -2526
rect 228 -2538 234 -2532
rect 228 -2544 234 -2538
rect 228 -2550 234 -2544
rect 228 -2556 234 -2550
rect 228 -2562 234 -2556
rect 228 -2568 234 -2562
rect 228 -2574 234 -2568
rect 228 -2580 234 -2574
rect 228 -2586 234 -2580
rect 228 -2592 234 -2586
rect 228 -2598 234 -2592
rect 228 -2604 234 -2598
rect 228 -2610 234 -2604
rect 228 -2616 234 -2610
rect 228 -2622 234 -2616
rect 228 -2628 234 -2622
rect 228 -2634 234 -2628
rect 228 -2640 234 -2634
rect 228 -2646 234 -2640
rect 228 -2652 234 -2646
rect 228 -2658 234 -2652
rect 228 -2664 234 -2658
rect 228 -2670 234 -2664
rect 228 -2676 234 -2670
rect 228 -2682 234 -2676
rect 228 -2688 234 -2682
rect 228 -2694 234 -2688
rect 228 -2700 234 -2694
rect 228 -2706 234 -2700
rect 228 -2712 234 -2706
rect 228 -2718 234 -2712
rect 228 -2724 234 -2718
rect 228 -2730 234 -2724
rect 228 -2736 234 -2730
rect 228 -2742 234 -2736
rect 228 -2748 234 -2742
rect 228 -2754 234 -2748
rect 228 -2760 234 -2754
rect 228 -2766 234 -2760
rect 228 -2772 234 -2766
rect 228 -2778 234 -2772
rect 228 -2784 234 -2778
rect 228 -2790 234 -2784
rect 228 -2796 234 -2790
rect 228 -2802 234 -2796
rect 228 -2808 234 -2802
rect 228 -2814 234 -2808
rect 228 -2820 234 -2814
rect 228 -2826 234 -2820
rect 228 -2832 234 -2826
rect 228 -2838 234 -2832
rect 228 -2844 234 -2838
rect 228 -2850 234 -2844
rect 228 -2856 234 -2850
rect 228 -2862 234 -2856
rect 228 -2868 234 -2862
rect 228 -2874 234 -2868
rect 228 -2880 234 -2874
rect 228 -2886 234 -2880
rect 228 -2892 234 -2886
rect 228 -2898 234 -2892
rect 228 -2904 234 -2898
rect 228 -2910 234 -2904
rect 228 -2916 234 -2910
rect 228 -2922 234 -2916
rect 228 -2928 234 -2922
rect 228 -2934 234 -2928
rect 228 -2940 234 -2934
rect 228 -2946 234 -2940
rect 228 -2952 234 -2946
rect 228 -2958 234 -2952
rect 228 -2964 234 -2958
rect 228 -2970 234 -2964
rect 228 -2976 234 -2970
rect 228 -2982 234 -2976
rect 228 -2988 234 -2982
rect 228 -2994 234 -2988
rect 228 -3000 234 -2994
rect 228 -3006 234 -3000
rect 228 -3012 234 -3006
rect 228 -3018 234 -3012
rect 234 -1596 240 -1590
rect 234 -1602 240 -1596
rect 234 -1608 240 -1602
rect 234 -1614 240 -1608
rect 234 -1620 240 -1614
rect 234 -1626 240 -1620
rect 234 -1632 240 -1626
rect 234 -1638 240 -1632
rect 234 -1644 240 -1638
rect 234 -1650 240 -1644
rect 234 -1656 240 -1650
rect 234 -1662 240 -1656
rect 234 -1668 240 -1662
rect 234 -1674 240 -1668
rect 234 -1680 240 -1674
rect 234 -1686 240 -1680
rect 234 -1692 240 -1686
rect 234 -1698 240 -1692
rect 234 -1704 240 -1698
rect 234 -1710 240 -1704
rect 234 -1716 240 -1710
rect 234 -1722 240 -1716
rect 234 -1728 240 -1722
rect 234 -1734 240 -1728
rect 234 -1740 240 -1734
rect 234 -1746 240 -1740
rect 234 -1752 240 -1746
rect 234 -1758 240 -1752
rect 234 -1764 240 -1758
rect 234 -1770 240 -1764
rect 234 -1776 240 -1770
rect 234 -1782 240 -1776
rect 234 -1788 240 -1782
rect 234 -1794 240 -1788
rect 234 -1800 240 -1794
rect 234 -1806 240 -1800
rect 234 -1812 240 -1806
rect 234 -1818 240 -1812
rect 234 -1824 240 -1818
rect 234 -1830 240 -1824
rect 234 -1836 240 -1830
rect 234 -1842 240 -1836
rect 234 -1848 240 -1842
rect 234 -1854 240 -1848
rect 234 -1860 240 -1854
rect 234 -1866 240 -1860
rect 234 -1872 240 -1866
rect 234 -1878 240 -1872
rect 234 -1884 240 -1878
rect 234 -1890 240 -1884
rect 234 -1896 240 -1890
rect 234 -1902 240 -1896
rect 234 -1908 240 -1902
rect 234 -1914 240 -1908
rect 234 -1920 240 -1914
rect 234 -1926 240 -1920
rect 234 -1932 240 -1926
rect 234 -1938 240 -1932
rect 234 -1944 240 -1938
rect 234 -1950 240 -1944
rect 234 -1956 240 -1950
rect 234 -1962 240 -1956
rect 234 -1968 240 -1962
rect 234 -1974 240 -1968
rect 234 -1980 240 -1974
rect 234 -1986 240 -1980
rect 234 -1992 240 -1986
rect 234 -1998 240 -1992
rect 234 -2004 240 -1998
rect 234 -2010 240 -2004
rect 234 -2016 240 -2010
rect 234 -2022 240 -2016
rect 234 -2028 240 -2022
rect 234 -2034 240 -2028
rect 234 -2040 240 -2034
rect 234 -2046 240 -2040
rect 234 -2052 240 -2046
rect 234 -2058 240 -2052
rect 234 -2064 240 -2058
rect 234 -2070 240 -2064
rect 234 -2076 240 -2070
rect 234 -2550 240 -2544
rect 234 -2556 240 -2550
rect 234 -2562 240 -2556
rect 234 -2568 240 -2562
rect 234 -2574 240 -2568
rect 234 -2580 240 -2574
rect 234 -2586 240 -2580
rect 234 -2592 240 -2586
rect 234 -2598 240 -2592
rect 234 -2604 240 -2598
rect 234 -2610 240 -2604
rect 234 -2616 240 -2610
rect 234 -2622 240 -2616
rect 234 -2628 240 -2622
rect 234 -2634 240 -2628
rect 234 -2640 240 -2634
rect 234 -2646 240 -2640
rect 234 -2652 240 -2646
rect 234 -2658 240 -2652
rect 234 -2664 240 -2658
rect 234 -2670 240 -2664
rect 234 -2676 240 -2670
rect 234 -2682 240 -2676
rect 234 -2688 240 -2682
rect 234 -2694 240 -2688
rect 234 -2700 240 -2694
rect 234 -2706 240 -2700
rect 234 -2712 240 -2706
rect 234 -2718 240 -2712
rect 234 -2724 240 -2718
rect 234 -2730 240 -2724
rect 234 -2736 240 -2730
rect 234 -2742 240 -2736
rect 234 -2748 240 -2742
rect 234 -2754 240 -2748
rect 234 -2760 240 -2754
rect 234 -2766 240 -2760
rect 234 -2772 240 -2766
rect 234 -2778 240 -2772
rect 234 -2784 240 -2778
rect 234 -2790 240 -2784
rect 234 -2796 240 -2790
rect 234 -2802 240 -2796
rect 234 -2808 240 -2802
rect 234 -2814 240 -2808
rect 234 -2820 240 -2814
rect 234 -2826 240 -2820
rect 234 -2832 240 -2826
rect 234 -2838 240 -2832
rect 234 -2844 240 -2838
rect 234 -2850 240 -2844
rect 234 -2856 240 -2850
rect 234 -2862 240 -2856
rect 234 -2868 240 -2862
rect 234 -2874 240 -2868
rect 234 -2880 240 -2874
rect 234 -2886 240 -2880
rect 234 -2892 240 -2886
rect 234 -2898 240 -2892
rect 234 -2904 240 -2898
rect 234 -2910 240 -2904
rect 234 -2916 240 -2910
rect 234 -2922 240 -2916
rect 234 -2928 240 -2922
rect 234 -2934 240 -2928
rect 234 -2940 240 -2934
rect 234 -2946 240 -2940
rect 234 -2952 240 -2946
rect 234 -2958 240 -2952
rect 234 -2964 240 -2958
rect 234 -2970 240 -2964
rect 234 -2976 240 -2970
rect 234 -2982 240 -2976
rect 234 -2988 240 -2982
rect 234 -2994 240 -2988
rect 234 -3000 240 -2994
rect 234 -3006 240 -3000
rect 234 -3012 240 -3006
rect 234 -3018 240 -3012
rect 234 -3024 240 -3018
rect 234 -3030 240 -3024
rect 240 -1590 246 -1584
rect 240 -1596 246 -1590
rect 240 -1602 246 -1596
rect 240 -1608 246 -1602
rect 240 -1614 246 -1608
rect 240 -1620 246 -1614
rect 240 -1626 246 -1620
rect 240 -1632 246 -1626
rect 240 -1638 246 -1632
rect 240 -1644 246 -1638
rect 240 -1650 246 -1644
rect 240 -1656 246 -1650
rect 240 -1662 246 -1656
rect 240 -1668 246 -1662
rect 240 -1674 246 -1668
rect 240 -1680 246 -1674
rect 240 -1686 246 -1680
rect 240 -1692 246 -1686
rect 240 -1698 246 -1692
rect 240 -1704 246 -1698
rect 240 -1710 246 -1704
rect 240 -1716 246 -1710
rect 240 -1722 246 -1716
rect 240 -1728 246 -1722
rect 240 -1734 246 -1728
rect 240 -1740 246 -1734
rect 240 -1746 246 -1740
rect 240 -1752 246 -1746
rect 240 -1758 246 -1752
rect 240 -1764 246 -1758
rect 240 -1770 246 -1764
rect 240 -1776 246 -1770
rect 240 -1782 246 -1776
rect 240 -1788 246 -1782
rect 240 -1794 246 -1788
rect 240 -1800 246 -1794
rect 240 -1806 246 -1800
rect 240 -1812 246 -1806
rect 240 -1818 246 -1812
rect 240 -1824 246 -1818
rect 240 -1830 246 -1824
rect 240 -1836 246 -1830
rect 240 -1842 246 -1836
rect 240 -1848 246 -1842
rect 240 -1854 246 -1848
rect 240 -1860 246 -1854
rect 240 -1866 246 -1860
rect 240 -1872 246 -1866
rect 240 -1878 246 -1872
rect 240 -1884 246 -1878
rect 240 -1890 246 -1884
rect 240 -1896 246 -1890
rect 240 -1902 246 -1896
rect 240 -1908 246 -1902
rect 240 -1914 246 -1908
rect 240 -1920 246 -1914
rect 240 -1926 246 -1920
rect 240 -1932 246 -1926
rect 240 -1938 246 -1932
rect 240 -1944 246 -1938
rect 240 -1950 246 -1944
rect 240 -1956 246 -1950
rect 240 -1962 246 -1956
rect 240 -1968 246 -1962
rect 240 -1974 246 -1968
rect 240 -1980 246 -1974
rect 240 -1986 246 -1980
rect 240 -1992 246 -1986
rect 240 -1998 246 -1992
rect 240 -2004 246 -1998
rect 240 -2010 246 -2004
rect 240 -2016 246 -2010
rect 240 -2022 246 -2016
rect 240 -2028 246 -2022
rect 240 -2034 246 -2028
rect 240 -2040 246 -2034
rect 240 -2046 246 -2040
rect 240 -2052 246 -2046
rect 240 -2574 246 -2568
rect 240 -2580 246 -2574
rect 240 -2586 246 -2580
rect 240 -2592 246 -2586
rect 240 -2598 246 -2592
rect 240 -2604 246 -2598
rect 240 -2610 246 -2604
rect 240 -2616 246 -2610
rect 240 -2622 246 -2616
rect 240 -2628 246 -2622
rect 240 -2634 246 -2628
rect 240 -2640 246 -2634
rect 240 -2646 246 -2640
rect 240 -2652 246 -2646
rect 240 -2658 246 -2652
rect 240 -2664 246 -2658
rect 240 -2670 246 -2664
rect 240 -2676 246 -2670
rect 240 -2682 246 -2676
rect 240 -2688 246 -2682
rect 240 -2694 246 -2688
rect 240 -2700 246 -2694
rect 240 -2706 246 -2700
rect 240 -2712 246 -2706
rect 240 -2718 246 -2712
rect 240 -2724 246 -2718
rect 240 -2730 246 -2724
rect 240 -2736 246 -2730
rect 240 -2742 246 -2736
rect 240 -2748 246 -2742
rect 240 -2754 246 -2748
rect 240 -2760 246 -2754
rect 240 -2766 246 -2760
rect 240 -2772 246 -2766
rect 240 -2778 246 -2772
rect 240 -2784 246 -2778
rect 240 -2790 246 -2784
rect 240 -2796 246 -2790
rect 240 -2802 246 -2796
rect 240 -2808 246 -2802
rect 240 -2814 246 -2808
rect 240 -2820 246 -2814
rect 240 -2826 246 -2820
rect 240 -2832 246 -2826
rect 240 -2838 246 -2832
rect 240 -2844 246 -2838
rect 240 -2850 246 -2844
rect 240 -2856 246 -2850
rect 240 -2862 246 -2856
rect 240 -2868 246 -2862
rect 240 -2874 246 -2868
rect 240 -2880 246 -2874
rect 240 -2886 246 -2880
rect 240 -2892 246 -2886
rect 240 -2898 246 -2892
rect 240 -2904 246 -2898
rect 240 -2910 246 -2904
rect 240 -2916 246 -2910
rect 240 -2922 246 -2916
rect 240 -2928 246 -2922
rect 240 -2934 246 -2928
rect 240 -2940 246 -2934
rect 240 -2946 246 -2940
rect 240 -2952 246 -2946
rect 240 -2958 246 -2952
rect 240 -2964 246 -2958
rect 240 -2970 246 -2964
rect 240 -2976 246 -2970
rect 240 -2982 246 -2976
rect 240 -2988 246 -2982
rect 240 -2994 246 -2988
rect 240 -3000 246 -2994
rect 240 -3006 246 -3000
rect 240 -3012 246 -3006
rect 240 -3018 246 -3012
rect 240 -3024 246 -3018
rect 240 -3030 246 -3024
rect 240 -3036 246 -3030
rect 246 -1584 252 -1578
rect 246 -1590 252 -1584
rect 246 -1596 252 -1590
rect 246 -1602 252 -1596
rect 246 -1608 252 -1602
rect 246 -1614 252 -1608
rect 246 -1620 252 -1614
rect 246 -1626 252 -1620
rect 246 -1632 252 -1626
rect 246 -1638 252 -1632
rect 246 -1644 252 -1638
rect 246 -1650 252 -1644
rect 246 -1656 252 -1650
rect 246 -1662 252 -1656
rect 246 -1668 252 -1662
rect 246 -1674 252 -1668
rect 246 -1680 252 -1674
rect 246 -1686 252 -1680
rect 246 -1692 252 -1686
rect 246 -1698 252 -1692
rect 246 -1704 252 -1698
rect 246 -1710 252 -1704
rect 246 -1716 252 -1710
rect 246 -1722 252 -1716
rect 246 -1728 252 -1722
rect 246 -1734 252 -1728
rect 246 -1740 252 -1734
rect 246 -1746 252 -1740
rect 246 -1752 252 -1746
rect 246 -1758 252 -1752
rect 246 -1764 252 -1758
rect 246 -1770 252 -1764
rect 246 -1776 252 -1770
rect 246 -1782 252 -1776
rect 246 -1788 252 -1782
rect 246 -1794 252 -1788
rect 246 -1800 252 -1794
rect 246 -1806 252 -1800
rect 246 -1812 252 -1806
rect 246 -1818 252 -1812
rect 246 -1824 252 -1818
rect 246 -1830 252 -1824
rect 246 -1836 252 -1830
rect 246 -1842 252 -1836
rect 246 -1848 252 -1842
rect 246 -1854 252 -1848
rect 246 -1860 252 -1854
rect 246 -1866 252 -1860
rect 246 -1872 252 -1866
rect 246 -1878 252 -1872
rect 246 -1884 252 -1878
rect 246 -1890 252 -1884
rect 246 -1896 252 -1890
rect 246 -1902 252 -1896
rect 246 -1908 252 -1902
rect 246 -1914 252 -1908
rect 246 -1920 252 -1914
rect 246 -1926 252 -1920
rect 246 -1932 252 -1926
rect 246 -1938 252 -1932
rect 246 -1944 252 -1938
rect 246 -1950 252 -1944
rect 246 -1956 252 -1950
rect 246 -1962 252 -1956
rect 246 -1968 252 -1962
rect 246 -1974 252 -1968
rect 246 -1980 252 -1974
rect 246 -1986 252 -1980
rect 246 -1992 252 -1986
rect 246 -1998 252 -1992
rect 246 -2004 252 -1998
rect 246 -2010 252 -2004
rect 246 -2016 252 -2010
rect 246 -2022 252 -2016
rect 246 -2028 252 -2022
rect 246 -2034 252 -2028
rect 246 -2592 252 -2586
rect 246 -2598 252 -2592
rect 246 -2604 252 -2598
rect 246 -2610 252 -2604
rect 246 -2616 252 -2610
rect 246 -2622 252 -2616
rect 246 -2628 252 -2622
rect 246 -2634 252 -2628
rect 246 -2640 252 -2634
rect 246 -2646 252 -2640
rect 246 -2652 252 -2646
rect 246 -2658 252 -2652
rect 246 -2664 252 -2658
rect 246 -2670 252 -2664
rect 246 -2676 252 -2670
rect 246 -2682 252 -2676
rect 246 -2688 252 -2682
rect 246 -2694 252 -2688
rect 246 -2700 252 -2694
rect 246 -2706 252 -2700
rect 246 -2712 252 -2706
rect 246 -2718 252 -2712
rect 246 -2724 252 -2718
rect 246 -2730 252 -2724
rect 246 -2736 252 -2730
rect 246 -2742 252 -2736
rect 246 -2748 252 -2742
rect 246 -2754 252 -2748
rect 246 -2760 252 -2754
rect 246 -2766 252 -2760
rect 246 -2772 252 -2766
rect 246 -2778 252 -2772
rect 246 -2784 252 -2778
rect 246 -2790 252 -2784
rect 246 -2796 252 -2790
rect 246 -2802 252 -2796
rect 246 -2808 252 -2802
rect 246 -2814 252 -2808
rect 246 -2820 252 -2814
rect 246 -2826 252 -2820
rect 246 -2832 252 -2826
rect 246 -2838 252 -2832
rect 246 -2844 252 -2838
rect 246 -2850 252 -2844
rect 246 -2856 252 -2850
rect 246 -2862 252 -2856
rect 246 -2868 252 -2862
rect 246 -2874 252 -2868
rect 246 -2880 252 -2874
rect 246 -2886 252 -2880
rect 246 -2892 252 -2886
rect 246 -2898 252 -2892
rect 246 -2904 252 -2898
rect 246 -2910 252 -2904
rect 246 -2916 252 -2910
rect 246 -2922 252 -2916
rect 246 -2928 252 -2922
rect 246 -2934 252 -2928
rect 246 -2940 252 -2934
rect 246 -2946 252 -2940
rect 246 -2952 252 -2946
rect 246 -2958 252 -2952
rect 246 -2964 252 -2958
rect 246 -2970 252 -2964
rect 246 -2976 252 -2970
rect 246 -2982 252 -2976
rect 246 -2988 252 -2982
rect 246 -2994 252 -2988
rect 246 -3000 252 -2994
rect 246 -3006 252 -3000
rect 246 -3012 252 -3006
rect 246 -3018 252 -3012
rect 246 -3024 252 -3018
rect 246 -3030 252 -3024
rect 246 -3036 252 -3030
rect 246 -3042 252 -3036
rect 252 -1572 258 -1566
rect 252 -1578 258 -1572
rect 252 -1584 258 -1578
rect 252 -1590 258 -1584
rect 252 -1596 258 -1590
rect 252 -1602 258 -1596
rect 252 -1608 258 -1602
rect 252 -1614 258 -1608
rect 252 -1620 258 -1614
rect 252 -1626 258 -1620
rect 252 -1632 258 -1626
rect 252 -1638 258 -1632
rect 252 -1644 258 -1638
rect 252 -1650 258 -1644
rect 252 -1656 258 -1650
rect 252 -1662 258 -1656
rect 252 -1668 258 -1662
rect 252 -1674 258 -1668
rect 252 -1680 258 -1674
rect 252 -1686 258 -1680
rect 252 -1692 258 -1686
rect 252 -1698 258 -1692
rect 252 -1704 258 -1698
rect 252 -1710 258 -1704
rect 252 -1716 258 -1710
rect 252 -1722 258 -1716
rect 252 -1728 258 -1722
rect 252 -1734 258 -1728
rect 252 -1740 258 -1734
rect 252 -1746 258 -1740
rect 252 -1752 258 -1746
rect 252 -1758 258 -1752
rect 252 -1764 258 -1758
rect 252 -1770 258 -1764
rect 252 -1776 258 -1770
rect 252 -1782 258 -1776
rect 252 -1788 258 -1782
rect 252 -1794 258 -1788
rect 252 -1800 258 -1794
rect 252 -1806 258 -1800
rect 252 -1812 258 -1806
rect 252 -1818 258 -1812
rect 252 -1824 258 -1818
rect 252 -1830 258 -1824
rect 252 -1836 258 -1830
rect 252 -1842 258 -1836
rect 252 -1848 258 -1842
rect 252 -1854 258 -1848
rect 252 -1860 258 -1854
rect 252 -1866 258 -1860
rect 252 -1872 258 -1866
rect 252 -1878 258 -1872
rect 252 -1884 258 -1878
rect 252 -1890 258 -1884
rect 252 -1896 258 -1890
rect 252 -1902 258 -1896
rect 252 -1908 258 -1902
rect 252 -1914 258 -1908
rect 252 -1920 258 -1914
rect 252 -1926 258 -1920
rect 252 -1932 258 -1926
rect 252 -1938 258 -1932
rect 252 -1944 258 -1938
rect 252 -1950 258 -1944
rect 252 -1956 258 -1950
rect 252 -1962 258 -1956
rect 252 -1968 258 -1962
rect 252 -1974 258 -1968
rect 252 -1980 258 -1974
rect 252 -1986 258 -1980
rect 252 -1992 258 -1986
rect 252 -1998 258 -1992
rect 252 -2004 258 -1998
rect 252 -2010 258 -2004
rect 252 -2616 258 -2610
rect 252 -2622 258 -2616
rect 252 -2628 258 -2622
rect 252 -2634 258 -2628
rect 252 -2640 258 -2634
rect 252 -2646 258 -2640
rect 252 -2652 258 -2646
rect 252 -2658 258 -2652
rect 252 -2664 258 -2658
rect 252 -2670 258 -2664
rect 252 -2676 258 -2670
rect 252 -2682 258 -2676
rect 252 -2688 258 -2682
rect 252 -2694 258 -2688
rect 252 -2700 258 -2694
rect 252 -2706 258 -2700
rect 252 -2712 258 -2706
rect 252 -2718 258 -2712
rect 252 -2724 258 -2718
rect 252 -2730 258 -2724
rect 252 -2736 258 -2730
rect 252 -2742 258 -2736
rect 252 -2748 258 -2742
rect 252 -2754 258 -2748
rect 252 -2760 258 -2754
rect 252 -2766 258 -2760
rect 252 -2772 258 -2766
rect 252 -2778 258 -2772
rect 252 -2784 258 -2778
rect 252 -2790 258 -2784
rect 252 -2796 258 -2790
rect 252 -2802 258 -2796
rect 252 -2808 258 -2802
rect 252 -2814 258 -2808
rect 252 -2820 258 -2814
rect 252 -2826 258 -2820
rect 252 -2832 258 -2826
rect 252 -2838 258 -2832
rect 252 -2844 258 -2838
rect 252 -2850 258 -2844
rect 252 -2856 258 -2850
rect 252 -2862 258 -2856
rect 252 -2868 258 -2862
rect 252 -2874 258 -2868
rect 252 -2880 258 -2874
rect 252 -2886 258 -2880
rect 252 -2892 258 -2886
rect 252 -2898 258 -2892
rect 252 -2904 258 -2898
rect 252 -2910 258 -2904
rect 252 -2916 258 -2910
rect 252 -2922 258 -2916
rect 252 -2928 258 -2922
rect 252 -2934 258 -2928
rect 252 -2940 258 -2934
rect 252 -2946 258 -2940
rect 252 -2952 258 -2946
rect 252 -2958 258 -2952
rect 252 -2964 258 -2958
rect 252 -2970 258 -2964
rect 252 -2976 258 -2970
rect 252 -2982 258 -2976
rect 252 -2988 258 -2982
rect 252 -2994 258 -2988
rect 252 -3000 258 -2994
rect 252 -3006 258 -3000
rect 252 -3012 258 -3006
rect 252 -3018 258 -3012
rect 252 -3024 258 -3018
rect 252 -3030 258 -3024
rect 252 -3036 258 -3030
rect 252 -3042 258 -3036
rect 252 -3048 258 -3042
rect 252 -3054 258 -3048
rect 258 -1566 264 -1560
rect 258 -1572 264 -1566
rect 258 -1578 264 -1572
rect 258 -1584 264 -1578
rect 258 -1590 264 -1584
rect 258 -1596 264 -1590
rect 258 -1602 264 -1596
rect 258 -1608 264 -1602
rect 258 -1614 264 -1608
rect 258 -1620 264 -1614
rect 258 -1626 264 -1620
rect 258 -1632 264 -1626
rect 258 -1638 264 -1632
rect 258 -1644 264 -1638
rect 258 -1650 264 -1644
rect 258 -1656 264 -1650
rect 258 -1662 264 -1656
rect 258 -1668 264 -1662
rect 258 -1674 264 -1668
rect 258 -1680 264 -1674
rect 258 -1686 264 -1680
rect 258 -1692 264 -1686
rect 258 -1698 264 -1692
rect 258 -1704 264 -1698
rect 258 -1710 264 -1704
rect 258 -1716 264 -1710
rect 258 -1722 264 -1716
rect 258 -1728 264 -1722
rect 258 -1734 264 -1728
rect 258 -1740 264 -1734
rect 258 -1746 264 -1740
rect 258 -1752 264 -1746
rect 258 -1758 264 -1752
rect 258 -1764 264 -1758
rect 258 -1770 264 -1764
rect 258 -1776 264 -1770
rect 258 -1782 264 -1776
rect 258 -1788 264 -1782
rect 258 -1794 264 -1788
rect 258 -1800 264 -1794
rect 258 -1806 264 -1800
rect 258 -1812 264 -1806
rect 258 -1818 264 -1812
rect 258 -1824 264 -1818
rect 258 -1830 264 -1824
rect 258 -1836 264 -1830
rect 258 -1842 264 -1836
rect 258 -1848 264 -1842
rect 258 -1854 264 -1848
rect 258 -1860 264 -1854
rect 258 -1866 264 -1860
rect 258 -1872 264 -1866
rect 258 -1878 264 -1872
rect 258 -1884 264 -1878
rect 258 -1890 264 -1884
rect 258 -1896 264 -1890
rect 258 -1902 264 -1896
rect 258 -1908 264 -1902
rect 258 -1914 264 -1908
rect 258 -1920 264 -1914
rect 258 -1926 264 -1920
rect 258 -1932 264 -1926
rect 258 -1938 264 -1932
rect 258 -1944 264 -1938
rect 258 -1950 264 -1944
rect 258 -1956 264 -1950
rect 258 -1962 264 -1956
rect 258 -1968 264 -1962
rect 258 -1974 264 -1968
rect 258 -1980 264 -1974
rect 258 -1986 264 -1980
rect 258 -1992 264 -1986
rect 258 -2634 264 -2628
rect 258 -2640 264 -2634
rect 258 -2646 264 -2640
rect 258 -2652 264 -2646
rect 258 -2658 264 -2652
rect 258 -2664 264 -2658
rect 258 -2670 264 -2664
rect 258 -2676 264 -2670
rect 258 -2682 264 -2676
rect 258 -2688 264 -2682
rect 258 -2694 264 -2688
rect 258 -2700 264 -2694
rect 258 -2706 264 -2700
rect 258 -2712 264 -2706
rect 258 -2718 264 -2712
rect 258 -2724 264 -2718
rect 258 -2730 264 -2724
rect 258 -2736 264 -2730
rect 258 -2742 264 -2736
rect 258 -2748 264 -2742
rect 258 -2754 264 -2748
rect 258 -2760 264 -2754
rect 258 -2766 264 -2760
rect 258 -2772 264 -2766
rect 258 -2778 264 -2772
rect 258 -2784 264 -2778
rect 258 -2790 264 -2784
rect 258 -2796 264 -2790
rect 258 -2802 264 -2796
rect 258 -2808 264 -2802
rect 258 -2814 264 -2808
rect 258 -2820 264 -2814
rect 258 -2826 264 -2820
rect 258 -2832 264 -2826
rect 258 -2838 264 -2832
rect 258 -2844 264 -2838
rect 258 -2850 264 -2844
rect 258 -2856 264 -2850
rect 258 -2862 264 -2856
rect 258 -2868 264 -2862
rect 258 -2874 264 -2868
rect 258 -2880 264 -2874
rect 258 -2886 264 -2880
rect 258 -2892 264 -2886
rect 258 -2898 264 -2892
rect 258 -2904 264 -2898
rect 258 -2910 264 -2904
rect 258 -2916 264 -2910
rect 258 -2922 264 -2916
rect 258 -2928 264 -2922
rect 258 -2934 264 -2928
rect 258 -2940 264 -2934
rect 258 -2946 264 -2940
rect 258 -2952 264 -2946
rect 258 -2958 264 -2952
rect 258 -2964 264 -2958
rect 258 -2970 264 -2964
rect 258 -2976 264 -2970
rect 258 -2982 264 -2976
rect 258 -2988 264 -2982
rect 258 -2994 264 -2988
rect 258 -3000 264 -2994
rect 258 -3006 264 -3000
rect 258 -3012 264 -3006
rect 258 -3018 264 -3012
rect 258 -3024 264 -3018
rect 258 -3030 264 -3024
rect 258 -3036 264 -3030
rect 258 -3042 264 -3036
rect 258 -3048 264 -3042
rect 258 -3054 264 -3048
rect 258 -3060 264 -3054
rect 264 -1560 270 -1554
rect 264 -1566 270 -1560
rect 264 -1572 270 -1566
rect 264 -1578 270 -1572
rect 264 -1584 270 -1578
rect 264 -1590 270 -1584
rect 264 -1596 270 -1590
rect 264 -1602 270 -1596
rect 264 -1608 270 -1602
rect 264 -1614 270 -1608
rect 264 -1620 270 -1614
rect 264 -1626 270 -1620
rect 264 -1632 270 -1626
rect 264 -1638 270 -1632
rect 264 -1644 270 -1638
rect 264 -1650 270 -1644
rect 264 -1656 270 -1650
rect 264 -1662 270 -1656
rect 264 -1668 270 -1662
rect 264 -1674 270 -1668
rect 264 -1680 270 -1674
rect 264 -1686 270 -1680
rect 264 -1692 270 -1686
rect 264 -1698 270 -1692
rect 264 -1704 270 -1698
rect 264 -1710 270 -1704
rect 264 -1716 270 -1710
rect 264 -1722 270 -1716
rect 264 -1728 270 -1722
rect 264 -1734 270 -1728
rect 264 -1740 270 -1734
rect 264 -1746 270 -1740
rect 264 -1752 270 -1746
rect 264 -1758 270 -1752
rect 264 -1764 270 -1758
rect 264 -1770 270 -1764
rect 264 -1776 270 -1770
rect 264 -1782 270 -1776
rect 264 -1788 270 -1782
rect 264 -1794 270 -1788
rect 264 -1800 270 -1794
rect 264 -1806 270 -1800
rect 264 -1812 270 -1806
rect 264 -1818 270 -1812
rect 264 -1824 270 -1818
rect 264 -1830 270 -1824
rect 264 -1836 270 -1830
rect 264 -1842 270 -1836
rect 264 -1848 270 -1842
rect 264 -1854 270 -1848
rect 264 -1860 270 -1854
rect 264 -1866 270 -1860
rect 264 -1872 270 -1866
rect 264 -1878 270 -1872
rect 264 -1884 270 -1878
rect 264 -1890 270 -1884
rect 264 -1896 270 -1890
rect 264 -1902 270 -1896
rect 264 -1908 270 -1902
rect 264 -1914 270 -1908
rect 264 -1920 270 -1914
rect 264 -1926 270 -1920
rect 264 -1932 270 -1926
rect 264 -1938 270 -1932
rect 264 -1944 270 -1938
rect 264 -1950 270 -1944
rect 264 -1956 270 -1950
rect 264 -1962 270 -1956
rect 264 -1968 270 -1962
rect 264 -1974 270 -1968
rect 264 -2652 270 -2646
rect 264 -2658 270 -2652
rect 264 -2664 270 -2658
rect 264 -2670 270 -2664
rect 264 -2676 270 -2670
rect 264 -2682 270 -2676
rect 264 -2688 270 -2682
rect 264 -2694 270 -2688
rect 264 -2700 270 -2694
rect 264 -2706 270 -2700
rect 264 -2712 270 -2706
rect 264 -2718 270 -2712
rect 264 -2724 270 -2718
rect 264 -2730 270 -2724
rect 264 -2736 270 -2730
rect 264 -2742 270 -2736
rect 264 -2748 270 -2742
rect 264 -2754 270 -2748
rect 264 -2760 270 -2754
rect 264 -2766 270 -2760
rect 264 -2772 270 -2766
rect 264 -2778 270 -2772
rect 264 -2784 270 -2778
rect 264 -2790 270 -2784
rect 264 -2796 270 -2790
rect 264 -2802 270 -2796
rect 264 -2808 270 -2802
rect 264 -2814 270 -2808
rect 264 -2820 270 -2814
rect 264 -2826 270 -2820
rect 264 -2832 270 -2826
rect 264 -2838 270 -2832
rect 264 -2844 270 -2838
rect 264 -2850 270 -2844
rect 264 -2856 270 -2850
rect 264 -2862 270 -2856
rect 264 -2868 270 -2862
rect 264 -2874 270 -2868
rect 264 -2880 270 -2874
rect 264 -2886 270 -2880
rect 264 -2892 270 -2886
rect 264 -2898 270 -2892
rect 264 -2904 270 -2898
rect 264 -2910 270 -2904
rect 264 -2916 270 -2910
rect 264 -2922 270 -2916
rect 264 -2928 270 -2922
rect 264 -2934 270 -2928
rect 264 -2940 270 -2934
rect 264 -2946 270 -2940
rect 264 -2952 270 -2946
rect 264 -2958 270 -2952
rect 264 -2964 270 -2958
rect 264 -2970 270 -2964
rect 264 -2976 270 -2970
rect 264 -2982 270 -2976
rect 264 -2988 270 -2982
rect 264 -2994 270 -2988
rect 264 -3000 270 -2994
rect 264 -3006 270 -3000
rect 264 -3012 270 -3006
rect 264 -3018 270 -3012
rect 264 -3024 270 -3018
rect 264 -3030 270 -3024
rect 264 -3036 270 -3030
rect 264 -3042 270 -3036
rect 264 -3048 270 -3042
rect 264 -3054 270 -3048
rect 264 -3060 270 -3054
rect 264 -3066 270 -3060
rect 270 -1554 276 -1548
rect 270 -1560 276 -1554
rect 270 -1566 276 -1560
rect 270 -1572 276 -1566
rect 270 -1578 276 -1572
rect 270 -1584 276 -1578
rect 270 -1590 276 -1584
rect 270 -1596 276 -1590
rect 270 -1602 276 -1596
rect 270 -1608 276 -1602
rect 270 -1614 276 -1608
rect 270 -1620 276 -1614
rect 270 -1626 276 -1620
rect 270 -1632 276 -1626
rect 270 -1638 276 -1632
rect 270 -1644 276 -1638
rect 270 -1650 276 -1644
rect 270 -1656 276 -1650
rect 270 -1662 276 -1656
rect 270 -1668 276 -1662
rect 270 -1674 276 -1668
rect 270 -1680 276 -1674
rect 270 -1686 276 -1680
rect 270 -1692 276 -1686
rect 270 -1698 276 -1692
rect 270 -1704 276 -1698
rect 270 -1710 276 -1704
rect 270 -1716 276 -1710
rect 270 -1722 276 -1716
rect 270 -1728 276 -1722
rect 270 -1734 276 -1728
rect 270 -1740 276 -1734
rect 270 -1746 276 -1740
rect 270 -1752 276 -1746
rect 270 -1758 276 -1752
rect 270 -1764 276 -1758
rect 270 -1770 276 -1764
rect 270 -1776 276 -1770
rect 270 -1782 276 -1776
rect 270 -1788 276 -1782
rect 270 -1794 276 -1788
rect 270 -1800 276 -1794
rect 270 -1806 276 -1800
rect 270 -1812 276 -1806
rect 270 -1818 276 -1812
rect 270 -1824 276 -1818
rect 270 -1830 276 -1824
rect 270 -1836 276 -1830
rect 270 -1842 276 -1836
rect 270 -1848 276 -1842
rect 270 -1854 276 -1848
rect 270 -1860 276 -1854
rect 270 -1866 276 -1860
rect 270 -1872 276 -1866
rect 270 -1878 276 -1872
rect 270 -1884 276 -1878
rect 270 -1890 276 -1884
rect 270 -1896 276 -1890
rect 270 -1902 276 -1896
rect 270 -1908 276 -1902
rect 270 -1914 276 -1908
rect 270 -1920 276 -1914
rect 270 -1926 276 -1920
rect 270 -1932 276 -1926
rect 270 -1938 276 -1932
rect 270 -1944 276 -1938
rect 270 -1950 276 -1944
rect 270 -1956 276 -1950
rect 270 -1962 276 -1956
rect 270 -2664 276 -2658
rect 270 -2670 276 -2664
rect 270 -2676 276 -2670
rect 270 -2682 276 -2676
rect 270 -2688 276 -2682
rect 270 -2694 276 -2688
rect 270 -2700 276 -2694
rect 270 -2706 276 -2700
rect 270 -2712 276 -2706
rect 270 -2718 276 -2712
rect 270 -2724 276 -2718
rect 270 -2730 276 -2724
rect 270 -2736 276 -2730
rect 270 -2742 276 -2736
rect 270 -2748 276 -2742
rect 270 -2754 276 -2748
rect 270 -2760 276 -2754
rect 270 -2766 276 -2760
rect 270 -2772 276 -2766
rect 270 -2778 276 -2772
rect 270 -2784 276 -2778
rect 270 -2790 276 -2784
rect 270 -2796 276 -2790
rect 270 -2802 276 -2796
rect 270 -2808 276 -2802
rect 270 -2814 276 -2808
rect 270 -2820 276 -2814
rect 270 -2826 276 -2820
rect 270 -2832 276 -2826
rect 270 -2838 276 -2832
rect 270 -2844 276 -2838
rect 270 -2850 276 -2844
rect 270 -2856 276 -2850
rect 270 -2862 276 -2856
rect 270 -2868 276 -2862
rect 270 -2874 276 -2868
rect 270 -2880 276 -2874
rect 270 -2886 276 -2880
rect 270 -2892 276 -2886
rect 270 -2898 276 -2892
rect 270 -2904 276 -2898
rect 270 -2910 276 -2904
rect 270 -2916 276 -2910
rect 270 -2922 276 -2916
rect 270 -2928 276 -2922
rect 270 -2934 276 -2928
rect 270 -2940 276 -2934
rect 270 -2946 276 -2940
rect 270 -2952 276 -2946
rect 270 -2958 276 -2952
rect 270 -2964 276 -2958
rect 270 -2970 276 -2964
rect 270 -2976 276 -2970
rect 270 -2982 276 -2976
rect 270 -2988 276 -2982
rect 270 -2994 276 -2988
rect 270 -3000 276 -2994
rect 270 -3006 276 -3000
rect 270 -3012 276 -3006
rect 270 -3018 276 -3012
rect 270 -3024 276 -3018
rect 270 -3030 276 -3024
rect 270 -3036 276 -3030
rect 270 -3042 276 -3036
rect 270 -3048 276 -3042
rect 270 -3054 276 -3048
rect 270 -3060 276 -3054
rect 270 -3066 276 -3060
rect 270 -3072 276 -3066
rect 270 -3078 276 -3072
rect 276 -1542 282 -1536
rect 276 -1548 282 -1542
rect 276 -1554 282 -1548
rect 276 -1560 282 -1554
rect 276 -1566 282 -1560
rect 276 -1572 282 -1566
rect 276 -1578 282 -1572
rect 276 -1584 282 -1578
rect 276 -1590 282 -1584
rect 276 -1596 282 -1590
rect 276 -1602 282 -1596
rect 276 -1608 282 -1602
rect 276 -1614 282 -1608
rect 276 -1620 282 -1614
rect 276 -1626 282 -1620
rect 276 -1632 282 -1626
rect 276 -1638 282 -1632
rect 276 -1644 282 -1638
rect 276 -1650 282 -1644
rect 276 -1656 282 -1650
rect 276 -1662 282 -1656
rect 276 -1668 282 -1662
rect 276 -1674 282 -1668
rect 276 -1680 282 -1674
rect 276 -1686 282 -1680
rect 276 -1692 282 -1686
rect 276 -1698 282 -1692
rect 276 -1704 282 -1698
rect 276 -1710 282 -1704
rect 276 -1716 282 -1710
rect 276 -1722 282 -1716
rect 276 -1728 282 -1722
rect 276 -1734 282 -1728
rect 276 -1740 282 -1734
rect 276 -1746 282 -1740
rect 276 -1752 282 -1746
rect 276 -1758 282 -1752
rect 276 -1764 282 -1758
rect 276 -1770 282 -1764
rect 276 -1776 282 -1770
rect 276 -1782 282 -1776
rect 276 -1788 282 -1782
rect 276 -1794 282 -1788
rect 276 -1800 282 -1794
rect 276 -1806 282 -1800
rect 276 -1812 282 -1806
rect 276 -1818 282 -1812
rect 276 -1824 282 -1818
rect 276 -1830 282 -1824
rect 276 -1836 282 -1830
rect 276 -1842 282 -1836
rect 276 -1848 282 -1842
rect 276 -1854 282 -1848
rect 276 -1860 282 -1854
rect 276 -1866 282 -1860
rect 276 -1872 282 -1866
rect 276 -1878 282 -1872
rect 276 -1884 282 -1878
rect 276 -1890 282 -1884
rect 276 -1896 282 -1890
rect 276 -1902 282 -1896
rect 276 -1908 282 -1902
rect 276 -1914 282 -1908
rect 276 -1920 282 -1914
rect 276 -1926 282 -1920
rect 276 -1932 282 -1926
rect 276 -1938 282 -1932
rect 276 -1944 282 -1938
rect 276 -2682 282 -2676
rect 276 -2688 282 -2682
rect 276 -2694 282 -2688
rect 276 -2700 282 -2694
rect 276 -2706 282 -2700
rect 276 -2712 282 -2706
rect 276 -2718 282 -2712
rect 276 -2724 282 -2718
rect 276 -2730 282 -2724
rect 276 -2736 282 -2730
rect 276 -2742 282 -2736
rect 276 -2748 282 -2742
rect 276 -2754 282 -2748
rect 276 -2760 282 -2754
rect 276 -2766 282 -2760
rect 276 -2772 282 -2766
rect 276 -2778 282 -2772
rect 276 -2784 282 -2778
rect 276 -2790 282 -2784
rect 276 -2796 282 -2790
rect 276 -2802 282 -2796
rect 276 -2808 282 -2802
rect 276 -2814 282 -2808
rect 276 -2820 282 -2814
rect 276 -2826 282 -2820
rect 276 -2832 282 -2826
rect 276 -2838 282 -2832
rect 276 -2844 282 -2838
rect 276 -2850 282 -2844
rect 276 -2856 282 -2850
rect 276 -2862 282 -2856
rect 276 -2868 282 -2862
rect 276 -2874 282 -2868
rect 276 -2880 282 -2874
rect 276 -2886 282 -2880
rect 276 -2892 282 -2886
rect 276 -2898 282 -2892
rect 276 -2904 282 -2898
rect 276 -2910 282 -2904
rect 276 -2916 282 -2910
rect 276 -2922 282 -2916
rect 276 -2928 282 -2922
rect 276 -2934 282 -2928
rect 276 -2940 282 -2934
rect 276 -2946 282 -2940
rect 276 -2952 282 -2946
rect 276 -2958 282 -2952
rect 276 -2964 282 -2958
rect 276 -2970 282 -2964
rect 276 -2976 282 -2970
rect 276 -2982 282 -2976
rect 276 -2988 282 -2982
rect 276 -2994 282 -2988
rect 276 -3000 282 -2994
rect 276 -3006 282 -3000
rect 276 -3012 282 -3006
rect 276 -3018 282 -3012
rect 276 -3024 282 -3018
rect 276 -3030 282 -3024
rect 276 -3036 282 -3030
rect 276 -3042 282 -3036
rect 276 -3048 282 -3042
rect 276 -3054 282 -3048
rect 276 -3060 282 -3054
rect 276 -3066 282 -3060
rect 276 -3072 282 -3066
rect 276 -3078 282 -3072
rect 276 -3084 282 -3078
rect 282 -1536 288 -1530
rect 282 -1542 288 -1536
rect 282 -1548 288 -1542
rect 282 -1554 288 -1548
rect 282 -1560 288 -1554
rect 282 -1566 288 -1560
rect 282 -1572 288 -1566
rect 282 -1578 288 -1572
rect 282 -1584 288 -1578
rect 282 -1590 288 -1584
rect 282 -1596 288 -1590
rect 282 -1602 288 -1596
rect 282 -1608 288 -1602
rect 282 -1614 288 -1608
rect 282 -1620 288 -1614
rect 282 -1626 288 -1620
rect 282 -1632 288 -1626
rect 282 -1638 288 -1632
rect 282 -1644 288 -1638
rect 282 -1650 288 -1644
rect 282 -1656 288 -1650
rect 282 -1662 288 -1656
rect 282 -1668 288 -1662
rect 282 -1674 288 -1668
rect 282 -1680 288 -1674
rect 282 -1686 288 -1680
rect 282 -1692 288 -1686
rect 282 -1698 288 -1692
rect 282 -1704 288 -1698
rect 282 -1710 288 -1704
rect 282 -1716 288 -1710
rect 282 -1722 288 -1716
rect 282 -1728 288 -1722
rect 282 -1734 288 -1728
rect 282 -1740 288 -1734
rect 282 -1746 288 -1740
rect 282 -1752 288 -1746
rect 282 -1758 288 -1752
rect 282 -1764 288 -1758
rect 282 -1770 288 -1764
rect 282 -1776 288 -1770
rect 282 -1782 288 -1776
rect 282 -1788 288 -1782
rect 282 -1794 288 -1788
rect 282 -1800 288 -1794
rect 282 -1806 288 -1800
rect 282 -1812 288 -1806
rect 282 -1818 288 -1812
rect 282 -1824 288 -1818
rect 282 -1830 288 -1824
rect 282 -1836 288 -1830
rect 282 -1842 288 -1836
rect 282 -1848 288 -1842
rect 282 -1854 288 -1848
rect 282 -1860 288 -1854
rect 282 -1866 288 -1860
rect 282 -1872 288 -1866
rect 282 -1878 288 -1872
rect 282 -1884 288 -1878
rect 282 -1890 288 -1884
rect 282 -1896 288 -1890
rect 282 -1902 288 -1896
rect 282 -1908 288 -1902
rect 282 -1914 288 -1908
rect 282 -1920 288 -1914
rect 282 -1926 288 -1920
rect 282 -2700 288 -2694
rect 282 -2706 288 -2700
rect 282 -2712 288 -2706
rect 282 -2718 288 -2712
rect 282 -2724 288 -2718
rect 282 -2730 288 -2724
rect 282 -2736 288 -2730
rect 282 -2742 288 -2736
rect 282 -2748 288 -2742
rect 282 -2754 288 -2748
rect 282 -2760 288 -2754
rect 282 -2766 288 -2760
rect 282 -2772 288 -2766
rect 282 -2778 288 -2772
rect 282 -2784 288 -2778
rect 282 -2790 288 -2784
rect 282 -2796 288 -2790
rect 282 -2802 288 -2796
rect 282 -2808 288 -2802
rect 282 -2814 288 -2808
rect 282 -2820 288 -2814
rect 282 -2826 288 -2820
rect 282 -2832 288 -2826
rect 282 -2838 288 -2832
rect 282 -2844 288 -2838
rect 282 -2850 288 -2844
rect 282 -2856 288 -2850
rect 282 -2862 288 -2856
rect 282 -2868 288 -2862
rect 282 -2874 288 -2868
rect 282 -2880 288 -2874
rect 282 -2886 288 -2880
rect 282 -2892 288 -2886
rect 282 -2898 288 -2892
rect 282 -2904 288 -2898
rect 282 -2910 288 -2904
rect 282 -2916 288 -2910
rect 282 -2922 288 -2916
rect 282 -2928 288 -2922
rect 282 -2934 288 -2928
rect 282 -2940 288 -2934
rect 282 -2946 288 -2940
rect 282 -2952 288 -2946
rect 282 -2958 288 -2952
rect 282 -2964 288 -2958
rect 282 -2970 288 -2964
rect 282 -2976 288 -2970
rect 282 -2982 288 -2976
rect 282 -2988 288 -2982
rect 282 -2994 288 -2988
rect 282 -3000 288 -2994
rect 282 -3006 288 -3000
rect 282 -3012 288 -3006
rect 282 -3018 288 -3012
rect 282 -3024 288 -3018
rect 282 -3030 288 -3024
rect 282 -3036 288 -3030
rect 282 -3042 288 -3036
rect 282 -3048 288 -3042
rect 282 -3054 288 -3048
rect 282 -3060 288 -3054
rect 282 -3066 288 -3060
rect 282 -3072 288 -3066
rect 282 -3078 288 -3072
rect 282 -3084 288 -3078
rect 282 -3090 288 -3084
rect 288 -1530 294 -1524
rect 288 -1536 294 -1530
rect 288 -1542 294 -1536
rect 288 -1548 294 -1542
rect 288 -1554 294 -1548
rect 288 -1560 294 -1554
rect 288 -1566 294 -1560
rect 288 -1572 294 -1566
rect 288 -1578 294 -1572
rect 288 -1584 294 -1578
rect 288 -1590 294 -1584
rect 288 -1596 294 -1590
rect 288 -1602 294 -1596
rect 288 -1608 294 -1602
rect 288 -1614 294 -1608
rect 288 -1620 294 -1614
rect 288 -1626 294 -1620
rect 288 -1632 294 -1626
rect 288 -1638 294 -1632
rect 288 -1644 294 -1638
rect 288 -1650 294 -1644
rect 288 -1656 294 -1650
rect 288 -1662 294 -1656
rect 288 -1668 294 -1662
rect 288 -1674 294 -1668
rect 288 -1680 294 -1674
rect 288 -1686 294 -1680
rect 288 -1692 294 -1686
rect 288 -1698 294 -1692
rect 288 -1704 294 -1698
rect 288 -1710 294 -1704
rect 288 -1716 294 -1710
rect 288 -1722 294 -1716
rect 288 -1728 294 -1722
rect 288 -1734 294 -1728
rect 288 -1740 294 -1734
rect 288 -1746 294 -1740
rect 288 -1752 294 -1746
rect 288 -1758 294 -1752
rect 288 -1764 294 -1758
rect 288 -1770 294 -1764
rect 288 -1776 294 -1770
rect 288 -1782 294 -1776
rect 288 -1788 294 -1782
rect 288 -1794 294 -1788
rect 288 -1800 294 -1794
rect 288 -1806 294 -1800
rect 288 -1812 294 -1806
rect 288 -1818 294 -1812
rect 288 -1824 294 -1818
rect 288 -1830 294 -1824
rect 288 -1836 294 -1830
rect 288 -1842 294 -1836
rect 288 -1848 294 -1842
rect 288 -1854 294 -1848
rect 288 -1860 294 -1854
rect 288 -1866 294 -1860
rect 288 -1872 294 -1866
rect 288 -1878 294 -1872
rect 288 -1884 294 -1878
rect 288 -1890 294 -1884
rect 288 -1896 294 -1890
rect 288 -1902 294 -1896
rect 288 -1908 294 -1902
rect 288 -1914 294 -1908
rect 288 -2712 294 -2706
rect 288 -2718 294 -2712
rect 288 -2724 294 -2718
rect 288 -2730 294 -2724
rect 288 -2736 294 -2730
rect 288 -2742 294 -2736
rect 288 -2748 294 -2742
rect 288 -2754 294 -2748
rect 288 -2760 294 -2754
rect 288 -2766 294 -2760
rect 288 -2772 294 -2766
rect 288 -2778 294 -2772
rect 288 -2784 294 -2778
rect 288 -2790 294 -2784
rect 288 -2796 294 -2790
rect 288 -2802 294 -2796
rect 288 -2808 294 -2802
rect 288 -2814 294 -2808
rect 288 -2820 294 -2814
rect 288 -2826 294 -2820
rect 288 -2832 294 -2826
rect 288 -2838 294 -2832
rect 288 -2844 294 -2838
rect 288 -2850 294 -2844
rect 288 -2856 294 -2850
rect 288 -2862 294 -2856
rect 288 -2868 294 -2862
rect 288 -2874 294 -2868
rect 288 -2880 294 -2874
rect 288 -2886 294 -2880
rect 288 -2892 294 -2886
rect 288 -2898 294 -2892
rect 288 -2904 294 -2898
rect 288 -2910 294 -2904
rect 288 -2916 294 -2910
rect 288 -2922 294 -2916
rect 288 -2928 294 -2922
rect 288 -2934 294 -2928
rect 288 -2940 294 -2934
rect 288 -2946 294 -2940
rect 288 -2952 294 -2946
rect 288 -2958 294 -2952
rect 288 -2964 294 -2958
rect 288 -2970 294 -2964
rect 288 -2976 294 -2970
rect 288 -2982 294 -2976
rect 288 -2988 294 -2982
rect 288 -2994 294 -2988
rect 288 -3000 294 -2994
rect 288 -3006 294 -3000
rect 288 -3012 294 -3006
rect 288 -3018 294 -3012
rect 288 -3024 294 -3018
rect 288 -3030 294 -3024
rect 288 -3036 294 -3030
rect 288 -3042 294 -3036
rect 288 -3048 294 -3042
rect 288 -3054 294 -3048
rect 288 -3060 294 -3054
rect 288 -3066 294 -3060
rect 288 -3072 294 -3066
rect 288 -3078 294 -3072
rect 288 -3084 294 -3078
rect 288 -3090 294 -3084
rect 288 -3096 294 -3090
rect 294 -1524 300 -1518
rect 294 -1530 300 -1524
rect 294 -1536 300 -1530
rect 294 -1542 300 -1536
rect 294 -1548 300 -1542
rect 294 -1554 300 -1548
rect 294 -1560 300 -1554
rect 294 -1566 300 -1560
rect 294 -1572 300 -1566
rect 294 -1578 300 -1572
rect 294 -1584 300 -1578
rect 294 -1590 300 -1584
rect 294 -1596 300 -1590
rect 294 -1602 300 -1596
rect 294 -1608 300 -1602
rect 294 -1614 300 -1608
rect 294 -1620 300 -1614
rect 294 -1626 300 -1620
rect 294 -1632 300 -1626
rect 294 -1638 300 -1632
rect 294 -1644 300 -1638
rect 294 -1650 300 -1644
rect 294 -1656 300 -1650
rect 294 -1662 300 -1656
rect 294 -1668 300 -1662
rect 294 -1674 300 -1668
rect 294 -1680 300 -1674
rect 294 -1686 300 -1680
rect 294 -1692 300 -1686
rect 294 -1698 300 -1692
rect 294 -1704 300 -1698
rect 294 -1710 300 -1704
rect 294 -1716 300 -1710
rect 294 -1722 300 -1716
rect 294 -1728 300 -1722
rect 294 -1734 300 -1728
rect 294 -1740 300 -1734
rect 294 -1746 300 -1740
rect 294 -1752 300 -1746
rect 294 -1758 300 -1752
rect 294 -1764 300 -1758
rect 294 -1770 300 -1764
rect 294 -1776 300 -1770
rect 294 -1782 300 -1776
rect 294 -1788 300 -1782
rect 294 -1794 300 -1788
rect 294 -1800 300 -1794
rect 294 -1806 300 -1800
rect 294 -1812 300 -1806
rect 294 -1818 300 -1812
rect 294 -1824 300 -1818
rect 294 -1830 300 -1824
rect 294 -1836 300 -1830
rect 294 -1842 300 -1836
rect 294 -1848 300 -1842
rect 294 -1854 300 -1848
rect 294 -1860 300 -1854
rect 294 -1866 300 -1860
rect 294 -1872 300 -1866
rect 294 -1878 300 -1872
rect 294 -1884 300 -1878
rect 294 -1890 300 -1884
rect 294 -1896 300 -1890
rect 294 -1902 300 -1896
rect 294 -2724 300 -2718
rect 294 -2730 300 -2724
rect 294 -2736 300 -2730
rect 294 -2742 300 -2736
rect 294 -2748 300 -2742
rect 294 -2754 300 -2748
rect 294 -2760 300 -2754
rect 294 -2766 300 -2760
rect 294 -2772 300 -2766
rect 294 -2778 300 -2772
rect 294 -2784 300 -2778
rect 294 -2790 300 -2784
rect 294 -2796 300 -2790
rect 294 -2802 300 -2796
rect 294 -2808 300 -2802
rect 294 -2814 300 -2808
rect 294 -2820 300 -2814
rect 294 -2826 300 -2820
rect 294 -2832 300 -2826
rect 294 -2838 300 -2832
rect 294 -2844 300 -2838
rect 294 -2850 300 -2844
rect 294 -2856 300 -2850
rect 294 -2862 300 -2856
rect 294 -2868 300 -2862
rect 294 -2874 300 -2868
rect 294 -2880 300 -2874
rect 294 -2886 300 -2880
rect 294 -2892 300 -2886
rect 294 -2898 300 -2892
rect 294 -2904 300 -2898
rect 294 -2910 300 -2904
rect 294 -2916 300 -2910
rect 294 -2922 300 -2916
rect 294 -2928 300 -2922
rect 294 -2934 300 -2928
rect 294 -2940 300 -2934
rect 294 -2946 300 -2940
rect 294 -2952 300 -2946
rect 294 -2958 300 -2952
rect 294 -2964 300 -2958
rect 294 -2970 300 -2964
rect 294 -2976 300 -2970
rect 294 -2982 300 -2976
rect 294 -2988 300 -2982
rect 294 -2994 300 -2988
rect 294 -3000 300 -2994
rect 294 -3006 300 -3000
rect 294 -3012 300 -3006
rect 294 -3018 300 -3012
rect 294 -3024 300 -3018
rect 294 -3030 300 -3024
rect 294 -3036 300 -3030
rect 294 -3042 300 -3036
rect 294 -3048 300 -3042
rect 294 -3054 300 -3048
rect 294 -3060 300 -3054
rect 294 -3066 300 -3060
rect 294 -3072 300 -3066
rect 294 -3078 300 -3072
rect 294 -3084 300 -3078
rect 294 -3090 300 -3084
rect 294 -3096 300 -3090
rect 294 -3102 300 -3096
rect 300 -1518 306 -1512
rect 300 -1524 306 -1518
rect 300 -1530 306 -1524
rect 300 -1536 306 -1530
rect 300 -1542 306 -1536
rect 300 -1548 306 -1542
rect 300 -1554 306 -1548
rect 300 -1560 306 -1554
rect 300 -1566 306 -1560
rect 300 -1572 306 -1566
rect 300 -1578 306 -1572
rect 300 -1584 306 -1578
rect 300 -1590 306 -1584
rect 300 -1596 306 -1590
rect 300 -1602 306 -1596
rect 300 -1608 306 -1602
rect 300 -1614 306 -1608
rect 300 -1620 306 -1614
rect 300 -1626 306 -1620
rect 300 -1632 306 -1626
rect 300 -1638 306 -1632
rect 300 -1644 306 -1638
rect 300 -1650 306 -1644
rect 300 -1656 306 -1650
rect 300 -1662 306 -1656
rect 300 -1668 306 -1662
rect 300 -1674 306 -1668
rect 300 -1680 306 -1674
rect 300 -1686 306 -1680
rect 300 -1692 306 -1686
rect 300 -1698 306 -1692
rect 300 -1704 306 -1698
rect 300 -1710 306 -1704
rect 300 -1716 306 -1710
rect 300 -1722 306 -1716
rect 300 -1728 306 -1722
rect 300 -1734 306 -1728
rect 300 -1740 306 -1734
rect 300 -1746 306 -1740
rect 300 -1752 306 -1746
rect 300 -1758 306 -1752
rect 300 -1764 306 -1758
rect 300 -1770 306 -1764
rect 300 -1776 306 -1770
rect 300 -1782 306 -1776
rect 300 -1788 306 -1782
rect 300 -1794 306 -1788
rect 300 -1800 306 -1794
rect 300 -1806 306 -1800
rect 300 -1812 306 -1806
rect 300 -1818 306 -1812
rect 300 -1824 306 -1818
rect 300 -1830 306 -1824
rect 300 -1836 306 -1830
rect 300 -1842 306 -1836
rect 300 -1848 306 -1842
rect 300 -1854 306 -1848
rect 300 -1860 306 -1854
rect 300 -1866 306 -1860
rect 300 -1872 306 -1866
rect 300 -1878 306 -1872
rect 300 -1884 306 -1878
rect 300 -1890 306 -1884
rect 300 -2736 306 -2730
rect 300 -2742 306 -2736
rect 300 -2748 306 -2742
rect 300 -2754 306 -2748
rect 300 -2760 306 -2754
rect 300 -2766 306 -2760
rect 300 -2772 306 -2766
rect 300 -2778 306 -2772
rect 300 -2784 306 -2778
rect 300 -2790 306 -2784
rect 300 -2796 306 -2790
rect 300 -2802 306 -2796
rect 300 -2808 306 -2802
rect 300 -2814 306 -2808
rect 300 -2820 306 -2814
rect 300 -2826 306 -2820
rect 300 -2832 306 -2826
rect 300 -2838 306 -2832
rect 300 -2844 306 -2838
rect 300 -2850 306 -2844
rect 300 -2856 306 -2850
rect 300 -2862 306 -2856
rect 300 -2868 306 -2862
rect 300 -2874 306 -2868
rect 300 -2880 306 -2874
rect 300 -2886 306 -2880
rect 300 -2892 306 -2886
rect 300 -2898 306 -2892
rect 300 -2904 306 -2898
rect 300 -2910 306 -2904
rect 300 -2916 306 -2910
rect 300 -2922 306 -2916
rect 300 -2928 306 -2922
rect 300 -2934 306 -2928
rect 300 -2940 306 -2934
rect 300 -2946 306 -2940
rect 300 -2952 306 -2946
rect 300 -2958 306 -2952
rect 300 -2964 306 -2958
rect 300 -2970 306 -2964
rect 300 -2976 306 -2970
rect 300 -2982 306 -2976
rect 300 -2988 306 -2982
rect 300 -2994 306 -2988
rect 300 -3000 306 -2994
rect 300 -3006 306 -3000
rect 300 -3012 306 -3006
rect 300 -3018 306 -3012
rect 300 -3024 306 -3018
rect 300 -3030 306 -3024
rect 300 -3036 306 -3030
rect 300 -3042 306 -3036
rect 300 -3048 306 -3042
rect 300 -3054 306 -3048
rect 300 -3060 306 -3054
rect 300 -3066 306 -3060
rect 300 -3072 306 -3066
rect 300 -3078 306 -3072
rect 300 -3084 306 -3078
rect 300 -3090 306 -3084
rect 300 -3096 306 -3090
rect 300 -3102 306 -3096
rect 300 -3108 306 -3102
rect 306 -1512 312 -1506
rect 306 -1518 312 -1512
rect 306 -1524 312 -1518
rect 306 -1530 312 -1524
rect 306 -1536 312 -1530
rect 306 -1542 312 -1536
rect 306 -1548 312 -1542
rect 306 -1554 312 -1548
rect 306 -1560 312 -1554
rect 306 -1566 312 -1560
rect 306 -1572 312 -1566
rect 306 -1578 312 -1572
rect 306 -1584 312 -1578
rect 306 -1590 312 -1584
rect 306 -1596 312 -1590
rect 306 -1602 312 -1596
rect 306 -1608 312 -1602
rect 306 -1614 312 -1608
rect 306 -1620 312 -1614
rect 306 -1626 312 -1620
rect 306 -1632 312 -1626
rect 306 -1638 312 -1632
rect 306 -1644 312 -1638
rect 306 -1650 312 -1644
rect 306 -1656 312 -1650
rect 306 -1662 312 -1656
rect 306 -1668 312 -1662
rect 306 -1674 312 -1668
rect 306 -1680 312 -1674
rect 306 -1686 312 -1680
rect 306 -1692 312 -1686
rect 306 -1698 312 -1692
rect 306 -1704 312 -1698
rect 306 -1710 312 -1704
rect 306 -1716 312 -1710
rect 306 -1722 312 -1716
rect 306 -1728 312 -1722
rect 306 -1734 312 -1728
rect 306 -1740 312 -1734
rect 306 -1746 312 -1740
rect 306 -1752 312 -1746
rect 306 -1758 312 -1752
rect 306 -1764 312 -1758
rect 306 -1770 312 -1764
rect 306 -1776 312 -1770
rect 306 -1782 312 -1776
rect 306 -1788 312 -1782
rect 306 -1794 312 -1788
rect 306 -1800 312 -1794
rect 306 -1806 312 -1800
rect 306 -1812 312 -1806
rect 306 -1818 312 -1812
rect 306 -1824 312 -1818
rect 306 -1830 312 -1824
rect 306 -1836 312 -1830
rect 306 -1842 312 -1836
rect 306 -1848 312 -1842
rect 306 -1854 312 -1848
rect 306 -1860 312 -1854
rect 306 -1866 312 -1860
rect 306 -1872 312 -1866
rect 306 -1878 312 -1872
rect 306 -2754 312 -2748
rect 306 -2760 312 -2754
rect 306 -2766 312 -2760
rect 306 -2772 312 -2766
rect 306 -2778 312 -2772
rect 306 -2784 312 -2778
rect 306 -2790 312 -2784
rect 306 -2796 312 -2790
rect 306 -2802 312 -2796
rect 306 -2808 312 -2802
rect 306 -2814 312 -2808
rect 306 -2820 312 -2814
rect 306 -2826 312 -2820
rect 306 -2832 312 -2826
rect 306 -2838 312 -2832
rect 306 -2844 312 -2838
rect 306 -2850 312 -2844
rect 306 -2856 312 -2850
rect 306 -2862 312 -2856
rect 306 -2868 312 -2862
rect 306 -2874 312 -2868
rect 306 -2880 312 -2874
rect 306 -2886 312 -2880
rect 306 -2892 312 -2886
rect 306 -2898 312 -2892
rect 306 -2904 312 -2898
rect 306 -2910 312 -2904
rect 306 -2916 312 -2910
rect 306 -2922 312 -2916
rect 306 -2928 312 -2922
rect 306 -2934 312 -2928
rect 306 -2940 312 -2934
rect 306 -2946 312 -2940
rect 306 -2952 312 -2946
rect 306 -2958 312 -2952
rect 306 -2964 312 -2958
rect 306 -2970 312 -2964
rect 306 -2976 312 -2970
rect 306 -2982 312 -2976
rect 306 -2988 312 -2982
rect 306 -2994 312 -2988
rect 306 -3000 312 -2994
rect 306 -3006 312 -3000
rect 306 -3012 312 -3006
rect 306 -3018 312 -3012
rect 306 -3024 312 -3018
rect 306 -3030 312 -3024
rect 306 -3036 312 -3030
rect 306 -3042 312 -3036
rect 306 -3048 312 -3042
rect 306 -3054 312 -3048
rect 306 -3060 312 -3054
rect 306 -3066 312 -3060
rect 306 -3072 312 -3066
rect 306 -3078 312 -3072
rect 306 -3084 312 -3078
rect 306 -3090 312 -3084
rect 306 -3096 312 -3090
rect 306 -3102 312 -3096
rect 306 -3108 312 -3102
rect 306 -3114 312 -3108
rect 306 -3120 312 -3114
rect 312 -1500 318 -1494
rect 312 -1506 318 -1500
rect 312 -1512 318 -1506
rect 312 -1518 318 -1512
rect 312 -1524 318 -1518
rect 312 -1530 318 -1524
rect 312 -1536 318 -1530
rect 312 -1542 318 -1536
rect 312 -1548 318 -1542
rect 312 -1554 318 -1548
rect 312 -1560 318 -1554
rect 312 -1566 318 -1560
rect 312 -1572 318 -1566
rect 312 -1578 318 -1572
rect 312 -1584 318 -1578
rect 312 -1590 318 -1584
rect 312 -1596 318 -1590
rect 312 -1602 318 -1596
rect 312 -1608 318 -1602
rect 312 -1614 318 -1608
rect 312 -1620 318 -1614
rect 312 -1626 318 -1620
rect 312 -1632 318 -1626
rect 312 -1638 318 -1632
rect 312 -1644 318 -1638
rect 312 -1650 318 -1644
rect 312 -1656 318 -1650
rect 312 -1662 318 -1656
rect 312 -1668 318 -1662
rect 312 -1674 318 -1668
rect 312 -1680 318 -1674
rect 312 -1686 318 -1680
rect 312 -1692 318 -1686
rect 312 -1698 318 -1692
rect 312 -1704 318 -1698
rect 312 -1710 318 -1704
rect 312 -1716 318 -1710
rect 312 -1722 318 -1716
rect 312 -1728 318 -1722
rect 312 -1734 318 -1728
rect 312 -1740 318 -1734
rect 312 -1746 318 -1740
rect 312 -1752 318 -1746
rect 312 -1758 318 -1752
rect 312 -1764 318 -1758
rect 312 -1770 318 -1764
rect 312 -1776 318 -1770
rect 312 -1782 318 -1776
rect 312 -1788 318 -1782
rect 312 -1794 318 -1788
rect 312 -1800 318 -1794
rect 312 -1806 318 -1800
rect 312 -1812 318 -1806
rect 312 -1818 318 -1812
rect 312 -1824 318 -1818
rect 312 -1830 318 -1824
rect 312 -1836 318 -1830
rect 312 -1842 318 -1836
rect 312 -1848 318 -1842
rect 312 -1854 318 -1848
rect 312 -1860 318 -1854
rect 312 -1866 318 -1860
rect 312 -2766 318 -2760
rect 312 -2772 318 -2766
rect 312 -2778 318 -2772
rect 312 -2784 318 -2778
rect 312 -2790 318 -2784
rect 312 -2796 318 -2790
rect 312 -2802 318 -2796
rect 312 -2808 318 -2802
rect 312 -2814 318 -2808
rect 312 -2820 318 -2814
rect 312 -2826 318 -2820
rect 312 -2832 318 -2826
rect 312 -2838 318 -2832
rect 312 -2844 318 -2838
rect 312 -2850 318 -2844
rect 312 -2856 318 -2850
rect 312 -2862 318 -2856
rect 312 -2868 318 -2862
rect 312 -2874 318 -2868
rect 312 -2880 318 -2874
rect 312 -2886 318 -2880
rect 312 -2892 318 -2886
rect 312 -2898 318 -2892
rect 312 -2904 318 -2898
rect 312 -2910 318 -2904
rect 312 -2916 318 -2910
rect 312 -2922 318 -2916
rect 312 -2928 318 -2922
rect 312 -2934 318 -2928
rect 312 -2940 318 -2934
rect 312 -2946 318 -2940
rect 312 -2952 318 -2946
rect 312 -2958 318 -2952
rect 312 -2964 318 -2958
rect 312 -2970 318 -2964
rect 312 -2976 318 -2970
rect 312 -2982 318 -2976
rect 312 -2988 318 -2982
rect 312 -2994 318 -2988
rect 312 -3000 318 -2994
rect 312 -3006 318 -3000
rect 312 -3012 318 -3006
rect 312 -3018 318 -3012
rect 312 -3024 318 -3018
rect 312 -3030 318 -3024
rect 312 -3036 318 -3030
rect 312 -3042 318 -3036
rect 312 -3048 318 -3042
rect 312 -3054 318 -3048
rect 312 -3060 318 -3054
rect 312 -3066 318 -3060
rect 312 -3072 318 -3066
rect 312 -3078 318 -3072
rect 312 -3084 318 -3078
rect 312 -3090 318 -3084
rect 312 -3096 318 -3090
rect 312 -3102 318 -3096
rect 312 -3108 318 -3102
rect 312 -3114 318 -3108
rect 312 -3120 318 -3114
rect 312 -3126 318 -3120
rect 318 -1494 324 -1488
rect 318 -1500 324 -1494
rect 318 -1506 324 -1500
rect 318 -1512 324 -1506
rect 318 -1518 324 -1512
rect 318 -1524 324 -1518
rect 318 -1530 324 -1524
rect 318 -1536 324 -1530
rect 318 -1542 324 -1536
rect 318 -1548 324 -1542
rect 318 -1554 324 -1548
rect 318 -1560 324 -1554
rect 318 -1566 324 -1560
rect 318 -1572 324 -1566
rect 318 -1578 324 -1572
rect 318 -1584 324 -1578
rect 318 -1590 324 -1584
rect 318 -1596 324 -1590
rect 318 -1602 324 -1596
rect 318 -1608 324 -1602
rect 318 -1614 324 -1608
rect 318 -1620 324 -1614
rect 318 -1626 324 -1620
rect 318 -1632 324 -1626
rect 318 -1638 324 -1632
rect 318 -1644 324 -1638
rect 318 -1650 324 -1644
rect 318 -1656 324 -1650
rect 318 -1662 324 -1656
rect 318 -1668 324 -1662
rect 318 -1674 324 -1668
rect 318 -1680 324 -1674
rect 318 -1686 324 -1680
rect 318 -1692 324 -1686
rect 318 -1698 324 -1692
rect 318 -1704 324 -1698
rect 318 -1710 324 -1704
rect 318 -1716 324 -1710
rect 318 -1722 324 -1716
rect 318 -1728 324 -1722
rect 318 -1734 324 -1728
rect 318 -1740 324 -1734
rect 318 -1746 324 -1740
rect 318 -1752 324 -1746
rect 318 -1758 324 -1752
rect 318 -1764 324 -1758
rect 318 -1770 324 -1764
rect 318 -1776 324 -1770
rect 318 -1782 324 -1776
rect 318 -1788 324 -1782
rect 318 -1794 324 -1788
rect 318 -1800 324 -1794
rect 318 -1806 324 -1800
rect 318 -1812 324 -1806
rect 318 -1818 324 -1812
rect 318 -1824 324 -1818
rect 318 -1830 324 -1824
rect 318 -1836 324 -1830
rect 318 -1842 324 -1836
rect 318 -1848 324 -1842
rect 318 -1854 324 -1848
rect 318 -2778 324 -2772
rect 318 -2784 324 -2778
rect 318 -2790 324 -2784
rect 318 -2796 324 -2790
rect 318 -2802 324 -2796
rect 318 -2808 324 -2802
rect 318 -2814 324 -2808
rect 318 -2820 324 -2814
rect 318 -2826 324 -2820
rect 318 -2832 324 -2826
rect 318 -2838 324 -2832
rect 318 -2844 324 -2838
rect 318 -2850 324 -2844
rect 318 -2856 324 -2850
rect 318 -2862 324 -2856
rect 318 -2868 324 -2862
rect 318 -2874 324 -2868
rect 318 -2880 324 -2874
rect 318 -2886 324 -2880
rect 318 -2892 324 -2886
rect 318 -2898 324 -2892
rect 318 -2904 324 -2898
rect 318 -2910 324 -2904
rect 318 -2916 324 -2910
rect 318 -2922 324 -2916
rect 318 -2928 324 -2922
rect 318 -2934 324 -2928
rect 318 -2940 324 -2934
rect 318 -2946 324 -2940
rect 318 -2952 324 -2946
rect 318 -2958 324 -2952
rect 318 -2964 324 -2958
rect 318 -2970 324 -2964
rect 318 -2976 324 -2970
rect 318 -2982 324 -2976
rect 318 -2988 324 -2982
rect 318 -2994 324 -2988
rect 318 -3000 324 -2994
rect 318 -3006 324 -3000
rect 318 -3012 324 -3006
rect 318 -3018 324 -3012
rect 318 -3024 324 -3018
rect 318 -3030 324 -3024
rect 318 -3036 324 -3030
rect 318 -3042 324 -3036
rect 318 -3048 324 -3042
rect 318 -3054 324 -3048
rect 318 -3060 324 -3054
rect 318 -3066 324 -3060
rect 318 -3072 324 -3066
rect 318 -3078 324 -3072
rect 318 -3084 324 -3078
rect 318 -3090 324 -3084
rect 318 -3096 324 -3090
rect 318 -3102 324 -3096
rect 318 -3108 324 -3102
rect 318 -3114 324 -3108
rect 318 -3120 324 -3114
rect 318 -3126 324 -3120
rect 318 -3132 324 -3126
rect 324 -1488 330 -1482
rect 324 -1494 330 -1488
rect 324 -1500 330 -1494
rect 324 -1506 330 -1500
rect 324 -1512 330 -1506
rect 324 -1518 330 -1512
rect 324 -1524 330 -1518
rect 324 -1530 330 -1524
rect 324 -1536 330 -1530
rect 324 -1542 330 -1536
rect 324 -1548 330 -1542
rect 324 -1554 330 -1548
rect 324 -1560 330 -1554
rect 324 -1566 330 -1560
rect 324 -1572 330 -1566
rect 324 -1578 330 -1572
rect 324 -1584 330 -1578
rect 324 -1590 330 -1584
rect 324 -1596 330 -1590
rect 324 -1602 330 -1596
rect 324 -1608 330 -1602
rect 324 -1614 330 -1608
rect 324 -1620 330 -1614
rect 324 -1626 330 -1620
rect 324 -1632 330 -1626
rect 324 -1638 330 -1632
rect 324 -1644 330 -1638
rect 324 -1650 330 -1644
rect 324 -1656 330 -1650
rect 324 -1662 330 -1656
rect 324 -1668 330 -1662
rect 324 -1674 330 -1668
rect 324 -1680 330 -1674
rect 324 -1686 330 -1680
rect 324 -1692 330 -1686
rect 324 -1698 330 -1692
rect 324 -1704 330 -1698
rect 324 -1710 330 -1704
rect 324 -1716 330 -1710
rect 324 -1722 330 -1716
rect 324 -1728 330 -1722
rect 324 -1734 330 -1728
rect 324 -1740 330 -1734
rect 324 -1746 330 -1740
rect 324 -1752 330 -1746
rect 324 -1758 330 -1752
rect 324 -1764 330 -1758
rect 324 -1770 330 -1764
rect 324 -1776 330 -1770
rect 324 -1782 330 -1776
rect 324 -1788 330 -1782
rect 324 -1794 330 -1788
rect 324 -1800 330 -1794
rect 324 -1806 330 -1800
rect 324 -1812 330 -1806
rect 324 -1818 330 -1812
rect 324 -1824 330 -1818
rect 324 -1830 330 -1824
rect 324 -1836 330 -1830
rect 324 -1842 330 -1836
rect 324 -2790 330 -2784
rect 324 -2796 330 -2790
rect 324 -2802 330 -2796
rect 324 -2808 330 -2802
rect 324 -2814 330 -2808
rect 324 -2820 330 -2814
rect 324 -2826 330 -2820
rect 324 -2832 330 -2826
rect 324 -2838 330 -2832
rect 324 -2844 330 -2838
rect 324 -2850 330 -2844
rect 324 -2856 330 -2850
rect 324 -2862 330 -2856
rect 324 -2868 330 -2862
rect 324 -2874 330 -2868
rect 324 -2880 330 -2874
rect 324 -2886 330 -2880
rect 324 -2892 330 -2886
rect 324 -2898 330 -2892
rect 324 -2904 330 -2898
rect 324 -2910 330 -2904
rect 324 -2916 330 -2910
rect 324 -2922 330 -2916
rect 324 -2928 330 -2922
rect 324 -2934 330 -2928
rect 324 -2940 330 -2934
rect 324 -2946 330 -2940
rect 324 -2952 330 -2946
rect 324 -2958 330 -2952
rect 324 -2964 330 -2958
rect 324 -2970 330 -2964
rect 324 -2976 330 -2970
rect 324 -2982 330 -2976
rect 324 -2988 330 -2982
rect 324 -2994 330 -2988
rect 324 -3000 330 -2994
rect 324 -3006 330 -3000
rect 324 -3012 330 -3006
rect 324 -3018 330 -3012
rect 324 -3024 330 -3018
rect 324 -3030 330 -3024
rect 324 -3036 330 -3030
rect 324 -3042 330 -3036
rect 324 -3048 330 -3042
rect 324 -3054 330 -3048
rect 324 -3060 330 -3054
rect 324 -3066 330 -3060
rect 324 -3072 330 -3066
rect 324 -3078 330 -3072
rect 324 -3084 330 -3078
rect 324 -3090 330 -3084
rect 324 -3096 330 -3090
rect 324 -3102 330 -3096
rect 324 -3108 330 -3102
rect 324 -3114 330 -3108
rect 324 -3120 330 -3114
rect 324 -3126 330 -3120
rect 324 -3132 330 -3126
rect 324 -3138 330 -3132
rect 330 -1482 336 -1476
rect 330 -1488 336 -1482
rect 330 -1494 336 -1488
rect 330 -1500 336 -1494
rect 330 -1506 336 -1500
rect 330 -1512 336 -1506
rect 330 -1518 336 -1512
rect 330 -1524 336 -1518
rect 330 -1530 336 -1524
rect 330 -1536 336 -1530
rect 330 -1542 336 -1536
rect 330 -1548 336 -1542
rect 330 -1554 336 -1548
rect 330 -1560 336 -1554
rect 330 -1566 336 -1560
rect 330 -1572 336 -1566
rect 330 -1578 336 -1572
rect 330 -1584 336 -1578
rect 330 -1590 336 -1584
rect 330 -1596 336 -1590
rect 330 -1602 336 -1596
rect 330 -1608 336 -1602
rect 330 -1614 336 -1608
rect 330 -1620 336 -1614
rect 330 -1626 336 -1620
rect 330 -1632 336 -1626
rect 330 -1638 336 -1632
rect 330 -1644 336 -1638
rect 330 -1650 336 -1644
rect 330 -1656 336 -1650
rect 330 -1662 336 -1656
rect 330 -1668 336 -1662
rect 330 -1674 336 -1668
rect 330 -1680 336 -1674
rect 330 -1686 336 -1680
rect 330 -1692 336 -1686
rect 330 -1698 336 -1692
rect 330 -1704 336 -1698
rect 330 -1710 336 -1704
rect 330 -1716 336 -1710
rect 330 -1722 336 -1716
rect 330 -1728 336 -1722
rect 330 -1734 336 -1728
rect 330 -1740 336 -1734
rect 330 -1746 336 -1740
rect 330 -1752 336 -1746
rect 330 -1758 336 -1752
rect 330 -1764 336 -1758
rect 330 -1770 336 -1764
rect 330 -1776 336 -1770
rect 330 -1782 336 -1776
rect 330 -1788 336 -1782
rect 330 -1794 336 -1788
rect 330 -1800 336 -1794
rect 330 -1806 336 -1800
rect 330 -1812 336 -1806
rect 330 -1818 336 -1812
rect 330 -1824 336 -1818
rect 330 -1830 336 -1824
rect 330 -2796 336 -2790
rect 330 -2802 336 -2796
rect 330 -2808 336 -2802
rect 330 -2814 336 -2808
rect 330 -2820 336 -2814
rect 330 -2826 336 -2820
rect 330 -2832 336 -2826
rect 330 -2838 336 -2832
rect 330 -2844 336 -2838
rect 330 -2850 336 -2844
rect 330 -2856 336 -2850
rect 330 -2862 336 -2856
rect 330 -2868 336 -2862
rect 330 -2874 336 -2868
rect 330 -2880 336 -2874
rect 330 -2886 336 -2880
rect 330 -2892 336 -2886
rect 330 -2898 336 -2892
rect 330 -2904 336 -2898
rect 330 -2910 336 -2904
rect 330 -2916 336 -2910
rect 330 -2922 336 -2916
rect 330 -2928 336 -2922
rect 330 -2934 336 -2928
rect 330 -2940 336 -2934
rect 330 -2946 336 -2940
rect 330 -2952 336 -2946
rect 330 -2958 336 -2952
rect 330 -2964 336 -2958
rect 330 -2970 336 -2964
rect 330 -2976 336 -2970
rect 330 -2982 336 -2976
rect 330 -2988 336 -2982
rect 330 -2994 336 -2988
rect 330 -3000 336 -2994
rect 330 -3006 336 -3000
rect 330 -3012 336 -3006
rect 330 -3018 336 -3012
rect 330 -3024 336 -3018
rect 330 -3030 336 -3024
rect 330 -3036 336 -3030
rect 330 -3042 336 -3036
rect 330 -3048 336 -3042
rect 330 -3054 336 -3048
rect 330 -3060 336 -3054
rect 330 -3066 336 -3060
rect 330 -3072 336 -3066
rect 330 -3078 336 -3072
rect 330 -3084 336 -3078
rect 330 -3090 336 -3084
rect 330 -3096 336 -3090
rect 330 -3102 336 -3096
rect 330 -3108 336 -3102
rect 330 -3114 336 -3108
rect 330 -3120 336 -3114
rect 330 -3126 336 -3120
rect 330 -3132 336 -3126
rect 330 -3138 336 -3132
rect 330 -3144 336 -3138
rect 336 -1476 342 -1470
rect 336 -1482 342 -1476
rect 336 -1488 342 -1482
rect 336 -1494 342 -1488
rect 336 -1500 342 -1494
rect 336 -1506 342 -1500
rect 336 -1512 342 -1506
rect 336 -1518 342 -1512
rect 336 -1524 342 -1518
rect 336 -1530 342 -1524
rect 336 -1536 342 -1530
rect 336 -1542 342 -1536
rect 336 -1548 342 -1542
rect 336 -1554 342 -1548
rect 336 -1560 342 -1554
rect 336 -1566 342 -1560
rect 336 -1572 342 -1566
rect 336 -1578 342 -1572
rect 336 -1584 342 -1578
rect 336 -1590 342 -1584
rect 336 -1596 342 -1590
rect 336 -1602 342 -1596
rect 336 -1608 342 -1602
rect 336 -1614 342 -1608
rect 336 -1620 342 -1614
rect 336 -1626 342 -1620
rect 336 -1632 342 -1626
rect 336 -1638 342 -1632
rect 336 -1644 342 -1638
rect 336 -1650 342 -1644
rect 336 -1656 342 -1650
rect 336 -1662 342 -1656
rect 336 -1668 342 -1662
rect 336 -1674 342 -1668
rect 336 -1680 342 -1674
rect 336 -1686 342 -1680
rect 336 -1692 342 -1686
rect 336 -1698 342 -1692
rect 336 -1704 342 -1698
rect 336 -1710 342 -1704
rect 336 -1716 342 -1710
rect 336 -1722 342 -1716
rect 336 -1728 342 -1722
rect 336 -1734 342 -1728
rect 336 -1740 342 -1734
rect 336 -1746 342 -1740
rect 336 -1752 342 -1746
rect 336 -1758 342 -1752
rect 336 -1764 342 -1758
rect 336 -1770 342 -1764
rect 336 -1776 342 -1770
rect 336 -1782 342 -1776
rect 336 -1788 342 -1782
rect 336 -1794 342 -1788
rect 336 -1800 342 -1794
rect 336 -1806 342 -1800
rect 336 -1812 342 -1806
rect 336 -1818 342 -1812
rect 336 -2808 342 -2802
rect 336 -2814 342 -2808
rect 336 -2820 342 -2814
rect 336 -2826 342 -2820
rect 336 -2832 342 -2826
rect 336 -2838 342 -2832
rect 336 -2844 342 -2838
rect 336 -2850 342 -2844
rect 336 -2856 342 -2850
rect 336 -2862 342 -2856
rect 336 -2868 342 -2862
rect 336 -2874 342 -2868
rect 336 -2880 342 -2874
rect 336 -2886 342 -2880
rect 336 -2892 342 -2886
rect 336 -2898 342 -2892
rect 336 -2904 342 -2898
rect 336 -2910 342 -2904
rect 336 -2916 342 -2910
rect 336 -2922 342 -2916
rect 336 -2928 342 -2922
rect 336 -2934 342 -2928
rect 336 -2940 342 -2934
rect 336 -2946 342 -2940
rect 336 -2952 342 -2946
rect 336 -2958 342 -2952
rect 336 -2964 342 -2958
rect 336 -2970 342 -2964
rect 336 -2976 342 -2970
rect 336 -2982 342 -2976
rect 336 -2988 342 -2982
rect 336 -2994 342 -2988
rect 336 -3000 342 -2994
rect 336 -3006 342 -3000
rect 336 -3012 342 -3006
rect 336 -3018 342 -3012
rect 336 -3024 342 -3018
rect 336 -3030 342 -3024
rect 336 -3036 342 -3030
rect 336 -3042 342 -3036
rect 336 -3048 342 -3042
rect 336 -3054 342 -3048
rect 336 -3060 342 -3054
rect 336 -3066 342 -3060
rect 336 -3072 342 -3066
rect 336 -3078 342 -3072
rect 336 -3084 342 -3078
rect 336 -3090 342 -3084
rect 336 -3096 342 -3090
rect 336 -3102 342 -3096
rect 336 -3108 342 -3102
rect 336 -3114 342 -3108
rect 336 -3120 342 -3114
rect 336 -3126 342 -3120
rect 336 -3132 342 -3126
rect 336 -3138 342 -3132
rect 336 -3144 342 -3138
rect 336 -3150 342 -3144
rect 342 -1470 348 -1464
rect 342 -1476 348 -1470
rect 342 -1482 348 -1476
rect 342 -1488 348 -1482
rect 342 -1494 348 -1488
rect 342 -1500 348 -1494
rect 342 -1506 348 -1500
rect 342 -1512 348 -1506
rect 342 -1518 348 -1512
rect 342 -1524 348 -1518
rect 342 -1530 348 -1524
rect 342 -1536 348 -1530
rect 342 -1542 348 -1536
rect 342 -1548 348 -1542
rect 342 -1554 348 -1548
rect 342 -1560 348 -1554
rect 342 -1566 348 -1560
rect 342 -1572 348 -1566
rect 342 -1578 348 -1572
rect 342 -1584 348 -1578
rect 342 -1590 348 -1584
rect 342 -1596 348 -1590
rect 342 -1602 348 -1596
rect 342 -1608 348 -1602
rect 342 -1614 348 -1608
rect 342 -1620 348 -1614
rect 342 -1626 348 -1620
rect 342 -1632 348 -1626
rect 342 -1638 348 -1632
rect 342 -1644 348 -1638
rect 342 -1650 348 -1644
rect 342 -1656 348 -1650
rect 342 -1662 348 -1656
rect 342 -1668 348 -1662
rect 342 -1674 348 -1668
rect 342 -1680 348 -1674
rect 342 -1686 348 -1680
rect 342 -1692 348 -1686
rect 342 -1698 348 -1692
rect 342 -1704 348 -1698
rect 342 -1710 348 -1704
rect 342 -1716 348 -1710
rect 342 -1722 348 -1716
rect 342 -1728 348 -1722
rect 342 -1734 348 -1728
rect 342 -1740 348 -1734
rect 342 -1746 348 -1740
rect 342 -1752 348 -1746
rect 342 -1758 348 -1752
rect 342 -1764 348 -1758
rect 342 -1770 348 -1764
rect 342 -1776 348 -1770
rect 342 -1782 348 -1776
rect 342 -1788 348 -1782
rect 342 -1794 348 -1788
rect 342 -1800 348 -1794
rect 342 -1806 348 -1800
rect 342 -2820 348 -2814
rect 342 -2826 348 -2820
rect 342 -2832 348 -2826
rect 342 -2838 348 -2832
rect 342 -2844 348 -2838
rect 342 -2850 348 -2844
rect 342 -2856 348 -2850
rect 342 -2862 348 -2856
rect 342 -2868 348 -2862
rect 342 -2874 348 -2868
rect 342 -2880 348 -2874
rect 342 -2886 348 -2880
rect 342 -2892 348 -2886
rect 342 -2898 348 -2892
rect 342 -2904 348 -2898
rect 342 -2910 348 -2904
rect 342 -2916 348 -2910
rect 342 -2922 348 -2916
rect 342 -2928 348 -2922
rect 342 -2934 348 -2928
rect 342 -2940 348 -2934
rect 342 -2946 348 -2940
rect 342 -2952 348 -2946
rect 342 -2958 348 -2952
rect 342 -2964 348 -2958
rect 342 -2970 348 -2964
rect 342 -2976 348 -2970
rect 342 -2982 348 -2976
rect 342 -2988 348 -2982
rect 342 -2994 348 -2988
rect 342 -3000 348 -2994
rect 342 -3006 348 -3000
rect 342 -3012 348 -3006
rect 342 -3018 348 -3012
rect 342 -3024 348 -3018
rect 342 -3030 348 -3024
rect 342 -3036 348 -3030
rect 342 -3042 348 -3036
rect 342 -3048 348 -3042
rect 342 -3054 348 -3048
rect 342 -3060 348 -3054
rect 342 -3066 348 -3060
rect 342 -3072 348 -3066
rect 342 -3078 348 -3072
rect 342 -3084 348 -3078
rect 342 -3090 348 -3084
rect 342 -3096 348 -3090
rect 342 -3102 348 -3096
rect 342 -3108 348 -3102
rect 342 -3114 348 -3108
rect 342 -3120 348 -3114
rect 342 -3126 348 -3120
rect 342 -3132 348 -3126
rect 342 -3138 348 -3132
rect 342 -3144 348 -3138
rect 342 -3150 348 -3144
rect 342 -3156 348 -3150
rect 348 -1464 354 -1458
rect 348 -1470 354 -1464
rect 348 -1476 354 -1470
rect 348 -1482 354 -1476
rect 348 -1488 354 -1482
rect 348 -1494 354 -1488
rect 348 -1500 354 -1494
rect 348 -1506 354 -1500
rect 348 -1512 354 -1506
rect 348 -1518 354 -1512
rect 348 -1524 354 -1518
rect 348 -1530 354 -1524
rect 348 -1536 354 -1530
rect 348 -1542 354 -1536
rect 348 -1548 354 -1542
rect 348 -1554 354 -1548
rect 348 -1560 354 -1554
rect 348 -1566 354 -1560
rect 348 -1572 354 -1566
rect 348 -1578 354 -1572
rect 348 -1584 354 -1578
rect 348 -1590 354 -1584
rect 348 -1596 354 -1590
rect 348 -1602 354 -1596
rect 348 -1608 354 -1602
rect 348 -1614 354 -1608
rect 348 -1620 354 -1614
rect 348 -1626 354 -1620
rect 348 -1632 354 -1626
rect 348 -1638 354 -1632
rect 348 -1644 354 -1638
rect 348 -1650 354 -1644
rect 348 -1656 354 -1650
rect 348 -1662 354 -1656
rect 348 -1668 354 -1662
rect 348 -1674 354 -1668
rect 348 -1680 354 -1674
rect 348 -1686 354 -1680
rect 348 -1692 354 -1686
rect 348 -1698 354 -1692
rect 348 -1704 354 -1698
rect 348 -1710 354 -1704
rect 348 -1716 354 -1710
rect 348 -1722 354 -1716
rect 348 -1728 354 -1722
rect 348 -1734 354 -1728
rect 348 -1740 354 -1734
rect 348 -1746 354 -1740
rect 348 -1752 354 -1746
rect 348 -1758 354 -1752
rect 348 -1764 354 -1758
rect 348 -1770 354 -1764
rect 348 -1776 354 -1770
rect 348 -1782 354 -1776
rect 348 -1788 354 -1782
rect 348 -1794 354 -1788
rect 348 -2832 354 -2826
rect 348 -2838 354 -2832
rect 348 -2844 354 -2838
rect 348 -2850 354 -2844
rect 348 -2856 354 -2850
rect 348 -2862 354 -2856
rect 348 -2868 354 -2862
rect 348 -2874 354 -2868
rect 348 -2880 354 -2874
rect 348 -2886 354 -2880
rect 348 -2892 354 -2886
rect 348 -2898 354 -2892
rect 348 -2904 354 -2898
rect 348 -2910 354 -2904
rect 348 -2916 354 -2910
rect 348 -2922 354 -2916
rect 348 -2928 354 -2922
rect 348 -2934 354 -2928
rect 348 -2940 354 -2934
rect 348 -2946 354 -2940
rect 348 -2952 354 -2946
rect 348 -2958 354 -2952
rect 348 -2964 354 -2958
rect 348 -2970 354 -2964
rect 348 -2976 354 -2970
rect 348 -2982 354 -2976
rect 348 -2988 354 -2982
rect 348 -2994 354 -2988
rect 348 -3000 354 -2994
rect 348 -3006 354 -3000
rect 348 -3012 354 -3006
rect 348 -3018 354 -3012
rect 348 -3024 354 -3018
rect 348 -3030 354 -3024
rect 348 -3036 354 -3030
rect 348 -3042 354 -3036
rect 348 -3048 354 -3042
rect 348 -3054 354 -3048
rect 348 -3060 354 -3054
rect 348 -3066 354 -3060
rect 348 -3072 354 -3066
rect 348 -3078 354 -3072
rect 348 -3084 354 -3078
rect 348 -3090 354 -3084
rect 348 -3096 354 -3090
rect 348 -3102 354 -3096
rect 348 -3108 354 -3102
rect 348 -3114 354 -3108
rect 348 -3120 354 -3114
rect 348 -3126 354 -3120
rect 348 -3132 354 -3126
rect 348 -3138 354 -3132
rect 348 -3144 354 -3138
rect 348 -3150 354 -3144
rect 348 -3156 354 -3150
rect 348 -3162 354 -3156
rect 354 -1458 360 -1452
rect 354 -1464 360 -1458
rect 354 -1470 360 -1464
rect 354 -1476 360 -1470
rect 354 -1482 360 -1476
rect 354 -1488 360 -1482
rect 354 -1494 360 -1488
rect 354 -1500 360 -1494
rect 354 -1506 360 -1500
rect 354 -1512 360 -1506
rect 354 -1518 360 -1512
rect 354 -1524 360 -1518
rect 354 -1530 360 -1524
rect 354 -1536 360 -1530
rect 354 -1542 360 -1536
rect 354 -1548 360 -1542
rect 354 -1554 360 -1548
rect 354 -1560 360 -1554
rect 354 -1566 360 -1560
rect 354 -1572 360 -1566
rect 354 -1578 360 -1572
rect 354 -1584 360 -1578
rect 354 -1590 360 -1584
rect 354 -1596 360 -1590
rect 354 -1602 360 -1596
rect 354 -1608 360 -1602
rect 354 -1614 360 -1608
rect 354 -1620 360 -1614
rect 354 -1626 360 -1620
rect 354 -1632 360 -1626
rect 354 -1638 360 -1632
rect 354 -1644 360 -1638
rect 354 -1650 360 -1644
rect 354 -1656 360 -1650
rect 354 -1662 360 -1656
rect 354 -1668 360 -1662
rect 354 -1674 360 -1668
rect 354 -1680 360 -1674
rect 354 -1686 360 -1680
rect 354 -1692 360 -1686
rect 354 -1698 360 -1692
rect 354 -1704 360 -1698
rect 354 -1710 360 -1704
rect 354 -1716 360 -1710
rect 354 -1722 360 -1716
rect 354 -1728 360 -1722
rect 354 -1734 360 -1728
rect 354 -1740 360 -1734
rect 354 -1746 360 -1740
rect 354 -1752 360 -1746
rect 354 -1758 360 -1752
rect 354 -1764 360 -1758
rect 354 -1770 360 -1764
rect 354 -1776 360 -1770
rect 354 -1782 360 -1776
rect 354 -1788 360 -1782
rect 354 -2838 360 -2832
rect 354 -2844 360 -2838
rect 354 -2850 360 -2844
rect 354 -2856 360 -2850
rect 354 -2862 360 -2856
rect 354 -2868 360 -2862
rect 354 -2874 360 -2868
rect 354 -2880 360 -2874
rect 354 -2886 360 -2880
rect 354 -2892 360 -2886
rect 354 -2898 360 -2892
rect 354 -2904 360 -2898
rect 354 -2910 360 -2904
rect 354 -2916 360 -2910
rect 354 -2922 360 -2916
rect 354 -2928 360 -2922
rect 354 -2934 360 -2928
rect 354 -2940 360 -2934
rect 354 -2946 360 -2940
rect 354 -2952 360 -2946
rect 354 -2958 360 -2952
rect 354 -2964 360 -2958
rect 354 -2970 360 -2964
rect 354 -2976 360 -2970
rect 354 -2982 360 -2976
rect 354 -2988 360 -2982
rect 354 -2994 360 -2988
rect 354 -3000 360 -2994
rect 354 -3006 360 -3000
rect 354 -3012 360 -3006
rect 354 -3018 360 -3012
rect 354 -3024 360 -3018
rect 354 -3030 360 -3024
rect 354 -3036 360 -3030
rect 354 -3042 360 -3036
rect 354 -3048 360 -3042
rect 354 -3054 360 -3048
rect 354 -3060 360 -3054
rect 354 -3066 360 -3060
rect 354 -3072 360 -3066
rect 354 -3078 360 -3072
rect 354 -3084 360 -3078
rect 354 -3090 360 -3084
rect 354 -3096 360 -3090
rect 354 -3102 360 -3096
rect 354 -3108 360 -3102
rect 354 -3114 360 -3108
rect 354 -3120 360 -3114
rect 354 -3126 360 -3120
rect 354 -3132 360 -3126
rect 354 -3138 360 -3132
rect 354 -3144 360 -3138
rect 354 -3150 360 -3144
rect 354 -3156 360 -3150
rect 354 -3162 360 -3156
rect 354 -3168 360 -3162
rect 360 -1452 366 -1446
rect 360 -1458 366 -1452
rect 360 -1464 366 -1458
rect 360 -1470 366 -1464
rect 360 -1476 366 -1470
rect 360 -1482 366 -1476
rect 360 -1488 366 -1482
rect 360 -1494 366 -1488
rect 360 -1500 366 -1494
rect 360 -1506 366 -1500
rect 360 -1512 366 -1506
rect 360 -1518 366 -1512
rect 360 -1524 366 -1518
rect 360 -1530 366 -1524
rect 360 -1536 366 -1530
rect 360 -1542 366 -1536
rect 360 -1548 366 -1542
rect 360 -1554 366 -1548
rect 360 -1560 366 -1554
rect 360 -1566 366 -1560
rect 360 -1572 366 -1566
rect 360 -1578 366 -1572
rect 360 -1584 366 -1578
rect 360 -1590 366 -1584
rect 360 -1596 366 -1590
rect 360 -1602 366 -1596
rect 360 -1608 366 -1602
rect 360 -1614 366 -1608
rect 360 -1620 366 -1614
rect 360 -1626 366 -1620
rect 360 -1632 366 -1626
rect 360 -1638 366 -1632
rect 360 -1644 366 -1638
rect 360 -1650 366 -1644
rect 360 -1656 366 -1650
rect 360 -1662 366 -1656
rect 360 -1668 366 -1662
rect 360 -1674 366 -1668
rect 360 -1680 366 -1674
rect 360 -1686 366 -1680
rect 360 -1692 366 -1686
rect 360 -1698 366 -1692
rect 360 -1704 366 -1698
rect 360 -1710 366 -1704
rect 360 -1716 366 -1710
rect 360 -1722 366 -1716
rect 360 -1728 366 -1722
rect 360 -1734 366 -1728
rect 360 -1740 366 -1734
rect 360 -1746 366 -1740
rect 360 -1752 366 -1746
rect 360 -1758 366 -1752
rect 360 -1764 366 -1758
rect 360 -1770 366 -1764
rect 360 -1776 366 -1770
rect 360 -2850 366 -2844
rect 360 -2856 366 -2850
rect 360 -2862 366 -2856
rect 360 -2868 366 -2862
rect 360 -2874 366 -2868
rect 360 -2880 366 -2874
rect 360 -2886 366 -2880
rect 360 -2892 366 -2886
rect 360 -2898 366 -2892
rect 360 -2904 366 -2898
rect 360 -2910 366 -2904
rect 360 -2916 366 -2910
rect 360 -2922 366 -2916
rect 360 -2928 366 -2922
rect 360 -2934 366 -2928
rect 360 -2940 366 -2934
rect 360 -2946 366 -2940
rect 360 -2952 366 -2946
rect 360 -2958 366 -2952
rect 360 -2964 366 -2958
rect 360 -2970 366 -2964
rect 360 -2976 366 -2970
rect 360 -2982 366 -2976
rect 360 -2988 366 -2982
rect 360 -2994 366 -2988
rect 360 -3000 366 -2994
rect 360 -3006 366 -3000
rect 360 -3012 366 -3006
rect 360 -3018 366 -3012
rect 360 -3024 366 -3018
rect 360 -3030 366 -3024
rect 360 -3036 366 -3030
rect 360 -3042 366 -3036
rect 360 -3048 366 -3042
rect 360 -3054 366 -3048
rect 360 -3060 366 -3054
rect 360 -3066 366 -3060
rect 360 -3072 366 -3066
rect 360 -3078 366 -3072
rect 360 -3084 366 -3078
rect 360 -3090 366 -3084
rect 360 -3096 366 -3090
rect 360 -3102 366 -3096
rect 360 -3108 366 -3102
rect 360 -3114 366 -3108
rect 360 -3120 366 -3114
rect 360 -3126 366 -3120
rect 360 -3132 366 -3126
rect 360 -3138 366 -3132
rect 360 -3144 366 -3138
rect 360 -3150 366 -3144
rect 360 -3156 366 -3150
rect 360 -3162 366 -3156
rect 360 -3168 366 -3162
rect 360 -3174 366 -3168
rect 366 -1446 372 -1440
rect 366 -1452 372 -1446
rect 366 -1458 372 -1452
rect 366 -1464 372 -1458
rect 366 -1470 372 -1464
rect 366 -1476 372 -1470
rect 366 -1482 372 -1476
rect 366 -1488 372 -1482
rect 366 -1494 372 -1488
rect 366 -1500 372 -1494
rect 366 -1506 372 -1500
rect 366 -1512 372 -1506
rect 366 -1518 372 -1512
rect 366 -1524 372 -1518
rect 366 -1530 372 -1524
rect 366 -1536 372 -1530
rect 366 -1542 372 -1536
rect 366 -1548 372 -1542
rect 366 -1554 372 -1548
rect 366 -1560 372 -1554
rect 366 -1566 372 -1560
rect 366 -1572 372 -1566
rect 366 -1578 372 -1572
rect 366 -1584 372 -1578
rect 366 -1590 372 -1584
rect 366 -1596 372 -1590
rect 366 -1602 372 -1596
rect 366 -1608 372 -1602
rect 366 -1614 372 -1608
rect 366 -1620 372 -1614
rect 366 -1626 372 -1620
rect 366 -1632 372 -1626
rect 366 -1638 372 -1632
rect 366 -1644 372 -1638
rect 366 -1650 372 -1644
rect 366 -1656 372 -1650
rect 366 -1662 372 -1656
rect 366 -1668 372 -1662
rect 366 -1674 372 -1668
rect 366 -1680 372 -1674
rect 366 -1686 372 -1680
rect 366 -1692 372 -1686
rect 366 -1698 372 -1692
rect 366 -1704 372 -1698
rect 366 -1710 372 -1704
rect 366 -1716 372 -1710
rect 366 -1722 372 -1716
rect 366 -1728 372 -1722
rect 366 -1734 372 -1728
rect 366 -1740 372 -1734
rect 366 -1746 372 -1740
rect 366 -1752 372 -1746
rect 366 -1758 372 -1752
rect 366 -1764 372 -1758
rect 366 -1770 372 -1764
rect 366 -2856 372 -2850
rect 366 -2862 372 -2856
rect 366 -2868 372 -2862
rect 366 -2874 372 -2868
rect 366 -2880 372 -2874
rect 366 -2886 372 -2880
rect 366 -2892 372 -2886
rect 366 -2898 372 -2892
rect 366 -2904 372 -2898
rect 366 -2910 372 -2904
rect 366 -2916 372 -2910
rect 366 -2922 372 -2916
rect 366 -2928 372 -2922
rect 366 -2934 372 -2928
rect 366 -2940 372 -2934
rect 366 -2946 372 -2940
rect 366 -2952 372 -2946
rect 366 -2958 372 -2952
rect 366 -2964 372 -2958
rect 366 -2970 372 -2964
rect 366 -2976 372 -2970
rect 366 -2982 372 -2976
rect 366 -2988 372 -2982
rect 366 -2994 372 -2988
rect 366 -3000 372 -2994
rect 366 -3006 372 -3000
rect 366 -3012 372 -3006
rect 366 -3018 372 -3012
rect 366 -3024 372 -3018
rect 366 -3030 372 -3024
rect 366 -3036 372 -3030
rect 366 -3042 372 -3036
rect 366 -3048 372 -3042
rect 366 -3054 372 -3048
rect 366 -3060 372 -3054
rect 366 -3066 372 -3060
rect 366 -3072 372 -3066
rect 366 -3078 372 -3072
rect 366 -3084 372 -3078
rect 366 -3090 372 -3084
rect 366 -3096 372 -3090
rect 366 -3102 372 -3096
rect 366 -3108 372 -3102
rect 366 -3114 372 -3108
rect 366 -3120 372 -3114
rect 366 -3126 372 -3120
rect 366 -3132 372 -3126
rect 366 -3138 372 -3132
rect 366 -3144 372 -3138
rect 366 -3150 372 -3144
rect 366 -3156 372 -3150
rect 366 -3162 372 -3156
rect 366 -3168 372 -3162
rect 366 -3174 372 -3168
rect 366 -3180 372 -3174
rect 372 -1440 378 -1434
rect 372 -1446 378 -1440
rect 372 -1452 378 -1446
rect 372 -1458 378 -1452
rect 372 -1464 378 -1458
rect 372 -1470 378 -1464
rect 372 -1476 378 -1470
rect 372 -1482 378 -1476
rect 372 -1488 378 -1482
rect 372 -1494 378 -1488
rect 372 -1500 378 -1494
rect 372 -1506 378 -1500
rect 372 -1512 378 -1506
rect 372 -1518 378 -1512
rect 372 -1524 378 -1518
rect 372 -1530 378 -1524
rect 372 -1536 378 -1530
rect 372 -1542 378 -1536
rect 372 -1548 378 -1542
rect 372 -1554 378 -1548
rect 372 -1560 378 -1554
rect 372 -1566 378 -1560
rect 372 -1572 378 -1566
rect 372 -1578 378 -1572
rect 372 -1584 378 -1578
rect 372 -1590 378 -1584
rect 372 -1596 378 -1590
rect 372 -1602 378 -1596
rect 372 -1608 378 -1602
rect 372 -1614 378 -1608
rect 372 -1620 378 -1614
rect 372 -1626 378 -1620
rect 372 -1632 378 -1626
rect 372 -1638 378 -1632
rect 372 -1644 378 -1638
rect 372 -1650 378 -1644
rect 372 -1656 378 -1650
rect 372 -1662 378 -1656
rect 372 -1668 378 -1662
rect 372 -1674 378 -1668
rect 372 -1680 378 -1674
rect 372 -1686 378 -1680
rect 372 -1692 378 -1686
rect 372 -1698 378 -1692
rect 372 -1704 378 -1698
rect 372 -1710 378 -1704
rect 372 -1716 378 -1710
rect 372 -1722 378 -1716
rect 372 -1728 378 -1722
rect 372 -1734 378 -1728
rect 372 -1740 378 -1734
rect 372 -1746 378 -1740
rect 372 -1752 378 -1746
rect 372 -1758 378 -1752
rect 372 -2868 378 -2862
rect 372 -2874 378 -2868
rect 372 -2880 378 -2874
rect 372 -2886 378 -2880
rect 372 -2892 378 -2886
rect 372 -2898 378 -2892
rect 372 -2904 378 -2898
rect 372 -2910 378 -2904
rect 372 -2916 378 -2910
rect 372 -2922 378 -2916
rect 372 -2928 378 -2922
rect 372 -2934 378 -2928
rect 372 -2940 378 -2934
rect 372 -2946 378 -2940
rect 372 -2952 378 -2946
rect 372 -2958 378 -2952
rect 372 -2964 378 -2958
rect 372 -2970 378 -2964
rect 372 -2976 378 -2970
rect 372 -2982 378 -2976
rect 372 -2988 378 -2982
rect 372 -2994 378 -2988
rect 372 -3000 378 -2994
rect 372 -3006 378 -3000
rect 372 -3012 378 -3006
rect 372 -3018 378 -3012
rect 372 -3024 378 -3018
rect 372 -3030 378 -3024
rect 372 -3036 378 -3030
rect 372 -3042 378 -3036
rect 372 -3048 378 -3042
rect 372 -3054 378 -3048
rect 372 -3060 378 -3054
rect 372 -3066 378 -3060
rect 372 -3072 378 -3066
rect 372 -3078 378 -3072
rect 372 -3084 378 -3078
rect 372 -3090 378 -3084
rect 372 -3096 378 -3090
rect 372 -3102 378 -3096
rect 372 -3108 378 -3102
rect 372 -3114 378 -3108
rect 372 -3120 378 -3114
rect 372 -3126 378 -3120
rect 372 -3132 378 -3126
rect 372 -3138 378 -3132
rect 372 -3144 378 -3138
rect 372 -3150 378 -3144
rect 372 -3156 378 -3150
rect 372 -3162 378 -3156
rect 372 -3168 378 -3162
rect 372 -3174 378 -3168
rect 372 -3180 378 -3174
rect 372 -3186 378 -3180
rect 378 -1434 384 -1428
rect 378 -1440 384 -1434
rect 378 -1446 384 -1440
rect 378 -1452 384 -1446
rect 378 -1458 384 -1452
rect 378 -1464 384 -1458
rect 378 -1470 384 -1464
rect 378 -1476 384 -1470
rect 378 -1482 384 -1476
rect 378 -1488 384 -1482
rect 378 -1494 384 -1488
rect 378 -1500 384 -1494
rect 378 -1506 384 -1500
rect 378 -1512 384 -1506
rect 378 -1518 384 -1512
rect 378 -1524 384 -1518
rect 378 -1530 384 -1524
rect 378 -1536 384 -1530
rect 378 -1542 384 -1536
rect 378 -1548 384 -1542
rect 378 -1554 384 -1548
rect 378 -1560 384 -1554
rect 378 -1566 384 -1560
rect 378 -1572 384 -1566
rect 378 -1578 384 -1572
rect 378 -1584 384 -1578
rect 378 -1590 384 -1584
rect 378 -1596 384 -1590
rect 378 -1602 384 -1596
rect 378 -1608 384 -1602
rect 378 -1614 384 -1608
rect 378 -1620 384 -1614
rect 378 -1626 384 -1620
rect 378 -1632 384 -1626
rect 378 -1638 384 -1632
rect 378 -1644 384 -1638
rect 378 -1650 384 -1644
rect 378 -1656 384 -1650
rect 378 -1662 384 -1656
rect 378 -1668 384 -1662
rect 378 -1674 384 -1668
rect 378 -1680 384 -1674
rect 378 -1686 384 -1680
rect 378 -1692 384 -1686
rect 378 -1698 384 -1692
rect 378 -1704 384 -1698
rect 378 -1710 384 -1704
rect 378 -1716 384 -1710
rect 378 -1722 384 -1716
rect 378 -1728 384 -1722
rect 378 -1734 384 -1728
rect 378 -1740 384 -1734
rect 378 -1746 384 -1740
rect 378 -1752 384 -1746
rect 378 -2880 384 -2874
rect 378 -2886 384 -2880
rect 378 -2892 384 -2886
rect 378 -2898 384 -2892
rect 378 -2904 384 -2898
rect 378 -2910 384 -2904
rect 378 -2916 384 -2910
rect 378 -2922 384 -2916
rect 378 -2928 384 -2922
rect 378 -2934 384 -2928
rect 378 -2940 384 -2934
rect 378 -2946 384 -2940
rect 378 -2952 384 -2946
rect 378 -2958 384 -2952
rect 378 -2964 384 -2958
rect 378 -2970 384 -2964
rect 378 -2976 384 -2970
rect 378 -2982 384 -2976
rect 378 -2988 384 -2982
rect 378 -2994 384 -2988
rect 378 -3000 384 -2994
rect 378 -3006 384 -3000
rect 378 -3012 384 -3006
rect 378 -3018 384 -3012
rect 378 -3024 384 -3018
rect 378 -3030 384 -3024
rect 378 -3036 384 -3030
rect 378 -3042 384 -3036
rect 378 -3048 384 -3042
rect 378 -3054 384 -3048
rect 378 -3060 384 -3054
rect 378 -3066 384 -3060
rect 378 -3072 384 -3066
rect 378 -3078 384 -3072
rect 378 -3084 384 -3078
rect 378 -3090 384 -3084
rect 378 -3096 384 -3090
rect 378 -3102 384 -3096
rect 378 -3108 384 -3102
rect 378 -3114 384 -3108
rect 378 -3120 384 -3114
rect 378 -3126 384 -3120
rect 378 -3132 384 -3126
rect 378 -3138 384 -3132
rect 378 -3144 384 -3138
rect 378 -3150 384 -3144
rect 378 -3156 384 -3150
rect 378 -3162 384 -3156
rect 378 -3168 384 -3162
rect 378 -3174 384 -3168
rect 378 -3180 384 -3174
rect 378 -3186 384 -3180
rect 378 -3192 384 -3186
rect 384 -1428 390 -1422
rect 384 -1434 390 -1428
rect 384 -1440 390 -1434
rect 384 -1446 390 -1440
rect 384 -1452 390 -1446
rect 384 -1458 390 -1452
rect 384 -1464 390 -1458
rect 384 -1470 390 -1464
rect 384 -1476 390 -1470
rect 384 -1482 390 -1476
rect 384 -1488 390 -1482
rect 384 -1494 390 -1488
rect 384 -1500 390 -1494
rect 384 -1506 390 -1500
rect 384 -1512 390 -1506
rect 384 -1518 390 -1512
rect 384 -1524 390 -1518
rect 384 -1530 390 -1524
rect 384 -1536 390 -1530
rect 384 -1542 390 -1536
rect 384 -1548 390 -1542
rect 384 -1554 390 -1548
rect 384 -1560 390 -1554
rect 384 -1566 390 -1560
rect 384 -1572 390 -1566
rect 384 -1578 390 -1572
rect 384 -1584 390 -1578
rect 384 -1590 390 -1584
rect 384 -1596 390 -1590
rect 384 -1602 390 -1596
rect 384 -1608 390 -1602
rect 384 -1614 390 -1608
rect 384 -1620 390 -1614
rect 384 -1626 390 -1620
rect 384 -1632 390 -1626
rect 384 -1638 390 -1632
rect 384 -1644 390 -1638
rect 384 -1650 390 -1644
rect 384 -1656 390 -1650
rect 384 -1662 390 -1656
rect 384 -1668 390 -1662
rect 384 -1674 390 -1668
rect 384 -1680 390 -1674
rect 384 -1686 390 -1680
rect 384 -1692 390 -1686
rect 384 -1698 390 -1692
rect 384 -1704 390 -1698
rect 384 -1710 390 -1704
rect 384 -1716 390 -1710
rect 384 -1722 390 -1716
rect 384 -1728 390 -1722
rect 384 -1734 390 -1728
rect 384 -1740 390 -1734
rect 384 -2886 390 -2880
rect 384 -2892 390 -2886
rect 384 -2898 390 -2892
rect 384 -2904 390 -2898
rect 384 -2910 390 -2904
rect 384 -2916 390 -2910
rect 384 -2922 390 -2916
rect 384 -2928 390 -2922
rect 384 -2934 390 -2928
rect 384 -2940 390 -2934
rect 384 -2946 390 -2940
rect 384 -2952 390 -2946
rect 384 -2958 390 -2952
rect 384 -2964 390 -2958
rect 384 -2970 390 -2964
rect 384 -2976 390 -2970
rect 384 -2982 390 -2976
rect 384 -2988 390 -2982
rect 384 -2994 390 -2988
rect 384 -3000 390 -2994
rect 384 -3006 390 -3000
rect 384 -3012 390 -3006
rect 384 -3018 390 -3012
rect 384 -3024 390 -3018
rect 384 -3030 390 -3024
rect 384 -3036 390 -3030
rect 384 -3042 390 -3036
rect 384 -3048 390 -3042
rect 384 -3054 390 -3048
rect 384 -3060 390 -3054
rect 384 -3066 390 -3060
rect 384 -3072 390 -3066
rect 384 -3078 390 -3072
rect 384 -3084 390 -3078
rect 384 -3090 390 -3084
rect 384 -3096 390 -3090
rect 384 -3102 390 -3096
rect 384 -3108 390 -3102
rect 384 -3114 390 -3108
rect 384 -3120 390 -3114
rect 384 -3126 390 -3120
rect 384 -3132 390 -3126
rect 384 -3138 390 -3132
rect 384 -3144 390 -3138
rect 384 -3150 390 -3144
rect 384 -3156 390 -3150
rect 384 -3162 390 -3156
rect 384 -3168 390 -3162
rect 384 -3174 390 -3168
rect 384 -3180 390 -3174
rect 384 -3186 390 -3180
rect 384 -3192 390 -3186
rect 384 -3198 390 -3192
rect 390 -1422 396 -1416
rect 390 -1428 396 -1422
rect 390 -1434 396 -1428
rect 390 -1440 396 -1434
rect 390 -1446 396 -1440
rect 390 -1452 396 -1446
rect 390 -1458 396 -1452
rect 390 -1464 396 -1458
rect 390 -1470 396 -1464
rect 390 -1476 396 -1470
rect 390 -1482 396 -1476
rect 390 -1488 396 -1482
rect 390 -1494 396 -1488
rect 390 -1500 396 -1494
rect 390 -1506 396 -1500
rect 390 -1512 396 -1506
rect 390 -1518 396 -1512
rect 390 -1524 396 -1518
rect 390 -1530 396 -1524
rect 390 -1536 396 -1530
rect 390 -1542 396 -1536
rect 390 -1548 396 -1542
rect 390 -1554 396 -1548
rect 390 -1560 396 -1554
rect 390 -1566 396 -1560
rect 390 -1572 396 -1566
rect 390 -1578 396 -1572
rect 390 -1584 396 -1578
rect 390 -1590 396 -1584
rect 390 -1596 396 -1590
rect 390 -1602 396 -1596
rect 390 -1608 396 -1602
rect 390 -1614 396 -1608
rect 390 -1620 396 -1614
rect 390 -1626 396 -1620
rect 390 -1632 396 -1626
rect 390 -1638 396 -1632
rect 390 -1644 396 -1638
rect 390 -1650 396 -1644
rect 390 -1656 396 -1650
rect 390 -1662 396 -1656
rect 390 -1668 396 -1662
rect 390 -1674 396 -1668
rect 390 -1680 396 -1674
rect 390 -1686 396 -1680
rect 390 -1692 396 -1686
rect 390 -1698 396 -1692
rect 390 -1704 396 -1698
rect 390 -1710 396 -1704
rect 390 -1716 396 -1710
rect 390 -1722 396 -1716
rect 390 -1728 396 -1722
rect 390 -1734 396 -1728
rect 390 -2892 396 -2886
rect 390 -2898 396 -2892
rect 390 -2904 396 -2898
rect 390 -2910 396 -2904
rect 390 -2916 396 -2910
rect 390 -2922 396 -2916
rect 390 -2928 396 -2922
rect 390 -2934 396 -2928
rect 390 -2940 396 -2934
rect 390 -2946 396 -2940
rect 390 -2952 396 -2946
rect 390 -2958 396 -2952
rect 390 -2964 396 -2958
rect 390 -2970 396 -2964
rect 390 -2976 396 -2970
rect 390 -2982 396 -2976
rect 390 -2988 396 -2982
rect 390 -2994 396 -2988
rect 390 -3000 396 -2994
rect 390 -3006 396 -3000
rect 390 -3012 396 -3006
rect 390 -3018 396 -3012
rect 390 -3024 396 -3018
rect 390 -3030 396 -3024
rect 390 -3036 396 -3030
rect 390 -3042 396 -3036
rect 390 -3048 396 -3042
rect 390 -3054 396 -3048
rect 390 -3060 396 -3054
rect 390 -3066 396 -3060
rect 390 -3072 396 -3066
rect 390 -3078 396 -3072
rect 390 -3084 396 -3078
rect 390 -3090 396 -3084
rect 390 -3096 396 -3090
rect 390 -3102 396 -3096
rect 390 -3108 396 -3102
rect 390 -3114 396 -3108
rect 390 -3120 396 -3114
rect 390 -3126 396 -3120
rect 390 -3132 396 -3126
rect 390 -3138 396 -3132
rect 390 -3144 396 -3138
rect 390 -3150 396 -3144
rect 390 -3156 396 -3150
rect 390 -3162 396 -3156
rect 390 -3168 396 -3162
rect 390 -3174 396 -3168
rect 390 -3180 396 -3174
rect 390 -3186 396 -3180
rect 390 -3192 396 -3186
rect 390 -3198 396 -3192
rect 390 -3204 396 -3198
rect 396 -1416 402 -1410
rect 396 -1422 402 -1416
rect 396 -1428 402 -1422
rect 396 -1434 402 -1428
rect 396 -1440 402 -1434
rect 396 -1446 402 -1440
rect 396 -1452 402 -1446
rect 396 -1458 402 -1452
rect 396 -1464 402 -1458
rect 396 -1470 402 -1464
rect 396 -1476 402 -1470
rect 396 -1482 402 -1476
rect 396 -1488 402 -1482
rect 396 -1494 402 -1488
rect 396 -1500 402 -1494
rect 396 -1506 402 -1500
rect 396 -1512 402 -1506
rect 396 -1518 402 -1512
rect 396 -1524 402 -1518
rect 396 -1530 402 -1524
rect 396 -1536 402 -1530
rect 396 -1542 402 -1536
rect 396 -1548 402 -1542
rect 396 -1554 402 -1548
rect 396 -1560 402 -1554
rect 396 -1566 402 -1560
rect 396 -1572 402 -1566
rect 396 -1578 402 -1572
rect 396 -1584 402 -1578
rect 396 -1590 402 -1584
rect 396 -1596 402 -1590
rect 396 -1602 402 -1596
rect 396 -1608 402 -1602
rect 396 -1614 402 -1608
rect 396 -1620 402 -1614
rect 396 -1626 402 -1620
rect 396 -1632 402 -1626
rect 396 -1638 402 -1632
rect 396 -1644 402 -1638
rect 396 -1650 402 -1644
rect 396 -1656 402 -1650
rect 396 -1662 402 -1656
rect 396 -1668 402 -1662
rect 396 -1674 402 -1668
rect 396 -1680 402 -1674
rect 396 -1686 402 -1680
rect 396 -1692 402 -1686
rect 396 -1698 402 -1692
rect 396 -1704 402 -1698
rect 396 -1710 402 -1704
rect 396 -1716 402 -1710
rect 396 -1722 402 -1716
rect 396 -2904 402 -2898
rect 396 -2910 402 -2904
rect 396 -2916 402 -2910
rect 396 -2922 402 -2916
rect 396 -2928 402 -2922
rect 396 -2934 402 -2928
rect 396 -2940 402 -2934
rect 396 -2946 402 -2940
rect 396 -2952 402 -2946
rect 396 -2958 402 -2952
rect 396 -2964 402 -2958
rect 396 -2970 402 -2964
rect 396 -2976 402 -2970
rect 396 -2982 402 -2976
rect 396 -2988 402 -2982
rect 396 -2994 402 -2988
rect 396 -3000 402 -2994
rect 396 -3006 402 -3000
rect 396 -3012 402 -3006
rect 396 -3018 402 -3012
rect 396 -3024 402 -3018
rect 396 -3030 402 -3024
rect 396 -3036 402 -3030
rect 396 -3042 402 -3036
rect 396 -3048 402 -3042
rect 396 -3054 402 -3048
rect 396 -3060 402 -3054
rect 396 -3066 402 -3060
rect 396 -3072 402 -3066
rect 396 -3078 402 -3072
rect 396 -3084 402 -3078
rect 396 -3090 402 -3084
rect 396 -3096 402 -3090
rect 396 -3102 402 -3096
rect 396 -3108 402 -3102
rect 396 -3114 402 -3108
rect 396 -3120 402 -3114
rect 396 -3126 402 -3120
rect 396 -3132 402 -3126
rect 396 -3138 402 -3132
rect 396 -3144 402 -3138
rect 396 -3150 402 -3144
rect 396 -3156 402 -3150
rect 396 -3162 402 -3156
rect 396 -3168 402 -3162
rect 396 -3174 402 -3168
rect 396 -3180 402 -3174
rect 396 -3186 402 -3180
rect 396 -3192 402 -3186
rect 396 -3198 402 -3192
rect 396 -3204 402 -3198
rect 396 -3210 402 -3204
rect 402 -1410 408 -1404
rect 402 -1416 408 -1410
rect 402 -1422 408 -1416
rect 402 -1428 408 -1422
rect 402 -1434 408 -1428
rect 402 -1440 408 -1434
rect 402 -1446 408 -1440
rect 402 -1452 408 -1446
rect 402 -1458 408 -1452
rect 402 -1464 408 -1458
rect 402 -1470 408 -1464
rect 402 -1476 408 -1470
rect 402 -1482 408 -1476
rect 402 -1488 408 -1482
rect 402 -1494 408 -1488
rect 402 -1500 408 -1494
rect 402 -1506 408 -1500
rect 402 -1512 408 -1506
rect 402 -1518 408 -1512
rect 402 -1524 408 -1518
rect 402 -1530 408 -1524
rect 402 -1536 408 -1530
rect 402 -1542 408 -1536
rect 402 -1548 408 -1542
rect 402 -1554 408 -1548
rect 402 -1560 408 -1554
rect 402 -1566 408 -1560
rect 402 -1572 408 -1566
rect 402 -1578 408 -1572
rect 402 -1584 408 -1578
rect 402 -1590 408 -1584
rect 402 -1596 408 -1590
rect 402 -1602 408 -1596
rect 402 -1608 408 -1602
rect 402 -1614 408 -1608
rect 402 -1620 408 -1614
rect 402 -1626 408 -1620
rect 402 -1632 408 -1626
rect 402 -1638 408 -1632
rect 402 -1644 408 -1638
rect 402 -1650 408 -1644
rect 402 -1656 408 -1650
rect 402 -1662 408 -1656
rect 402 -1668 408 -1662
rect 402 -1674 408 -1668
rect 402 -1680 408 -1674
rect 402 -1686 408 -1680
rect 402 -1692 408 -1686
rect 402 -1698 408 -1692
rect 402 -1704 408 -1698
rect 402 -1710 408 -1704
rect 402 -1716 408 -1710
rect 402 -2910 408 -2904
rect 402 -2916 408 -2910
rect 402 -2922 408 -2916
rect 402 -2928 408 -2922
rect 402 -2934 408 -2928
rect 402 -2940 408 -2934
rect 402 -2946 408 -2940
rect 402 -2952 408 -2946
rect 402 -2958 408 -2952
rect 402 -2964 408 -2958
rect 402 -2970 408 -2964
rect 402 -2976 408 -2970
rect 402 -2982 408 -2976
rect 402 -2988 408 -2982
rect 402 -2994 408 -2988
rect 402 -3000 408 -2994
rect 402 -3006 408 -3000
rect 402 -3012 408 -3006
rect 402 -3018 408 -3012
rect 402 -3024 408 -3018
rect 402 -3030 408 -3024
rect 402 -3036 408 -3030
rect 402 -3042 408 -3036
rect 402 -3048 408 -3042
rect 402 -3054 408 -3048
rect 402 -3060 408 -3054
rect 402 -3066 408 -3060
rect 402 -3072 408 -3066
rect 402 -3078 408 -3072
rect 402 -3084 408 -3078
rect 402 -3090 408 -3084
rect 402 -3096 408 -3090
rect 402 -3102 408 -3096
rect 402 -3108 408 -3102
rect 402 -3114 408 -3108
rect 402 -3120 408 -3114
rect 402 -3126 408 -3120
rect 402 -3132 408 -3126
rect 402 -3138 408 -3132
rect 402 -3144 408 -3138
rect 402 -3150 408 -3144
rect 402 -3156 408 -3150
rect 402 -3162 408 -3156
rect 402 -3168 408 -3162
rect 402 -3174 408 -3168
rect 402 -3180 408 -3174
rect 402 -3186 408 -3180
rect 402 -3192 408 -3186
rect 402 -3198 408 -3192
rect 402 -3204 408 -3198
rect 402 -3210 408 -3204
rect 402 -3216 408 -3210
rect 408 -1410 414 -1404
rect 408 -1416 414 -1410
rect 408 -1422 414 -1416
rect 408 -1428 414 -1422
rect 408 -1434 414 -1428
rect 408 -1440 414 -1434
rect 408 -1446 414 -1440
rect 408 -1452 414 -1446
rect 408 -1458 414 -1452
rect 408 -1464 414 -1458
rect 408 -1470 414 -1464
rect 408 -1476 414 -1470
rect 408 -1482 414 -1476
rect 408 -1488 414 -1482
rect 408 -1494 414 -1488
rect 408 -1500 414 -1494
rect 408 -1506 414 -1500
rect 408 -1512 414 -1506
rect 408 -1518 414 -1512
rect 408 -1524 414 -1518
rect 408 -1530 414 -1524
rect 408 -1536 414 -1530
rect 408 -1542 414 -1536
rect 408 -1548 414 -1542
rect 408 -1554 414 -1548
rect 408 -1560 414 -1554
rect 408 -1566 414 -1560
rect 408 -1572 414 -1566
rect 408 -1578 414 -1572
rect 408 -1584 414 -1578
rect 408 -1590 414 -1584
rect 408 -1596 414 -1590
rect 408 -1602 414 -1596
rect 408 -1608 414 -1602
rect 408 -1614 414 -1608
rect 408 -1620 414 -1614
rect 408 -1626 414 -1620
rect 408 -1632 414 -1626
rect 408 -1638 414 -1632
rect 408 -1644 414 -1638
rect 408 -1650 414 -1644
rect 408 -1656 414 -1650
rect 408 -1662 414 -1656
rect 408 -1668 414 -1662
rect 408 -1674 414 -1668
rect 408 -1680 414 -1674
rect 408 -1686 414 -1680
rect 408 -1692 414 -1686
rect 408 -1698 414 -1692
rect 408 -1704 414 -1698
rect 408 -1710 414 -1704
rect 408 -2922 414 -2916
rect 408 -2928 414 -2922
rect 408 -2934 414 -2928
rect 408 -2940 414 -2934
rect 408 -2946 414 -2940
rect 408 -2952 414 -2946
rect 408 -2958 414 -2952
rect 408 -2964 414 -2958
rect 408 -2970 414 -2964
rect 408 -2976 414 -2970
rect 408 -2982 414 -2976
rect 408 -2988 414 -2982
rect 408 -2994 414 -2988
rect 408 -3000 414 -2994
rect 408 -3006 414 -3000
rect 408 -3012 414 -3006
rect 408 -3018 414 -3012
rect 408 -3024 414 -3018
rect 408 -3030 414 -3024
rect 408 -3036 414 -3030
rect 408 -3042 414 -3036
rect 408 -3048 414 -3042
rect 408 -3054 414 -3048
rect 408 -3060 414 -3054
rect 408 -3066 414 -3060
rect 408 -3072 414 -3066
rect 408 -3078 414 -3072
rect 408 -3084 414 -3078
rect 408 -3090 414 -3084
rect 408 -3096 414 -3090
rect 408 -3102 414 -3096
rect 408 -3108 414 -3102
rect 408 -3114 414 -3108
rect 408 -3120 414 -3114
rect 408 -3126 414 -3120
rect 408 -3132 414 -3126
rect 408 -3138 414 -3132
rect 408 -3144 414 -3138
rect 408 -3150 414 -3144
rect 408 -3156 414 -3150
rect 408 -3162 414 -3156
rect 408 -3168 414 -3162
rect 408 -3174 414 -3168
rect 408 -3180 414 -3174
rect 408 -3186 414 -3180
rect 408 -3192 414 -3186
rect 408 -3198 414 -3192
rect 408 -3204 414 -3198
rect 408 -3210 414 -3204
rect 408 -3216 414 -3210
rect 408 -3222 414 -3216
rect 414 -1404 420 -1398
rect 414 -1410 420 -1404
rect 414 -1416 420 -1410
rect 414 -1422 420 -1416
rect 414 -1428 420 -1422
rect 414 -1434 420 -1428
rect 414 -1440 420 -1434
rect 414 -1446 420 -1440
rect 414 -1452 420 -1446
rect 414 -1458 420 -1452
rect 414 -1464 420 -1458
rect 414 -1470 420 -1464
rect 414 -1476 420 -1470
rect 414 -1482 420 -1476
rect 414 -1488 420 -1482
rect 414 -1494 420 -1488
rect 414 -1500 420 -1494
rect 414 -1506 420 -1500
rect 414 -1512 420 -1506
rect 414 -1518 420 -1512
rect 414 -1524 420 -1518
rect 414 -1530 420 -1524
rect 414 -1536 420 -1530
rect 414 -1542 420 -1536
rect 414 -1548 420 -1542
rect 414 -1554 420 -1548
rect 414 -1560 420 -1554
rect 414 -1566 420 -1560
rect 414 -1572 420 -1566
rect 414 -1578 420 -1572
rect 414 -1584 420 -1578
rect 414 -1590 420 -1584
rect 414 -1596 420 -1590
rect 414 -1602 420 -1596
rect 414 -1608 420 -1602
rect 414 -1614 420 -1608
rect 414 -1620 420 -1614
rect 414 -1626 420 -1620
rect 414 -1632 420 -1626
rect 414 -1638 420 -1632
rect 414 -1644 420 -1638
rect 414 -1650 420 -1644
rect 414 -1656 420 -1650
rect 414 -1662 420 -1656
rect 414 -1668 420 -1662
rect 414 -1674 420 -1668
rect 414 -1680 420 -1674
rect 414 -1686 420 -1680
rect 414 -1692 420 -1686
rect 414 -1698 420 -1692
rect 414 -2928 420 -2922
rect 414 -2934 420 -2928
rect 414 -2940 420 -2934
rect 414 -2946 420 -2940
rect 414 -2952 420 -2946
rect 414 -2958 420 -2952
rect 414 -2964 420 -2958
rect 414 -2970 420 -2964
rect 414 -2976 420 -2970
rect 414 -2982 420 -2976
rect 414 -2988 420 -2982
rect 414 -2994 420 -2988
rect 414 -3000 420 -2994
rect 414 -3006 420 -3000
rect 414 -3012 420 -3006
rect 414 -3018 420 -3012
rect 414 -3024 420 -3018
rect 414 -3030 420 -3024
rect 414 -3036 420 -3030
rect 414 -3042 420 -3036
rect 414 -3048 420 -3042
rect 414 -3054 420 -3048
rect 414 -3060 420 -3054
rect 414 -3066 420 -3060
rect 414 -3072 420 -3066
rect 414 -3078 420 -3072
rect 414 -3084 420 -3078
rect 414 -3090 420 -3084
rect 414 -3096 420 -3090
rect 414 -3102 420 -3096
rect 414 -3108 420 -3102
rect 414 -3114 420 -3108
rect 414 -3120 420 -3114
rect 414 -3126 420 -3120
rect 414 -3132 420 -3126
rect 414 -3138 420 -3132
rect 414 -3144 420 -3138
rect 414 -3150 420 -3144
rect 414 -3156 420 -3150
rect 414 -3162 420 -3156
rect 414 -3168 420 -3162
rect 414 -3174 420 -3168
rect 414 -3180 420 -3174
rect 414 -3186 420 -3180
rect 414 -3192 420 -3186
rect 414 -3198 420 -3192
rect 414 -3204 420 -3198
rect 414 -3210 420 -3204
rect 414 -3216 420 -3210
rect 414 -3222 420 -3216
rect 420 -1398 426 -1392
rect 420 -1404 426 -1398
rect 420 -1410 426 -1404
rect 420 -1416 426 -1410
rect 420 -1422 426 -1416
rect 420 -1428 426 -1422
rect 420 -1434 426 -1428
rect 420 -1440 426 -1434
rect 420 -1446 426 -1440
rect 420 -1452 426 -1446
rect 420 -1458 426 -1452
rect 420 -1464 426 -1458
rect 420 -1470 426 -1464
rect 420 -1476 426 -1470
rect 420 -1482 426 -1476
rect 420 -1488 426 -1482
rect 420 -1494 426 -1488
rect 420 -1500 426 -1494
rect 420 -1506 426 -1500
rect 420 -1512 426 -1506
rect 420 -1518 426 -1512
rect 420 -1524 426 -1518
rect 420 -1530 426 -1524
rect 420 -1536 426 -1530
rect 420 -1542 426 -1536
rect 420 -1548 426 -1542
rect 420 -1554 426 -1548
rect 420 -1560 426 -1554
rect 420 -1566 426 -1560
rect 420 -1572 426 -1566
rect 420 -1578 426 -1572
rect 420 -1584 426 -1578
rect 420 -1590 426 -1584
rect 420 -1596 426 -1590
rect 420 -1602 426 -1596
rect 420 -1608 426 -1602
rect 420 -1614 426 -1608
rect 420 -1620 426 -1614
rect 420 -1626 426 -1620
rect 420 -1632 426 -1626
rect 420 -1638 426 -1632
rect 420 -1644 426 -1638
rect 420 -1650 426 -1644
rect 420 -1656 426 -1650
rect 420 -1662 426 -1656
rect 420 -1668 426 -1662
rect 420 -1674 426 -1668
rect 420 -1680 426 -1674
rect 420 -1686 426 -1680
rect 420 -1692 426 -1686
rect 420 -2934 426 -2928
rect 420 -2940 426 -2934
rect 420 -2946 426 -2940
rect 420 -2952 426 -2946
rect 420 -2958 426 -2952
rect 420 -2964 426 -2958
rect 420 -2970 426 -2964
rect 420 -2976 426 -2970
rect 420 -2982 426 -2976
rect 420 -2988 426 -2982
rect 420 -2994 426 -2988
rect 420 -3000 426 -2994
rect 420 -3006 426 -3000
rect 420 -3012 426 -3006
rect 420 -3018 426 -3012
rect 420 -3024 426 -3018
rect 420 -3030 426 -3024
rect 420 -3036 426 -3030
rect 420 -3042 426 -3036
rect 420 -3048 426 -3042
rect 420 -3054 426 -3048
rect 420 -3060 426 -3054
rect 420 -3066 426 -3060
rect 420 -3072 426 -3066
rect 420 -3078 426 -3072
rect 420 -3084 426 -3078
rect 420 -3090 426 -3084
rect 420 -3096 426 -3090
rect 420 -3102 426 -3096
rect 420 -3108 426 -3102
rect 420 -3114 426 -3108
rect 420 -3120 426 -3114
rect 420 -3126 426 -3120
rect 420 -3132 426 -3126
rect 420 -3138 426 -3132
rect 420 -3144 426 -3138
rect 420 -3150 426 -3144
rect 420 -3156 426 -3150
rect 420 -3162 426 -3156
rect 420 -3168 426 -3162
rect 420 -3174 426 -3168
rect 420 -3180 426 -3174
rect 420 -3186 426 -3180
rect 420 -3192 426 -3186
rect 420 -3198 426 -3192
rect 420 -3204 426 -3198
rect 420 -3210 426 -3204
rect 420 -3216 426 -3210
rect 420 -3222 426 -3216
rect 420 -3228 426 -3222
rect 426 -1392 432 -1386
rect 426 -1398 432 -1392
rect 426 -1404 432 -1398
rect 426 -1410 432 -1404
rect 426 -1416 432 -1410
rect 426 -1422 432 -1416
rect 426 -1428 432 -1422
rect 426 -1434 432 -1428
rect 426 -1440 432 -1434
rect 426 -1446 432 -1440
rect 426 -1452 432 -1446
rect 426 -1458 432 -1452
rect 426 -1464 432 -1458
rect 426 -1470 432 -1464
rect 426 -1476 432 -1470
rect 426 -1482 432 -1476
rect 426 -1488 432 -1482
rect 426 -1494 432 -1488
rect 426 -1500 432 -1494
rect 426 -1506 432 -1500
rect 426 -1512 432 -1506
rect 426 -1518 432 -1512
rect 426 -1524 432 -1518
rect 426 -1530 432 -1524
rect 426 -1536 432 -1530
rect 426 -1542 432 -1536
rect 426 -1548 432 -1542
rect 426 -1554 432 -1548
rect 426 -1560 432 -1554
rect 426 -1566 432 -1560
rect 426 -1572 432 -1566
rect 426 -1578 432 -1572
rect 426 -1584 432 -1578
rect 426 -1590 432 -1584
rect 426 -1596 432 -1590
rect 426 -1602 432 -1596
rect 426 -1608 432 -1602
rect 426 -1614 432 -1608
rect 426 -1620 432 -1614
rect 426 -1626 432 -1620
rect 426 -1632 432 -1626
rect 426 -1638 432 -1632
rect 426 -1644 432 -1638
rect 426 -1650 432 -1644
rect 426 -1656 432 -1650
rect 426 -1662 432 -1656
rect 426 -1668 432 -1662
rect 426 -1674 432 -1668
rect 426 -1680 432 -1674
rect 426 -1686 432 -1680
rect 426 -2940 432 -2934
rect 426 -2946 432 -2940
rect 426 -2952 432 -2946
rect 426 -2958 432 -2952
rect 426 -2964 432 -2958
rect 426 -2970 432 -2964
rect 426 -2976 432 -2970
rect 426 -2982 432 -2976
rect 426 -2988 432 -2982
rect 426 -2994 432 -2988
rect 426 -3000 432 -2994
rect 426 -3006 432 -3000
rect 426 -3012 432 -3006
rect 426 -3018 432 -3012
rect 426 -3024 432 -3018
rect 426 -3030 432 -3024
rect 426 -3036 432 -3030
rect 426 -3042 432 -3036
rect 426 -3048 432 -3042
rect 426 -3054 432 -3048
rect 426 -3060 432 -3054
rect 426 -3066 432 -3060
rect 426 -3072 432 -3066
rect 426 -3078 432 -3072
rect 426 -3084 432 -3078
rect 426 -3090 432 -3084
rect 426 -3096 432 -3090
rect 426 -3102 432 -3096
rect 426 -3108 432 -3102
rect 426 -3114 432 -3108
rect 426 -3120 432 -3114
rect 426 -3126 432 -3120
rect 426 -3132 432 -3126
rect 426 -3138 432 -3132
rect 426 -3144 432 -3138
rect 426 -3150 432 -3144
rect 426 -3156 432 -3150
rect 426 -3162 432 -3156
rect 426 -3168 432 -3162
rect 426 -3174 432 -3168
rect 426 -3180 432 -3174
rect 426 -3186 432 -3180
rect 426 -3192 432 -3186
rect 426 -3198 432 -3192
rect 426 -3204 432 -3198
rect 426 -3210 432 -3204
rect 426 -3216 432 -3210
rect 426 -3222 432 -3216
rect 426 -3228 432 -3222
rect 426 -3234 432 -3228
rect 432 -1386 438 -1380
rect 432 -1392 438 -1386
rect 432 -1398 438 -1392
rect 432 -1404 438 -1398
rect 432 -1410 438 -1404
rect 432 -1416 438 -1410
rect 432 -1422 438 -1416
rect 432 -1428 438 -1422
rect 432 -1434 438 -1428
rect 432 -1440 438 -1434
rect 432 -1446 438 -1440
rect 432 -1452 438 -1446
rect 432 -1458 438 -1452
rect 432 -1464 438 -1458
rect 432 -1470 438 -1464
rect 432 -1476 438 -1470
rect 432 -1482 438 -1476
rect 432 -1488 438 -1482
rect 432 -1494 438 -1488
rect 432 -1500 438 -1494
rect 432 -1506 438 -1500
rect 432 -1512 438 -1506
rect 432 -1518 438 -1512
rect 432 -1524 438 -1518
rect 432 -1530 438 -1524
rect 432 -1536 438 -1530
rect 432 -1542 438 -1536
rect 432 -1548 438 -1542
rect 432 -1554 438 -1548
rect 432 -1560 438 -1554
rect 432 -1566 438 -1560
rect 432 -1572 438 -1566
rect 432 -1578 438 -1572
rect 432 -1584 438 -1578
rect 432 -1590 438 -1584
rect 432 -1596 438 -1590
rect 432 -1602 438 -1596
rect 432 -1608 438 -1602
rect 432 -1614 438 -1608
rect 432 -1620 438 -1614
rect 432 -1626 438 -1620
rect 432 -1632 438 -1626
rect 432 -1638 438 -1632
rect 432 -1644 438 -1638
rect 432 -1650 438 -1644
rect 432 -1656 438 -1650
rect 432 -1662 438 -1656
rect 432 -1668 438 -1662
rect 432 -1674 438 -1668
rect 432 -2952 438 -2946
rect 432 -2958 438 -2952
rect 432 -2964 438 -2958
rect 432 -2970 438 -2964
rect 432 -2976 438 -2970
rect 432 -2982 438 -2976
rect 432 -2988 438 -2982
rect 432 -2994 438 -2988
rect 432 -3000 438 -2994
rect 432 -3006 438 -3000
rect 432 -3012 438 -3006
rect 432 -3018 438 -3012
rect 432 -3024 438 -3018
rect 432 -3030 438 -3024
rect 432 -3036 438 -3030
rect 432 -3042 438 -3036
rect 432 -3048 438 -3042
rect 432 -3054 438 -3048
rect 432 -3060 438 -3054
rect 432 -3066 438 -3060
rect 432 -3072 438 -3066
rect 432 -3078 438 -3072
rect 432 -3084 438 -3078
rect 432 -3090 438 -3084
rect 432 -3096 438 -3090
rect 432 -3102 438 -3096
rect 432 -3108 438 -3102
rect 432 -3114 438 -3108
rect 432 -3120 438 -3114
rect 432 -3126 438 -3120
rect 432 -3132 438 -3126
rect 432 -3138 438 -3132
rect 432 -3144 438 -3138
rect 432 -3150 438 -3144
rect 432 -3156 438 -3150
rect 432 -3162 438 -3156
rect 432 -3168 438 -3162
rect 432 -3174 438 -3168
rect 432 -3180 438 -3174
rect 432 -3186 438 -3180
rect 432 -3192 438 -3186
rect 432 -3198 438 -3192
rect 432 -3204 438 -3198
rect 432 -3210 438 -3204
rect 432 -3216 438 -3210
rect 432 -3222 438 -3216
rect 432 -3228 438 -3222
rect 432 -3234 438 -3228
rect 432 -3240 438 -3234
rect 438 -1380 444 -1374
rect 438 -1386 444 -1380
rect 438 -1392 444 -1386
rect 438 -1398 444 -1392
rect 438 -1404 444 -1398
rect 438 -1410 444 -1404
rect 438 -1416 444 -1410
rect 438 -1422 444 -1416
rect 438 -1428 444 -1422
rect 438 -1434 444 -1428
rect 438 -1440 444 -1434
rect 438 -1446 444 -1440
rect 438 -1452 444 -1446
rect 438 -1458 444 -1452
rect 438 -1464 444 -1458
rect 438 -1470 444 -1464
rect 438 -1476 444 -1470
rect 438 -1482 444 -1476
rect 438 -1488 444 -1482
rect 438 -1494 444 -1488
rect 438 -1500 444 -1494
rect 438 -1506 444 -1500
rect 438 -1512 444 -1506
rect 438 -1518 444 -1512
rect 438 -1524 444 -1518
rect 438 -1530 444 -1524
rect 438 -1536 444 -1530
rect 438 -1542 444 -1536
rect 438 -1548 444 -1542
rect 438 -1554 444 -1548
rect 438 -1560 444 -1554
rect 438 -1566 444 -1560
rect 438 -1572 444 -1566
rect 438 -1578 444 -1572
rect 438 -1584 444 -1578
rect 438 -1590 444 -1584
rect 438 -1596 444 -1590
rect 438 -1602 444 -1596
rect 438 -1608 444 -1602
rect 438 -1614 444 -1608
rect 438 -1620 444 -1614
rect 438 -1626 444 -1620
rect 438 -1632 444 -1626
rect 438 -1638 444 -1632
rect 438 -1644 444 -1638
rect 438 -1650 444 -1644
rect 438 -1656 444 -1650
rect 438 -1662 444 -1656
rect 438 -1668 444 -1662
rect 438 -2958 444 -2952
rect 438 -2964 444 -2958
rect 438 -2970 444 -2964
rect 438 -2976 444 -2970
rect 438 -2982 444 -2976
rect 438 -2988 444 -2982
rect 438 -2994 444 -2988
rect 438 -3000 444 -2994
rect 438 -3006 444 -3000
rect 438 -3012 444 -3006
rect 438 -3018 444 -3012
rect 438 -3024 444 -3018
rect 438 -3030 444 -3024
rect 438 -3036 444 -3030
rect 438 -3042 444 -3036
rect 438 -3048 444 -3042
rect 438 -3054 444 -3048
rect 438 -3060 444 -3054
rect 438 -3066 444 -3060
rect 438 -3072 444 -3066
rect 438 -3078 444 -3072
rect 438 -3084 444 -3078
rect 438 -3090 444 -3084
rect 438 -3096 444 -3090
rect 438 -3102 444 -3096
rect 438 -3108 444 -3102
rect 438 -3114 444 -3108
rect 438 -3120 444 -3114
rect 438 -3126 444 -3120
rect 438 -3132 444 -3126
rect 438 -3138 444 -3132
rect 438 -3144 444 -3138
rect 438 -3150 444 -3144
rect 438 -3156 444 -3150
rect 438 -3162 444 -3156
rect 438 -3168 444 -3162
rect 438 -3174 444 -3168
rect 438 -3180 444 -3174
rect 438 -3186 444 -3180
rect 438 -3192 444 -3186
rect 438 -3198 444 -3192
rect 438 -3204 444 -3198
rect 438 -3210 444 -3204
rect 438 -3216 444 -3210
rect 438 -3222 444 -3216
rect 438 -3228 444 -3222
rect 438 -3234 444 -3228
rect 438 -3240 444 -3234
rect 438 -3246 444 -3240
rect 444 -1374 450 -1368
rect 444 -1380 450 -1374
rect 444 -1386 450 -1380
rect 444 -1392 450 -1386
rect 444 -1398 450 -1392
rect 444 -1404 450 -1398
rect 444 -1410 450 -1404
rect 444 -1416 450 -1410
rect 444 -1422 450 -1416
rect 444 -1428 450 -1422
rect 444 -1434 450 -1428
rect 444 -1440 450 -1434
rect 444 -1446 450 -1440
rect 444 -1452 450 -1446
rect 444 -1458 450 -1452
rect 444 -1464 450 -1458
rect 444 -1470 450 -1464
rect 444 -1476 450 -1470
rect 444 -1482 450 -1476
rect 444 -1488 450 -1482
rect 444 -1494 450 -1488
rect 444 -1500 450 -1494
rect 444 -1506 450 -1500
rect 444 -1512 450 -1506
rect 444 -1518 450 -1512
rect 444 -1524 450 -1518
rect 444 -1530 450 -1524
rect 444 -1536 450 -1530
rect 444 -1542 450 -1536
rect 444 -1548 450 -1542
rect 444 -1554 450 -1548
rect 444 -1560 450 -1554
rect 444 -1566 450 -1560
rect 444 -1572 450 -1566
rect 444 -1578 450 -1572
rect 444 -1584 450 -1578
rect 444 -1590 450 -1584
rect 444 -1596 450 -1590
rect 444 -1602 450 -1596
rect 444 -1608 450 -1602
rect 444 -1614 450 -1608
rect 444 -1620 450 -1614
rect 444 -1626 450 -1620
rect 444 -1632 450 -1626
rect 444 -1638 450 -1632
rect 444 -1644 450 -1638
rect 444 -1650 450 -1644
rect 444 -1656 450 -1650
rect 444 -1662 450 -1656
rect 444 -2964 450 -2958
rect 444 -2970 450 -2964
rect 444 -2976 450 -2970
rect 444 -2982 450 -2976
rect 444 -2988 450 -2982
rect 444 -2994 450 -2988
rect 444 -3000 450 -2994
rect 444 -3006 450 -3000
rect 444 -3012 450 -3006
rect 444 -3018 450 -3012
rect 444 -3024 450 -3018
rect 444 -3030 450 -3024
rect 444 -3036 450 -3030
rect 444 -3042 450 -3036
rect 444 -3048 450 -3042
rect 444 -3054 450 -3048
rect 444 -3060 450 -3054
rect 444 -3066 450 -3060
rect 444 -3072 450 -3066
rect 444 -3078 450 -3072
rect 444 -3084 450 -3078
rect 444 -3090 450 -3084
rect 444 -3096 450 -3090
rect 444 -3102 450 -3096
rect 444 -3108 450 -3102
rect 444 -3114 450 -3108
rect 444 -3120 450 -3114
rect 444 -3126 450 -3120
rect 444 -3132 450 -3126
rect 444 -3138 450 -3132
rect 444 -3144 450 -3138
rect 444 -3150 450 -3144
rect 444 -3156 450 -3150
rect 444 -3162 450 -3156
rect 444 -3168 450 -3162
rect 444 -3174 450 -3168
rect 444 -3180 450 -3174
rect 444 -3186 450 -3180
rect 444 -3192 450 -3186
rect 444 -3198 450 -3192
rect 444 -3204 450 -3198
rect 444 -3210 450 -3204
rect 444 -3216 450 -3210
rect 444 -3222 450 -3216
rect 444 -3228 450 -3222
rect 444 -3234 450 -3228
rect 444 -3240 450 -3234
rect 444 -3246 450 -3240
rect 444 -3252 450 -3246
rect 450 -1374 456 -1368
rect 450 -1380 456 -1374
rect 450 -1386 456 -1380
rect 450 -1392 456 -1386
rect 450 -1398 456 -1392
rect 450 -1404 456 -1398
rect 450 -1410 456 -1404
rect 450 -1416 456 -1410
rect 450 -1422 456 -1416
rect 450 -1428 456 -1422
rect 450 -1434 456 -1428
rect 450 -1440 456 -1434
rect 450 -1446 456 -1440
rect 450 -1452 456 -1446
rect 450 -1458 456 -1452
rect 450 -1464 456 -1458
rect 450 -1470 456 -1464
rect 450 -1476 456 -1470
rect 450 -1482 456 -1476
rect 450 -1488 456 -1482
rect 450 -1494 456 -1488
rect 450 -1500 456 -1494
rect 450 -1506 456 -1500
rect 450 -1512 456 -1506
rect 450 -1518 456 -1512
rect 450 -1524 456 -1518
rect 450 -1530 456 -1524
rect 450 -1536 456 -1530
rect 450 -1542 456 -1536
rect 450 -1548 456 -1542
rect 450 -1554 456 -1548
rect 450 -1560 456 -1554
rect 450 -1566 456 -1560
rect 450 -1572 456 -1566
rect 450 -1578 456 -1572
rect 450 -1584 456 -1578
rect 450 -1590 456 -1584
rect 450 -1596 456 -1590
rect 450 -1602 456 -1596
rect 450 -1608 456 -1602
rect 450 -1614 456 -1608
rect 450 -1620 456 -1614
rect 450 -1626 456 -1620
rect 450 -1632 456 -1626
rect 450 -1638 456 -1632
rect 450 -1644 456 -1638
rect 450 -1650 456 -1644
rect 450 -1656 456 -1650
rect 450 -2970 456 -2964
rect 450 -2976 456 -2970
rect 450 -2982 456 -2976
rect 450 -2988 456 -2982
rect 450 -2994 456 -2988
rect 450 -3000 456 -2994
rect 450 -3006 456 -3000
rect 450 -3012 456 -3006
rect 450 -3018 456 -3012
rect 450 -3024 456 -3018
rect 450 -3030 456 -3024
rect 450 -3036 456 -3030
rect 450 -3042 456 -3036
rect 450 -3048 456 -3042
rect 450 -3054 456 -3048
rect 450 -3060 456 -3054
rect 450 -3066 456 -3060
rect 450 -3072 456 -3066
rect 450 -3078 456 -3072
rect 450 -3084 456 -3078
rect 450 -3090 456 -3084
rect 450 -3096 456 -3090
rect 450 -3102 456 -3096
rect 450 -3108 456 -3102
rect 450 -3114 456 -3108
rect 450 -3120 456 -3114
rect 450 -3126 456 -3120
rect 450 -3132 456 -3126
rect 450 -3138 456 -3132
rect 450 -3144 456 -3138
rect 450 -3150 456 -3144
rect 450 -3156 456 -3150
rect 450 -3162 456 -3156
rect 450 -3168 456 -3162
rect 450 -3174 456 -3168
rect 450 -3180 456 -3174
rect 450 -3186 456 -3180
rect 450 -3192 456 -3186
rect 450 -3198 456 -3192
rect 450 -3204 456 -3198
rect 450 -3210 456 -3204
rect 450 -3216 456 -3210
rect 450 -3222 456 -3216
rect 450 -3228 456 -3222
rect 450 -3234 456 -3228
rect 450 -3240 456 -3234
rect 450 -3246 456 -3240
rect 450 -3252 456 -3246
rect 456 -1368 462 -1362
rect 456 -1374 462 -1368
rect 456 -1380 462 -1374
rect 456 -1386 462 -1380
rect 456 -1392 462 -1386
rect 456 -1398 462 -1392
rect 456 -1404 462 -1398
rect 456 -1410 462 -1404
rect 456 -1416 462 -1410
rect 456 -1422 462 -1416
rect 456 -1428 462 -1422
rect 456 -1434 462 -1428
rect 456 -1440 462 -1434
rect 456 -1446 462 -1440
rect 456 -1452 462 -1446
rect 456 -1458 462 -1452
rect 456 -1464 462 -1458
rect 456 -1470 462 -1464
rect 456 -1476 462 -1470
rect 456 -1482 462 -1476
rect 456 -1488 462 -1482
rect 456 -1494 462 -1488
rect 456 -1500 462 -1494
rect 456 -1506 462 -1500
rect 456 -1512 462 -1506
rect 456 -1518 462 -1512
rect 456 -1524 462 -1518
rect 456 -1530 462 -1524
rect 456 -1536 462 -1530
rect 456 -1542 462 -1536
rect 456 -1548 462 -1542
rect 456 -1554 462 -1548
rect 456 -1560 462 -1554
rect 456 -1566 462 -1560
rect 456 -1572 462 -1566
rect 456 -1578 462 -1572
rect 456 -1584 462 -1578
rect 456 -1590 462 -1584
rect 456 -1596 462 -1590
rect 456 -1602 462 -1596
rect 456 -1608 462 -1602
rect 456 -1614 462 -1608
rect 456 -1620 462 -1614
rect 456 -1626 462 -1620
rect 456 -1632 462 -1626
rect 456 -1638 462 -1632
rect 456 -1644 462 -1638
rect 456 -1650 462 -1644
rect 456 -2976 462 -2970
rect 456 -2982 462 -2976
rect 456 -2988 462 -2982
rect 456 -2994 462 -2988
rect 456 -3000 462 -2994
rect 456 -3006 462 -3000
rect 456 -3012 462 -3006
rect 456 -3018 462 -3012
rect 456 -3024 462 -3018
rect 456 -3030 462 -3024
rect 456 -3036 462 -3030
rect 456 -3042 462 -3036
rect 456 -3048 462 -3042
rect 456 -3054 462 -3048
rect 456 -3060 462 -3054
rect 456 -3066 462 -3060
rect 456 -3072 462 -3066
rect 456 -3078 462 -3072
rect 456 -3084 462 -3078
rect 456 -3090 462 -3084
rect 456 -3096 462 -3090
rect 456 -3102 462 -3096
rect 456 -3108 462 -3102
rect 456 -3114 462 -3108
rect 456 -3120 462 -3114
rect 456 -3126 462 -3120
rect 456 -3132 462 -3126
rect 456 -3138 462 -3132
rect 456 -3144 462 -3138
rect 456 -3150 462 -3144
rect 456 -3156 462 -3150
rect 456 -3162 462 -3156
rect 456 -3168 462 -3162
rect 456 -3174 462 -3168
rect 456 -3180 462 -3174
rect 456 -3186 462 -3180
rect 456 -3192 462 -3186
rect 456 -3198 462 -3192
rect 456 -3204 462 -3198
rect 456 -3210 462 -3204
rect 456 -3216 462 -3210
rect 456 -3222 462 -3216
rect 456 -3228 462 -3222
rect 456 -3234 462 -3228
rect 456 -3240 462 -3234
rect 456 -3246 462 -3240
rect 456 -3252 462 -3246
rect 456 -3258 462 -3252
rect 462 -1362 468 -1356
rect 462 -1368 468 -1362
rect 462 -1374 468 -1368
rect 462 -1380 468 -1374
rect 462 -1386 468 -1380
rect 462 -1392 468 -1386
rect 462 -1398 468 -1392
rect 462 -1404 468 -1398
rect 462 -1410 468 -1404
rect 462 -1416 468 -1410
rect 462 -1422 468 -1416
rect 462 -1428 468 -1422
rect 462 -1434 468 -1428
rect 462 -1440 468 -1434
rect 462 -1446 468 -1440
rect 462 -1452 468 -1446
rect 462 -1458 468 -1452
rect 462 -1464 468 -1458
rect 462 -1470 468 -1464
rect 462 -1476 468 -1470
rect 462 -1482 468 -1476
rect 462 -1488 468 -1482
rect 462 -1494 468 -1488
rect 462 -1500 468 -1494
rect 462 -1506 468 -1500
rect 462 -1512 468 -1506
rect 462 -1518 468 -1512
rect 462 -1524 468 -1518
rect 462 -1530 468 -1524
rect 462 -1536 468 -1530
rect 462 -1542 468 -1536
rect 462 -1548 468 -1542
rect 462 -1554 468 -1548
rect 462 -1560 468 -1554
rect 462 -1566 468 -1560
rect 462 -1572 468 -1566
rect 462 -1578 468 -1572
rect 462 -1584 468 -1578
rect 462 -1590 468 -1584
rect 462 -1596 468 -1590
rect 462 -1602 468 -1596
rect 462 -1608 468 -1602
rect 462 -1614 468 -1608
rect 462 -1620 468 -1614
rect 462 -1626 468 -1620
rect 462 -1632 468 -1626
rect 462 -1638 468 -1632
rect 462 -1644 468 -1638
rect 462 -2988 468 -2982
rect 462 -2994 468 -2988
rect 462 -3000 468 -2994
rect 462 -3006 468 -3000
rect 462 -3012 468 -3006
rect 462 -3018 468 -3012
rect 462 -3024 468 -3018
rect 462 -3030 468 -3024
rect 462 -3036 468 -3030
rect 462 -3042 468 -3036
rect 462 -3048 468 -3042
rect 462 -3054 468 -3048
rect 462 -3060 468 -3054
rect 462 -3066 468 -3060
rect 462 -3072 468 -3066
rect 462 -3078 468 -3072
rect 462 -3084 468 -3078
rect 462 -3090 468 -3084
rect 462 -3096 468 -3090
rect 462 -3102 468 -3096
rect 462 -3108 468 -3102
rect 462 -3114 468 -3108
rect 462 -3120 468 -3114
rect 462 -3126 468 -3120
rect 462 -3132 468 -3126
rect 462 -3138 468 -3132
rect 462 -3144 468 -3138
rect 462 -3150 468 -3144
rect 462 -3156 468 -3150
rect 462 -3162 468 -3156
rect 462 -3168 468 -3162
rect 462 -3174 468 -3168
rect 462 -3180 468 -3174
rect 462 -3186 468 -3180
rect 462 -3192 468 -3186
rect 462 -3198 468 -3192
rect 462 -3204 468 -3198
rect 462 -3210 468 -3204
rect 462 -3216 468 -3210
rect 462 -3222 468 -3216
rect 462 -3228 468 -3222
rect 462 -3234 468 -3228
rect 462 -3240 468 -3234
rect 462 -3246 468 -3240
rect 462 -3252 468 -3246
rect 462 -3258 468 -3252
rect 462 -3264 468 -3258
rect 468 -1356 474 -1350
rect 468 -1362 474 -1356
rect 468 -1368 474 -1362
rect 468 -1374 474 -1368
rect 468 -1380 474 -1374
rect 468 -1386 474 -1380
rect 468 -1392 474 -1386
rect 468 -1398 474 -1392
rect 468 -1404 474 -1398
rect 468 -1410 474 -1404
rect 468 -1416 474 -1410
rect 468 -1422 474 -1416
rect 468 -1428 474 -1422
rect 468 -1434 474 -1428
rect 468 -1440 474 -1434
rect 468 -1446 474 -1440
rect 468 -1452 474 -1446
rect 468 -1458 474 -1452
rect 468 -1464 474 -1458
rect 468 -1470 474 -1464
rect 468 -1476 474 -1470
rect 468 -1482 474 -1476
rect 468 -1488 474 -1482
rect 468 -1494 474 -1488
rect 468 -1500 474 -1494
rect 468 -1506 474 -1500
rect 468 -1512 474 -1506
rect 468 -1518 474 -1512
rect 468 -1524 474 -1518
rect 468 -1530 474 -1524
rect 468 -1536 474 -1530
rect 468 -1542 474 -1536
rect 468 -1548 474 -1542
rect 468 -1554 474 -1548
rect 468 -1560 474 -1554
rect 468 -1566 474 -1560
rect 468 -1572 474 -1566
rect 468 -1578 474 -1572
rect 468 -1584 474 -1578
rect 468 -1590 474 -1584
rect 468 -1596 474 -1590
rect 468 -1602 474 -1596
rect 468 -1608 474 -1602
rect 468 -1614 474 -1608
rect 468 -1620 474 -1614
rect 468 -1626 474 -1620
rect 468 -1632 474 -1626
rect 468 -2994 474 -2988
rect 468 -3000 474 -2994
rect 468 -3006 474 -3000
rect 468 -3012 474 -3006
rect 468 -3018 474 -3012
rect 468 -3024 474 -3018
rect 468 -3030 474 -3024
rect 468 -3036 474 -3030
rect 468 -3042 474 -3036
rect 468 -3048 474 -3042
rect 468 -3054 474 -3048
rect 468 -3060 474 -3054
rect 468 -3066 474 -3060
rect 468 -3072 474 -3066
rect 468 -3078 474 -3072
rect 468 -3084 474 -3078
rect 468 -3090 474 -3084
rect 468 -3096 474 -3090
rect 468 -3102 474 -3096
rect 468 -3108 474 -3102
rect 468 -3114 474 -3108
rect 468 -3120 474 -3114
rect 468 -3126 474 -3120
rect 468 -3132 474 -3126
rect 468 -3138 474 -3132
rect 468 -3144 474 -3138
rect 468 -3150 474 -3144
rect 468 -3156 474 -3150
rect 468 -3162 474 -3156
rect 468 -3168 474 -3162
rect 468 -3174 474 -3168
rect 468 -3180 474 -3174
rect 468 -3186 474 -3180
rect 468 -3192 474 -3186
rect 468 -3198 474 -3192
rect 468 -3204 474 -3198
rect 468 -3210 474 -3204
rect 468 -3216 474 -3210
rect 468 -3222 474 -3216
rect 468 -3228 474 -3222
rect 468 -3234 474 -3228
rect 468 -3240 474 -3234
rect 468 -3246 474 -3240
rect 468 -3252 474 -3246
rect 468 -3258 474 -3252
rect 468 -3264 474 -3258
rect 468 -3270 474 -3264
rect 474 -1356 480 -1350
rect 474 -1362 480 -1356
rect 474 -1368 480 -1362
rect 474 -1374 480 -1368
rect 474 -1380 480 -1374
rect 474 -1386 480 -1380
rect 474 -1392 480 -1386
rect 474 -1398 480 -1392
rect 474 -1404 480 -1398
rect 474 -1410 480 -1404
rect 474 -1416 480 -1410
rect 474 -1422 480 -1416
rect 474 -1428 480 -1422
rect 474 -1434 480 -1428
rect 474 -1440 480 -1434
rect 474 -1446 480 -1440
rect 474 -1452 480 -1446
rect 474 -1458 480 -1452
rect 474 -1464 480 -1458
rect 474 -1470 480 -1464
rect 474 -1476 480 -1470
rect 474 -1482 480 -1476
rect 474 -1488 480 -1482
rect 474 -1494 480 -1488
rect 474 -1500 480 -1494
rect 474 -1506 480 -1500
rect 474 -1512 480 -1506
rect 474 -1518 480 -1512
rect 474 -1524 480 -1518
rect 474 -1530 480 -1524
rect 474 -1536 480 -1530
rect 474 -1542 480 -1536
rect 474 -1548 480 -1542
rect 474 -1554 480 -1548
rect 474 -1560 480 -1554
rect 474 -1566 480 -1560
rect 474 -1572 480 -1566
rect 474 -1578 480 -1572
rect 474 -1584 480 -1578
rect 474 -1590 480 -1584
rect 474 -1596 480 -1590
rect 474 -1602 480 -1596
rect 474 -1608 480 -1602
rect 474 -1614 480 -1608
rect 474 -1620 480 -1614
rect 474 -1626 480 -1620
rect 474 -3000 480 -2994
rect 474 -3006 480 -3000
rect 474 -3012 480 -3006
rect 474 -3018 480 -3012
rect 474 -3024 480 -3018
rect 474 -3030 480 -3024
rect 474 -3036 480 -3030
rect 474 -3042 480 -3036
rect 474 -3048 480 -3042
rect 474 -3054 480 -3048
rect 474 -3060 480 -3054
rect 474 -3066 480 -3060
rect 474 -3072 480 -3066
rect 474 -3078 480 -3072
rect 474 -3084 480 -3078
rect 474 -3090 480 -3084
rect 474 -3096 480 -3090
rect 474 -3102 480 -3096
rect 474 -3108 480 -3102
rect 474 -3114 480 -3108
rect 474 -3120 480 -3114
rect 474 -3126 480 -3120
rect 474 -3132 480 -3126
rect 474 -3138 480 -3132
rect 474 -3144 480 -3138
rect 474 -3150 480 -3144
rect 474 -3156 480 -3150
rect 474 -3162 480 -3156
rect 474 -3168 480 -3162
rect 474 -3174 480 -3168
rect 474 -3180 480 -3174
rect 474 -3186 480 -3180
rect 474 -3192 480 -3186
rect 474 -3198 480 -3192
rect 474 -3204 480 -3198
rect 474 -3210 480 -3204
rect 474 -3216 480 -3210
rect 474 -3222 480 -3216
rect 474 -3228 480 -3222
rect 474 -3234 480 -3228
rect 474 -3240 480 -3234
rect 474 -3246 480 -3240
rect 474 -3252 480 -3246
rect 474 -3258 480 -3252
rect 474 -3264 480 -3258
rect 474 -3270 480 -3264
rect 474 -3276 480 -3270
rect 480 -1350 486 -1344
rect 480 -1356 486 -1350
rect 480 -1362 486 -1356
rect 480 -1368 486 -1362
rect 480 -1374 486 -1368
rect 480 -1380 486 -1374
rect 480 -1386 486 -1380
rect 480 -1392 486 -1386
rect 480 -1398 486 -1392
rect 480 -1404 486 -1398
rect 480 -1410 486 -1404
rect 480 -1416 486 -1410
rect 480 -1422 486 -1416
rect 480 -1428 486 -1422
rect 480 -1434 486 -1428
rect 480 -1440 486 -1434
rect 480 -1446 486 -1440
rect 480 -1452 486 -1446
rect 480 -1458 486 -1452
rect 480 -1464 486 -1458
rect 480 -1470 486 -1464
rect 480 -1476 486 -1470
rect 480 -1482 486 -1476
rect 480 -1488 486 -1482
rect 480 -1494 486 -1488
rect 480 -1500 486 -1494
rect 480 -1506 486 -1500
rect 480 -1512 486 -1506
rect 480 -1518 486 -1512
rect 480 -1524 486 -1518
rect 480 -1530 486 -1524
rect 480 -1536 486 -1530
rect 480 -1542 486 -1536
rect 480 -1548 486 -1542
rect 480 -1554 486 -1548
rect 480 -1560 486 -1554
rect 480 -1566 486 -1560
rect 480 -1572 486 -1566
rect 480 -1578 486 -1572
rect 480 -1584 486 -1578
rect 480 -1590 486 -1584
rect 480 -1596 486 -1590
rect 480 -1602 486 -1596
rect 480 -1608 486 -1602
rect 480 -1614 486 -1608
rect 480 -1620 486 -1614
rect 480 -3006 486 -3000
rect 480 -3012 486 -3006
rect 480 -3018 486 -3012
rect 480 -3024 486 -3018
rect 480 -3030 486 -3024
rect 480 -3036 486 -3030
rect 480 -3042 486 -3036
rect 480 -3048 486 -3042
rect 480 -3054 486 -3048
rect 480 -3060 486 -3054
rect 480 -3066 486 -3060
rect 480 -3072 486 -3066
rect 480 -3078 486 -3072
rect 480 -3084 486 -3078
rect 480 -3090 486 -3084
rect 480 -3096 486 -3090
rect 480 -3102 486 -3096
rect 480 -3108 486 -3102
rect 480 -3114 486 -3108
rect 480 -3120 486 -3114
rect 480 -3126 486 -3120
rect 480 -3132 486 -3126
rect 480 -3138 486 -3132
rect 480 -3144 486 -3138
rect 480 -3150 486 -3144
rect 480 -3156 486 -3150
rect 480 -3162 486 -3156
rect 480 -3168 486 -3162
rect 480 -3174 486 -3168
rect 480 -3180 486 -3174
rect 480 -3186 486 -3180
rect 480 -3192 486 -3186
rect 480 -3198 486 -3192
rect 480 -3204 486 -3198
rect 480 -3210 486 -3204
rect 480 -3216 486 -3210
rect 480 -3222 486 -3216
rect 480 -3228 486 -3222
rect 480 -3234 486 -3228
rect 480 -3240 486 -3234
rect 480 -3246 486 -3240
rect 480 -3252 486 -3246
rect 480 -3258 486 -3252
rect 480 -3264 486 -3258
rect 480 -3270 486 -3264
rect 480 -3276 486 -3270
rect 486 -1344 492 -1338
rect 486 -1350 492 -1344
rect 486 -1356 492 -1350
rect 486 -1362 492 -1356
rect 486 -1368 492 -1362
rect 486 -1374 492 -1368
rect 486 -1380 492 -1374
rect 486 -1386 492 -1380
rect 486 -1392 492 -1386
rect 486 -1398 492 -1392
rect 486 -1404 492 -1398
rect 486 -1410 492 -1404
rect 486 -1416 492 -1410
rect 486 -1422 492 -1416
rect 486 -1428 492 -1422
rect 486 -1434 492 -1428
rect 486 -1440 492 -1434
rect 486 -1446 492 -1440
rect 486 -1452 492 -1446
rect 486 -1458 492 -1452
rect 486 -1464 492 -1458
rect 486 -1470 492 -1464
rect 486 -1476 492 -1470
rect 486 -1482 492 -1476
rect 486 -1488 492 -1482
rect 486 -1494 492 -1488
rect 486 -1500 492 -1494
rect 486 -1506 492 -1500
rect 486 -1512 492 -1506
rect 486 -1518 492 -1512
rect 486 -1524 492 -1518
rect 486 -1530 492 -1524
rect 486 -1536 492 -1530
rect 486 -1542 492 -1536
rect 486 -1548 492 -1542
rect 486 -1554 492 -1548
rect 486 -1560 492 -1554
rect 486 -1566 492 -1560
rect 486 -1572 492 -1566
rect 486 -1578 492 -1572
rect 486 -1584 492 -1578
rect 486 -1590 492 -1584
rect 486 -1596 492 -1590
rect 486 -1602 492 -1596
rect 486 -1608 492 -1602
rect 486 -1614 492 -1608
rect 486 -3012 492 -3006
rect 486 -3018 492 -3012
rect 486 -3024 492 -3018
rect 486 -3030 492 -3024
rect 486 -3036 492 -3030
rect 486 -3042 492 -3036
rect 486 -3048 492 -3042
rect 486 -3054 492 -3048
rect 486 -3060 492 -3054
rect 486 -3066 492 -3060
rect 486 -3072 492 -3066
rect 486 -3078 492 -3072
rect 486 -3084 492 -3078
rect 486 -3090 492 -3084
rect 486 -3096 492 -3090
rect 486 -3102 492 -3096
rect 486 -3108 492 -3102
rect 486 -3114 492 -3108
rect 486 -3120 492 -3114
rect 486 -3126 492 -3120
rect 486 -3132 492 -3126
rect 486 -3138 492 -3132
rect 486 -3144 492 -3138
rect 486 -3150 492 -3144
rect 486 -3156 492 -3150
rect 486 -3162 492 -3156
rect 486 -3168 492 -3162
rect 486 -3174 492 -3168
rect 486 -3180 492 -3174
rect 486 -3186 492 -3180
rect 486 -3192 492 -3186
rect 486 -3198 492 -3192
rect 486 -3204 492 -3198
rect 486 -3210 492 -3204
rect 486 -3216 492 -3210
rect 486 -3222 492 -3216
rect 486 -3228 492 -3222
rect 486 -3234 492 -3228
rect 486 -3240 492 -3234
rect 486 -3246 492 -3240
rect 486 -3252 492 -3246
rect 486 -3258 492 -3252
rect 486 -3264 492 -3258
rect 486 -3270 492 -3264
rect 486 -3276 492 -3270
rect 486 -3282 492 -3276
rect 492 -1338 498 -1332
rect 492 -1344 498 -1338
rect 492 -1350 498 -1344
rect 492 -1356 498 -1350
rect 492 -1362 498 -1356
rect 492 -1368 498 -1362
rect 492 -1374 498 -1368
rect 492 -1380 498 -1374
rect 492 -1386 498 -1380
rect 492 -1392 498 -1386
rect 492 -1398 498 -1392
rect 492 -1404 498 -1398
rect 492 -1410 498 -1404
rect 492 -1416 498 -1410
rect 492 -1422 498 -1416
rect 492 -1428 498 -1422
rect 492 -1434 498 -1428
rect 492 -1440 498 -1434
rect 492 -1446 498 -1440
rect 492 -1452 498 -1446
rect 492 -1458 498 -1452
rect 492 -1464 498 -1458
rect 492 -1470 498 -1464
rect 492 -1476 498 -1470
rect 492 -1482 498 -1476
rect 492 -1488 498 -1482
rect 492 -1494 498 -1488
rect 492 -1500 498 -1494
rect 492 -1506 498 -1500
rect 492 -1512 498 -1506
rect 492 -1518 498 -1512
rect 492 -1524 498 -1518
rect 492 -1530 498 -1524
rect 492 -1536 498 -1530
rect 492 -1542 498 -1536
rect 492 -1548 498 -1542
rect 492 -1554 498 -1548
rect 492 -1560 498 -1554
rect 492 -1566 498 -1560
rect 492 -1572 498 -1566
rect 492 -1578 498 -1572
rect 492 -1584 498 -1578
rect 492 -1590 498 -1584
rect 492 -1596 498 -1590
rect 492 -1602 498 -1596
rect 492 -1608 498 -1602
rect 492 -3018 498 -3012
rect 492 -3024 498 -3018
rect 492 -3030 498 -3024
rect 492 -3036 498 -3030
rect 492 -3042 498 -3036
rect 492 -3048 498 -3042
rect 492 -3054 498 -3048
rect 492 -3060 498 -3054
rect 492 -3066 498 -3060
rect 492 -3072 498 -3066
rect 492 -3078 498 -3072
rect 492 -3084 498 -3078
rect 492 -3090 498 -3084
rect 492 -3096 498 -3090
rect 492 -3102 498 -3096
rect 492 -3108 498 -3102
rect 492 -3114 498 -3108
rect 492 -3120 498 -3114
rect 492 -3126 498 -3120
rect 492 -3132 498 -3126
rect 492 -3138 498 -3132
rect 492 -3144 498 -3138
rect 492 -3150 498 -3144
rect 492 -3156 498 -3150
rect 492 -3162 498 -3156
rect 492 -3168 498 -3162
rect 492 -3174 498 -3168
rect 492 -3180 498 -3174
rect 492 -3186 498 -3180
rect 492 -3192 498 -3186
rect 492 -3198 498 -3192
rect 492 -3204 498 -3198
rect 492 -3210 498 -3204
rect 492 -3216 498 -3210
rect 492 -3222 498 -3216
rect 492 -3228 498 -3222
rect 492 -3234 498 -3228
rect 492 -3240 498 -3234
rect 492 -3246 498 -3240
rect 492 -3252 498 -3246
rect 492 -3258 498 -3252
rect 492 -3264 498 -3258
rect 492 -3270 498 -3264
rect 492 -3276 498 -3270
rect 492 -3282 498 -3276
rect 492 -3288 498 -3282
rect 498 -1338 504 -1332
rect 498 -1344 504 -1338
rect 498 -1350 504 -1344
rect 498 -1356 504 -1350
rect 498 -1362 504 -1356
rect 498 -1368 504 -1362
rect 498 -1374 504 -1368
rect 498 -1380 504 -1374
rect 498 -1386 504 -1380
rect 498 -1392 504 -1386
rect 498 -1398 504 -1392
rect 498 -1404 504 -1398
rect 498 -1410 504 -1404
rect 498 -1416 504 -1410
rect 498 -1422 504 -1416
rect 498 -1428 504 -1422
rect 498 -1434 504 -1428
rect 498 -1440 504 -1434
rect 498 -1446 504 -1440
rect 498 -1452 504 -1446
rect 498 -1458 504 -1452
rect 498 -1464 504 -1458
rect 498 -1470 504 -1464
rect 498 -1476 504 -1470
rect 498 -1482 504 -1476
rect 498 -1488 504 -1482
rect 498 -1494 504 -1488
rect 498 -1500 504 -1494
rect 498 -1506 504 -1500
rect 498 -1512 504 -1506
rect 498 -1518 504 -1512
rect 498 -1524 504 -1518
rect 498 -1530 504 -1524
rect 498 -1536 504 -1530
rect 498 -1542 504 -1536
rect 498 -1548 504 -1542
rect 498 -1554 504 -1548
rect 498 -1560 504 -1554
rect 498 -1566 504 -1560
rect 498 -1572 504 -1566
rect 498 -1578 504 -1572
rect 498 -1584 504 -1578
rect 498 -1590 504 -1584
rect 498 -1596 504 -1590
rect 498 -1602 504 -1596
rect 498 -3024 504 -3018
rect 498 -3030 504 -3024
rect 498 -3036 504 -3030
rect 498 -3042 504 -3036
rect 498 -3048 504 -3042
rect 498 -3054 504 -3048
rect 498 -3060 504 -3054
rect 498 -3066 504 -3060
rect 498 -3072 504 -3066
rect 498 -3078 504 -3072
rect 498 -3084 504 -3078
rect 498 -3090 504 -3084
rect 498 -3096 504 -3090
rect 498 -3102 504 -3096
rect 498 -3108 504 -3102
rect 498 -3114 504 -3108
rect 498 -3120 504 -3114
rect 498 -3126 504 -3120
rect 498 -3132 504 -3126
rect 498 -3138 504 -3132
rect 498 -3144 504 -3138
rect 498 -3150 504 -3144
rect 498 -3156 504 -3150
rect 498 -3162 504 -3156
rect 498 -3168 504 -3162
rect 498 -3174 504 -3168
rect 498 -3180 504 -3174
rect 498 -3186 504 -3180
rect 498 -3192 504 -3186
rect 498 -3198 504 -3192
rect 498 -3204 504 -3198
rect 498 -3210 504 -3204
rect 498 -3216 504 -3210
rect 498 -3222 504 -3216
rect 498 -3228 504 -3222
rect 498 -3234 504 -3228
rect 498 -3240 504 -3234
rect 498 -3246 504 -3240
rect 498 -3252 504 -3246
rect 498 -3258 504 -3252
rect 498 -3264 504 -3258
rect 498 -3270 504 -3264
rect 498 -3276 504 -3270
rect 498 -3282 504 -3276
rect 498 -3288 504 -3282
rect 498 -3294 504 -3288
rect 504 -1332 510 -1326
rect 504 -1338 510 -1332
rect 504 -1344 510 -1338
rect 504 -1350 510 -1344
rect 504 -1356 510 -1350
rect 504 -1362 510 -1356
rect 504 -1368 510 -1362
rect 504 -1374 510 -1368
rect 504 -1380 510 -1374
rect 504 -1386 510 -1380
rect 504 -1392 510 -1386
rect 504 -1398 510 -1392
rect 504 -1404 510 -1398
rect 504 -1410 510 -1404
rect 504 -1416 510 -1410
rect 504 -1422 510 -1416
rect 504 -1428 510 -1422
rect 504 -1434 510 -1428
rect 504 -1440 510 -1434
rect 504 -1446 510 -1440
rect 504 -1452 510 -1446
rect 504 -1458 510 -1452
rect 504 -1464 510 -1458
rect 504 -1470 510 -1464
rect 504 -1476 510 -1470
rect 504 -1482 510 -1476
rect 504 -1488 510 -1482
rect 504 -1494 510 -1488
rect 504 -1500 510 -1494
rect 504 -1506 510 -1500
rect 504 -1512 510 -1506
rect 504 -1518 510 -1512
rect 504 -1524 510 -1518
rect 504 -1530 510 -1524
rect 504 -1536 510 -1530
rect 504 -1542 510 -1536
rect 504 -1548 510 -1542
rect 504 -1554 510 -1548
rect 504 -1560 510 -1554
rect 504 -1566 510 -1560
rect 504 -1572 510 -1566
rect 504 -1578 510 -1572
rect 504 -1584 510 -1578
rect 504 -1590 510 -1584
rect 504 -1596 510 -1590
rect 504 -3030 510 -3024
rect 504 -3036 510 -3030
rect 504 -3042 510 -3036
rect 504 -3048 510 -3042
rect 504 -3054 510 -3048
rect 504 -3060 510 -3054
rect 504 -3066 510 -3060
rect 504 -3072 510 -3066
rect 504 -3078 510 -3072
rect 504 -3084 510 -3078
rect 504 -3090 510 -3084
rect 504 -3096 510 -3090
rect 504 -3102 510 -3096
rect 504 -3108 510 -3102
rect 504 -3114 510 -3108
rect 504 -3120 510 -3114
rect 504 -3126 510 -3120
rect 504 -3132 510 -3126
rect 504 -3138 510 -3132
rect 504 -3144 510 -3138
rect 504 -3150 510 -3144
rect 504 -3156 510 -3150
rect 504 -3162 510 -3156
rect 504 -3168 510 -3162
rect 504 -3174 510 -3168
rect 504 -3180 510 -3174
rect 504 -3186 510 -3180
rect 504 -3192 510 -3186
rect 504 -3198 510 -3192
rect 504 -3204 510 -3198
rect 504 -3210 510 -3204
rect 504 -3216 510 -3210
rect 504 -3222 510 -3216
rect 504 -3228 510 -3222
rect 504 -3234 510 -3228
rect 504 -3240 510 -3234
rect 504 -3246 510 -3240
rect 504 -3252 510 -3246
rect 504 -3258 510 -3252
rect 504 -3264 510 -3258
rect 504 -3270 510 -3264
rect 504 -3276 510 -3270
rect 504 -3282 510 -3276
rect 504 -3288 510 -3282
rect 504 -3294 510 -3288
rect 510 -1326 516 -1320
rect 510 -1332 516 -1326
rect 510 -1338 516 -1332
rect 510 -1344 516 -1338
rect 510 -1350 516 -1344
rect 510 -1356 516 -1350
rect 510 -1362 516 -1356
rect 510 -1368 516 -1362
rect 510 -1374 516 -1368
rect 510 -1380 516 -1374
rect 510 -1386 516 -1380
rect 510 -1392 516 -1386
rect 510 -1398 516 -1392
rect 510 -1404 516 -1398
rect 510 -1410 516 -1404
rect 510 -1416 516 -1410
rect 510 -1422 516 -1416
rect 510 -1428 516 -1422
rect 510 -1434 516 -1428
rect 510 -1440 516 -1434
rect 510 -1446 516 -1440
rect 510 -1452 516 -1446
rect 510 -1458 516 -1452
rect 510 -1464 516 -1458
rect 510 -1470 516 -1464
rect 510 -1476 516 -1470
rect 510 -1482 516 -1476
rect 510 -1488 516 -1482
rect 510 -1494 516 -1488
rect 510 -1500 516 -1494
rect 510 -1506 516 -1500
rect 510 -1512 516 -1506
rect 510 -1518 516 -1512
rect 510 -1524 516 -1518
rect 510 -1530 516 -1524
rect 510 -1536 516 -1530
rect 510 -1542 516 -1536
rect 510 -1548 516 -1542
rect 510 -1554 516 -1548
rect 510 -1560 516 -1554
rect 510 -1566 516 -1560
rect 510 -1572 516 -1566
rect 510 -1578 516 -1572
rect 510 -1584 516 -1578
rect 510 -1590 516 -1584
rect 510 -3036 516 -3030
rect 510 -3042 516 -3036
rect 510 -3048 516 -3042
rect 510 -3054 516 -3048
rect 510 -3060 516 -3054
rect 510 -3066 516 -3060
rect 510 -3072 516 -3066
rect 510 -3078 516 -3072
rect 510 -3084 516 -3078
rect 510 -3090 516 -3084
rect 510 -3096 516 -3090
rect 510 -3102 516 -3096
rect 510 -3108 516 -3102
rect 510 -3114 516 -3108
rect 510 -3120 516 -3114
rect 510 -3126 516 -3120
rect 510 -3132 516 -3126
rect 510 -3138 516 -3132
rect 510 -3144 516 -3138
rect 510 -3150 516 -3144
rect 510 -3156 516 -3150
rect 510 -3162 516 -3156
rect 510 -3168 516 -3162
rect 510 -3174 516 -3168
rect 510 -3180 516 -3174
rect 510 -3186 516 -3180
rect 510 -3192 516 -3186
rect 510 -3198 516 -3192
rect 510 -3204 516 -3198
rect 510 -3210 516 -3204
rect 510 -3216 516 -3210
rect 510 -3222 516 -3216
rect 510 -3228 516 -3222
rect 510 -3234 516 -3228
rect 510 -3240 516 -3234
rect 510 -3246 516 -3240
rect 510 -3252 516 -3246
rect 510 -3258 516 -3252
rect 510 -3264 516 -3258
rect 510 -3270 516 -3264
rect 510 -3276 516 -3270
rect 510 -3282 516 -3276
rect 510 -3288 516 -3282
rect 510 -3294 516 -3288
rect 510 -3300 516 -3294
rect 516 -1320 522 -1314
rect 516 -1326 522 -1320
rect 516 -1332 522 -1326
rect 516 -1338 522 -1332
rect 516 -1344 522 -1338
rect 516 -1350 522 -1344
rect 516 -1356 522 -1350
rect 516 -1362 522 -1356
rect 516 -1368 522 -1362
rect 516 -1374 522 -1368
rect 516 -1380 522 -1374
rect 516 -1386 522 -1380
rect 516 -1392 522 -1386
rect 516 -1398 522 -1392
rect 516 -1404 522 -1398
rect 516 -1410 522 -1404
rect 516 -1416 522 -1410
rect 516 -1422 522 -1416
rect 516 -1428 522 -1422
rect 516 -1434 522 -1428
rect 516 -1440 522 -1434
rect 516 -1446 522 -1440
rect 516 -1452 522 -1446
rect 516 -1458 522 -1452
rect 516 -1464 522 -1458
rect 516 -1470 522 -1464
rect 516 -1476 522 -1470
rect 516 -1482 522 -1476
rect 516 -1488 522 -1482
rect 516 -1494 522 -1488
rect 516 -1500 522 -1494
rect 516 -1506 522 -1500
rect 516 -1512 522 -1506
rect 516 -1518 522 -1512
rect 516 -1524 522 -1518
rect 516 -1530 522 -1524
rect 516 -1536 522 -1530
rect 516 -1542 522 -1536
rect 516 -1548 522 -1542
rect 516 -1554 522 -1548
rect 516 -1560 522 -1554
rect 516 -1566 522 -1560
rect 516 -1572 522 -1566
rect 516 -1578 522 -1572
rect 516 -1584 522 -1578
rect 516 -3042 522 -3036
rect 516 -3048 522 -3042
rect 516 -3054 522 -3048
rect 516 -3060 522 -3054
rect 516 -3066 522 -3060
rect 516 -3072 522 -3066
rect 516 -3078 522 -3072
rect 516 -3084 522 -3078
rect 516 -3090 522 -3084
rect 516 -3096 522 -3090
rect 516 -3102 522 -3096
rect 516 -3108 522 -3102
rect 516 -3114 522 -3108
rect 516 -3120 522 -3114
rect 516 -3126 522 -3120
rect 516 -3132 522 -3126
rect 516 -3138 522 -3132
rect 516 -3144 522 -3138
rect 516 -3150 522 -3144
rect 516 -3156 522 -3150
rect 516 -3162 522 -3156
rect 516 -3168 522 -3162
rect 516 -3174 522 -3168
rect 516 -3180 522 -3174
rect 516 -3186 522 -3180
rect 516 -3192 522 -3186
rect 516 -3198 522 -3192
rect 516 -3204 522 -3198
rect 516 -3210 522 -3204
rect 516 -3216 522 -3210
rect 516 -3222 522 -3216
rect 516 -3228 522 -3222
rect 516 -3234 522 -3228
rect 516 -3240 522 -3234
rect 516 -3246 522 -3240
rect 516 -3252 522 -3246
rect 516 -3258 522 -3252
rect 516 -3264 522 -3258
rect 516 -3270 522 -3264
rect 516 -3276 522 -3270
rect 516 -3282 522 -3276
rect 516 -3288 522 -3282
rect 516 -3294 522 -3288
rect 516 -3300 522 -3294
rect 516 -3306 522 -3300
rect 522 -1320 528 -1314
rect 522 -1326 528 -1320
rect 522 -1332 528 -1326
rect 522 -1338 528 -1332
rect 522 -1344 528 -1338
rect 522 -1350 528 -1344
rect 522 -1356 528 -1350
rect 522 -1362 528 -1356
rect 522 -1368 528 -1362
rect 522 -1374 528 -1368
rect 522 -1380 528 -1374
rect 522 -1386 528 -1380
rect 522 -1392 528 -1386
rect 522 -1398 528 -1392
rect 522 -1404 528 -1398
rect 522 -1410 528 -1404
rect 522 -1416 528 -1410
rect 522 -1422 528 -1416
rect 522 -1428 528 -1422
rect 522 -1434 528 -1428
rect 522 -1440 528 -1434
rect 522 -1446 528 -1440
rect 522 -1452 528 -1446
rect 522 -1458 528 -1452
rect 522 -1464 528 -1458
rect 522 -1470 528 -1464
rect 522 -1476 528 -1470
rect 522 -1482 528 -1476
rect 522 -1488 528 -1482
rect 522 -1494 528 -1488
rect 522 -1500 528 -1494
rect 522 -1506 528 -1500
rect 522 -1512 528 -1506
rect 522 -1518 528 -1512
rect 522 -1524 528 -1518
rect 522 -1530 528 -1524
rect 522 -1536 528 -1530
rect 522 -1542 528 -1536
rect 522 -1548 528 -1542
rect 522 -1554 528 -1548
rect 522 -1560 528 -1554
rect 522 -1566 528 -1560
rect 522 -1572 528 -1566
rect 522 -1578 528 -1572
rect 522 -3048 528 -3042
rect 522 -3054 528 -3048
rect 522 -3060 528 -3054
rect 522 -3066 528 -3060
rect 522 -3072 528 -3066
rect 522 -3078 528 -3072
rect 522 -3084 528 -3078
rect 522 -3090 528 -3084
rect 522 -3096 528 -3090
rect 522 -3102 528 -3096
rect 522 -3108 528 -3102
rect 522 -3114 528 -3108
rect 522 -3120 528 -3114
rect 522 -3126 528 -3120
rect 522 -3132 528 -3126
rect 522 -3138 528 -3132
rect 522 -3144 528 -3138
rect 522 -3150 528 -3144
rect 522 -3156 528 -3150
rect 522 -3162 528 -3156
rect 522 -3168 528 -3162
rect 522 -3174 528 -3168
rect 522 -3180 528 -3174
rect 522 -3186 528 -3180
rect 522 -3192 528 -3186
rect 522 -3198 528 -3192
rect 522 -3204 528 -3198
rect 522 -3210 528 -3204
rect 522 -3216 528 -3210
rect 522 -3222 528 -3216
rect 522 -3228 528 -3222
rect 522 -3234 528 -3228
rect 522 -3240 528 -3234
rect 522 -3246 528 -3240
rect 522 -3252 528 -3246
rect 522 -3258 528 -3252
rect 522 -3264 528 -3258
rect 522 -3270 528 -3264
rect 522 -3276 528 -3270
rect 522 -3282 528 -3276
rect 522 -3288 528 -3282
rect 522 -3294 528 -3288
rect 522 -3300 528 -3294
rect 522 -3306 528 -3300
rect 528 -1314 534 -1308
rect 528 -1320 534 -1314
rect 528 -1326 534 -1320
rect 528 -1332 534 -1326
rect 528 -1338 534 -1332
rect 528 -1344 534 -1338
rect 528 -1350 534 -1344
rect 528 -1356 534 -1350
rect 528 -1362 534 -1356
rect 528 -1368 534 -1362
rect 528 -1374 534 -1368
rect 528 -1380 534 -1374
rect 528 -1386 534 -1380
rect 528 -1392 534 -1386
rect 528 -1398 534 -1392
rect 528 -1404 534 -1398
rect 528 -1410 534 -1404
rect 528 -1416 534 -1410
rect 528 -1422 534 -1416
rect 528 -1428 534 -1422
rect 528 -1434 534 -1428
rect 528 -1440 534 -1434
rect 528 -1446 534 -1440
rect 528 -1452 534 -1446
rect 528 -1458 534 -1452
rect 528 -1464 534 -1458
rect 528 -1470 534 -1464
rect 528 -1476 534 -1470
rect 528 -1482 534 -1476
rect 528 -1488 534 -1482
rect 528 -1494 534 -1488
rect 528 -1500 534 -1494
rect 528 -1506 534 -1500
rect 528 -1512 534 -1506
rect 528 -1518 534 -1512
rect 528 -1524 534 -1518
rect 528 -1530 534 -1524
rect 528 -1536 534 -1530
rect 528 -1542 534 -1536
rect 528 -1548 534 -1542
rect 528 -1554 534 -1548
rect 528 -1560 534 -1554
rect 528 -1566 534 -1560
rect 528 -1572 534 -1566
rect 528 -3054 534 -3048
rect 528 -3060 534 -3054
rect 528 -3066 534 -3060
rect 528 -3072 534 -3066
rect 528 -3078 534 -3072
rect 528 -3084 534 -3078
rect 528 -3090 534 -3084
rect 528 -3096 534 -3090
rect 528 -3102 534 -3096
rect 528 -3108 534 -3102
rect 528 -3114 534 -3108
rect 528 -3120 534 -3114
rect 528 -3126 534 -3120
rect 528 -3132 534 -3126
rect 528 -3138 534 -3132
rect 528 -3144 534 -3138
rect 528 -3150 534 -3144
rect 528 -3156 534 -3150
rect 528 -3162 534 -3156
rect 528 -3168 534 -3162
rect 528 -3174 534 -3168
rect 528 -3180 534 -3174
rect 528 -3186 534 -3180
rect 528 -3192 534 -3186
rect 528 -3198 534 -3192
rect 528 -3204 534 -3198
rect 528 -3210 534 -3204
rect 528 -3216 534 -3210
rect 528 -3222 534 -3216
rect 528 -3228 534 -3222
rect 528 -3234 534 -3228
rect 528 -3240 534 -3234
rect 528 -3246 534 -3240
rect 528 -3252 534 -3246
rect 528 -3258 534 -3252
rect 528 -3264 534 -3258
rect 528 -3270 534 -3264
rect 528 -3276 534 -3270
rect 528 -3282 534 -3276
rect 528 -3288 534 -3282
rect 528 -3294 534 -3288
rect 528 -3300 534 -3294
rect 528 -3306 534 -3300
rect 528 -3312 534 -3306
rect 534 -1308 540 -1302
rect 534 -1314 540 -1308
rect 534 -1320 540 -1314
rect 534 -1326 540 -1320
rect 534 -1332 540 -1326
rect 534 -1338 540 -1332
rect 534 -1344 540 -1338
rect 534 -1350 540 -1344
rect 534 -1356 540 -1350
rect 534 -1362 540 -1356
rect 534 -1368 540 -1362
rect 534 -1374 540 -1368
rect 534 -1380 540 -1374
rect 534 -1386 540 -1380
rect 534 -1392 540 -1386
rect 534 -1398 540 -1392
rect 534 -1404 540 -1398
rect 534 -1410 540 -1404
rect 534 -1416 540 -1410
rect 534 -1422 540 -1416
rect 534 -1428 540 -1422
rect 534 -1434 540 -1428
rect 534 -1440 540 -1434
rect 534 -1446 540 -1440
rect 534 -1452 540 -1446
rect 534 -1458 540 -1452
rect 534 -1464 540 -1458
rect 534 -1470 540 -1464
rect 534 -1476 540 -1470
rect 534 -1482 540 -1476
rect 534 -1488 540 -1482
rect 534 -1494 540 -1488
rect 534 -1500 540 -1494
rect 534 -1506 540 -1500
rect 534 -1512 540 -1506
rect 534 -1518 540 -1512
rect 534 -1524 540 -1518
rect 534 -1530 540 -1524
rect 534 -1536 540 -1530
rect 534 -1542 540 -1536
rect 534 -1548 540 -1542
rect 534 -1554 540 -1548
rect 534 -1560 540 -1554
rect 534 -1566 540 -1560
rect 534 -3060 540 -3054
rect 534 -3066 540 -3060
rect 534 -3072 540 -3066
rect 534 -3078 540 -3072
rect 534 -3084 540 -3078
rect 534 -3090 540 -3084
rect 534 -3096 540 -3090
rect 534 -3102 540 -3096
rect 534 -3108 540 -3102
rect 534 -3114 540 -3108
rect 534 -3120 540 -3114
rect 534 -3126 540 -3120
rect 534 -3132 540 -3126
rect 534 -3138 540 -3132
rect 534 -3144 540 -3138
rect 534 -3150 540 -3144
rect 534 -3156 540 -3150
rect 534 -3162 540 -3156
rect 534 -3168 540 -3162
rect 534 -3174 540 -3168
rect 534 -3180 540 -3174
rect 534 -3186 540 -3180
rect 534 -3192 540 -3186
rect 534 -3198 540 -3192
rect 534 -3204 540 -3198
rect 534 -3210 540 -3204
rect 534 -3216 540 -3210
rect 534 -3222 540 -3216
rect 534 -3228 540 -3222
rect 534 -3234 540 -3228
rect 534 -3240 540 -3234
rect 534 -3246 540 -3240
rect 534 -3252 540 -3246
rect 534 -3258 540 -3252
rect 534 -3264 540 -3258
rect 534 -3270 540 -3264
rect 534 -3276 540 -3270
rect 534 -3282 540 -3276
rect 534 -3288 540 -3282
rect 534 -3294 540 -3288
rect 534 -3300 540 -3294
rect 534 -3306 540 -3300
rect 534 -3312 540 -3306
rect 534 -3318 540 -3312
rect 540 -1308 546 -1302
rect 540 -1314 546 -1308
rect 540 -1320 546 -1314
rect 540 -1326 546 -1320
rect 540 -1332 546 -1326
rect 540 -1338 546 -1332
rect 540 -1344 546 -1338
rect 540 -1350 546 -1344
rect 540 -1356 546 -1350
rect 540 -1362 546 -1356
rect 540 -1368 546 -1362
rect 540 -1374 546 -1368
rect 540 -1380 546 -1374
rect 540 -1386 546 -1380
rect 540 -1392 546 -1386
rect 540 -1398 546 -1392
rect 540 -1404 546 -1398
rect 540 -1410 546 -1404
rect 540 -1416 546 -1410
rect 540 -1422 546 -1416
rect 540 -1428 546 -1422
rect 540 -1434 546 -1428
rect 540 -1440 546 -1434
rect 540 -1446 546 -1440
rect 540 -1452 546 -1446
rect 540 -1458 546 -1452
rect 540 -1464 546 -1458
rect 540 -1470 546 -1464
rect 540 -1476 546 -1470
rect 540 -1482 546 -1476
rect 540 -1488 546 -1482
rect 540 -1494 546 -1488
rect 540 -1500 546 -1494
rect 540 -1506 546 -1500
rect 540 -1512 546 -1506
rect 540 -1518 546 -1512
rect 540 -1524 546 -1518
rect 540 -1530 546 -1524
rect 540 -1536 546 -1530
rect 540 -1542 546 -1536
rect 540 -1548 546 -1542
rect 540 -1554 546 -1548
rect 540 -1560 546 -1554
rect 540 -1566 546 -1560
rect 540 -3066 546 -3060
rect 540 -3072 546 -3066
rect 540 -3078 546 -3072
rect 540 -3084 546 -3078
rect 540 -3090 546 -3084
rect 540 -3096 546 -3090
rect 540 -3102 546 -3096
rect 540 -3108 546 -3102
rect 540 -3114 546 -3108
rect 540 -3120 546 -3114
rect 540 -3126 546 -3120
rect 540 -3132 546 -3126
rect 540 -3138 546 -3132
rect 540 -3144 546 -3138
rect 540 -3150 546 -3144
rect 540 -3156 546 -3150
rect 540 -3162 546 -3156
rect 540 -3168 546 -3162
rect 540 -3174 546 -3168
rect 540 -3180 546 -3174
rect 540 -3186 546 -3180
rect 540 -3192 546 -3186
rect 540 -3198 546 -3192
rect 540 -3204 546 -3198
rect 540 -3210 546 -3204
rect 540 -3216 546 -3210
rect 540 -3222 546 -3216
rect 540 -3228 546 -3222
rect 540 -3234 546 -3228
rect 540 -3240 546 -3234
rect 540 -3246 546 -3240
rect 540 -3252 546 -3246
rect 540 -3258 546 -3252
rect 540 -3264 546 -3258
rect 540 -3270 546 -3264
rect 540 -3276 546 -3270
rect 540 -3282 546 -3276
rect 540 -3288 546 -3282
rect 540 -3294 546 -3288
rect 540 -3300 546 -3294
rect 540 -3306 546 -3300
rect 540 -3312 546 -3306
rect 540 -3318 546 -3312
rect 540 -3324 546 -3318
rect 546 -1302 552 -1296
rect 546 -1308 552 -1302
rect 546 -1314 552 -1308
rect 546 -1320 552 -1314
rect 546 -1326 552 -1320
rect 546 -1332 552 -1326
rect 546 -1338 552 -1332
rect 546 -1344 552 -1338
rect 546 -1350 552 -1344
rect 546 -1356 552 -1350
rect 546 -1362 552 -1356
rect 546 -1368 552 -1362
rect 546 -1374 552 -1368
rect 546 -1380 552 -1374
rect 546 -1386 552 -1380
rect 546 -1392 552 -1386
rect 546 -1398 552 -1392
rect 546 -1404 552 -1398
rect 546 -1410 552 -1404
rect 546 -1416 552 -1410
rect 546 -1422 552 -1416
rect 546 -1428 552 -1422
rect 546 -1434 552 -1428
rect 546 -1440 552 -1434
rect 546 -1446 552 -1440
rect 546 -1452 552 -1446
rect 546 -1458 552 -1452
rect 546 -1464 552 -1458
rect 546 -1470 552 -1464
rect 546 -1476 552 -1470
rect 546 -1482 552 -1476
rect 546 -1488 552 -1482
rect 546 -1494 552 -1488
rect 546 -1500 552 -1494
rect 546 -1506 552 -1500
rect 546 -1512 552 -1506
rect 546 -1518 552 -1512
rect 546 -1524 552 -1518
rect 546 -1530 552 -1524
rect 546 -1536 552 -1530
rect 546 -1542 552 -1536
rect 546 -1548 552 -1542
rect 546 -1554 552 -1548
rect 546 -1560 552 -1554
rect 546 -3066 552 -3060
rect 546 -3072 552 -3066
rect 546 -3078 552 -3072
rect 546 -3084 552 -3078
rect 546 -3090 552 -3084
rect 546 -3096 552 -3090
rect 546 -3102 552 -3096
rect 546 -3108 552 -3102
rect 546 -3114 552 -3108
rect 546 -3120 552 -3114
rect 546 -3126 552 -3120
rect 546 -3132 552 -3126
rect 546 -3138 552 -3132
rect 546 -3144 552 -3138
rect 546 -3150 552 -3144
rect 546 -3156 552 -3150
rect 546 -3162 552 -3156
rect 546 -3168 552 -3162
rect 546 -3174 552 -3168
rect 546 -3180 552 -3174
rect 546 -3186 552 -3180
rect 546 -3192 552 -3186
rect 546 -3198 552 -3192
rect 546 -3204 552 -3198
rect 546 -3210 552 -3204
rect 546 -3216 552 -3210
rect 546 -3222 552 -3216
rect 546 -3228 552 -3222
rect 546 -3234 552 -3228
rect 546 -3240 552 -3234
rect 546 -3246 552 -3240
rect 546 -3252 552 -3246
rect 546 -3258 552 -3252
rect 546 -3264 552 -3258
rect 546 -3270 552 -3264
rect 546 -3276 552 -3270
rect 546 -3282 552 -3276
rect 546 -3288 552 -3282
rect 546 -3294 552 -3288
rect 546 -3300 552 -3294
rect 546 -3306 552 -3300
rect 546 -3312 552 -3306
rect 546 -3318 552 -3312
rect 546 -3324 552 -3318
rect 552 -1296 558 -1290
rect 552 -1302 558 -1296
rect 552 -1308 558 -1302
rect 552 -1314 558 -1308
rect 552 -1320 558 -1314
rect 552 -1326 558 -1320
rect 552 -1332 558 -1326
rect 552 -1338 558 -1332
rect 552 -1344 558 -1338
rect 552 -1350 558 -1344
rect 552 -1356 558 -1350
rect 552 -1362 558 -1356
rect 552 -1368 558 -1362
rect 552 -1374 558 -1368
rect 552 -1380 558 -1374
rect 552 -1386 558 -1380
rect 552 -1392 558 -1386
rect 552 -1398 558 -1392
rect 552 -1404 558 -1398
rect 552 -1410 558 -1404
rect 552 -1416 558 -1410
rect 552 -1422 558 -1416
rect 552 -1428 558 -1422
rect 552 -1434 558 -1428
rect 552 -1440 558 -1434
rect 552 -1446 558 -1440
rect 552 -1452 558 -1446
rect 552 -1458 558 -1452
rect 552 -1464 558 -1458
rect 552 -1470 558 -1464
rect 552 -1476 558 -1470
rect 552 -1482 558 -1476
rect 552 -1488 558 -1482
rect 552 -1494 558 -1488
rect 552 -1500 558 -1494
rect 552 -1506 558 -1500
rect 552 -1512 558 -1506
rect 552 -1518 558 -1512
rect 552 -1524 558 -1518
rect 552 -1530 558 -1524
rect 552 -1536 558 -1530
rect 552 -1542 558 -1536
rect 552 -1548 558 -1542
rect 552 -1554 558 -1548
rect 552 -3072 558 -3066
rect 552 -3078 558 -3072
rect 552 -3084 558 -3078
rect 552 -3090 558 -3084
rect 552 -3096 558 -3090
rect 552 -3102 558 -3096
rect 552 -3108 558 -3102
rect 552 -3114 558 -3108
rect 552 -3120 558 -3114
rect 552 -3126 558 -3120
rect 552 -3132 558 -3126
rect 552 -3138 558 -3132
rect 552 -3144 558 -3138
rect 552 -3150 558 -3144
rect 552 -3156 558 -3150
rect 552 -3162 558 -3156
rect 552 -3168 558 -3162
rect 552 -3174 558 -3168
rect 552 -3180 558 -3174
rect 552 -3186 558 -3180
rect 552 -3192 558 -3186
rect 552 -3198 558 -3192
rect 552 -3204 558 -3198
rect 552 -3210 558 -3204
rect 552 -3216 558 -3210
rect 552 -3222 558 -3216
rect 552 -3228 558 -3222
rect 552 -3234 558 -3228
rect 552 -3240 558 -3234
rect 552 -3246 558 -3240
rect 552 -3252 558 -3246
rect 552 -3258 558 -3252
rect 552 -3264 558 -3258
rect 552 -3270 558 -3264
rect 552 -3276 558 -3270
rect 552 -3282 558 -3276
rect 552 -3288 558 -3282
rect 552 -3294 558 -3288
rect 552 -3300 558 -3294
rect 552 -3306 558 -3300
rect 552 -3312 558 -3306
rect 552 -3318 558 -3312
rect 552 -3324 558 -3318
rect 552 -3330 558 -3324
rect 558 -1296 564 -1290
rect 558 -1302 564 -1296
rect 558 -1308 564 -1302
rect 558 -1314 564 -1308
rect 558 -1320 564 -1314
rect 558 -1326 564 -1320
rect 558 -1332 564 -1326
rect 558 -1338 564 -1332
rect 558 -1344 564 -1338
rect 558 -1350 564 -1344
rect 558 -1356 564 -1350
rect 558 -1362 564 -1356
rect 558 -1368 564 -1362
rect 558 -1374 564 -1368
rect 558 -1380 564 -1374
rect 558 -1386 564 -1380
rect 558 -1392 564 -1386
rect 558 -1398 564 -1392
rect 558 -1404 564 -1398
rect 558 -1410 564 -1404
rect 558 -1416 564 -1410
rect 558 -1422 564 -1416
rect 558 -1428 564 -1422
rect 558 -1434 564 -1428
rect 558 -1440 564 -1434
rect 558 -1446 564 -1440
rect 558 -1452 564 -1446
rect 558 -1458 564 -1452
rect 558 -1464 564 -1458
rect 558 -1470 564 -1464
rect 558 -1476 564 -1470
rect 558 -1482 564 -1476
rect 558 -1488 564 -1482
rect 558 -1494 564 -1488
rect 558 -1500 564 -1494
rect 558 -1506 564 -1500
rect 558 -1512 564 -1506
rect 558 -1518 564 -1512
rect 558 -1524 564 -1518
rect 558 -1530 564 -1524
rect 558 -1536 564 -1530
rect 558 -1542 564 -1536
rect 558 -1548 564 -1542
rect 558 -3078 564 -3072
rect 558 -3084 564 -3078
rect 558 -3090 564 -3084
rect 558 -3096 564 -3090
rect 558 -3102 564 -3096
rect 558 -3108 564 -3102
rect 558 -3114 564 -3108
rect 558 -3120 564 -3114
rect 558 -3126 564 -3120
rect 558 -3132 564 -3126
rect 558 -3138 564 -3132
rect 558 -3144 564 -3138
rect 558 -3150 564 -3144
rect 558 -3156 564 -3150
rect 558 -3162 564 -3156
rect 558 -3168 564 -3162
rect 558 -3174 564 -3168
rect 558 -3180 564 -3174
rect 558 -3186 564 -3180
rect 558 -3192 564 -3186
rect 558 -3198 564 -3192
rect 558 -3204 564 -3198
rect 558 -3210 564 -3204
rect 558 -3216 564 -3210
rect 558 -3222 564 -3216
rect 558 -3228 564 -3222
rect 558 -3234 564 -3228
rect 558 -3240 564 -3234
rect 558 -3246 564 -3240
rect 558 -3252 564 -3246
rect 558 -3258 564 -3252
rect 558 -3264 564 -3258
rect 558 -3270 564 -3264
rect 558 -3276 564 -3270
rect 558 -3282 564 -3276
rect 558 -3288 564 -3282
rect 558 -3294 564 -3288
rect 558 -3300 564 -3294
rect 558 -3306 564 -3300
rect 558 -3312 564 -3306
rect 558 -3318 564 -3312
rect 558 -3324 564 -3318
rect 558 -3330 564 -3324
rect 564 -1290 570 -1284
rect 564 -1296 570 -1290
rect 564 -1302 570 -1296
rect 564 -1308 570 -1302
rect 564 -1314 570 -1308
rect 564 -1320 570 -1314
rect 564 -1326 570 -1320
rect 564 -1332 570 -1326
rect 564 -1338 570 -1332
rect 564 -1344 570 -1338
rect 564 -1350 570 -1344
rect 564 -1356 570 -1350
rect 564 -1362 570 -1356
rect 564 -1368 570 -1362
rect 564 -1374 570 -1368
rect 564 -1380 570 -1374
rect 564 -1386 570 -1380
rect 564 -1392 570 -1386
rect 564 -1398 570 -1392
rect 564 -1404 570 -1398
rect 564 -1410 570 -1404
rect 564 -1416 570 -1410
rect 564 -1422 570 -1416
rect 564 -1428 570 -1422
rect 564 -1434 570 -1428
rect 564 -1440 570 -1434
rect 564 -1446 570 -1440
rect 564 -1452 570 -1446
rect 564 -1458 570 -1452
rect 564 -1464 570 -1458
rect 564 -1470 570 -1464
rect 564 -1476 570 -1470
rect 564 -1482 570 -1476
rect 564 -1488 570 -1482
rect 564 -1494 570 -1488
rect 564 -1500 570 -1494
rect 564 -1506 570 -1500
rect 564 -1512 570 -1506
rect 564 -1518 570 -1512
rect 564 -1524 570 -1518
rect 564 -1530 570 -1524
rect 564 -1536 570 -1530
rect 564 -1542 570 -1536
rect 564 -3084 570 -3078
rect 564 -3090 570 -3084
rect 564 -3096 570 -3090
rect 564 -3102 570 -3096
rect 564 -3108 570 -3102
rect 564 -3114 570 -3108
rect 564 -3120 570 -3114
rect 564 -3126 570 -3120
rect 564 -3132 570 -3126
rect 564 -3138 570 -3132
rect 564 -3144 570 -3138
rect 564 -3150 570 -3144
rect 564 -3156 570 -3150
rect 564 -3162 570 -3156
rect 564 -3168 570 -3162
rect 564 -3174 570 -3168
rect 564 -3180 570 -3174
rect 564 -3186 570 -3180
rect 564 -3192 570 -3186
rect 564 -3198 570 -3192
rect 564 -3204 570 -3198
rect 564 -3210 570 -3204
rect 564 -3216 570 -3210
rect 564 -3222 570 -3216
rect 564 -3228 570 -3222
rect 564 -3234 570 -3228
rect 564 -3240 570 -3234
rect 564 -3246 570 -3240
rect 564 -3252 570 -3246
rect 564 -3258 570 -3252
rect 564 -3264 570 -3258
rect 564 -3270 570 -3264
rect 564 -3276 570 -3270
rect 564 -3282 570 -3276
rect 564 -3288 570 -3282
rect 564 -3294 570 -3288
rect 564 -3300 570 -3294
rect 564 -3306 570 -3300
rect 564 -3312 570 -3306
rect 564 -3318 570 -3312
rect 564 -3324 570 -3318
rect 564 -3330 570 -3324
rect 564 -3336 570 -3330
rect 570 -1290 576 -1284
rect 570 -1296 576 -1290
rect 570 -1302 576 -1296
rect 570 -1308 576 -1302
rect 570 -1314 576 -1308
rect 570 -1320 576 -1314
rect 570 -1326 576 -1320
rect 570 -1332 576 -1326
rect 570 -1338 576 -1332
rect 570 -1344 576 -1338
rect 570 -1350 576 -1344
rect 570 -1356 576 -1350
rect 570 -1362 576 -1356
rect 570 -1368 576 -1362
rect 570 -1374 576 -1368
rect 570 -1380 576 -1374
rect 570 -1386 576 -1380
rect 570 -1392 576 -1386
rect 570 -1398 576 -1392
rect 570 -1404 576 -1398
rect 570 -1410 576 -1404
rect 570 -1416 576 -1410
rect 570 -1422 576 -1416
rect 570 -1428 576 -1422
rect 570 -1434 576 -1428
rect 570 -1440 576 -1434
rect 570 -1446 576 -1440
rect 570 -1452 576 -1446
rect 570 -1458 576 -1452
rect 570 -1464 576 -1458
rect 570 -1470 576 -1464
rect 570 -1476 576 -1470
rect 570 -1482 576 -1476
rect 570 -1488 576 -1482
rect 570 -1494 576 -1488
rect 570 -1500 576 -1494
rect 570 -1506 576 -1500
rect 570 -1512 576 -1506
rect 570 -1518 576 -1512
rect 570 -1524 576 -1518
rect 570 -1530 576 -1524
rect 570 -1536 576 -1530
rect 570 -3090 576 -3084
rect 570 -3096 576 -3090
rect 570 -3102 576 -3096
rect 570 -3108 576 -3102
rect 570 -3114 576 -3108
rect 570 -3120 576 -3114
rect 570 -3126 576 -3120
rect 570 -3132 576 -3126
rect 570 -3138 576 -3132
rect 570 -3144 576 -3138
rect 570 -3150 576 -3144
rect 570 -3156 576 -3150
rect 570 -3162 576 -3156
rect 570 -3168 576 -3162
rect 570 -3174 576 -3168
rect 570 -3180 576 -3174
rect 570 -3186 576 -3180
rect 570 -3192 576 -3186
rect 570 -3198 576 -3192
rect 570 -3204 576 -3198
rect 570 -3210 576 -3204
rect 570 -3216 576 -3210
rect 570 -3222 576 -3216
rect 570 -3228 576 -3222
rect 570 -3234 576 -3228
rect 570 -3240 576 -3234
rect 570 -3246 576 -3240
rect 570 -3252 576 -3246
rect 570 -3258 576 -3252
rect 570 -3264 576 -3258
rect 570 -3270 576 -3264
rect 570 -3276 576 -3270
rect 570 -3282 576 -3276
rect 570 -3288 576 -3282
rect 570 -3294 576 -3288
rect 570 -3300 576 -3294
rect 570 -3306 576 -3300
rect 570 -3312 576 -3306
rect 570 -3318 576 -3312
rect 570 -3324 576 -3318
rect 570 -3330 576 -3324
rect 570 -3336 576 -3330
rect 570 -3342 576 -3336
rect 576 -1284 582 -1278
rect 576 -1290 582 -1284
rect 576 -1296 582 -1290
rect 576 -1302 582 -1296
rect 576 -1308 582 -1302
rect 576 -1314 582 -1308
rect 576 -1320 582 -1314
rect 576 -1326 582 -1320
rect 576 -1332 582 -1326
rect 576 -1338 582 -1332
rect 576 -1344 582 -1338
rect 576 -1350 582 -1344
rect 576 -1356 582 -1350
rect 576 -1362 582 -1356
rect 576 -1368 582 -1362
rect 576 -1374 582 -1368
rect 576 -1380 582 -1374
rect 576 -1386 582 -1380
rect 576 -1392 582 -1386
rect 576 -1398 582 -1392
rect 576 -1404 582 -1398
rect 576 -1410 582 -1404
rect 576 -1416 582 -1410
rect 576 -1422 582 -1416
rect 576 -1428 582 -1422
rect 576 -1434 582 -1428
rect 576 -1440 582 -1434
rect 576 -1446 582 -1440
rect 576 -1452 582 -1446
rect 576 -1458 582 -1452
rect 576 -1464 582 -1458
rect 576 -1470 582 -1464
rect 576 -1476 582 -1470
rect 576 -1482 582 -1476
rect 576 -1488 582 -1482
rect 576 -1494 582 -1488
rect 576 -1500 582 -1494
rect 576 -1506 582 -1500
rect 576 -1512 582 -1506
rect 576 -1518 582 -1512
rect 576 -1524 582 -1518
rect 576 -1530 582 -1524
rect 576 -3096 582 -3090
rect 576 -3102 582 -3096
rect 576 -3108 582 -3102
rect 576 -3114 582 -3108
rect 576 -3120 582 -3114
rect 576 -3126 582 -3120
rect 576 -3132 582 -3126
rect 576 -3138 582 -3132
rect 576 -3144 582 -3138
rect 576 -3150 582 -3144
rect 576 -3156 582 -3150
rect 576 -3162 582 -3156
rect 576 -3168 582 -3162
rect 576 -3174 582 -3168
rect 576 -3180 582 -3174
rect 576 -3186 582 -3180
rect 576 -3192 582 -3186
rect 576 -3198 582 -3192
rect 576 -3204 582 -3198
rect 576 -3210 582 -3204
rect 576 -3216 582 -3210
rect 576 -3222 582 -3216
rect 576 -3228 582 -3222
rect 576 -3234 582 -3228
rect 576 -3240 582 -3234
rect 576 -3246 582 -3240
rect 576 -3252 582 -3246
rect 576 -3258 582 -3252
rect 576 -3264 582 -3258
rect 576 -3270 582 -3264
rect 576 -3276 582 -3270
rect 576 -3282 582 -3276
rect 576 -3288 582 -3282
rect 576 -3294 582 -3288
rect 576 -3300 582 -3294
rect 576 -3306 582 -3300
rect 576 -3312 582 -3306
rect 576 -3318 582 -3312
rect 576 -3324 582 -3318
rect 576 -3330 582 -3324
rect 576 -3336 582 -3330
rect 576 -3342 582 -3336
rect 582 -1278 588 -1272
rect 582 -1284 588 -1278
rect 582 -1290 588 -1284
rect 582 -1296 588 -1290
rect 582 -1302 588 -1296
rect 582 -1308 588 -1302
rect 582 -1314 588 -1308
rect 582 -1320 588 -1314
rect 582 -1326 588 -1320
rect 582 -1332 588 -1326
rect 582 -1338 588 -1332
rect 582 -1344 588 -1338
rect 582 -1350 588 -1344
rect 582 -1356 588 -1350
rect 582 -1362 588 -1356
rect 582 -1368 588 -1362
rect 582 -1374 588 -1368
rect 582 -1380 588 -1374
rect 582 -1386 588 -1380
rect 582 -1392 588 -1386
rect 582 -1398 588 -1392
rect 582 -1404 588 -1398
rect 582 -1410 588 -1404
rect 582 -1416 588 -1410
rect 582 -1422 588 -1416
rect 582 -1428 588 -1422
rect 582 -1434 588 -1428
rect 582 -1440 588 -1434
rect 582 -1446 588 -1440
rect 582 -1452 588 -1446
rect 582 -1458 588 -1452
rect 582 -1464 588 -1458
rect 582 -1470 588 -1464
rect 582 -1476 588 -1470
rect 582 -1482 588 -1476
rect 582 -1488 588 -1482
rect 582 -1494 588 -1488
rect 582 -1500 588 -1494
rect 582 -1506 588 -1500
rect 582 -1512 588 -1506
rect 582 -1518 588 -1512
rect 582 -1524 588 -1518
rect 582 -1530 588 -1524
rect 582 -3102 588 -3096
rect 582 -3108 588 -3102
rect 582 -3114 588 -3108
rect 582 -3120 588 -3114
rect 582 -3126 588 -3120
rect 582 -3132 588 -3126
rect 582 -3138 588 -3132
rect 582 -3144 588 -3138
rect 582 -3150 588 -3144
rect 582 -3156 588 -3150
rect 582 -3162 588 -3156
rect 582 -3168 588 -3162
rect 582 -3174 588 -3168
rect 582 -3180 588 -3174
rect 582 -3186 588 -3180
rect 582 -3192 588 -3186
rect 582 -3198 588 -3192
rect 582 -3204 588 -3198
rect 582 -3210 588 -3204
rect 582 -3216 588 -3210
rect 582 -3222 588 -3216
rect 582 -3228 588 -3222
rect 582 -3234 588 -3228
rect 582 -3240 588 -3234
rect 582 -3246 588 -3240
rect 582 -3252 588 -3246
rect 582 -3258 588 -3252
rect 582 -3264 588 -3258
rect 582 -3270 588 -3264
rect 582 -3276 588 -3270
rect 582 -3282 588 -3276
rect 582 -3288 588 -3282
rect 582 -3294 588 -3288
rect 582 -3300 588 -3294
rect 582 -3306 588 -3300
rect 582 -3312 588 -3306
rect 582 -3318 588 -3312
rect 582 -3324 588 -3318
rect 582 -3330 588 -3324
rect 582 -3336 588 -3330
rect 582 -3342 588 -3336
rect 582 -3348 588 -3342
rect 588 -1278 594 -1272
rect 588 -1284 594 -1278
rect 588 -1290 594 -1284
rect 588 -1296 594 -1290
rect 588 -1302 594 -1296
rect 588 -1308 594 -1302
rect 588 -1314 594 -1308
rect 588 -1320 594 -1314
rect 588 -1326 594 -1320
rect 588 -1332 594 -1326
rect 588 -1338 594 -1332
rect 588 -1344 594 -1338
rect 588 -1350 594 -1344
rect 588 -1356 594 -1350
rect 588 -1362 594 -1356
rect 588 -1368 594 -1362
rect 588 -1374 594 -1368
rect 588 -1380 594 -1374
rect 588 -1386 594 -1380
rect 588 -1392 594 -1386
rect 588 -1398 594 -1392
rect 588 -1404 594 -1398
rect 588 -1410 594 -1404
rect 588 -1416 594 -1410
rect 588 -1422 594 -1416
rect 588 -1428 594 -1422
rect 588 -1434 594 -1428
rect 588 -1440 594 -1434
rect 588 -1446 594 -1440
rect 588 -1452 594 -1446
rect 588 -1458 594 -1452
rect 588 -1464 594 -1458
rect 588 -1470 594 -1464
rect 588 -1476 594 -1470
rect 588 -1482 594 -1476
rect 588 -1488 594 -1482
rect 588 -1494 594 -1488
rect 588 -1500 594 -1494
rect 588 -1506 594 -1500
rect 588 -1512 594 -1506
rect 588 -1518 594 -1512
rect 588 -1524 594 -1518
rect 588 -3102 594 -3096
rect 588 -3108 594 -3102
rect 588 -3114 594 -3108
rect 588 -3120 594 -3114
rect 588 -3126 594 -3120
rect 588 -3132 594 -3126
rect 588 -3138 594 -3132
rect 588 -3144 594 -3138
rect 588 -3150 594 -3144
rect 588 -3156 594 -3150
rect 588 -3162 594 -3156
rect 588 -3168 594 -3162
rect 588 -3174 594 -3168
rect 588 -3180 594 -3174
rect 588 -3186 594 -3180
rect 588 -3192 594 -3186
rect 588 -3198 594 -3192
rect 588 -3204 594 -3198
rect 588 -3210 594 -3204
rect 588 -3216 594 -3210
rect 588 -3222 594 -3216
rect 588 -3228 594 -3222
rect 588 -3234 594 -3228
rect 588 -3240 594 -3234
rect 588 -3246 594 -3240
rect 588 -3252 594 -3246
rect 588 -3258 594 -3252
rect 588 -3264 594 -3258
rect 588 -3270 594 -3264
rect 588 -3276 594 -3270
rect 588 -3282 594 -3276
rect 588 -3288 594 -3282
rect 588 -3294 594 -3288
rect 588 -3300 594 -3294
rect 588 -3306 594 -3300
rect 588 -3312 594 -3306
rect 588 -3318 594 -3312
rect 588 -3324 594 -3318
rect 588 -3330 594 -3324
rect 588 -3336 594 -3330
rect 588 -3342 594 -3336
rect 588 -3348 594 -3342
rect 588 -3354 594 -3348
rect 594 -1272 600 -1266
rect 594 -1278 600 -1272
rect 594 -1284 600 -1278
rect 594 -1290 600 -1284
rect 594 -1296 600 -1290
rect 594 -1302 600 -1296
rect 594 -1308 600 -1302
rect 594 -1314 600 -1308
rect 594 -1320 600 -1314
rect 594 -1326 600 -1320
rect 594 -1332 600 -1326
rect 594 -1338 600 -1332
rect 594 -1344 600 -1338
rect 594 -1350 600 -1344
rect 594 -1356 600 -1350
rect 594 -1362 600 -1356
rect 594 -1368 600 -1362
rect 594 -1374 600 -1368
rect 594 -1380 600 -1374
rect 594 -1386 600 -1380
rect 594 -1392 600 -1386
rect 594 -1398 600 -1392
rect 594 -1404 600 -1398
rect 594 -1410 600 -1404
rect 594 -1416 600 -1410
rect 594 -1422 600 -1416
rect 594 -1428 600 -1422
rect 594 -1434 600 -1428
rect 594 -1440 600 -1434
rect 594 -1446 600 -1440
rect 594 -1452 600 -1446
rect 594 -1458 600 -1452
rect 594 -1464 600 -1458
rect 594 -1470 600 -1464
rect 594 -1476 600 -1470
rect 594 -1482 600 -1476
rect 594 -1488 600 -1482
rect 594 -1494 600 -1488
rect 594 -1500 600 -1494
rect 594 -1506 600 -1500
rect 594 -1512 600 -1506
rect 594 -1518 600 -1512
rect 594 -3108 600 -3102
rect 594 -3114 600 -3108
rect 594 -3120 600 -3114
rect 594 -3126 600 -3120
rect 594 -3132 600 -3126
rect 594 -3138 600 -3132
rect 594 -3144 600 -3138
rect 594 -3150 600 -3144
rect 594 -3156 600 -3150
rect 594 -3162 600 -3156
rect 594 -3168 600 -3162
rect 594 -3174 600 -3168
rect 594 -3180 600 -3174
rect 594 -3186 600 -3180
rect 594 -3192 600 -3186
rect 594 -3198 600 -3192
rect 594 -3204 600 -3198
rect 594 -3210 600 -3204
rect 594 -3216 600 -3210
rect 594 -3222 600 -3216
rect 594 -3228 600 -3222
rect 594 -3234 600 -3228
rect 594 -3240 600 -3234
rect 594 -3246 600 -3240
rect 594 -3252 600 -3246
rect 594 -3258 600 -3252
rect 594 -3264 600 -3258
rect 594 -3270 600 -3264
rect 594 -3276 600 -3270
rect 594 -3282 600 -3276
rect 594 -3288 600 -3282
rect 594 -3294 600 -3288
rect 594 -3300 600 -3294
rect 594 -3306 600 -3300
rect 594 -3312 600 -3306
rect 594 -3318 600 -3312
rect 594 -3324 600 -3318
rect 594 -3330 600 -3324
rect 594 -3336 600 -3330
rect 594 -3342 600 -3336
rect 594 -3348 600 -3342
rect 594 -3354 600 -3348
rect 600 -1266 606 -1260
rect 600 -1272 606 -1266
rect 600 -1278 606 -1272
rect 600 -1284 606 -1278
rect 600 -1290 606 -1284
rect 600 -1296 606 -1290
rect 600 -1302 606 -1296
rect 600 -1308 606 -1302
rect 600 -1314 606 -1308
rect 600 -1320 606 -1314
rect 600 -1326 606 -1320
rect 600 -1332 606 -1326
rect 600 -1338 606 -1332
rect 600 -1344 606 -1338
rect 600 -1350 606 -1344
rect 600 -1356 606 -1350
rect 600 -1362 606 -1356
rect 600 -1368 606 -1362
rect 600 -1374 606 -1368
rect 600 -1380 606 -1374
rect 600 -1386 606 -1380
rect 600 -1392 606 -1386
rect 600 -1398 606 -1392
rect 600 -1404 606 -1398
rect 600 -1410 606 -1404
rect 600 -1416 606 -1410
rect 600 -1422 606 -1416
rect 600 -1428 606 -1422
rect 600 -1434 606 -1428
rect 600 -1440 606 -1434
rect 600 -1446 606 -1440
rect 600 -1452 606 -1446
rect 600 -1458 606 -1452
rect 600 -1464 606 -1458
rect 600 -1470 606 -1464
rect 600 -1476 606 -1470
rect 600 -1482 606 -1476
rect 600 -1488 606 -1482
rect 600 -1494 606 -1488
rect 600 -1500 606 -1494
rect 600 -1506 606 -1500
rect 600 -1512 606 -1506
rect 600 -3114 606 -3108
rect 600 -3120 606 -3114
rect 600 -3126 606 -3120
rect 600 -3132 606 -3126
rect 600 -3138 606 -3132
rect 600 -3144 606 -3138
rect 600 -3150 606 -3144
rect 600 -3156 606 -3150
rect 600 -3162 606 -3156
rect 600 -3168 606 -3162
rect 600 -3174 606 -3168
rect 600 -3180 606 -3174
rect 600 -3186 606 -3180
rect 600 -3192 606 -3186
rect 600 -3198 606 -3192
rect 600 -3204 606 -3198
rect 600 -3210 606 -3204
rect 600 -3216 606 -3210
rect 600 -3222 606 -3216
rect 600 -3228 606 -3222
rect 600 -3234 606 -3228
rect 600 -3240 606 -3234
rect 600 -3246 606 -3240
rect 600 -3252 606 -3246
rect 600 -3258 606 -3252
rect 600 -3264 606 -3258
rect 600 -3270 606 -3264
rect 600 -3276 606 -3270
rect 600 -3282 606 -3276
rect 600 -3288 606 -3282
rect 600 -3294 606 -3288
rect 600 -3300 606 -3294
rect 600 -3306 606 -3300
rect 600 -3312 606 -3306
rect 600 -3318 606 -3312
rect 600 -3324 606 -3318
rect 600 -3330 606 -3324
rect 600 -3336 606 -3330
rect 600 -3342 606 -3336
rect 600 -3348 606 -3342
rect 600 -3354 606 -3348
rect 600 -3360 606 -3354
rect 606 -1266 612 -1260
rect 606 -1272 612 -1266
rect 606 -1278 612 -1272
rect 606 -1284 612 -1278
rect 606 -1290 612 -1284
rect 606 -1296 612 -1290
rect 606 -1302 612 -1296
rect 606 -1308 612 -1302
rect 606 -1314 612 -1308
rect 606 -1320 612 -1314
rect 606 -1326 612 -1320
rect 606 -1332 612 -1326
rect 606 -1338 612 -1332
rect 606 -1344 612 -1338
rect 606 -1350 612 -1344
rect 606 -1356 612 -1350
rect 606 -1362 612 -1356
rect 606 -1368 612 -1362
rect 606 -1374 612 -1368
rect 606 -1380 612 -1374
rect 606 -1386 612 -1380
rect 606 -1392 612 -1386
rect 606 -1398 612 -1392
rect 606 -1404 612 -1398
rect 606 -1410 612 -1404
rect 606 -1416 612 -1410
rect 606 -1422 612 -1416
rect 606 -1428 612 -1422
rect 606 -1434 612 -1428
rect 606 -1440 612 -1434
rect 606 -1446 612 -1440
rect 606 -1452 612 -1446
rect 606 -1458 612 -1452
rect 606 -1464 612 -1458
rect 606 -1470 612 -1464
rect 606 -1476 612 -1470
rect 606 -1482 612 -1476
rect 606 -1488 612 -1482
rect 606 -1494 612 -1488
rect 606 -1500 612 -1494
rect 606 -1506 612 -1500
rect 606 -3120 612 -3114
rect 606 -3126 612 -3120
rect 606 -3132 612 -3126
rect 606 -3138 612 -3132
rect 606 -3144 612 -3138
rect 606 -3150 612 -3144
rect 606 -3156 612 -3150
rect 606 -3162 612 -3156
rect 606 -3168 612 -3162
rect 606 -3174 612 -3168
rect 606 -3180 612 -3174
rect 606 -3186 612 -3180
rect 606 -3192 612 -3186
rect 606 -3198 612 -3192
rect 606 -3204 612 -3198
rect 606 -3210 612 -3204
rect 606 -3216 612 -3210
rect 606 -3222 612 -3216
rect 606 -3228 612 -3222
rect 606 -3234 612 -3228
rect 606 -3240 612 -3234
rect 606 -3246 612 -3240
rect 606 -3252 612 -3246
rect 606 -3258 612 -3252
rect 606 -3264 612 -3258
rect 606 -3270 612 -3264
rect 606 -3276 612 -3270
rect 606 -3282 612 -3276
rect 606 -3288 612 -3282
rect 606 -3294 612 -3288
rect 606 -3300 612 -3294
rect 606 -3306 612 -3300
rect 606 -3312 612 -3306
rect 606 -3318 612 -3312
rect 606 -3324 612 -3318
rect 606 -3330 612 -3324
rect 606 -3336 612 -3330
rect 606 -3342 612 -3336
rect 606 -3348 612 -3342
rect 606 -3354 612 -3348
rect 606 -3360 612 -3354
rect 612 -1260 618 -1254
rect 612 -1266 618 -1260
rect 612 -1272 618 -1266
rect 612 -1278 618 -1272
rect 612 -1284 618 -1278
rect 612 -1290 618 -1284
rect 612 -1296 618 -1290
rect 612 -1302 618 -1296
rect 612 -1308 618 -1302
rect 612 -1314 618 -1308
rect 612 -1320 618 -1314
rect 612 -1326 618 -1320
rect 612 -1332 618 -1326
rect 612 -1338 618 -1332
rect 612 -1344 618 -1338
rect 612 -1350 618 -1344
rect 612 -1356 618 -1350
rect 612 -1362 618 -1356
rect 612 -1368 618 -1362
rect 612 -1374 618 -1368
rect 612 -1380 618 -1374
rect 612 -1386 618 -1380
rect 612 -1392 618 -1386
rect 612 -1398 618 -1392
rect 612 -1404 618 -1398
rect 612 -1410 618 -1404
rect 612 -1416 618 -1410
rect 612 -1422 618 -1416
rect 612 -1428 618 -1422
rect 612 -1434 618 -1428
rect 612 -1440 618 -1434
rect 612 -1446 618 -1440
rect 612 -1452 618 -1446
rect 612 -1458 618 -1452
rect 612 -1464 618 -1458
rect 612 -1470 618 -1464
rect 612 -1476 618 -1470
rect 612 -1482 618 -1476
rect 612 -1488 618 -1482
rect 612 -1494 618 -1488
rect 612 -1500 618 -1494
rect 612 -1506 618 -1500
rect 612 -3126 618 -3120
rect 612 -3132 618 -3126
rect 612 -3138 618 -3132
rect 612 -3144 618 -3138
rect 612 -3150 618 -3144
rect 612 -3156 618 -3150
rect 612 -3162 618 -3156
rect 612 -3168 618 -3162
rect 612 -3174 618 -3168
rect 612 -3180 618 -3174
rect 612 -3186 618 -3180
rect 612 -3192 618 -3186
rect 612 -3198 618 -3192
rect 612 -3204 618 -3198
rect 612 -3210 618 -3204
rect 612 -3216 618 -3210
rect 612 -3222 618 -3216
rect 612 -3228 618 -3222
rect 612 -3234 618 -3228
rect 612 -3240 618 -3234
rect 612 -3246 618 -3240
rect 612 -3252 618 -3246
rect 612 -3258 618 -3252
rect 612 -3264 618 -3258
rect 612 -3270 618 -3264
rect 612 -3276 618 -3270
rect 612 -3282 618 -3276
rect 612 -3288 618 -3282
rect 612 -3294 618 -3288
rect 612 -3300 618 -3294
rect 612 -3306 618 -3300
rect 612 -3312 618 -3306
rect 612 -3318 618 -3312
rect 612 -3324 618 -3318
rect 612 -3330 618 -3324
rect 612 -3336 618 -3330
rect 612 -3342 618 -3336
rect 612 -3348 618 -3342
rect 612 -3354 618 -3348
rect 612 -3360 618 -3354
rect 612 -3366 618 -3360
rect 618 -1260 624 -1254
rect 618 -1266 624 -1260
rect 618 -1272 624 -1266
rect 618 -1278 624 -1272
rect 618 -1284 624 -1278
rect 618 -1290 624 -1284
rect 618 -1296 624 -1290
rect 618 -1302 624 -1296
rect 618 -1308 624 -1302
rect 618 -1314 624 -1308
rect 618 -1320 624 -1314
rect 618 -1326 624 -1320
rect 618 -1332 624 -1326
rect 618 -1338 624 -1332
rect 618 -1344 624 -1338
rect 618 -1350 624 -1344
rect 618 -1356 624 -1350
rect 618 -1362 624 -1356
rect 618 -1368 624 -1362
rect 618 -1374 624 -1368
rect 618 -1380 624 -1374
rect 618 -1386 624 -1380
rect 618 -1392 624 -1386
rect 618 -1398 624 -1392
rect 618 -1404 624 -1398
rect 618 -1410 624 -1404
rect 618 -1416 624 -1410
rect 618 -1422 624 -1416
rect 618 -1428 624 -1422
rect 618 -1434 624 -1428
rect 618 -1440 624 -1434
rect 618 -1446 624 -1440
rect 618 -1452 624 -1446
rect 618 -1458 624 -1452
rect 618 -1464 624 -1458
rect 618 -1470 624 -1464
rect 618 -1476 624 -1470
rect 618 -1482 624 -1476
rect 618 -1488 624 -1482
rect 618 -1494 624 -1488
rect 618 -1500 624 -1494
rect 618 -3126 624 -3120
rect 618 -3132 624 -3126
rect 618 -3138 624 -3132
rect 618 -3144 624 -3138
rect 618 -3150 624 -3144
rect 618 -3156 624 -3150
rect 618 -3162 624 -3156
rect 618 -3168 624 -3162
rect 618 -3174 624 -3168
rect 618 -3180 624 -3174
rect 618 -3186 624 -3180
rect 618 -3192 624 -3186
rect 618 -3198 624 -3192
rect 618 -3204 624 -3198
rect 618 -3210 624 -3204
rect 618 -3216 624 -3210
rect 618 -3222 624 -3216
rect 618 -3228 624 -3222
rect 618 -3234 624 -3228
rect 618 -3240 624 -3234
rect 618 -3246 624 -3240
rect 618 -3252 624 -3246
rect 618 -3258 624 -3252
rect 618 -3264 624 -3258
rect 618 -3270 624 -3264
rect 618 -3276 624 -3270
rect 618 -3282 624 -3276
rect 618 -3288 624 -3282
rect 618 -3294 624 -3288
rect 618 -3300 624 -3294
rect 618 -3306 624 -3300
rect 618 -3312 624 -3306
rect 618 -3318 624 -3312
rect 618 -3324 624 -3318
rect 618 -3330 624 -3324
rect 618 -3336 624 -3330
rect 618 -3342 624 -3336
rect 618 -3348 624 -3342
rect 618 -3354 624 -3348
rect 618 -3360 624 -3354
rect 618 -3366 624 -3360
rect 618 -3372 624 -3366
rect 624 -1254 630 -1248
rect 624 -1260 630 -1254
rect 624 -1266 630 -1260
rect 624 -1272 630 -1266
rect 624 -1278 630 -1272
rect 624 -1284 630 -1278
rect 624 -1290 630 -1284
rect 624 -1296 630 -1290
rect 624 -1302 630 -1296
rect 624 -1308 630 -1302
rect 624 -1314 630 -1308
rect 624 -1320 630 -1314
rect 624 -1326 630 -1320
rect 624 -1332 630 -1326
rect 624 -1338 630 -1332
rect 624 -1344 630 -1338
rect 624 -1350 630 -1344
rect 624 -1356 630 -1350
rect 624 -1362 630 -1356
rect 624 -1368 630 -1362
rect 624 -1374 630 -1368
rect 624 -1380 630 -1374
rect 624 -1386 630 -1380
rect 624 -1392 630 -1386
rect 624 -1398 630 -1392
rect 624 -1404 630 -1398
rect 624 -1410 630 -1404
rect 624 -1416 630 -1410
rect 624 -1422 630 -1416
rect 624 -1428 630 -1422
rect 624 -1434 630 -1428
rect 624 -1440 630 -1434
rect 624 -1446 630 -1440
rect 624 -1452 630 -1446
rect 624 -1458 630 -1452
rect 624 -1464 630 -1458
rect 624 -1470 630 -1464
rect 624 -1476 630 -1470
rect 624 -1482 630 -1476
rect 624 -1488 630 -1482
rect 624 -1494 630 -1488
rect 624 -3132 630 -3126
rect 624 -3138 630 -3132
rect 624 -3144 630 -3138
rect 624 -3150 630 -3144
rect 624 -3156 630 -3150
rect 624 -3162 630 -3156
rect 624 -3168 630 -3162
rect 624 -3174 630 -3168
rect 624 -3180 630 -3174
rect 624 -3186 630 -3180
rect 624 -3192 630 -3186
rect 624 -3198 630 -3192
rect 624 -3204 630 -3198
rect 624 -3210 630 -3204
rect 624 -3216 630 -3210
rect 624 -3222 630 -3216
rect 624 -3228 630 -3222
rect 624 -3234 630 -3228
rect 624 -3240 630 -3234
rect 624 -3246 630 -3240
rect 624 -3252 630 -3246
rect 624 -3258 630 -3252
rect 624 -3264 630 -3258
rect 624 -3270 630 -3264
rect 624 -3276 630 -3270
rect 624 -3282 630 -3276
rect 624 -3288 630 -3282
rect 624 -3294 630 -3288
rect 624 -3300 630 -3294
rect 624 -3306 630 -3300
rect 624 -3312 630 -3306
rect 624 -3318 630 -3312
rect 624 -3324 630 -3318
rect 624 -3330 630 -3324
rect 624 -3336 630 -3330
rect 624 -3342 630 -3336
rect 624 -3348 630 -3342
rect 624 -3354 630 -3348
rect 624 -3360 630 -3354
rect 624 -3366 630 -3360
rect 624 -3372 630 -3366
rect 630 -1254 636 -1248
rect 630 -1260 636 -1254
rect 630 -1266 636 -1260
rect 630 -1272 636 -1266
rect 630 -1278 636 -1272
rect 630 -1284 636 -1278
rect 630 -1290 636 -1284
rect 630 -1296 636 -1290
rect 630 -1302 636 -1296
rect 630 -1308 636 -1302
rect 630 -1314 636 -1308
rect 630 -1320 636 -1314
rect 630 -1326 636 -1320
rect 630 -1332 636 -1326
rect 630 -1338 636 -1332
rect 630 -1344 636 -1338
rect 630 -1350 636 -1344
rect 630 -1356 636 -1350
rect 630 -1362 636 -1356
rect 630 -1368 636 -1362
rect 630 -1374 636 -1368
rect 630 -1380 636 -1374
rect 630 -1386 636 -1380
rect 630 -1392 636 -1386
rect 630 -1398 636 -1392
rect 630 -1404 636 -1398
rect 630 -1410 636 -1404
rect 630 -1416 636 -1410
rect 630 -1422 636 -1416
rect 630 -1428 636 -1422
rect 630 -1434 636 -1428
rect 630 -1440 636 -1434
rect 630 -1446 636 -1440
rect 630 -1452 636 -1446
rect 630 -1458 636 -1452
rect 630 -1464 636 -1458
rect 630 -1470 636 -1464
rect 630 -1476 636 -1470
rect 630 -1482 636 -1476
rect 630 -1488 636 -1482
rect 630 -1494 636 -1488
rect 630 -3138 636 -3132
rect 630 -3144 636 -3138
rect 630 -3150 636 -3144
rect 630 -3156 636 -3150
rect 630 -3162 636 -3156
rect 630 -3168 636 -3162
rect 630 -3174 636 -3168
rect 630 -3180 636 -3174
rect 630 -3186 636 -3180
rect 630 -3192 636 -3186
rect 630 -3198 636 -3192
rect 630 -3204 636 -3198
rect 630 -3210 636 -3204
rect 630 -3216 636 -3210
rect 630 -3222 636 -3216
rect 630 -3228 636 -3222
rect 630 -3234 636 -3228
rect 630 -3240 636 -3234
rect 630 -3246 636 -3240
rect 630 -3252 636 -3246
rect 630 -3258 636 -3252
rect 630 -3264 636 -3258
rect 630 -3270 636 -3264
rect 630 -3276 636 -3270
rect 630 -3282 636 -3276
rect 630 -3288 636 -3282
rect 630 -3294 636 -3288
rect 630 -3300 636 -3294
rect 630 -3306 636 -3300
rect 630 -3312 636 -3306
rect 630 -3318 636 -3312
rect 630 -3324 636 -3318
rect 630 -3330 636 -3324
rect 630 -3336 636 -3330
rect 630 -3342 636 -3336
rect 630 -3348 636 -3342
rect 630 -3354 636 -3348
rect 630 -3360 636 -3354
rect 630 -3366 636 -3360
rect 630 -3372 636 -3366
rect 630 -3378 636 -3372
rect 636 -1248 642 -1242
rect 636 -1254 642 -1248
rect 636 -1260 642 -1254
rect 636 -1266 642 -1260
rect 636 -1272 642 -1266
rect 636 -1278 642 -1272
rect 636 -1284 642 -1278
rect 636 -1290 642 -1284
rect 636 -1296 642 -1290
rect 636 -1302 642 -1296
rect 636 -1308 642 -1302
rect 636 -1314 642 -1308
rect 636 -1320 642 -1314
rect 636 -1326 642 -1320
rect 636 -1332 642 -1326
rect 636 -1338 642 -1332
rect 636 -1344 642 -1338
rect 636 -1350 642 -1344
rect 636 -1356 642 -1350
rect 636 -1362 642 -1356
rect 636 -1368 642 -1362
rect 636 -1374 642 -1368
rect 636 -1380 642 -1374
rect 636 -1386 642 -1380
rect 636 -1392 642 -1386
rect 636 -1398 642 -1392
rect 636 -1404 642 -1398
rect 636 -1410 642 -1404
rect 636 -1416 642 -1410
rect 636 -1422 642 -1416
rect 636 -1428 642 -1422
rect 636 -1434 642 -1428
rect 636 -1440 642 -1434
rect 636 -1446 642 -1440
rect 636 -1452 642 -1446
rect 636 -1458 642 -1452
rect 636 -1464 642 -1458
rect 636 -1470 642 -1464
rect 636 -1476 642 -1470
rect 636 -1482 642 -1476
rect 636 -1488 642 -1482
rect 636 -3144 642 -3138
rect 636 -3150 642 -3144
rect 636 -3156 642 -3150
rect 636 -3162 642 -3156
rect 636 -3168 642 -3162
rect 636 -3174 642 -3168
rect 636 -3180 642 -3174
rect 636 -3186 642 -3180
rect 636 -3192 642 -3186
rect 636 -3198 642 -3192
rect 636 -3204 642 -3198
rect 636 -3210 642 -3204
rect 636 -3216 642 -3210
rect 636 -3222 642 -3216
rect 636 -3228 642 -3222
rect 636 -3234 642 -3228
rect 636 -3240 642 -3234
rect 636 -3246 642 -3240
rect 636 -3252 642 -3246
rect 636 -3258 642 -3252
rect 636 -3264 642 -3258
rect 636 -3270 642 -3264
rect 636 -3276 642 -3270
rect 636 -3282 642 -3276
rect 636 -3288 642 -3282
rect 636 -3294 642 -3288
rect 636 -3300 642 -3294
rect 636 -3306 642 -3300
rect 636 -3312 642 -3306
rect 636 -3318 642 -3312
rect 636 -3324 642 -3318
rect 636 -3330 642 -3324
rect 636 -3336 642 -3330
rect 636 -3342 642 -3336
rect 636 -3348 642 -3342
rect 636 -3354 642 -3348
rect 636 -3360 642 -3354
rect 636 -3366 642 -3360
rect 636 -3372 642 -3366
rect 636 -3378 642 -3372
rect 642 -1248 648 -1242
rect 642 -1254 648 -1248
rect 642 -1260 648 -1254
rect 642 -1266 648 -1260
rect 642 -1272 648 -1266
rect 642 -1278 648 -1272
rect 642 -1284 648 -1278
rect 642 -1290 648 -1284
rect 642 -1296 648 -1290
rect 642 -1302 648 -1296
rect 642 -1308 648 -1302
rect 642 -1314 648 -1308
rect 642 -1320 648 -1314
rect 642 -1326 648 -1320
rect 642 -1332 648 -1326
rect 642 -1338 648 -1332
rect 642 -1344 648 -1338
rect 642 -1350 648 -1344
rect 642 -1356 648 -1350
rect 642 -1362 648 -1356
rect 642 -1368 648 -1362
rect 642 -1374 648 -1368
rect 642 -1380 648 -1374
rect 642 -1386 648 -1380
rect 642 -1392 648 -1386
rect 642 -1398 648 -1392
rect 642 -1404 648 -1398
rect 642 -1410 648 -1404
rect 642 -1416 648 -1410
rect 642 -1422 648 -1416
rect 642 -1428 648 -1422
rect 642 -1434 648 -1428
rect 642 -1440 648 -1434
rect 642 -1446 648 -1440
rect 642 -1452 648 -1446
rect 642 -1458 648 -1452
rect 642 -1464 648 -1458
rect 642 -1470 648 -1464
rect 642 -1476 648 -1470
rect 642 -1482 648 -1476
rect 642 -3144 648 -3138
rect 642 -3150 648 -3144
rect 642 -3156 648 -3150
rect 642 -3162 648 -3156
rect 642 -3168 648 -3162
rect 642 -3174 648 -3168
rect 642 -3180 648 -3174
rect 642 -3186 648 -3180
rect 642 -3192 648 -3186
rect 642 -3198 648 -3192
rect 642 -3204 648 -3198
rect 642 -3210 648 -3204
rect 642 -3216 648 -3210
rect 642 -3222 648 -3216
rect 642 -3228 648 -3222
rect 642 -3234 648 -3228
rect 642 -3240 648 -3234
rect 642 -3246 648 -3240
rect 642 -3252 648 -3246
rect 642 -3258 648 -3252
rect 642 -3264 648 -3258
rect 642 -3270 648 -3264
rect 642 -3276 648 -3270
rect 642 -3282 648 -3276
rect 642 -3288 648 -3282
rect 642 -3294 648 -3288
rect 642 -3300 648 -3294
rect 642 -3306 648 -3300
rect 642 -3312 648 -3306
rect 642 -3318 648 -3312
rect 642 -3324 648 -3318
rect 642 -3330 648 -3324
rect 642 -3336 648 -3330
rect 642 -3342 648 -3336
rect 642 -3348 648 -3342
rect 642 -3354 648 -3348
rect 642 -3360 648 -3354
rect 642 -3366 648 -3360
rect 642 -3372 648 -3366
rect 642 -3378 648 -3372
rect 642 -3384 648 -3378
rect 648 -1242 654 -1236
rect 648 -1248 654 -1242
rect 648 -1254 654 -1248
rect 648 -1260 654 -1254
rect 648 -1266 654 -1260
rect 648 -1272 654 -1266
rect 648 -1278 654 -1272
rect 648 -1284 654 -1278
rect 648 -1290 654 -1284
rect 648 -1296 654 -1290
rect 648 -1302 654 -1296
rect 648 -1308 654 -1302
rect 648 -1314 654 -1308
rect 648 -1320 654 -1314
rect 648 -1326 654 -1320
rect 648 -1332 654 -1326
rect 648 -1338 654 -1332
rect 648 -1344 654 -1338
rect 648 -1350 654 -1344
rect 648 -1356 654 -1350
rect 648 -1362 654 -1356
rect 648 -1368 654 -1362
rect 648 -1374 654 -1368
rect 648 -1380 654 -1374
rect 648 -1386 654 -1380
rect 648 -1392 654 -1386
rect 648 -1398 654 -1392
rect 648 -1404 654 -1398
rect 648 -1410 654 -1404
rect 648 -1416 654 -1410
rect 648 -1422 654 -1416
rect 648 -1428 654 -1422
rect 648 -1434 654 -1428
rect 648 -1440 654 -1434
rect 648 -1446 654 -1440
rect 648 -1452 654 -1446
rect 648 -1458 654 -1452
rect 648 -1464 654 -1458
rect 648 -1470 654 -1464
rect 648 -1476 654 -1470
rect 648 -3150 654 -3144
rect 648 -3156 654 -3150
rect 648 -3162 654 -3156
rect 648 -3168 654 -3162
rect 648 -3174 654 -3168
rect 648 -3180 654 -3174
rect 648 -3186 654 -3180
rect 648 -3192 654 -3186
rect 648 -3198 654 -3192
rect 648 -3204 654 -3198
rect 648 -3210 654 -3204
rect 648 -3216 654 -3210
rect 648 -3222 654 -3216
rect 648 -3228 654 -3222
rect 648 -3234 654 -3228
rect 648 -3240 654 -3234
rect 648 -3246 654 -3240
rect 648 -3252 654 -3246
rect 648 -3258 654 -3252
rect 648 -3264 654 -3258
rect 648 -3270 654 -3264
rect 648 -3276 654 -3270
rect 648 -3282 654 -3276
rect 648 -3288 654 -3282
rect 648 -3294 654 -3288
rect 648 -3300 654 -3294
rect 648 -3306 654 -3300
rect 648 -3312 654 -3306
rect 648 -3318 654 -3312
rect 648 -3324 654 -3318
rect 648 -3330 654 -3324
rect 648 -3336 654 -3330
rect 648 -3342 654 -3336
rect 648 -3348 654 -3342
rect 648 -3354 654 -3348
rect 648 -3360 654 -3354
rect 648 -3366 654 -3360
rect 648 -3372 654 -3366
rect 648 -3378 654 -3372
rect 648 -3384 654 -3378
rect 654 -1242 660 -1236
rect 654 -1248 660 -1242
rect 654 -1254 660 -1248
rect 654 -1260 660 -1254
rect 654 -1266 660 -1260
rect 654 -1272 660 -1266
rect 654 -1278 660 -1272
rect 654 -1284 660 -1278
rect 654 -1290 660 -1284
rect 654 -1296 660 -1290
rect 654 -1302 660 -1296
rect 654 -1308 660 -1302
rect 654 -1314 660 -1308
rect 654 -1320 660 -1314
rect 654 -1326 660 -1320
rect 654 -1332 660 -1326
rect 654 -1338 660 -1332
rect 654 -1344 660 -1338
rect 654 -1350 660 -1344
rect 654 -1356 660 -1350
rect 654 -1362 660 -1356
rect 654 -1368 660 -1362
rect 654 -1374 660 -1368
rect 654 -1380 660 -1374
rect 654 -1386 660 -1380
rect 654 -1392 660 -1386
rect 654 -1398 660 -1392
rect 654 -1404 660 -1398
rect 654 -1410 660 -1404
rect 654 -1416 660 -1410
rect 654 -1422 660 -1416
rect 654 -1428 660 -1422
rect 654 -1434 660 -1428
rect 654 -1440 660 -1434
rect 654 -1446 660 -1440
rect 654 -1452 660 -1446
rect 654 -1458 660 -1452
rect 654 -1464 660 -1458
rect 654 -1470 660 -1464
rect 654 -1476 660 -1470
rect 654 -3156 660 -3150
rect 654 -3162 660 -3156
rect 654 -3168 660 -3162
rect 654 -3174 660 -3168
rect 654 -3180 660 -3174
rect 654 -3186 660 -3180
rect 654 -3192 660 -3186
rect 654 -3198 660 -3192
rect 654 -3204 660 -3198
rect 654 -3210 660 -3204
rect 654 -3216 660 -3210
rect 654 -3222 660 -3216
rect 654 -3228 660 -3222
rect 654 -3234 660 -3228
rect 654 -3240 660 -3234
rect 654 -3246 660 -3240
rect 654 -3252 660 -3246
rect 654 -3258 660 -3252
rect 654 -3264 660 -3258
rect 654 -3270 660 -3264
rect 654 -3276 660 -3270
rect 654 -3282 660 -3276
rect 654 -3288 660 -3282
rect 654 -3294 660 -3288
rect 654 -3300 660 -3294
rect 654 -3306 660 -3300
rect 654 -3312 660 -3306
rect 654 -3318 660 -3312
rect 654 -3324 660 -3318
rect 654 -3330 660 -3324
rect 654 -3336 660 -3330
rect 654 -3342 660 -3336
rect 654 -3348 660 -3342
rect 654 -3354 660 -3348
rect 654 -3360 660 -3354
rect 654 -3366 660 -3360
rect 654 -3372 660 -3366
rect 654 -3378 660 -3372
rect 654 -3384 660 -3378
rect 654 -3390 660 -3384
rect 660 -1236 666 -1230
rect 660 -1242 666 -1236
rect 660 -1248 666 -1242
rect 660 -1254 666 -1248
rect 660 -1260 666 -1254
rect 660 -1266 666 -1260
rect 660 -1272 666 -1266
rect 660 -1278 666 -1272
rect 660 -1284 666 -1278
rect 660 -1290 666 -1284
rect 660 -1296 666 -1290
rect 660 -1302 666 -1296
rect 660 -1308 666 -1302
rect 660 -1314 666 -1308
rect 660 -1320 666 -1314
rect 660 -1326 666 -1320
rect 660 -1332 666 -1326
rect 660 -1338 666 -1332
rect 660 -1344 666 -1338
rect 660 -1350 666 -1344
rect 660 -1356 666 -1350
rect 660 -1362 666 -1356
rect 660 -1368 666 -1362
rect 660 -1374 666 -1368
rect 660 -1380 666 -1374
rect 660 -1386 666 -1380
rect 660 -1392 666 -1386
rect 660 -1398 666 -1392
rect 660 -1404 666 -1398
rect 660 -1410 666 -1404
rect 660 -1416 666 -1410
rect 660 -1422 666 -1416
rect 660 -1428 666 -1422
rect 660 -1434 666 -1428
rect 660 -1440 666 -1434
rect 660 -1446 666 -1440
rect 660 -1452 666 -1446
rect 660 -1458 666 -1452
rect 660 -1464 666 -1458
rect 660 -1470 666 -1464
rect 660 -3156 666 -3150
rect 660 -3162 666 -3156
rect 660 -3168 666 -3162
rect 660 -3174 666 -3168
rect 660 -3180 666 -3174
rect 660 -3186 666 -3180
rect 660 -3192 666 -3186
rect 660 -3198 666 -3192
rect 660 -3204 666 -3198
rect 660 -3210 666 -3204
rect 660 -3216 666 -3210
rect 660 -3222 666 -3216
rect 660 -3228 666 -3222
rect 660 -3234 666 -3228
rect 660 -3240 666 -3234
rect 660 -3246 666 -3240
rect 660 -3252 666 -3246
rect 660 -3258 666 -3252
rect 660 -3264 666 -3258
rect 660 -3270 666 -3264
rect 660 -3276 666 -3270
rect 660 -3282 666 -3276
rect 660 -3288 666 -3282
rect 660 -3294 666 -3288
rect 660 -3300 666 -3294
rect 660 -3306 666 -3300
rect 660 -3312 666 -3306
rect 660 -3318 666 -3312
rect 660 -3324 666 -3318
rect 660 -3330 666 -3324
rect 660 -3336 666 -3330
rect 660 -3342 666 -3336
rect 660 -3348 666 -3342
rect 660 -3354 666 -3348
rect 660 -3360 666 -3354
rect 660 -3366 666 -3360
rect 660 -3372 666 -3366
rect 660 -3378 666 -3372
rect 660 -3384 666 -3378
rect 660 -3390 666 -3384
rect 666 -1236 672 -1230
rect 666 -1242 672 -1236
rect 666 -1248 672 -1242
rect 666 -1254 672 -1248
rect 666 -1260 672 -1254
rect 666 -1266 672 -1260
rect 666 -1272 672 -1266
rect 666 -1278 672 -1272
rect 666 -1284 672 -1278
rect 666 -1290 672 -1284
rect 666 -1296 672 -1290
rect 666 -1302 672 -1296
rect 666 -1308 672 -1302
rect 666 -1314 672 -1308
rect 666 -1320 672 -1314
rect 666 -1326 672 -1320
rect 666 -1332 672 -1326
rect 666 -1338 672 -1332
rect 666 -1344 672 -1338
rect 666 -1350 672 -1344
rect 666 -1356 672 -1350
rect 666 -1362 672 -1356
rect 666 -1368 672 -1362
rect 666 -1374 672 -1368
rect 666 -1380 672 -1374
rect 666 -1386 672 -1380
rect 666 -1392 672 -1386
rect 666 -1398 672 -1392
rect 666 -1404 672 -1398
rect 666 -1410 672 -1404
rect 666 -1416 672 -1410
rect 666 -1422 672 -1416
rect 666 -1428 672 -1422
rect 666 -1434 672 -1428
rect 666 -1440 672 -1434
rect 666 -1446 672 -1440
rect 666 -1452 672 -1446
rect 666 -1458 672 -1452
rect 666 -1464 672 -1458
rect 666 -1470 672 -1464
rect 666 -3162 672 -3156
rect 666 -3168 672 -3162
rect 666 -3174 672 -3168
rect 666 -3180 672 -3174
rect 666 -3186 672 -3180
rect 666 -3192 672 -3186
rect 666 -3198 672 -3192
rect 666 -3204 672 -3198
rect 666 -3210 672 -3204
rect 666 -3216 672 -3210
rect 666 -3222 672 -3216
rect 666 -3228 672 -3222
rect 666 -3234 672 -3228
rect 666 -3240 672 -3234
rect 666 -3246 672 -3240
rect 666 -3252 672 -3246
rect 666 -3258 672 -3252
rect 666 -3264 672 -3258
rect 666 -3270 672 -3264
rect 666 -3276 672 -3270
rect 666 -3282 672 -3276
rect 666 -3288 672 -3282
rect 666 -3294 672 -3288
rect 666 -3300 672 -3294
rect 666 -3306 672 -3300
rect 666 -3312 672 -3306
rect 666 -3318 672 -3312
rect 666 -3324 672 -3318
rect 666 -3330 672 -3324
rect 666 -3336 672 -3330
rect 666 -3342 672 -3336
rect 666 -3348 672 -3342
rect 666 -3354 672 -3348
rect 666 -3360 672 -3354
rect 666 -3366 672 -3360
rect 666 -3372 672 -3366
rect 666 -3378 672 -3372
rect 666 -3384 672 -3378
rect 666 -3390 672 -3384
rect 666 -3396 672 -3390
rect 672 -1230 678 -1224
rect 672 -1236 678 -1230
rect 672 -1242 678 -1236
rect 672 -1248 678 -1242
rect 672 -1254 678 -1248
rect 672 -1260 678 -1254
rect 672 -1266 678 -1260
rect 672 -1272 678 -1266
rect 672 -1278 678 -1272
rect 672 -1284 678 -1278
rect 672 -1290 678 -1284
rect 672 -1296 678 -1290
rect 672 -1302 678 -1296
rect 672 -1308 678 -1302
rect 672 -1314 678 -1308
rect 672 -1320 678 -1314
rect 672 -1326 678 -1320
rect 672 -1332 678 -1326
rect 672 -1338 678 -1332
rect 672 -1344 678 -1338
rect 672 -1350 678 -1344
rect 672 -1356 678 -1350
rect 672 -1362 678 -1356
rect 672 -1368 678 -1362
rect 672 -1374 678 -1368
rect 672 -1380 678 -1374
rect 672 -1386 678 -1380
rect 672 -1392 678 -1386
rect 672 -1398 678 -1392
rect 672 -1404 678 -1398
rect 672 -1410 678 -1404
rect 672 -1416 678 -1410
rect 672 -1422 678 -1416
rect 672 -1428 678 -1422
rect 672 -1434 678 -1428
rect 672 -1440 678 -1434
rect 672 -1446 678 -1440
rect 672 -1452 678 -1446
rect 672 -1458 678 -1452
rect 672 -1464 678 -1458
rect 672 -3168 678 -3162
rect 672 -3174 678 -3168
rect 672 -3180 678 -3174
rect 672 -3186 678 -3180
rect 672 -3192 678 -3186
rect 672 -3198 678 -3192
rect 672 -3204 678 -3198
rect 672 -3210 678 -3204
rect 672 -3216 678 -3210
rect 672 -3222 678 -3216
rect 672 -3228 678 -3222
rect 672 -3234 678 -3228
rect 672 -3240 678 -3234
rect 672 -3246 678 -3240
rect 672 -3252 678 -3246
rect 672 -3258 678 -3252
rect 672 -3264 678 -3258
rect 672 -3270 678 -3264
rect 672 -3276 678 -3270
rect 672 -3282 678 -3276
rect 672 -3288 678 -3282
rect 672 -3294 678 -3288
rect 672 -3300 678 -3294
rect 672 -3306 678 -3300
rect 672 -3312 678 -3306
rect 672 -3318 678 -3312
rect 672 -3324 678 -3318
rect 672 -3330 678 -3324
rect 672 -3336 678 -3330
rect 672 -3342 678 -3336
rect 672 -3348 678 -3342
rect 672 -3354 678 -3348
rect 672 -3360 678 -3354
rect 672 -3366 678 -3360
rect 672 -3372 678 -3366
rect 672 -3378 678 -3372
rect 672 -3384 678 -3378
rect 672 -3390 678 -3384
rect 672 -3396 678 -3390
rect 672 -3402 678 -3396
rect 678 -1230 684 -1224
rect 678 -1236 684 -1230
rect 678 -1242 684 -1236
rect 678 -1248 684 -1242
rect 678 -1254 684 -1248
rect 678 -1260 684 -1254
rect 678 -1266 684 -1260
rect 678 -1272 684 -1266
rect 678 -1278 684 -1272
rect 678 -1284 684 -1278
rect 678 -1290 684 -1284
rect 678 -1296 684 -1290
rect 678 -1302 684 -1296
rect 678 -1308 684 -1302
rect 678 -1314 684 -1308
rect 678 -1320 684 -1314
rect 678 -1326 684 -1320
rect 678 -1332 684 -1326
rect 678 -1338 684 -1332
rect 678 -1344 684 -1338
rect 678 -1350 684 -1344
rect 678 -1356 684 -1350
rect 678 -1362 684 -1356
rect 678 -1368 684 -1362
rect 678 -1374 684 -1368
rect 678 -1380 684 -1374
rect 678 -1386 684 -1380
rect 678 -1392 684 -1386
rect 678 -1398 684 -1392
rect 678 -1404 684 -1398
rect 678 -1410 684 -1404
rect 678 -1416 684 -1410
rect 678 -1422 684 -1416
rect 678 -1428 684 -1422
rect 678 -1434 684 -1428
rect 678 -1440 684 -1434
rect 678 -1446 684 -1440
rect 678 -1452 684 -1446
rect 678 -1458 684 -1452
rect 678 -3168 684 -3162
rect 678 -3174 684 -3168
rect 678 -3180 684 -3174
rect 678 -3186 684 -3180
rect 678 -3192 684 -3186
rect 678 -3198 684 -3192
rect 678 -3204 684 -3198
rect 678 -3210 684 -3204
rect 678 -3216 684 -3210
rect 678 -3222 684 -3216
rect 678 -3228 684 -3222
rect 678 -3234 684 -3228
rect 678 -3240 684 -3234
rect 678 -3246 684 -3240
rect 678 -3252 684 -3246
rect 678 -3258 684 -3252
rect 678 -3264 684 -3258
rect 678 -3270 684 -3264
rect 678 -3276 684 -3270
rect 678 -3282 684 -3276
rect 678 -3288 684 -3282
rect 678 -3294 684 -3288
rect 678 -3300 684 -3294
rect 678 -3306 684 -3300
rect 678 -3312 684 -3306
rect 678 -3318 684 -3312
rect 678 -3324 684 -3318
rect 678 -3330 684 -3324
rect 678 -3336 684 -3330
rect 678 -3342 684 -3336
rect 678 -3348 684 -3342
rect 678 -3354 684 -3348
rect 678 -3360 684 -3354
rect 678 -3366 684 -3360
rect 678 -3372 684 -3366
rect 678 -3378 684 -3372
rect 678 -3384 684 -3378
rect 678 -3390 684 -3384
rect 678 -3396 684 -3390
rect 678 -3402 684 -3396
rect 684 -1224 690 -1218
rect 684 -1230 690 -1224
rect 684 -1236 690 -1230
rect 684 -1242 690 -1236
rect 684 -1248 690 -1242
rect 684 -1254 690 -1248
rect 684 -1260 690 -1254
rect 684 -1266 690 -1260
rect 684 -1272 690 -1266
rect 684 -1278 690 -1272
rect 684 -1284 690 -1278
rect 684 -1290 690 -1284
rect 684 -1296 690 -1290
rect 684 -1302 690 -1296
rect 684 -1308 690 -1302
rect 684 -1314 690 -1308
rect 684 -1320 690 -1314
rect 684 -1326 690 -1320
rect 684 -1332 690 -1326
rect 684 -1338 690 -1332
rect 684 -1344 690 -1338
rect 684 -1350 690 -1344
rect 684 -1356 690 -1350
rect 684 -1362 690 -1356
rect 684 -1368 690 -1362
rect 684 -1374 690 -1368
rect 684 -1380 690 -1374
rect 684 -1386 690 -1380
rect 684 -1392 690 -1386
rect 684 -1398 690 -1392
rect 684 -1404 690 -1398
rect 684 -1410 690 -1404
rect 684 -1416 690 -1410
rect 684 -1422 690 -1416
rect 684 -1428 690 -1422
rect 684 -1434 690 -1428
rect 684 -1440 690 -1434
rect 684 -1446 690 -1440
rect 684 -1452 690 -1446
rect 684 -1458 690 -1452
rect 684 -3174 690 -3168
rect 684 -3180 690 -3174
rect 684 -3186 690 -3180
rect 684 -3192 690 -3186
rect 684 -3198 690 -3192
rect 684 -3204 690 -3198
rect 684 -3210 690 -3204
rect 684 -3216 690 -3210
rect 684 -3222 690 -3216
rect 684 -3228 690 -3222
rect 684 -3234 690 -3228
rect 684 -3240 690 -3234
rect 684 -3246 690 -3240
rect 684 -3252 690 -3246
rect 684 -3258 690 -3252
rect 684 -3264 690 -3258
rect 684 -3270 690 -3264
rect 684 -3276 690 -3270
rect 684 -3282 690 -3276
rect 684 -3288 690 -3282
rect 684 -3294 690 -3288
rect 684 -3300 690 -3294
rect 684 -3306 690 -3300
rect 684 -3312 690 -3306
rect 684 -3318 690 -3312
rect 684 -3324 690 -3318
rect 684 -3330 690 -3324
rect 684 -3336 690 -3330
rect 684 -3342 690 -3336
rect 684 -3348 690 -3342
rect 684 -3354 690 -3348
rect 684 -3360 690 -3354
rect 684 -3366 690 -3360
rect 684 -3372 690 -3366
rect 684 -3378 690 -3372
rect 684 -3384 690 -3378
rect 684 -3390 690 -3384
rect 684 -3396 690 -3390
rect 684 -3402 690 -3396
rect 684 -3408 690 -3402
rect 690 -1224 696 -1218
rect 690 -1230 696 -1224
rect 690 -1236 696 -1230
rect 690 -1242 696 -1236
rect 690 -1248 696 -1242
rect 690 -1254 696 -1248
rect 690 -1260 696 -1254
rect 690 -1266 696 -1260
rect 690 -1272 696 -1266
rect 690 -1278 696 -1272
rect 690 -1284 696 -1278
rect 690 -1290 696 -1284
rect 690 -1296 696 -1290
rect 690 -1302 696 -1296
rect 690 -1308 696 -1302
rect 690 -1314 696 -1308
rect 690 -1320 696 -1314
rect 690 -1326 696 -1320
rect 690 -1332 696 -1326
rect 690 -1338 696 -1332
rect 690 -1344 696 -1338
rect 690 -1350 696 -1344
rect 690 -1356 696 -1350
rect 690 -1362 696 -1356
rect 690 -1368 696 -1362
rect 690 -1374 696 -1368
rect 690 -1380 696 -1374
rect 690 -1386 696 -1380
rect 690 -1392 696 -1386
rect 690 -1398 696 -1392
rect 690 -1404 696 -1398
rect 690 -1410 696 -1404
rect 690 -1416 696 -1410
rect 690 -1422 696 -1416
rect 690 -1428 696 -1422
rect 690 -1434 696 -1428
rect 690 -1440 696 -1434
rect 690 -1446 696 -1440
rect 690 -1452 696 -1446
rect 690 -3180 696 -3174
rect 690 -3186 696 -3180
rect 690 -3192 696 -3186
rect 690 -3198 696 -3192
rect 690 -3204 696 -3198
rect 690 -3210 696 -3204
rect 690 -3216 696 -3210
rect 690 -3222 696 -3216
rect 690 -3228 696 -3222
rect 690 -3234 696 -3228
rect 690 -3240 696 -3234
rect 690 -3246 696 -3240
rect 690 -3252 696 -3246
rect 690 -3258 696 -3252
rect 690 -3264 696 -3258
rect 690 -3270 696 -3264
rect 690 -3276 696 -3270
rect 690 -3282 696 -3276
rect 690 -3288 696 -3282
rect 690 -3294 696 -3288
rect 690 -3300 696 -3294
rect 690 -3306 696 -3300
rect 690 -3312 696 -3306
rect 690 -3318 696 -3312
rect 690 -3324 696 -3318
rect 690 -3330 696 -3324
rect 690 -3336 696 -3330
rect 690 -3342 696 -3336
rect 690 -3348 696 -3342
rect 690 -3354 696 -3348
rect 690 -3360 696 -3354
rect 690 -3366 696 -3360
rect 690 -3372 696 -3366
rect 690 -3378 696 -3372
rect 690 -3384 696 -3378
rect 690 -3390 696 -3384
rect 690 -3396 696 -3390
rect 690 -3402 696 -3396
rect 690 -3408 696 -3402
rect 696 -1218 702 -1212
rect 696 -1224 702 -1218
rect 696 -1230 702 -1224
rect 696 -1236 702 -1230
rect 696 -1242 702 -1236
rect 696 -1248 702 -1242
rect 696 -1254 702 -1248
rect 696 -1260 702 -1254
rect 696 -1266 702 -1260
rect 696 -1272 702 -1266
rect 696 -1278 702 -1272
rect 696 -1284 702 -1278
rect 696 -1290 702 -1284
rect 696 -1296 702 -1290
rect 696 -1302 702 -1296
rect 696 -1308 702 -1302
rect 696 -1314 702 -1308
rect 696 -1320 702 -1314
rect 696 -1326 702 -1320
rect 696 -1332 702 -1326
rect 696 -1338 702 -1332
rect 696 -1344 702 -1338
rect 696 -1350 702 -1344
rect 696 -1356 702 -1350
rect 696 -1362 702 -1356
rect 696 -1368 702 -1362
rect 696 -1374 702 -1368
rect 696 -1380 702 -1374
rect 696 -1386 702 -1380
rect 696 -1392 702 -1386
rect 696 -1398 702 -1392
rect 696 -1404 702 -1398
rect 696 -1410 702 -1404
rect 696 -1416 702 -1410
rect 696 -1422 702 -1416
rect 696 -1428 702 -1422
rect 696 -1434 702 -1428
rect 696 -1440 702 -1434
rect 696 -1446 702 -1440
rect 696 -3180 702 -3174
rect 696 -3186 702 -3180
rect 696 -3192 702 -3186
rect 696 -3198 702 -3192
rect 696 -3204 702 -3198
rect 696 -3210 702 -3204
rect 696 -3216 702 -3210
rect 696 -3222 702 -3216
rect 696 -3228 702 -3222
rect 696 -3234 702 -3228
rect 696 -3240 702 -3234
rect 696 -3246 702 -3240
rect 696 -3252 702 -3246
rect 696 -3258 702 -3252
rect 696 -3264 702 -3258
rect 696 -3270 702 -3264
rect 696 -3276 702 -3270
rect 696 -3282 702 -3276
rect 696 -3288 702 -3282
rect 696 -3294 702 -3288
rect 696 -3300 702 -3294
rect 696 -3306 702 -3300
rect 696 -3312 702 -3306
rect 696 -3318 702 -3312
rect 696 -3324 702 -3318
rect 696 -3330 702 -3324
rect 696 -3336 702 -3330
rect 696 -3342 702 -3336
rect 696 -3348 702 -3342
rect 696 -3354 702 -3348
rect 696 -3360 702 -3354
rect 696 -3366 702 -3360
rect 696 -3372 702 -3366
rect 696 -3378 702 -3372
rect 696 -3384 702 -3378
rect 696 -3390 702 -3384
rect 696 -3396 702 -3390
rect 696 -3402 702 -3396
rect 696 -3408 702 -3402
rect 696 -3414 702 -3408
rect 702 -1218 708 -1212
rect 702 -1224 708 -1218
rect 702 -1230 708 -1224
rect 702 -1236 708 -1230
rect 702 -1242 708 -1236
rect 702 -1248 708 -1242
rect 702 -1254 708 -1248
rect 702 -1260 708 -1254
rect 702 -1266 708 -1260
rect 702 -1272 708 -1266
rect 702 -1278 708 -1272
rect 702 -1284 708 -1278
rect 702 -1290 708 -1284
rect 702 -1296 708 -1290
rect 702 -1302 708 -1296
rect 702 -1308 708 -1302
rect 702 -1314 708 -1308
rect 702 -1320 708 -1314
rect 702 -1326 708 -1320
rect 702 -1332 708 -1326
rect 702 -1338 708 -1332
rect 702 -1344 708 -1338
rect 702 -1350 708 -1344
rect 702 -1356 708 -1350
rect 702 -1362 708 -1356
rect 702 -1368 708 -1362
rect 702 -1374 708 -1368
rect 702 -1380 708 -1374
rect 702 -1386 708 -1380
rect 702 -1392 708 -1386
rect 702 -1398 708 -1392
rect 702 -1404 708 -1398
rect 702 -1410 708 -1404
rect 702 -1416 708 -1410
rect 702 -1422 708 -1416
rect 702 -1428 708 -1422
rect 702 -1434 708 -1428
rect 702 -1440 708 -1434
rect 702 -1446 708 -1440
rect 702 -3186 708 -3180
rect 702 -3192 708 -3186
rect 702 -3198 708 -3192
rect 702 -3204 708 -3198
rect 702 -3210 708 -3204
rect 702 -3216 708 -3210
rect 702 -3222 708 -3216
rect 702 -3228 708 -3222
rect 702 -3234 708 -3228
rect 702 -3240 708 -3234
rect 702 -3246 708 -3240
rect 702 -3252 708 -3246
rect 702 -3258 708 -3252
rect 702 -3264 708 -3258
rect 702 -3270 708 -3264
rect 702 -3276 708 -3270
rect 702 -3282 708 -3276
rect 702 -3288 708 -3282
rect 702 -3294 708 -3288
rect 702 -3300 708 -3294
rect 702 -3306 708 -3300
rect 702 -3312 708 -3306
rect 702 -3318 708 -3312
rect 702 -3324 708 -3318
rect 702 -3330 708 -3324
rect 702 -3336 708 -3330
rect 702 -3342 708 -3336
rect 702 -3348 708 -3342
rect 702 -3354 708 -3348
rect 702 -3360 708 -3354
rect 702 -3366 708 -3360
rect 702 -3372 708 -3366
rect 702 -3378 708 -3372
rect 702 -3384 708 -3378
rect 702 -3390 708 -3384
rect 702 -3396 708 -3390
rect 702 -3402 708 -3396
rect 702 -3408 708 -3402
rect 702 -3414 708 -3408
rect 708 -1212 714 -1206
rect 708 -1218 714 -1212
rect 708 -1224 714 -1218
rect 708 -1230 714 -1224
rect 708 -1236 714 -1230
rect 708 -1242 714 -1236
rect 708 -1248 714 -1242
rect 708 -1254 714 -1248
rect 708 -1260 714 -1254
rect 708 -1266 714 -1260
rect 708 -1272 714 -1266
rect 708 -1278 714 -1272
rect 708 -1284 714 -1278
rect 708 -1290 714 -1284
rect 708 -1296 714 -1290
rect 708 -1302 714 -1296
rect 708 -1308 714 -1302
rect 708 -1314 714 -1308
rect 708 -1320 714 -1314
rect 708 -1326 714 -1320
rect 708 -1332 714 -1326
rect 708 -1338 714 -1332
rect 708 -1344 714 -1338
rect 708 -1350 714 -1344
rect 708 -1356 714 -1350
rect 708 -1362 714 -1356
rect 708 -1368 714 -1362
rect 708 -1374 714 -1368
rect 708 -1380 714 -1374
rect 708 -1386 714 -1380
rect 708 -1392 714 -1386
rect 708 -1398 714 -1392
rect 708 -1404 714 -1398
rect 708 -1410 714 -1404
rect 708 -1416 714 -1410
rect 708 -1422 714 -1416
rect 708 -1428 714 -1422
rect 708 -1434 714 -1428
rect 708 -1440 714 -1434
rect 708 -3186 714 -3180
rect 708 -3192 714 -3186
rect 708 -3198 714 -3192
rect 708 -3204 714 -3198
rect 708 -3210 714 -3204
rect 708 -3216 714 -3210
rect 708 -3222 714 -3216
rect 708 -3228 714 -3222
rect 708 -3234 714 -3228
rect 708 -3240 714 -3234
rect 708 -3246 714 -3240
rect 708 -3252 714 -3246
rect 708 -3258 714 -3252
rect 708 -3264 714 -3258
rect 708 -3270 714 -3264
rect 708 -3276 714 -3270
rect 708 -3282 714 -3276
rect 708 -3288 714 -3282
rect 708 -3294 714 -3288
rect 708 -3300 714 -3294
rect 708 -3306 714 -3300
rect 708 -3312 714 -3306
rect 708 -3318 714 -3312
rect 708 -3324 714 -3318
rect 708 -3330 714 -3324
rect 708 -3336 714 -3330
rect 708 -3342 714 -3336
rect 708 -3348 714 -3342
rect 708 -3354 714 -3348
rect 708 -3360 714 -3354
rect 708 -3366 714 -3360
rect 708 -3372 714 -3366
rect 708 -3378 714 -3372
rect 708 -3384 714 -3378
rect 708 -3390 714 -3384
rect 708 -3396 714 -3390
rect 708 -3402 714 -3396
rect 708 -3408 714 -3402
rect 708 -3414 714 -3408
rect 708 -3420 714 -3414
rect 714 -1212 720 -1206
rect 714 -1218 720 -1212
rect 714 -1224 720 -1218
rect 714 -1230 720 -1224
rect 714 -1236 720 -1230
rect 714 -1242 720 -1236
rect 714 -1248 720 -1242
rect 714 -1254 720 -1248
rect 714 -1260 720 -1254
rect 714 -1266 720 -1260
rect 714 -1272 720 -1266
rect 714 -1278 720 -1272
rect 714 -1284 720 -1278
rect 714 -1290 720 -1284
rect 714 -1296 720 -1290
rect 714 -1302 720 -1296
rect 714 -1308 720 -1302
rect 714 -1314 720 -1308
rect 714 -1320 720 -1314
rect 714 -1326 720 -1320
rect 714 -1332 720 -1326
rect 714 -1338 720 -1332
rect 714 -1344 720 -1338
rect 714 -1350 720 -1344
rect 714 -1356 720 -1350
rect 714 -1362 720 -1356
rect 714 -1368 720 -1362
rect 714 -1374 720 -1368
rect 714 -1380 720 -1374
rect 714 -1386 720 -1380
rect 714 -1392 720 -1386
rect 714 -1398 720 -1392
rect 714 -1404 720 -1398
rect 714 -1410 720 -1404
rect 714 -1416 720 -1410
rect 714 -1422 720 -1416
rect 714 -1428 720 -1422
rect 714 -1434 720 -1428
rect 714 -1440 720 -1434
rect 714 -3192 720 -3186
rect 714 -3198 720 -3192
rect 714 -3204 720 -3198
rect 714 -3210 720 -3204
rect 714 -3216 720 -3210
rect 714 -3222 720 -3216
rect 714 -3228 720 -3222
rect 714 -3234 720 -3228
rect 714 -3240 720 -3234
rect 714 -3246 720 -3240
rect 714 -3252 720 -3246
rect 714 -3258 720 -3252
rect 714 -3264 720 -3258
rect 714 -3270 720 -3264
rect 714 -3276 720 -3270
rect 714 -3282 720 -3276
rect 714 -3288 720 -3282
rect 714 -3294 720 -3288
rect 714 -3300 720 -3294
rect 714 -3306 720 -3300
rect 714 -3312 720 -3306
rect 714 -3318 720 -3312
rect 714 -3324 720 -3318
rect 714 -3330 720 -3324
rect 714 -3336 720 -3330
rect 714 -3342 720 -3336
rect 714 -3348 720 -3342
rect 714 -3354 720 -3348
rect 714 -3360 720 -3354
rect 714 -3366 720 -3360
rect 714 -3372 720 -3366
rect 714 -3378 720 -3372
rect 714 -3384 720 -3378
rect 714 -3390 720 -3384
rect 714 -3396 720 -3390
rect 720 -1206 726 -1200
rect 720 -1212 726 -1206
rect 720 -1218 726 -1212
rect 720 -1224 726 -1218
rect 720 -1230 726 -1224
rect 720 -1236 726 -1230
rect 720 -1242 726 -1236
rect 720 -1248 726 -1242
rect 720 -1254 726 -1248
rect 720 -1260 726 -1254
rect 720 -1266 726 -1260
rect 720 -1272 726 -1266
rect 720 -1278 726 -1272
rect 720 -1284 726 -1278
rect 720 -1290 726 -1284
rect 720 -1296 726 -1290
rect 720 -1302 726 -1296
rect 720 -1308 726 -1302
rect 720 -1314 726 -1308
rect 720 -1320 726 -1314
rect 720 -1326 726 -1320
rect 720 -1332 726 -1326
rect 720 -1338 726 -1332
rect 720 -1344 726 -1338
rect 720 -1350 726 -1344
rect 720 -1356 726 -1350
rect 720 -1362 726 -1356
rect 720 -1368 726 -1362
rect 720 -1374 726 -1368
rect 720 -1380 726 -1374
rect 720 -1386 726 -1380
rect 720 -1392 726 -1386
rect 720 -1398 726 -1392
rect 720 -1404 726 -1398
rect 720 -1410 726 -1404
rect 720 -1416 726 -1410
rect 720 -1422 726 -1416
rect 720 -1428 726 -1422
rect 720 -1434 726 -1428
rect 720 -3192 726 -3186
rect 720 -3198 726 -3192
rect 720 -3204 726 -3198
rect 720 -3210 726 -3204
rect 720 -3216 726 -3210
rect 720 -3222 726 -3216
rect 720 -3228 726 -3222
rect 720 -3234 726 -3228
rect 720 -3240 726 -3234
rect 720 -3246 726 -3240
rect 720 -3252 726 -3246
rect 720 -3258 726 -3252
rect 720 -3264 726 -3258
rect 720 -3270 726 -3264
rect 720 -3276 726 -3270
rect 720 -3282 726 -3276
rect 720 -3288 726 -3282
rect 720 -3294 726 -3288
rect 720 -3300 726 -3294
rect 720 -3306 726 -3300
rect 720 -3312 726 -3306
rect 720 -3318 726 -3312
rect 720 -3324 726 -3318
rect 720 -3330 726 -3324
rect 720 -3336 726 -3330
rect 720 -3342 726 -3336
rect 720 -3348 726 -3342
rect 726 -1206 732 -1200
rect 726 -1212 732 -1206
rect 726 -1218 732 -1212
rect 726 -1224 732 -1218
rect 726 -1230 732 -1224
rect 726 -1236 732 -1230
rect 726 -1242 732 -1236
rect 726 -1248 732 -1242
rect 726 -1254 732 -1248
rect 726 -1260 732 -1254
rect 726 -1266 732 -1260
rect 726 -1272 732 -1266
rect 726 -1278 732 -1272
rect 726 -1284 732 -1278
rect 726 -1290 732 -1284
rect 726 -1296 732 -1290
rect 726 -1302 732 -1296
rect 726 -1308 732 -1302
rect 726 -1314 732 -1308
rect 726 -1320 732 -1314
rect 726 -1326 732 -1320
rect 726 -1332 732 -1326
rect 726 -1338 732 -1332
rect 726 -1344 732 -1338
rect 726 -1350 732 -1344
rect 726 -1356 732 -1350
rect 726 -1362 732 -1356
rect 726 -1368 732 -1362
rect 726 -1374 732 -1368
rect 726 -1380 732 -1374
rect 726 -1386 732 -1380
rect 726 -1392 732 -1386
rect 726 -1398 732 -1392
rect 726 -1404 732 -1398
rect 726 -1410 732 -1404
rect 726 -1416 732 -1410
rect 726 -1422 732 -1416
rect 726 -1428 732 -1422
rect 726 -1434 732 -1428
rect 726 -3198 732 -3192
rect 726 -3204 732 -3198
rect 726 -3210 732 -3204
rect 726 -3216 732 -3210
rect 726 -3222 732 -3216
rect 726 -3228 732 -3222
rect 726 -3234 732 -3228
rect 726 -3240 732 -3234
rect 726 -3246 732 -3240
rect 726 -3252 732 -3246
rect 726 -3258 732 -3252
rect 726 -3264 732 -3258
rect 726 -3270 732 -3264
rect 726 -3276 732 -3270
rect 726 -3282 732 -3276
rect 726 -3288 732 -3282
rect 726 -3294 732 -3288
rect 726 -3300 732 -3294
rect 732 -1200 738 -1194
rect 732 -1206 738 -1200
rect 732 -1212 738 -1206
rect 732 -1218 738 -1212
rect 732 -1224 738 -1218
rect 732 -1230 738 -1224
rect 732 -1236 738 -1230
rect 732 -1242 738 -1236
rect 732 -1248 738 -1242
rect 732 -1254 738 -1248
rect 732 -1260 738 -1254
rect 732 -1266 738 -1260
rect 732 -1272 738 -1266
rect 732 -1278 738 -1272
rect 732 -1284 738 -1278
rect 732 -1290 738 -1284
rect 732 -1296 738 -1290
rect 732 -1302 738 -1296
rect 732 -1308 738 -1302
rect 732 -1314 738 -1308
rect 732 -1320 738 -1314
rect 732 -1326 738 -1320
rect 732 -1332 738 -1326
rect 732 -1338 738 -1332
rect 732 -1344 738 -1338
rect 732 -1350 738 -1344
rect 732 -1356 738 -1350
rect 732 -1362 738 -1356
rect 732 -1368 738 -1362
rect 732 -1374 738 -1368
rect 732 -1380 738 -1374
rect 732 -1386 738 -1380
rect 732 -1392 738 -1386
rect 732 -1398 738 -1392
rect 732 -1404 738 -1398
rect 732 -1410 738 -1404
rect 732 -1416 738 -1410
rect 732 -1422 738 -1416
rect 732 -1428 738 -1422
rect 732 -3198 738 -3192
rect 732 -3204 738 -3198
rect 732 -3210 738 -3204
rect 732 -3216 738 -3210
rect 732 -3222 738 -3216
rect 732 -3228 738 -3222
rect 732 -3234 738 -3228
rect 732 -3240 738 -3234
rect 732 -3246 738 -3240
rect 738 -1200 744 -1194
rect 738 -1206 744 -1200
rect 738 -1212 744 -1206
rect 738 -1218 744 -1212
rect 738 -1224 744 -1218
rect 738 -1230 744 -1224
rect 738 -1236 744 -1230
rect 738 -1242 744 -1236
rect 738 -1248 744 -1242
rect 738 -1254 744 -1248
rect 738 -1260 744 -1254
rect 738 -1266 744 -1260
rect 738 -1272 744 -1266
rect 738 -1278 744 -1272
rect 738 -1284 744 -1278
rect 738 -1290 744 -1284
rect 738 -1296 744 -1290
rect 738 -1302 744 -1296
rect 738 -1308 744 -1302
rect 738 -1314 744 -1308
rect 738 -1320 744 -1314
rect 738 -1326 744 -1320
rect 738 -1332 744 -1326
rect 738 -1338 744 -1332
rect 738 -1344 744 -1338
rect 738 -1350 744 -1344
rect 738 -1356 744 -1350
rect 738 -1362 744 -1356
rect 738 -1368 744 -1362
rect 738 -1374 744 -1368
rect 738 -1380 744 -1374
rect 738 -1386 744 -1380
rect 738 -1392 744 -1386
rect 738 -1398 744 -1392
rect 738 -1404 744 -1398
rect 738 -1410 744 -1404
rect 738 -1416 744 -1410
rect 738 -1422 744 -1416
rect 744 -1200 750 -1194
rect 744 -1206 750 -1200
rect 744 -1212 750 -1206
rect 744 -1218 750 -1212
rect 744 -1224 750 -1218
rect 744 -1230 750 -1224
rect 744 -1236 750 -1230
rect 744 -1242 750 -1236
rect 744 -1248 750 -1242
rect 744 -1254 750 -1248
rect 744 -1260 750 -1254
rect 744 -1266 750 -1260
rect 744 -1272 750 -1266
rect 744 -1278 750 -1272
rect 744 -1284 750 -1278
rect 744 -1290 750 -1284
rect 744 -1296 750 -1290
rect 744 -1302 750 -1296
rect 744 -1308 750 -1302
rect 744 -1314 750 -1308
rect 744 -1320 750 -1314
rect 744 -1326 750 -1320
rect 744 -1332 750 -1326
rect 744 -1338 750 -1332
rect 744 -1344 750 -1338
rect 744 -1350 750 -1344
rect 744 -1356 750 -1350
rect 744 -1362 750 -1356
rect 744 -1368 750 -1362
rect 744 -1374 750 -1368
rect 744 -1380 750 -1374
rect 744 -1386 750 -1380
rect 744 -1392 750 -1386
rect 744 -1398 750 -1392
rect 744 -1404 750 -1398
rect 744 -1410 750 -1404
rect 744 -1416 750 -1410
rect 744 -1422 750 -1416
rect 750 -1194 756 -1188
rect 750 -1200 756 -1194
rect 750 -1206 756 -1200
rect 750 -1212 756 -1206
rect 750 -1218 756 -1212
rect 750 -1224 756 -1218
rect 750 -1230 756 -1224
rect 750 -1236 756 -1230
rect 750 -1242 756 -1236
rect 750 -1248 756 -1242
rect 750 -1254 756 -1248
rect 750 -1260 756 -1254
rect 750 -1266 756 -1260
rect 750 -1272 756 -1266
rect 750 -1278 756 -1272
rect 750 -1284 756 -1278
rect 750 -1290 756 -1284
rect 750 -1296 756 -1290
rect 750 -1302 756 -1296
rect 750 -1308 756 -1302
rect 750 -1314 756 -1308
rect 750 -1320 756 -1314
rect 750 -1326 756 -1320
rect 750 -1332 756 -1326
rect 750 -1338 756 -1332
rect 750 -1344 756 -1338
rect 750 -1350 756 -1344
rect 750 -1356 756 -1350
rect 750 -1362 756 -1356
rect 750 -1368 756 -1362
rect 750 -1374 756 -1368
rect 750 -1380 756 -1374
rect 750 -1386 756 -1380
rect 750 -1392 756 -1386
rect 750 -1398 756 -1392
rect 750 -1404 756 -1398
rect 750 -1410 756 -1404
rect 750 -1416 756 -1410
rect 756 -1194 762 -1188
rect 756 -1200 762 -1194
rect 756 -1206 762 -1200
rect 756 -1212 762 -1206
rect 756 -1218 762 -1212
rect 756 -1224 762 -1218
rect 756 -1230 762 -1224
rect 756 -1236 762 -1230
rect 756 -1242 762 -1236
rect 756 -1248 762 -1242
rect 756 -1254 762 -1248
rect 756 -1260 762 -1254
rect 756 -1266 762 -1260
rect 756 -1272 762 -1266
rect 756 -1278 762 -1272
rect 756 -1284 762 -1278
rect 756 -1290 762 -1284
rect 756 -1296 762 -1290
rect 756 -1302 762 -1296
rect 756 -1308 762 -1302
rect 756 -1314 762 -1308
rect 756 -1320 762 -1314
rect 756 -1326 762 -1320
rect 756 -1332 762 -1326
rect 756 -1338 762 -1332
rect 756 -1344 762 -1338
rect 756 -1350 762 -1344
rect 756 -1356 762 -1350
rect 756 -1362 762 -1356
rect 756 -1368 762 -1362
rect 756 -1374 762 -1368
rect 756 -1380 762 -1374
rect 756 -1386 762 -1380
rect 756 -1392 762 -1386
rect 756 -1398 762 -1392
rect 756 -1404 762 -1398
rect 756 -1410 762 -1404
rect 756 -1416 762 -1410
rect 762 -1188 768 -1182
rect 762 -1194 768 -1188
rect 762 -1200 768 -1194
rect 762 -1206 768 -1200
rect 762 -1212 768 -1206
rect 762 -1218 768 -1212
rect 762 -1224 768 -1218
rect 762 -1230 768 -1224
rect 762 -1236 768 -1230
rect 762 -1242 768 -1236
rect 762 -1248 768 -1242
rect 762 -1254 768 -1248
rect 762 -1260 768 -1254
rect 762 -1266 768 -1260
rect 762 -1272 768 -1266
rect 762 -1278 768 -1272
rect 762 -1284 768 -1278
rect 762 -1290 768 -1284
rect 762 -1296 768 -1290
rect 762 -1302 768 -1296
rect 762 -1308 768 -1302
rect 762 -1314 768 -1308
rect 762 -1320 768 -1314
rect 762 -1326 768 -1320
rect 762 -1332 768 -1326
rect 762 -1338 768 -1332
rect 762 -1344 768 -1338
rect 762 -1350 768 -1344
rect 762 -1356 768 -1350
rect 762 -1362 768 -1356
rect 762 -1368 768 -1362
rect 762 -1374 768 -1368
rect 762 -1380 768 -1374
rect 762 -1386 768 -1380
rect 762 -1392 768 -1386
rect 762 -1398 768 -1392
rect 762 -1404 768 -1398
rect 762 -1410 768 -1404
rect 762 -3414 768 -3408
rect 768 -1188 774 -1182
rect 768 -1194 774 -1188
rect 768 -1200 774 -1194
rect 768 -1206 774 -1200
rect 768 -1212 774 -1206
rect 768 -1218 774 -1212
rect 768 -1224 774 -1218
rect 768 -1230 774 -1224
rect 768 -1236 774 -1230
rect 768 -1242 774 -1236
rect 768 -1248 774 -1242
rect 768 -1254 774 -1248
rect 768 -1260 774 -1254
rect 768 -1266 774 -1260
rect 768 -1272 774 -1266
rect 768 -1278 774 -1272
rect 768 -1284 774 -1278
rect 768 -1290 774 -1284
rect 768 -1296 774 -1290
rect 768 -1302 774 -1296
rect 768 -1308 774 -1302
rect 768 -1314 774 -1308
rect 768 -1320 774 -1314
rect 768 -1326 774 -1320
rect 768 -1332 774 -1326
rect 768 -1338 774 -1332
rect 768 -1344 774 -1338
rect 768 -1350 774 -1344
rect 768 -1356 774 -1350
rect 768 -1362 774 -1356
rect 768 -1368 774 -1362
rect 768 -1374 774 -1368
rect 768 -1380 774 -1374
rect 768 -1386 774 -1380
rect 768 -1392 774 -1386
rect 768 -1398 774 -1392
rect 768 -1404 774 -1398
rect 768 -1410 774 -1404
rect 768 -3384 774 -3378
rect 768 -3390 774 -3384
rect 768 -3396 774 -3390
rect 768 -3402 774 -3396
rect 774 -1188 780 -1182
rect 774 -1194 780 -1188
rect 774 -1200 780 -1194
rect 774 -1206 780 -1200
rect 774 -1212 780 -1206
rect 774 -1218 780 -1212
rect 774 -1224 780 -1218
rect 774 -1230 780 -1224
rect 774 -1236 780 -1230
rect 774 -1242 780 -1236
rect 774 -1248 780 -1242
rect 774 -1254 780 -1248
rect 774 -1260 780 -1254
rect 774 -1266 780 -1260
rect 774 -1272 780 -1266
rect 774 -1278 780 -1272
rect 774 -1284 780 -1278
rect 774 -1290 780 -1284
rect 774 -1296 780 -1290
rect 774 -1302 780 -1296
rect 774 -1308 780 -1302
rect 774 -1314 780 -1308
rect 774 -1320 780 -1314
rect 774 -1326 780 -1320
rect 774 -1332 780 -1326
rect 774 -1338 780 -1332
rect 774 -1344 780 -1338
rect 774 -1350 780 -1344
rect 774 -1356 780 -1350
rect 774 -1362 780 -1356
rect 774 -1368 780 -1362
rect 774 -1374 780 -1368
rect 774 -1380 780 -1374
rect 774 -1386 780 -1380
rect 774 -1392 780 -1386
rect 774 -1398 780 -1392
rect 774 -1404 780 -1398
rect 774 -3354 780 -3348
rect 774 -3360 780 -3354
rect 774 -3366 780 -3360
rect 774 -3372 780 -3366
rect 774 -3378 780 -3372
rect 774 -3384 780 -3378
rect 774 -3390 780 -3384
rect 780 -1182 786 -1176
rect 780 -1188 786 -1182
rect 780 -1194 786 -1188
rect 780 -1200 786 -1194
rect 780 -1206 786 -1200
rect 780 -1212 786 -1206
rect 780 -1218 786 -1212
rect 780 -1224 786 -1218
rect 780 -1230 786 -1224
rect 780 -1236 786 -1230
rect 780 -1242 786 -1236
rect 780 -1248 786 -1242
rect 780 -1254 786 -1248
rect 780 -1260 786 -1254
rect 780 -1266 786 -1260
rect 780 -1272 786 -1266
rect 780 -1278 786 -1272
rect 780 -1284 786 -1278
rect 780 -1290 786 -1284
rect 780 -1296 786 -1290
rect 780 -1302 786 -1296
rect 780 -1308 786 -1302
rect 780 -1314 786 -1308
rect 780 -1320 786 -1314
rect 780 -1326 786 -1320
rect 780 -1332 786 -1326
rect 780 -1338 786 -1332
rect 780 -1344 786 -1338
rect 780 -1350 786 -1344
rect 780 -1356 786 -1350
rect 780 -1362 786 -1356
rect 780 -1368 786 -1362
rect 780 -1374 786 -1368
rect 780 -1380 786 -1374
rect 780 -1386 786 -1380
rect 780 -1392 786 -1386
rect 780 -1398 786 -1392
rect 780 -1404 786 -1398
rect 780 -3318 786 -3312
rect 780 -3324 786 -3318
rect 780 -3330 786 -3324
rect 780 -3336 786 -3330
rect 780 -3342 786 -3336
rect 780 -3348 786 -3342
rect 780 -3354 786 -3348
rect 780 -3360 786 -3354
rect 780 -3366 786 -3360
rect 780 -3372 786 -3366
rect 780 -3378 786 -3372
rect 786 -1182 792 -1176
rect 786 -1188 792 -1182
rect 786 -1194 792 -1188
rect 786 -1200 792 -1194
rect 786 -1206 792 -1200
rect 786 -1212 792 -1206
rect 786 -1218 792 -1212
rect 786 -1224 792 -1218
rect 786 -1230 792 -1224
rect 786 -1236 792 -1230
rect 786 -1242 792 -1236
rect 786 -1248 792 -1242
rect 786 -1254 792 -1248
rect 786 -1260 792 -1254
rect 786 -1266 792 -1260
rect 786 -1272 792 -1266
rect 786 -1278 792 -1272
rect 786 -1284 792 -1278
rect 786 -1290 792 -1284
rect 786 -1296 792 -1290
rect 786 -1302 792 -1296
rect 786 -1308 792 -1302
rect 786 -1314 792 -1308
rect 786 -1320 792 -1314
rect 786 -1326 792 -1320
rect 786 -1332 792 -1326
rect 786 -1338 792 -1332
rect 786 -1344 792 -1338
rect 786 -1350 792 -1344
rect 786 -1356 792 -1350
rect 786 -1362 792 -1356
rect 786 -1368 792 -1362
rect 786 -1374 792 -1368
rect 786 -1380 792 -1374
rect 786 -1386 792 -1380
rect 786 -1392 792 -1386
rect 786 -1398 792 -1392
rect 786 -3288 792 -3282
rect 786 -3294 792 -3288
rect 786 -3300 792 -3294
rect 786 -3306 792 -3300
rect 786 -3312 792 -3306
rect 786 -3318 792 -3312
rect 786 -3324 792 -3318
rect 786 -3330 792 -3324
rect 786 -3336 792 -3330
rect 786 -3342 792 -3336
rect 786 -3348 792 -3342
rect 786 -3354 792 -3348
rect 786 -3360 792 -3354
rect 786 -3366 792 -3360
rect 792 -1176 798 -1170
rect 792 -1182 798 -1176
rect 792 -1188 798 -1182
rect 792 -1194 798 -1188
rect 792 -1200 798 -1194
rect 792 -1206 798 -1200
rect 792 -1212 798 -1206
rect 792 -1218 798 -1212
rect 792 -1224 798 -1218
rect 792 -1230 798 -1224
rect 792 -1236 798 -1230
rect 792 -1242 798 -1236
rect 792 -1248 798 -1242
rect 792 -1254 798 -1248
rect 792 -1260 798 -1254
rect 792 -1266 798 -1260
rect 792 -1272 798 -1266
rect 792 -1278 798 -1272
rect 792 -1284 798 -1278
rect 792 -1290 798 -1284
rect 792 -1296 798 -1290
rect 792 -1302 798 -1296
rect 792 -1308 798 -1302
rect 792 -1314 798 -1308
rect 792 -1320 798 -1314
rect 792 -1326 798 -1320
rect 792 -1332 798 -1326
rect 792 -1338 798 -1332
rect 792 -1344 798 -1338
rect 792 -1350 798 -1344
rect 792 -1356 798 -1350
rect 792 -1362 798 -1356
rect 792 -1368 798 -1362
rect 792 -1374 798 -1368
rect 792 -1380 798 -1374
rect 792 -1386 798 -1380
rect 792 -1392 798 -1386
rect 792 -1398 798 -1392
rect 792 -3258 798 -3252
rect 792 -3264 798 -3258
rect 792 -3270 798 -3264
rect 792 -3276 798 -3270
rect 792 -3282 798 -3276
rect 792 -3288 798 -3282
rect 792 -3294 798 -3288
rect 792 -3300 798 -3294
rect 792 -3306 798 -3300
rect 792 -3312 798 -3306
rect 792 -3318 798 -3312
rect 792 -3324 798 -3318
rect 792 -3330 798 -3324
rect 792 -3336 798 -3330
rect 792 -3342 798 -3336
rect 792 -3348 798 -3342
rect 792 -3354 798 -3348
rect 798 -1176 804 -1170
rect 798 -1182 804 -1176
rect 798 -1188 804 -1182
rect 798 -1194 804 -1188
rect 798 -1200 804 -1194
rect 798 -1206 804 -1200
rect 798 -1212 804 -1206
rect 798 -1218 804 -1212
rect 798 -1224 804 -1218
rect 798 -1230 804 -1224
rect 798 -1236 804 -1230
rect 798 -1242 804 -1236
rect 798 -1248 804 -1242
rect 798 -1254 804 -1248
rect 798 -1260 804 -1254
rect 798 -1266 804 -1260
rect 798 -1272 804 -1266
rect 798 -1278 804 -1272
rect 798 -1284 804 -1278
rect 798 -1290 804 -1284
rect 798 -1296 804 -1290
rect 798 -1302 804 -1296
rect 798 -1308 804 -1302
rect 798 -1314 804 -1308
rect 798 -1320 804 -1314
rect 798 -1326 804 -1320
rect 798 -1332 804 -1326
rect 798 -1338 804 -1332
rect 798 -1344 804 -1338
rect 798 -1350 804 -1344
rect 798 -1356 804 -1350
rect 798 -1362 804 -1356
rect 798 -1368 804 -1362
rect 798 -1374 804 -1368
rect 798 -1380 804 -1374
rect 798 -1386 804 -1380
rect 798 -1392 804 -1386
rect 798 -1398 804 -1392
rect 798 -3228 804 -3222
rect 798 -3234 804 -3228
rect 798 -3240 804 -3234
rect 798 -3246 804 -3240
rect 798 -3252 804 -3246
rect 798 -3258 804 -3252
rect 798 -3264 804 -3258
rect 798 -3270 804 -3264
rect 798 -3276 804 -3270
rect 798 -3282 804 -3276
rect 798 -3288 804 -3282
rect 798 -3294 804 -3288
rect 798 -3300 804 -3294
rect 798 -3306 804 -3300
rect 798 -3312 804 -3306
rect 798 -3318 804 -3312
rect 798 -3324 804 -3318
rect 798 -3330 804 -3324
rect 798 -3336 804 -3330
rect 798 -3342 804 -3336
rect 804 -1176 810 -1170
rect 804 -1182 810 -1176
rect 804 -1188 810 -1182
rect 804 -1194 810 -1188
rect 804 -1200 810 -1194
rect 804 -1206 810 -1200
rect 804 -1212 810 -1206
rect 804 -1218 810 -1212
rect 804 -1224 810 -1218
rect 804 -1230 810 -1224
rect 804 -1236 810 -1230
rect 804 -1242 810 -1236
rect 804 -1248 810 -1242
rect 804 -1254 810 -1248
rect 804 -1260 810 -1254
rect 804 -1266 810 -1260
rect 804 -1272 810 -1266
rect 804 -1278 810 -1272
rect 804 -1284 810 -1278
rect 804 -1290 810 -1284
rect 804 -1296 810 -1290
rect 804 -1302 810 -1296
rect 804 -1308 810 -1302
rect 804 -1314 810 -1308
rect 804 -1320 810 -1314
rect 804 -1326 810 -1320
rect 804 -1332 810 -1326
rect 804 -1338 810 -1332
rect 804 -1344 810 -1338
rect 804 -1350 810 -1344
rect 804 -1356 810 -1350
rect 804 -1362 810 -1356
rect 804 -1368 810 -1362
rect 804 -1374 810 -1368
rect 804 -1380 810 -1374
rect 804 -1386 810 -1380
rect 804 -1392 810 -1386
rect 804 -3198 810 -3192
rect 804 -3204 810 -3198
rect 804 -3210 810 -3204
rect 804 -3216 810 -3210
rect 804 -3222 810 -3216
rect 804 -3228 810 -3222
rect 804 -3234 810 -3228
rect 804 -3240 810 -3234
rect 804 -3246 810 -3240
rect 804 -3252 810 -3246
rect 804 -3258 810 -3252
rect 804 -3264 810 -3258
rect 804 -3270 810 -3264
rect 804 -3276 810 -3270
rect 804 -3282 810 -3276
rect 804 -3288 810 -3282
rect 804 -3294 810 -3288
rect 804 -3300 810 -3294
rect 804 -3306 810 -3300
rect 804 -3312 810 -3306
rect 804 -3318 810 -3312
rect 804 -3324 810 -3318
rect 804 -3330 810 -3324
rect 810 -1170 816 -1164
rect 810 -1176 816 -1170
rect 810 -1182 816 -1176
rect 810 -1188 816 -1182
rect 810 -1194 816 -1188
rect 810 -1200 816 -1194
rect 810 -1206 816 -1200
rect 810 -1212 816 -1206
rect 810 -1218 816 -1212
rect 810 -1224 816 -1218
rect 810 -1230 816 -1224
rect 810 -1236 816 -1230
rect 810 -1242 816 -1236
rect 810 -1248 816 -1242
rect 810 -1254 816 -1248
rect 810 -1260 816 -1254
rect 810 -1266 816 -1260
rect 810 -1272 816 -1266
rect 810 -1278 816 -1272
rect 810 -1284 816 -1278
rect 810 -1290 816 -1284
rect 810 -1296 816 -1290
rect 810 -1302 816 -1296
rect 810 -1308 816 -1302
rect 810 -1314 816 -1308
rect 810 -1320 816 -1314
rect 810 -1326 816 -1320
rect 810 -1332 816 -1326
rect 810 -1338 816 -1332
rect 810 -1344 816 -1338
rect 810 -1350 816 -1344
rect 810 -1356 816 -1350
rect 810 -1362 816 -1356
rect 810 -1368 816 -1362
rect 810 -1374 816 -1368
rect 810 -1380 816 -1374
rect 810 -1386 816 -1380
rect 810 -1392 816 -1386
rect 810 -3162 816 -3156
rect 810 -3168 816 -3162
rect 810 -3174 816 -3168
rect 810 -3180 816 -3174
rect 810 -3186 816 -3180
rect 810 -3192 816 -3186
rect 810 -3198 816 -3192
rect 810 -3204 816 -3198
rect 810 -3210 816 -3204
rect 810 -3216 816 -3210
rect 810 -3222 816 -3216
rect 810 -3228 816 -3222
rect 810 -3234 816 -3228
rect 810 -3240 816 -3234
rect 810 -3246 816 -3240
rect 810 -3252 816 -3246
rect 810 -3258 816 -3252
rect 810 -3264 816 -3258
rect 810 -3270 816 -3264
rect 810 -3276 816 -3270
rect 810 -3282 816 -3276
rect 810 -3288 816 -3282
rect 810 -3294 816 -3288
rect 810 -3300 816 -3294
rect 810 -3306 816 -3300
rect 810 -3312 816 -3306
rect 810 -3318 816 -3312
rect 816 -1170 822 -1164
rect 816 -1176 822 -1170
rect 816 -1182 822 -1176
rect 816 -1188 822 -1182
rect 816 -1194 822 -1188
rect 816 -1200 822 -1194
rect 816 -1206 822 -1200
rect 816 -1212 822 -1206
rect 816 -1218 822 -1212
rect 816 -1224 822 -1218
rect 816 -1230 822 -1224
rect 816 -1236 822 -1230
rect 816 -1242 822 -1236
rect 816 -1248 822 -1242
rect 816 -1254 822 -1248
rect 816 -1260 822 -1254
rect 816 -1266 822 -1260
rect 816 -1272 822 -1266
rect 816 -1278 822 -1272
rect 816 -1284 822 -1278
rect 816 -1290 822 -1284
rect 816 -1296 822 -1290
rect 816 -1302 822 -1296
rect 816 -1308 822 -1302
rect 816 -1314 822 -1308
rect 816 -1320 822 -1314
rect 816 -1326 822 -1320
rect 816 -1332 822 -1326
rect 816 -1338 822 -1332
rect 816 -1344 822 -1338
rect 816 -1350 822 -1344
rect 816 -1356 822 -1350
rect 816 -1362 822 -1356
rect 816 -1368 822 -1362
rect 816 -1374 822 -1368
rect 816 -1380 822 -1374
rect 816 -1386 822 -1380
rect 816 -3132 822 -3126
rect 816 -3138 822 -3132
rect 816 -3144 822 -3138
rect 816 -3150 822 -3144
rect 816 -3156 822 -3150
rect 816 -3162 822 -3156
rect 816 -3168 822 -3162
rect 816 -3174 822 -3168
rect 816 -3180 822 -3174
rect 816 -3186 822 -3180
rect 816 -3192 822 -3186
rect 816 -3198 822 -3192
rect 816 -3204 822 -3198
rect 816 -3210 822 -3204
rect 816 -3216 822 -3210
rect 816 -3222 822 -3216
rect 816 -3228 822 -3222
rect 816 -3234 822 -3228
rect 816 -3240 822 -3234
rect 816 -3246 822 -3240
rect 816 -3252 822 -3246
rect 816 -3258 822 -3252
rect 816 -3264 822 -3258
rect 816 -3270 822 -3264
rect 816 -3276 822 -3270
rect 816 -3282 822 -3276
rect 816 -3288 822 -3282
rect 816 -3294 822 -3288
rect 816 -3300 822 -3294
rect 822 -1170 828 -1164
rect 822 -1176 828 -1170
rect 822 -1182 828 -1176
rect 822 -1188 828 -1182
rect 822 -1194 828 -1188
rect 822 -1200 828 -1194
rect 822 -1206 828 -1200
rect 822 -1212 828 -1206
rect 822 -1218 828 -1212
rect 822 -1224 828 -1218
rect 822 -1230 828 -1224
rect 822 -1236 828 -1230
rect 822 -1242 828 -1236
rect 822 -1248 828 -1242
rect 822 -1254 828 -1248
rect 822 -1260 828 -1254
rect 822 -1266 828 -1260
rect 822 -1272 828 -1266
rect 822 -1278 828 -1272
rect 822 -1284 828 -1278
rect 822 -1290 828 -1284
rect 822 -1296 828 -1290
rect 822 -1302 828 -1296
rect 822 -1308 828 -1302
rect 822 -1314 828 -1308
rect 822 -1320 828 -1314
rect 822 -1326 828 -1320
rect 822 -1332 828 -1326
rect 822 -1338 828 -1332
rect 822 -1344 828 -1338
rect 822 -1350 828 -1344
rect 822 -1356 828 -1350
rect 822 -1362 828 -1356
rect 822 -1368 828 -1362
rect 822 -1374 828 -1368
rect 822 -1380 828 -1374
rect 822 -1386 828 -1380
rect 822 -3108 828 -3102
rect 822 -3114 828 -3108
rect 822 -3120 828 -3114
rect 822 -3126 828 -3120
rect 822 -3132 828 -3126
rect 822 -3138 828 -3132
rect 822 -3144 828 -3138
rect 822 -3150 828 -3144
rect 822 -3156 828 -3150
rect 822 -3162 828 -3156
rect 822 -3168 828 -3162
rect 822 -3174 828 -3168
rect 822 -3180 828 -3174
rect 822 -3186 828 -3180
rect 822 -3192 828 -3186
rect 822 -3198 828 -3192
rect 822 -3204 828 -3198
rect 822 -3210 828 -3204
rect 822 -3216 828 -3210
rect 822 -3222 828 -3216
rect 822 -3228 828 -3222
rect 822 -3234 828 -3228
rect 822 -3240 828 -3234
rect 822 -3246 828 -3240
rect 822 -3252 828 -3246
rect 822 -3258 828 -3252
rect 822 -3264 828 -3258
rect 822 -3270 828 -3264
rect 822 -3276 828 -3270
rect 822 -3282 828 -3276
rect 822 -3288 828 -3282
rect 822 -3456 828 -3450
rect 828 -1164 834 -1158
rect 828 -1170 834 -1164
rect 828 -1176 834 -1170
rect 828 -1182 834 -1176
rect 828 -1188 834 -1182
rect 828 -1194 834 -1188
rect 828 -1200 834 -1194
rect 828 -1206 834 -1200
rect 828 -1212 834 -1206
rect 828 -1218 834 -1212
rect 828 -1224 834 -1218
rect 828 -1230 834 -1224
rect 828 -1236 834 -1230
rect 828 -1242 834 -1236
rect 828 -1248 834 -1242
rect 828 -1254 834 -1248
rect 828 -1260 834 -1254
rect 828 -1266 834 -1260
rect 828 -1272 834 -1266
rect 828 -1278 834 -1272
rect 828 -1284 834 -1278
rect 828 -1290 834 -1284
rect 828 -1296 834 -1290
rect 828 -1302 834 -1296
rect 828 -1308 834 -1302
rect 828 -1314 834 -1308
rect 828 -1320 834 -1314
rect 828 -1326 834 -1320
rect 828 -1332 834 -1326
rect 828 -1338 834 -1332
rect 828 -1344 834 -1338
rect 828 -1350 834 -1344
rect 828 -1356 834 -1350
rect 828 -1362 834 -1356
rect 828 -1368 834 -1362
rect 828 -1374 834 -1368
rect 828 -1380 834 -1374
rect 828 -3078 834 -3072
rect 828 -3084 834 -3078
rect 828 -3090 834 -3084
rect 828 -3096 834 -3090
rect 828 -3102 834 -3096
rect 828 -3108 834 -3102
rect 828 -3114 834 -3108
rect 828 -3120 834 -3114
rect 828 -3126 834 -3120
rect 828 -3132 834 -3126
rect 828 -3138 834 -3132
rect 828 -3144 834 -3138
rect 828 -3150 834 -3144
rect 828 -3156 834 -3150
rect 828 -3162 834 -3156
rect 828 -3168 834 -3162
rect 828 -3174 834 -3168
rect 828 -3180 834 -3174
rect 828 -3186 834 -3180
rect 828 -3192 834 -3186
rect 828 -3198 834 -3192
rect 828 -3204 834 -3198
rect 828 -3210 834 -3204
rect 828 -3216 834 -3210
rect 828 -3222 834 -3216
rect 828 -3228 834 -3222
rect 828 -3234 834 -3228
rect 828 -3240 834 -3234
rect 828 -3246 834 -3240
rect 828 -3252 834 -3246
rect 828 -3258 834 -3252
rect 828 -3264 834 -3258
rect 828 -3270 834 -3264
rect 828 -3276 834 -3270
rect 828 -3444 834 -3438
rect 828 -3450 834 -3444
rect 834 -1164 840 -1158
rect 834 -1170 840 -1164
rect 834 -1176 840 -1170
rect 834 -1182 840 -1176
rect 834 -1188 840 -1182
rect 834 -1194 840 -1188
rect 834 -1200 840 -1194
rect 834 -1206 840 -1200
rect 834 -1212 840 -1206
rect 834 -1218 840 -1212
rect 834 -1224 840 -1218
rect 834 -1230 840 -1224
rect 834 -1236 840 -1230
rect 834 -1242 840 -1236
rect 834 -1248 840 -1242
rect 834 -1254 840 -1248
rect 834 -1260 840 -1254
rect 834 -1266 840 -1260
rect 834 -1272 840 -1266
rect 834 -1278 840 -1272
rect 834 -1284 840 -1278
rect 834 -1290 840 -1284
rect 834 -1296 840 -1290
rect 834 -1302 840 -1296
rect 834 -1308 840 -1302
rect 834 -1314 840 -1308
rect 834 -1320 840 -1314
rect 834 -1326 840 -1320
rect 834 -1332 840 -1326
rect 834 -1338 840 -1332
rect 834 -1344 840 -1338
rect 834 -1350 840 -1344
rect 834 -1356 840 -1350
rect 834 -1362 840 -1356
rect 834 -1368 840 -1362
rect 834 -1374 840 -1368
rect 834 -1380 840 -1374
rect 834 -3048 840 -3042
rect 834 -3054 840 -3048
rect 834 -3060 840 -3054
rect 834 -3066 840 -3060
rect 834 -3072 840 -3066
rect 834 -3078 840 -3072
rect 834 -3084 840 -3078
rect 834 -3090 840 -3084
rect 834 -3096 840 -3090
rect 834 -3102 840 -3096
rect 834 -3108 840 -3102
rect 834 -3114 840 -3108
rect 834 -3120 840 -3114
rect 834 -3126 840 -3120
rect 834 -3132 840 -3126
rect 834 -3138 840 -3132
rect 834 -3144 840 -3138
rect 834 -3150 840 -3144
rect 834 -3156 840 -3150
rect 834 -3162 840 -3156
rect 834 -3168 840 -3162
rect 834 -3174 840 -3168
rect 834 -3180 840 -3174
rect 834 -3186 840 -3180
rect 834 -3192 840 -3186
rect 834 -3198 840 -3192
rect 834 -3204 840 -3198
rect 834 -3210 840 -3204
rect 834 -3216 840 -3210
rect 834 -3222 840 -3216
rect 834 -3228 840 -3222
rect 834 -3234 840 -3228
rect 834 -3240 840 -3234
rect 834 -3246 840 -3240
rect 834 -3252 840 -3246
rect 834 -3258 840 -3252
rect 834 -3264 840 -3258
rect 834 -3432 840 -3426
rect 834 -3438 840 -3432
rect 834 -3444 840 -3438
rect 834 -3450 840 -3444
rect 840 -1164 846 -1158
rect 840 -1170 846 -1164
rect 840 -1176 846 -1170
rect 840 -1182 846 -1176
rect 840 -1188 846 -1182
rect 840 -1194 846 -1188
rect 840 -1200 846 -1194
rect 840 -1206 846 -1200
rect 840 -1212 846 -1206
rect 840 -1218 846 -1212
rect 840 -1224 846 -1218
rect 840 -1230 846 -1224
rect 840 -1236 846 -1230
rect 840 -1242 846 -1236
rect 840 -1248 846 -1242
rect 840 -1254 846 -1248
rect 840 -1260 846 -1254
rect 840 -1266 846 -1260
rect 840 -1272 846 -1266
rect 840 -1278 846 -1272
rect 840 -1284 846 -1278
rect 840 -1290 846 -1284
rect 840 -1296 846 -1290
rect 840 -1302 846 -1296
rect 840 -1308 846 -1302
rect 840 -1314 846 -1308
rect 840 -1320 846 -1314
rect 840 -1326 846 -1320
rect 840 -1332 846 -1326
rect 840 -1338 846 -1332
rect 840 -1344 846 -1338
rect 840 -1350 846 -1344
rect 840 -1356 846 -1350
rect 840 -1362 846 -1356
rect 840 -1368 846 -1362
rect 840 -1374 846 -1368
rect 840 -1380 846 -1374
rect 840 -3018 846 -3012
rect 840 -3024 846 -3018
rect 840 -3030 846 -3024
rect 840 -3036 846 -3030
rect 840 -3042 846 -3036
rect 840 -3048 846 -3042
rect 840 -3054 846 -3048
rect 840 -3060 846 -3054
rect 840 -3066 846 -3060
rect 840 -3072 846 -3066
rect 840 -3078 846 -3072
rect 840 -3084 846 -3078
rect 840 -3090 846 -3084
rect 840 -3096 846 -3090
rect 840 -3102 846 -3096
rect 840 -3108 846 -3102
rect 840 -3114 846 -3108
rect 840 -3120 846 -3114
rect 840 -3126 846 -3120
rect 840 -3132 846 -3126
rect 840 -3138 846 -3132
rect 840 -3144 846 -3138
rect 840 -3150 846 -3144
rect 840 -3156 846 -3150
rect 840 -3162 846 -3156
rect 840 -3168 846 -3162
rect 840 -3174 846 -3168
rect 840 -3180 846 -3174
rect 840 -3186 846 -3180
rect 840 -3192 846 -3186
rect 840 -3198 846 -3192
rect 840 -3204 846 -3198
rect 840 -3210 846 -3204
rect 840 -3216 846 -3210
rect 840 -3222 846 -3216
rect 840 -3228 846 -3222
rect 840 -3234 846 -3228
rect 840 -3240 846 -3234
rect 840 -3246 846 -3240
rect 840 -3252 846 -3246
rect 840 -3420 846 -3414
rect 840 -3426 846 -3420
rect 840 -3432 846 -3426
rect 840 -3438 846 -3432
rect 840 -3444 846 -3438
rect 846 -1158 852 -1152
rect 846 -1164 852 -1158
rect 846 -1170 852 -1164
rect 846 -1176 852 -1170
rect 846 -1182 852 -1176
rect 846 -1188 852 -1182
rect 846 -1194 852 -1188
rect 846 -1200 852 -1194
rect 846 -1206 852 -1200
rect 846 -1212 852 -1206
rect 846 -1218 852 -1212
rect 846 -1224 852 -1218
rect 846 -1230 852 -1224
rect 846 -1236 852 -1230
rect 846 -1242 852 -1236
rect 846 -1248 852 -1242
rect 846 -1254 852 -1248
rect 846 -1260 852 -1254
rect 846 -1266 852 -1260
rect 846 -1272 852 -1266
rect 846 -1278 852 -1272
rect 846 -1284 852 -1278
rect 846 -1290 852 -1284
rect 846 -1296 852 -1290
rect 846 -1302 852 -1296
rect 846 -1308 852 -1302
rect 846 -1314 852 -1308
rect 846 -1320 852 -1314
rect 846 -1326 852 -1320
rect 846 -1332 852 -1326
rect 846 -1338 852 -1332
rect 846 -1344 852 -1338
rect 846 -1350 852 -1344
rect 846 -1356 852 -1350
rect 846 -1362 852 -1356
rect 846 -1368 852 -1362
rect 846 -1374 852 -1368
rect 846 -2994 852 -2988
rect 846 -3000 852 -2994
rect 846 -3006 852 -3000
rect 846 -3012 852 -3006
rect 846 -3018 852 -3012
rect 846 -3024 852 -3018
rect 846 -3030 852 -3024
rect 846 -3036 852 -3030
rect 846 -3042 852 -3036
rect 846 -3048 852 -3042
rect 846 -3054 852 -3048
rect 846 -3060 852 -3054
rect 846 -3066 852 -3060
rect 846 -3072 852 -3066
rect 846 -3078 852 -3072
rect 846 -3084 852 -3078
rect 846 -3090 852 -3084
rect 846 -3096 852 -3090
rect 846 -3102 852 -3096
rect 846 -3108 852 -3102
rect 846 -3114 852 -3108
rect 846 -3120 852 -3114
rect 846 -3126 852 -3120
rect 846 -3132 852 -3126
rect 846 -3138 852 -3132
rect 846 -3144 852 -3138
rect 846 -3150 852 -3144
rect 846 -3156 852 -3150
rect 846 -3162 852 -3156
rect 846 -3168 852 -3162
rect 846 -3174 852 -3168
rect 846 -3180 852 -3174
rect 846 -3186 852 -3180
rect 846 -3192 852 -3186
rect 846 -3198 852 -3192
rect 846 -3204 852 -3198
rect 846 -3210 852 -3204
rect 846 -3216 852 -3210
rect 846 -3222 852 -3216
rect 846 -3228 852 -3222
rect 846 -3234 852 -3228
rect 846 -3240 852 -3234
rect 846 -3408 852 -3402
rect 846 -3414 852 -3408
rect 846 -3420 852 -3414
rect 846 -3426 852 -3420
rect 846 -3432 852 -3426
rect 846 -3438 852 -3432
rect 852 -1158 858 -1152
rect 852 -1164 858 -1158
rect 852 -1170 858 -1164
rect 852 -1176 858 -1170
rect 852 -1182 858 -1176
rect 852 -1188 858 -1182
rect 852 -1194 858 -1188
rect 852 -1200 858 -1194
rect 852 -1206 858 -1200
rect 852 -1212 858 -1206
rect 852 -1218 858 -1212
rect 852 -1224 858 -1218
rect 852 -1230 858 -1224
rect 852 -1236 858 -1230
rect 852 -1242 858 -1236
rect 852 -1248 858 -1242
rect 852 -1254 858 -1248
rect 852 -1260 858 -1254
rect 852 -1266 858 -1260
rect 852 -1272 858 -1266
rect 852 -1278 858 -1272
rect 852 -1284 858 -1278
rect 852 -1290 858 -1284
rect 852 -1296 858 -1290
rect 852 -1302 858 -1296
rect 852 -1308 858 -1302
rect 852 -1314 858 -1308
rect 852 -1320 858 -1314
rect 852 -1326 858 -1320
rect 852 -1332 858 -1326
rect 852 -1338 858 -1332
rect 852 -1344 858 -1338
rect 852 -1350 858 -1344
rect 852 -1356 858 -1350
rect 852 -1362 858 -1356
rect 852 -1368 858 -1362
rect 852 -1374 858 -1368
rect 852 -2964 858 -2958
rect 852 -2970 858 -2964
rect 852 -2976 858 -2970
rect 852 -2982 858 -2976
rect 852 -2988 858 -2982
rect 852 -2994 858 -2988
rect 852 -3000 858 -2994
rect 852 -3006 858 -3000
rect 852 -3012 858 -3006
rect 852 -3018 858 -3012
rect 852 -3024 858 -3018
rect 852 -3030 858 -3024
rect 852 -3036 858 -3030
rect 852 -3042 858 -3036
rect 852 -3048 858 -3042
rect 852 -3054 858 -3048
rect 852 -3060 858 -3054
rect 852 -3066 858 -3060
rect 852 -3072 858 -3066
rect 852 -3078 858 -3072
rect 852 -3084 858 -3078
rect 852 -3090 858 -3084
rect 852 -3096 858 -3090
rect 852 -3102 858 -3096
rect 852 -3108 858 -3102
rect 852 -3114 858 -3108
rect 852 -3120 858 -3114
rect 852 -3126 858 -3120
rect 852 -3132 858 -3126
rect 852 -3138 858 -3132
rect 852 -3144 858 -3138
rect 852 -3150 858 -3144
rect 852 -3156 858 -3150
rect 852 -3162 858 -3156
rect 852 -3168 858 -3162
rect 852 -3174 858 -3168
rect 852 -3180 858 -3174
rect 852 -3186 858 -3180
rect 852 -3192 858 -3186
rect 852 -3198 858 -3192
rect 852 -3204 858 -3198
rect 852 -3210 858 -3204
rect 852 -3216 858 -3210
rect 852 -3222 858 -3216
rect 852 -3228 858 -3222
rect 852 -3396 858 -3390
rect 852 -3402 858 -3396
rect 852 -3408 858 -3402
rect 852 -3414 858 -3408
rect 852 -3420 858 -3414
rect 852 -3426 858 -3420
rect 852 -3432 858 -3426
rect 852 -3438 858 -3432
rect 858 -1158 864 -1152
rect 858 -1164 864 -1158
rect 858 -1170 864 -1164
rect 858 -1176 864 -1170
rect 858 -1182 864 -1176
rect 858 -1188 864 -1182
rect 858 -1194 864 -1188
rect 858 -1200 864 -1194
rect 858 -1206 864 -1200
rect 858 -1212 864 -1206
rect 858 -1218 864 -1212
rect 858 -1224 864 -1218
rect 858 -1230 864 -1224
rect 858 -1236 864 -1230
rect 858 -1242 864 -1236
rect 858 -1248 864 -1242
rect 858 -1254 864 -1248
rect 858 -1260 864 -1254
rect 858 -1266 864 -1260
rect 858 -1272 864 -1266
rect 858 -1278 864 -1272
rect 858 -1284 864 -1278
rect 858 -1290 864 -1284
rect 858 -1296 864 -1290
rect 858 -1302 864 -1296
rect 858 -1308 864 -1302
rect 858 -1314 864 -1308
rect 858 -1320 864 -1314
rect 858 -1326 864 -1320
rect 858 -1332 864 -1326
rect 858 -1338 864 -1332
rect 858 -1344 864 -1338
rect 858 -1350 864 -1344
rect 858 -1356 864 -1350
rect 858 -1362 864 -1356
rect 858 -1368 864 -1362
rect 858 -2940 864 -2934
rect 858 -2946 864 -2940
rect 858 -2952 864 -2946
rect 858 -2958 864 -2952
rect 858 -2964 864 -2958
rect 858 -2970 864 -2964
rect 858 -2976 864 -2970
rect 858 -2982 864 -2976
rect 858 -2988 864 -2982
rect 858 -2994 864 -2988
rect 858 -3000 864 -2994
rect 858 -3006 864 -3000
rect 858 -3012 864 -3006
rect 858 -3018 864 -3012
rect 858 -3024 864 -3018
rect 858 -3030 864 -3024
rect 858 -3036 864 -3030
rect 858 -3042 864 -3036
rect 858 -3048 864 -3042
rect 858 -3054 864 -3048
rect 858 -3060 864 -3054
rect 858 -3066 864 -3060
rect 858 -3072 864 -3066
rect 858 -3078 864 -3072
rect 858 -3084 864 -3078
rect 858 -3090 864 -3084
rect 858 -3096 864 -3090
rect 858 -3102 864 -3096
rect 858 -3108 864 -3102
rect 858 -3114 864 -3108
rect 858 -3120 864 -3114
rect 858 -3126 864 -3120
rect 858 -3132 864 -3126
rect 858 -3138 864 -3132
rect 858 -3144 864 -3138
rect 858 -3150 864 -3144
rect 858 -3156 864 -3150
rect 858 -3162 864 -3156
rect 858 -3168 864 -3162
rect 858 -3174 864 -3168
rect 858 -3180 864 -3174
rect 858 -3186 864 -3180
rect 858 -3192 864 -3186
rect 858 -3198 864 -3192
rect 858 -3204 864 -3198
rect 858 -3210 864 -3204
rect 858 -3216 864 -3210
rect 858 -3384 864 -3378
rect 858 -3390 864 -3384
rect 858 -3396 864 -3390
rect 858 -3402 864 -3396
rect 858 -3408 864 -3402
rect 858 -3414 864 -3408
rect 858 -3420 864 -3414
rect 858 -3426 864 -3420
rect 858 -3432 864 -3426
rect 864 -1152 870 -1146
rect 864 -1158 870 -1152
rect 864 -1164 870 -1158
rect 864 -1170 870 -1164
rect 864 -1176 870 -1170
rect 864 -1182 870 -1176
rect 864 -1188 870 -1182
rect 864 -1194 870 -1188
rect 864 -1200 870 -1194
rect 864 -1206 870 -1200
rect 864 -1212 870 -1206
rect 864 -1218 870 -1212
rect 864 -1224 870 -1218
rect 864 -1230 870 -1224
rect 864 -1236 870 -1230
rect 864 -1242 870 -1236
rect 864 -1248 870 -1242
rect 864 -1254 870 -1248
rect 864 -1260 870 -1254
rect 864 -1266 870 -1260
rect 864 -1272 870 -1266
rect 864 -1278 870 -1272
rect 864 -1284 870 -1278
rect 864 -1290 870 -1284
rect 864 -1296 870 -1290
rect 864 -1302 870 -1296
rect 864 -1308 870 -1302
rect 864 -1314 870 -1308
rect 864 -1320 870 -1314
rect 864 -1326 870 -1320
rect 864 -1332 870 -1326
rect 864 -1338 870 -1332
rect 864 -1344 870 -1338
rect 864 -1350 870 -1344
rect 864 -1356 870 -1350
rect 864 -1362 870 -1356
rect 864 -1368 870 -1362
rect 864 -2910 870 -2904
rect 864 -2916 870 -2910
rect 864 -2922 870 -2916
rect 864 -2928 870 -2922
rect 864 -2934 870 -2928
rect 864 -2940 870 -2934
rect 864 -2946 870 -2940
rect 864 -2952 870 -2946
rect 864 -2958 870 -2952
rect 864 -2964 870 -2958
rect 864 -2970 870 -2964
rect 864 -2976 870 -2970
rect 864 -2982 870 -2976
rect 864 -2988 870 -2982
rect 864 -2994 870 -2988
rect 864 -3000 870 -2994
rect 864 -3006 870 -3000
rect 864 -3012 870 -3006
rect 864 -3018 870 -3012
rect 864 -3024 870 -3018
rect 864 -3030 870 -3024
rect 864 -3036 870 -3030
rect 864 -3042 870 -3036
rect 864 -3048 870 -3042
rect 864 -3054 870 -3048
rect 864 -3060 870 -3054
rect 864 -3066 870 -3060
rect 864 -3072 870 -3066
rect 864 -3078 870 -3072
rect 864 -3084 870 -3078
rect 864 -3090 870 -3084
rect 864 -3096 870 -3090
rect 864 -3102 870 -3096
rect 864 -3108 870 -3102
rect 864 -3114 870 -3108
rect 864 -3120 870 -3114
rect 864 -3126 870 -3120
rect 864 -3132 870 -3126
rect 864 -3138 870 -3132
rect 864 -3144 870 -3138
rect 864 -3150 870 -3144
rect 864 -3156 870 -3150
rect 864 -3162 870 -3156
rect 864 -3168 870 -3162
rect 864 -3174 870 -3168
rect 864 -3180 870 -3174
rect 864 -3186 870 -3180
rect 864 -3192 870 -3186
rect 864 -3198 870 -3192
rect 864 -3204 870 -3198
rect 864 -3378 870 -3372
rect 864 -3384 870 -3378
rect 864 -3390 870 -3384
rect 864 -3396 870 -3390
rect 864 -3402 870 -3396
rect 864 -3408 870 -3402
rect 864 -3414 870 -3408
rect 864 -3420 870 -3414
rect 864 -3426 870 -3420
rect 864 -3432 870 -3426
rect 870 -1152 876 -1146
rect 870 -1158 876 -1152
rect 870 -1164 876 -1158
rect 870 -1170 876 -1164
rect 870 -1176 876 -1170
rect 870 -1182 876 -1176
rect 870 -1188 876 -1182
rect 870 -1194 876 -1188
rect 870 -1200 876 -1194
rect 870 -1206 876 -1200
rect 870 -1212 876 -1206
rect 870 -1218 876 -1212
rect 870 -1224 876 -1218
rect 870 -1230 876 -1224
rect 870 -1236 876 -1230
rect 870 -1242 876 -1236
rect 870 -1248 876 -1242
rect 870 -1254 876 -1248
rect 870 -1260 876 -1254
rect 870 -1266 876 -1260
rect 870 -1272 876 -1266
rect 870 -1278 876 -1272
rect 870 -1284 876 -1278
rect 870 -1290 876 -1284
rect 870 -1296 876 -1290
rect 870 -1302 876 -1296
rect 870 -1308 876 -1302
rect 870 -1314 876 -1308
rect 870 -1320 876 -1314
rect 870 -1326 876 -1320
rect 870 -1332 876 -1326
rect 870 -1338 876 -1332
rect 870 -1344 876 -1338
rect 870 -1350 876 -1344
rect 870 -1356 876 -1350
rect 870 -1362 876 -1356
rect 870 -1368 876 -1362
rect 870 -2886 876 -2880
rect 870 -2892 876 -2886
rect 870 -2898 876 -2892
rect 870 -2904 876 -2898
rect 870 -2910 876 -2904
rect 870 -2916 876 -2910
rect 870 -2922 876 -2916
rect 870 -2928 876 -2922
rect 870 -2934 876 -2928
rect 870 -2940 876 -2934
rect 870 -2946 876 -2940
rect 870 -2952 876 -2946
rect 870 -2958 876 -2952
rect 870 -2964 876 -2958
rect 870 -2970 876 -2964
rect 870 -2976 876 -2970
rect 870 -2982 876 -2976
rect 870 -2988 876 -2982
rect 870 -2994 876 -2988
rect 870 -3000 876 -2994
rect 870 -3006 876 -3000
rect 870 -3012 876 -3006
rect 870 -3018 876 -3012
rect 870 -3024 876 -3018
rect 870 -3030 876 -3024
rect 870 -3036 876 -3030
rect 870 -3042 876 -3036
rect 870 -3048 876 -3042
rect 870 -3054 876 -3048
rect 870 -3060 876 -3054
rect 870 -3066 876 -3060
rect 870 -3072 876 -3066
rect 870 -3078 876 -3072
rect 870 -3084 876 -3078
rect 870 -3090 876 -3084
rect 870 -3096 876 -3090
rect 870 -3102 876 -3096
rect 870 -3108 876 -3102
rect 870 -3114 876 -3108
rect 870 -3120 876 -3114
rect 870 -3126 876 -3120
rect 870 -3132 876 -3126
rect 870 -3138 876 -3132
rect 870 -3144 876 -3138
rect 870 -3150 876 -3144
rect 870 -3156 876 -3150
rect 870 -3162 876 -3156
rect 870 -3168 876 -3162
rect 870 -3174 876 -3168
rect 870 -3180 876 -3174
rect 870 -3186 876 -3180
rect 870 -3192 876 -3186
rect 870 -3366 876 -3360
rect 870 -3372 876 -3366
rect 870 -3378 876 -3372
rect 870 -3384 876 -3378
rect 870 -3390 876 -3384
rect 870 -3396 876 -3390
rect 870 -3402 876 -3396
rect 870 -3408 876 -3402
rect 870 -3414 876 -3408
rect 870 -3420 876 -3414
rect 870 -3426 876 -3420
rect 876 -1152 882 -1146
rect 876 -1158 882 -1152
rect 876 -1164 882 -1158
rect 876 -1170 882 -1164
rect 876 -1176 882 -1170
rect 876 -1182 882 -1176
rect 876 -1188 882 -1182
rect 876 -1194 882 -1188
rect 876 -1200 882 -1194
rect 876 -1206 882 -1200
rect 876 -1212 882 -1206
rect 876 -1218 882 -1212
rect 876 -1224 882 -1218
rect 876 -1230 882 -1224
rect 876 -1236 882 -1230
rect 876 -1242 882 -1236
rect 876 -1248 882 -1242
rect 876 -1254 882 -1248
rect 876 -1260 882 -1254
rect 876 -1266 882 -1260
rect 876 -1272 882 -1266
rect 876 -1278 882 -1272
rect 876 -1284 882 -1278
rect 876 -1290 882 -1284
rect 876 -1296 882 -1290
rect 876 -1302 882 -1296
rect 876 -1308 882 -1302
rect 876 -1314 882 -1308
rect 876 -1320 882 -1314
rect 876 -1326 882 -1320
rect 876 -1332 882 -1326
rect 876 -1338 882 -1332
rect 876 -1344 882 -1338
rect 876 -1350 882 -1344
rect 876 -1356 882 -1350
rect 876 -1362 882 -1356
rect 876 -2862 882 -2856
rect 876 -2868 882 -2862
rect 876 -2874 882 -2868
rect 876 -2880 882 -2874
rect 876 -2886 882 -2880
rect 876 -2892 882 -2886
rect 876 -2898 882 -2892
rect 876 -2904 882 -2898
rect 876 -2910 882 -2904
rect 876 -2916 882 -2910
rect 876 -2922 882 -2916
rect 876 -2928 882 -2922
rect 876 -2934 882 -2928
rect 876 -2940 882 -2934
rect 876 -2946 882 -2940
rect 876 -2952 882 -2946
rect 876 -2958 882 -2952
rect 876 -2964 882 -2958
rect 876 -2970 882 -2964
rect 876 -2976 882 -2970
rect 876 -2982 882 -2976
rect 876 -2988 882 -2982
rect 876 -2994 882 -2988
rect 876 -3000 882 -2994
rect 876 -3006 882 -3000
rect 876 -3012 882 -3006
rect 876 -3018 882 -3012
rect 876 -3024 882 -3018
rect 876 -3030 882 -3024
rect 876 -3036 882 -3030
rect 876 -3042 882 -3036
rect 876 -3048 882 -3042
rect 876 -3054 882 -3048
rect 876 -3060 882 -3054
rect 876 -3066 882 -3060
rect 876 -3072 882 -3066
rect 876 -3078 882 -3072
rect 876 -3084 882 -3078
rect 876 -3090 882 -3084
rect 876 -3096 882 -3090
rect 876 -3102 882 -3096
rect 876 -3108 882 -3102
rect 876 -3114 882 -3108
rect 876 -3120 882 -3114
rect 876 -3126 882 -3120
rect 876 -3132 882 -3126
rect 876 -3138 882 -3132
rect 876 -3144 882 -3138
rect 876 -3150 882 -3144
rect 876 -3156 882 -3150
rect 876 -3162 882 -3156
rect 876 -3168 882 -3162
rect 876 -3174 882 -3168
rect 876 -3180 882 -3174
rect 876 -3360 882 -3354
rect 876 -3366 882 -3360
rect 876 -3372 882 -3366
rect 876 -3378 882 -3372
rect 876 -3384 882 -3378
rect 876 -3390 882 -3384
rect 876 -3396 882 -3390
rect 876 -3402 882 -3396
rect 876 -3408 882 -3402
rect 876 -3414 882 -3408
rect 876 -3420 882 -3414
rect 882 -1152 888 -1146
rect 882 -1158 888 -1152
rect 882 -1164 888 -1158
rect 882 -1170 888 -1164
rect 882 -1176 888 -1170
rect 882 -1182 888 -1176
rect 882 -1188 888 -1182
rect 882 -1194 888 -1188
rect 882 -1200 888 -1194
rect 882 -1206 888 -1200
rect 882 -1212 888 -1206
rect 882 -1218 888 -1212
rect 882 -1224 888 -1218
rect 882 -1230 888 -1224
rect 882 -1236 888 -1230
rect 882 -1242 888 -1236
rect 882 -1248 888 -1242
rect 882 -1254 888 -1248
rect 882 -1260 888 -1254
rect 882 -1266 888 -1260
rect 882 -1272 888 -1266
rect 882 -1278 888 -1272
rect 882 -1284 888 -1278
rect 882 -1290 888 -1284
rect 882 -1296 888 -1290
rect 882 -1302 888 -1296
rect 882 -1308 888 -1302
rect 882 -1314 888 -1308
rect 882 -1320 888 -1314
rect 882 -1326 888 -1320
rect 882 -1332 888 -1326
rect 882 -1338 888 -1332
rect 882 -1344 888 -1338
rect 882 -1350 888 -1344
rect 882 -1356 888 -1350
rect 882 -1362 888 -1356
rect 882 -2838 888 -2832
rect 882 -2844 888 -2838
rect 882 -2850 888 -2844
rect 882 -2856 888 -2850
rect 882 -2862 888 -2856
rect 882 -2868 888 -2862
rect 882 -2874 888 -2868
rect 882 -2880 888 -2874
rect 882 -2886 888 -2880
rect 882 -2892 888 -2886
rect 882 -2898 888 -2892
rect 882 -2904 888 -2898
rect 882 -2910 888 -2904
rect 882 -2916 888 -2910
rect 882 -2922 888 -2916
rect 882 -2928 888 -2922
rect 882 -2934 888 -2928
rect 882 -2940 888 -2934
rect 882 -2946 888 -2940
rect 882 -2952 888 -2946
rect 882 -2958 888 -2952
rect 882 -2964 888 -2958
rect 882 -2970 888 -2964
rect 882 -2976 888 -2970
rect 882 -2982 888 -2976
rect 882 -2988 888 -2982
rect 882 -2994 888 -2988
rect 882 -3000 888 -2994
rect 882 -3006 888 -3000
rect 882 -3012 888 -3006
rect 882 -3018 888 -3012
rect 882 -3024 888 -3018
rect 882 -3030 888 -3024
rect 882 -3036 888 -3030
rect 882 -3042 888 -3036
rect 882 -3048 888 -3042
rect 882 -3054 888 -3048
rect 882 -3060 888 -3054
rect 882 -3066 888 -3060
rect 882 -3072 888 -3066
rect 882 -3078 888 -3072
rect 882 -3084 888 -3078
rect 882 -3090 888 -3084
rect 882 -3096 888 -3090
rect 882 -3102 888 -3096
rect 882 -3108 888 -3102
rect 882 -3114 888 -3108
rect 882 -3120 888 -3114
rect 882 -3126 888 -3120
rect 882 -3132 888 -3126
rect 882 -3138 888 -3132
rect 882 -3144 888 -3138
rect 882 -3150 888 -3144
rect 882 -3156 888 -3150
rect 882 -3162 888 -3156
rect 882 -3168 888 -3162
rect 882 -3348 888 -3342
rect 882 -3354 888 -3348
rect 882 -3360 888 -3354
rect 882 -3366 888 -3360
rect 882 -3372 888 -3366
rect 882 -3378 888 -3372
rect 882 -3384 888 -3378
rect 882 -3390 888 -3384
rect 882 -3396 888 -3390
rect 882 -3402 888 -3396
rect 882 -3408 888 -3402
rect 882 -3414 888 -3408
rect 882 -3420 888 -3414
rect 888 -1146 894 -1140
rect 888 -1152 894 -1146
rect 888 -1158 894 -1152
rect 888 -1164 894 -1158
rect 888 -1170 894 -1164
rect 888 -1176 894 -1170
rect 888 -1182 894 -1176
rect 888 -1188 894 -1182
rect 888 -1194 894 -1188
rect 888 -1200 894 -1194
rect 888 -1206 894 -1200
rect 888 -1212 894 -1206
rect 888 -1218 894 -1212
rect 888 -1224 894 -1218
rect 888 -1230 894 -1224
rect 888 -1236 894 -1230
rect 888 -1242 894 -1236
rect 888 -1248 894 -1242
rect 888 -1254 894 -1248
rect 888 -1260 894 -1254
rect 888 -1266 894 -1260
rect 888 -1272 894 -1266
rect 888 -1278 894 -1272
rect 888 -1284 894 -1278
rect 888 -1290 894 -1284
rect 888 -1296 894 -1290
rect 888 -1302 894 -1296
rect 888 -1308 894 -1302
rect 888 -1314 894 -1308
rect 888 -1320 894 -1314
rect 888 -1326 894 -1320
rect 888 -1332 894 -1326
rect 888 -1338 894 -1332
rect 888 -1344 894 -1338
rect 888 -1350 894 -1344
rect 888 -1356 894 -1350
rect 888 -1362 894 -1356
rect 888 -2814 894 -2808
rect 888 -2820 894 -2814
rect 888 -2826 894 -2820
rect 888 -2832 894 -2826
rect 888 -2838 894 -2832
rect 888 -2844 894 -2838
rect 888 -2850 894 -2844
rect 888 -2856 894 -2850
rect 888 -2862 894 -2856
rect 888 -2868 894 -2862
rect 888 -2874 894 -2868
rect 888 -2880 894 -2874
rect 888 -2886 894 -2880
rect 888 -2892 894 -2886
rect 888 -2898 894 -2892
rect 888 -2904 894 -2898
rect 888 -2910 894 -2904
rect 888 -2916 894 -2910
rect 888 -2922 894 -2916
rect 888 -2928 894 -2922
rect 888 -2934 894 -2928
rect 888 -2940 894 -2934
rect 888 -2946 894 -2940
rect 888 -2952 894 -2946
rect 888 -2958 894 -2952
rect 888 -2964 894 -2958
rect 888 -2970 894 -2964
rect 888 -2976 894 -2970
rect 888 -2982 894 -2976
rect 888 -2988 894 -2982
rect 888 -2994 894 -2988
rect 888 -3000 894 -2994
rect 888 -3006 894 -3000
rect 888 -3012 894 -3006
rect 888 -3018 894 -3012
rect 888 -3024 894 -3018
rect 888 -3030 894 -3024
rect 888 -3036 894 -3030
rect 888 -3042 894 -3036
rect 888 -3048 894 -3042
rect 888 -3054 894 -3048
rect 888 -3060 894 -3054
rect 888 -3066 894 -3060
rect 888 -3072 894 -3066
rect 888 -3078 894 -3072
rect 888 -3084 894 -3078
rect 888 -3090 894 -3084
rect 888 -3096 894 -3090
rect 888 -3102 894 -3096
rect 888 -3108 894 -3102
rect 888 -3114 894 -3108
rect 888 -3120 894 -3114
rect 888 -3126 894 -3120
rect 888 -3132 894 -3126
rect 888 -3138 894 -3132
rect 888 -3144 894 -3138
rect 888 -3150 894 -3144
rect 888 -3156 894 -3150
rect 888 -3342 894 -3336
rect 888 -3348 894 -3342
rect 888 -3354 894 -3348
rect 888 -3360 894 -3354
rect 888 -3366 894 -3360
rect 888 -3372 894 -3366
rect 888 -3378 894 -3372
rect 888 -3384 894 -3378
rect 888 -3390 894 -3384
rect 888 -3396 894 -3390
rect 888 -3402 894 -3396
rect 888 -3408 894 -3402
rect 888 -3414 894 -3408
rect 894 -1146 900 -1140
rect 894 -1152 900 -1146
rect 894 -1158 900 -1152
rect 894 -1164 900 -1158
rect 894 -1170 900 -1164
rect 894 -1176 900 -1170
rect 894 -1182 900 -1176
rect 894 -1188 900 -1182
rect 894 -1194 900 -1188
rect 894 -1200 900 -1194
rect 894 -1206 900 -1200
rect 894 -1212 900 -1206
rect 894 -1218 900 -1212
rect 894 -1224 900 -1218
rect 894 -1230 900 -1224
rect 894 -1236 900 -1230
rect 894 -1242 900 -1236
rect 894 -1248 900 -1242
rect 894 -1254 900 -1248
rect 894 -1260 900 -1254
rect 894 -1266 900 -1260
rect 894 -1272 900 -1266
rect 894 -1278 900 -1272
rect 894 -1284 900 -1278
rect 894 -1290 900 -1284
rect 894 -1296 900 -1290
rect 894 -1302 900 -1296
rect 894 -1308 900 -1302
rect 894 -1314 900 -1308
rect 894 -1320 900 -1314
rect 894 -1326 900 -1320
rect 894 -1332 900 -1326
rect 894 -1338 900 -1332
rect 894 -1344 900 -1338
rect 894 -1350 900 -1344
rect 894 -1356 900 -1350
rect 894 -2790 900 -2784
rect 894 -2796 900 -2790
rect 894 -2802 900 -2796
rect 894 -2808 900 -2802
rect 894 -2814 900 -2808
rect 894 -2820 900 -2814
rect 894 -2826 900 -2820
rect 894 -2832 900 -2826
rect 894 -2838 900 -2832
rect 894 -2844 900 -2838
rect 894 -2850 900 -2844
rect 894 -2856 900 -2850
rect 894 -2862 900 -2856
rect 894 -2868 900 -2862
rect 894 -2874 900 -2868
rect 894 -2880 900 -2874
rect 894 -2886 900 -2880
rect 894 -2892 900 -2886
rect 894 -2898 900 -2892
rect 894 -2904 900 -2898
rect 894 -2910 900 -2904
rect 894 -2916 900 -2910
rect 894 -2922 900 -2916
rect 894 -2928 900 -2922
rect 894 -2934 900 -2928
rect 894 -2940 900 -2934
rect 894 -2946 900 -2940
rect 894 -2952 900 -2946
rect 894 -2958 900 -2952
rect 894 -2964 900 -2958
rect 894 -2970 900 -2964
rect 894 -2976 900 -2970
rect 894 -2982 900 -2976
rect 894 -2988 900 -2982
rect 894 -2994 900 -2988
rect 894 -3000 900 -2994
rect 894 -3006 900 -3000
rect 894 -3012 900 -3006
rect 894 -3018 900 -3012
rect 894 -3024 900 -3018
rect 894 -3030 900 -3024
rect 894 -3036 900 -3030
rect 894 -3042 900 -3036
rect 894 -3048 900 -3042
rect 894 -3054 900 -3048
rect 894 -3060 900 -3054
rect 894 -3066 900 -3060
rect 894 -3072 900 -3066
rect 894 -3078 900 -3072
rect 894 -3084 900 -3078
rect 894 -3090 900 -3084
rect 894 -3096 900 -3090
rect 894 -3102 900 -3096
rect 894 -3108 900 -3102
rect 894 -3114 900 -3108
rect 894 -3120 900 -3114
rect 894 -3126 900 -3120
rect 894 -3132 900 -3126
rect 894 -3138 900 -3132
rect 894 -3144 900 -3138
rect 894 -3336 900 -3330
rect 894 -3342 900 -3336
rect 894 -3348 900 -3342
rect 894 -3354 900 -3348
rect 894 -3360 900 -3354
rect 894 -3366 900 -3360
rect 894 -3372 900 -3366
rect 894 -3378 900 -3372
rect 894 -3384 900 -3378
rect 894 -3390 900 -3384
rect 894 -3396 900 -3390
rect 894 -3402 900 -3396
rect 894 -3408 900 -3402
rect 894 -3480 900 -3474
rect 900 -1146 906 -1140
rect 900 -1152 906 -1146
rect 900 -1158 906 -1152
rect 900 -1164 906 -1158
rect 900 -1170 906 -1164
rect 900 -1176 906 -1170
rect 900 -1182 906 -1176
rect 900 -1188 906 -1182
rect 900 -1194 906 -1188
rect 900 -1200 906 -1194
rect 900 -1206 906 -1200
rect 900 -1212 906 -1206
rect 900 -1218 906 -1212
rect 900 -1224 906 -1218
rect 900 -1230 906 -1224
rect 900 -1236 906 -1230
rect 900 -1242 906 -1236
rect 900 -1248 906 -1242
rect 900 -1254 906 -1248
rect 900 -1260 906 -1254
rect 900 -1266 906 -1260
rect 900 -1272 906 -1266
rect 900 -1278 906 -1272
rect 900 -1284 906 -1278
rect 900 -1290 906 -1284
rect 900 -1296 906 -1290
rect 900 -1302 906 -1296
rect 900 -1308 906 -1302
rect 900 -1314 906 -1308
rect 900 -1320 906 -1314
rect 900 -1326 906 -1320
rect 900 -1332 906 -1326
rect 900 -1338 906 -1332
rect 900 -1344 906 -1338
rect 900 -1350 906 -1344
rect 900 -1356 906 -1350
rect 900 -2766 906 -2760
rect 900 -2772 906 -2766
rect 900 -2778 906 -2772
rect 900 -2784 906 -2778
rect 900 -2790 906 -2784
rect 900 -2796 906 -2790
rect 900 -2802 906 -2796
rect 900 -2808 906 -2802
rect 900 -2814 906 -2808
rect 900 -2820 906 -2814
rect 900 -2826 906 -2820
rect 900 -2832 906 -2826
rect 900 -2838 906 -2832
rect 900 -2844 906 -2838
rect 900 -2850 906 -2844
rect 900 -2856 906 -2850
rect 900 -2862 906 -2856
rect 900 -2868 906 -2862
rect 900 -2874 906 -2868
rect 900 -2880 906 -2874
rect 900 -2886 906 -2880
rect 900 -2892 906 -2886
rect 900 -2898 906 -2892
rect 900 -2904 906 -2898
rect 900 -2910 906 -2904
rect 900 -2916 906 -2910
rect 900 -2922 906 -2916
rect 900 -2928 906 -2922
rect 900 -2934 906 -2928
rect 900 -2940 906 -2934
rect 900 -2946 906 -2940
rect 900 -2952 906 -2946
rect 900 -2958 906 -2952
rect 900 -2964 906 -2958
rect 900 -2970 906 -2964
rect 900 -2976 906 -2970
rect 900 -2982 906 -2976
rect 900 -2988 906 -2982
rect 900 -2994 906 -2988
rect 900 -3000 906 -2994
rect 900 -3006 906 -3000
rect 900 -3012 906 -3006
rect 900 -3018 906 -3012
rect 900 -3024 906 -3018
rect 900 -3030 906 -3024
rect 900 -3036 906 -3030
rect 900 -3042 906 -3036
rect 900 -3048 906 -3042
rect 900 -3054 906 -3048
rect 900 -3060 906 -3054
rect 900 -3066 906 -3060
rect 900 -3072 906 -3066
rect 900 -3078 906 -3072
rect 900 -3084 906 -3078
rect 900 -3090 906 -3084
rect 900 -3096 906 -3090
rect 900 -3102 906 -3096
rect 900 -3108 906 -3102
rect 900 -3114 906 -3108
rect 900 -3120 906 -3114
rect 900 -3126 906 -3120
rect 900 -3132 906 -3126
rect 900 -3330 906 -3324
rect 900 -3336 906 -3330
rect 900 -3342 906 -3336
rect 900 -3348 906 -3342
rect 900 -3354 906 -3348
rect 900 -3360 906 -3354
rect 900 -3366 906 -3360
rect 900 -3372 906 -3366
rect 900 -3378 906 -3372
rect 900 -3384 906 -3378
rect 900 -3390 906 -3384
rect 900 -3396 906 -3390
rect 900 -3402 906 -3396
rect 900 -3408 906 -3402
rect 900 -3474 906 -3468
rect 900 -3480 906 -3474
rect 906 -1140 912 -1134
rect 906 -1146 912 -1140
rect 906 -1152 912 -1146
rect 906 -1158 912 -1152
rect 906 -1164 912 -1158
rect 906 -1170 912 -1164
rect 906 -1176 912 -1170
rect 906 -1182 912 -1176
rect 906 -1188 912 -1182
rect 906 -1194 912 -1188
rect 906 -1200 912 -1194
rect 906 -1206 912 -1200
rect 906 -1212 912 -1206
rect 906 -1218 912 -1212
rect 906 -1224 912 -1218
rect 906 -1230 912 -1224
rect 906 -1236 912 -1230
rect 906 -1242 912 -1236
rect 906 -1248 912 -1242
rect 906 -1254 912 -1248
rect 906 -1260 912 -1254
rect 906 -1266 912 -1260
rect 906 -1272 912 -1266
rect 906 -1278 912 -1272
rect 906 -1284 912 -1278
rect 906 -1290 912 -1284
rect 906 -1296 912 -1290
rect 906 -1302 912 -1296
rect 906 -1308 912 -1302
rect 906 -1314 912 -1308
rect 906 -1320 912 -1314
rect 906 -1326 912 -1320
rect 906 -1332 912 -1326
rect 906 -1338 912 -1332
rect 906 -1344 912 -1338
rect 906 -1350 912 -1344
rect 906 -1356 912 -1350
rect 906 -2748 912 -2742
rect 906 -2754 912 -2748
rect 906 -2760 912 -2754
rect 906 -2766 912 -2760
rect 906 -2772 912 -2766
rect 906 -2778 912 -2772
rect 906 -2784 912 -2778
rect 906 -2790 912 -2784
rect 906 -2796 912 -2790
rect 906 -2802 912 -2796
rect 906 -2808 912 -2802
rect 906 -2814 912 -2808
rect 906 -2820 912 -2814
rect 906 -2826 912 -2820
rect 906 -2832 912 -2826
rect 906 -2838 912 -2832
rect 906 -2844 912 -2838
rect 906 -2850 912 -2844
rect 906 -2856 912 -2850
rect 906 -2862 912 -2856
rect 906 -2868 912 -2862
rect 906 -2874 912 -2868
rect 906 -2880 912 -2874
rect 906 -2886 912 -2880
rect 906 -2892 912 -2886
rect 906 -2898 912 -2892
rect 906 -2904 912 -2898
rect 906 -2910 912 -2904
rect 906 -2916 912 -2910
rect 906 -2922 912 -2916
rect 906 -2928 912 -2922
rect 906 -2934 912 -2928
rect 906 -2940 912 -2934
rect 906 -2946 912 -2940
rect 906 -2952 912 -2946
rect 906 -2958 912 -2952
rect 906 -2964 912 -2958
rect 906 -2970 912 -2964
rect 906 -2976 912 -2970
rect 906 -2982 912 -2976
rect 906 -2988 912 -2982
rect 906 -2994 912 -2988
rect 906 -3000 912 -2994
rect 906 -3006 912 -3000
rect 906 -3012 912 -3006
rect 906 -3018 912 -3012
rect 906 -3024 912 -3018
rect 906 -3030 912 -3024
rect 906 -3036 912 -3030
rect 906 -3042 912 -3036
rect 906 -3048 912 -3042
rect 906 -3054 912 -3048
rect 906 -3060 912 -3054
rect 906 -3066 912 -3060
rect 906 -3072 912 -3066
rect 906 -3078 912 -3072
rect 906 -3084 912 -3078
rect 906 -3090 912 -3084
rect 906 -3096 912 -3090
rect 906 -3102 912 -3096
rect 906 -3108 912 -3102
rect 906 -3114 912 -3108
rect 906 -3120 912 -3114
rect 906 -3324 912 -3318
rect 906 -3330 912 -3324
rect 906 -3336 912 -3330
rect 906 -3342 912 -3336
rect 906 -3348 912 -3342
rect 906 -3354 912 -3348
rect 906 -3360 912 -3354
rect 906 -3366 912 -3360
rect 906 -3372 912 -3366
rect 906 -3378 912 -3372
rect 906 -3384 912 -3378
rect 906 -3390 912 -3384
rect 906 -3396 912 -3390
rect 906 -3402 912 -3396
rect 906 -3468 912 -3462
rect 906 -3474 912 -3468
rect 906 -3480 912 -3474
rect 912 -1140 918 -1134
rect 912 -1146 918 -1140
rect 912 -1152 918 -1146
rect 912 -1158 918 -1152
rect 912 -1164 918 -1158
rect 912 -1170 918 -1164
rect 912 -1176 918 -1170
rect 912 -1182 918 -1176
rect 912 -1188 918 -1182
rect 912 -1194 918 -1188
rect 912 -1200 918 -1194
rect 912 -1206 918 -1200
rect 912 -1212 918 -1206
rect 912 -1218 918 -1212
rect 912 -1224 918 -1218
rect 912 -1230 918 -1224
rect 912 -1236 918 -1230
rect 912 -1242 918 -1236
rect 912 -1248 918 -1242
rect 912 -1254 918 -1248
rect 912 -1260 918 -1254
rect 912 -1266 918 -1260
rect 912 -1272 918 -1266
rect 912 -1278 918 -1272
rect 912 -1284 918 -1278
rect 912 -1290 918 -1284
rect 912 -1296 918 -1290
rect 912 -1302 918 -1296
rect 912 -1308 918 -1302
rect 912 -1314 918 -1308
rect 912 -1320 918 -1314
rect 912 -1326 918 -1320
rect 912 -1332 918 -1326
rect 912 -1338 918 -1332
rect 912 -1344 918 -1338
rect 912 -1350 918 -1344
rect 912 -2724 918 -2718
rect 912 -2730 918 -2724
rect 912 -2736 918 -2730
rect 912 -2742 918 -2736
rect 912 -2748 918 -2742
rect 912 -2754 918 -2748
rect 912 -2760 918 -2754
rect 912 -2766 918 -2760
rect 912 -2772 918 -2766
rect 912 -2778 918 -2772
rect 912 -2784 918 -2778
rect 912 -2790 918 -2784
rect 912 -2796 918 -2790
rect 912 -2802 918 -2796
rect 912 -2808 918 -2802
rect 912 -2814 918 -2808
rect 912 -2820 918 -2814
rect 912 -2826 918 -2820
rect 912 -2832 918 -2826
rect 912 -2838 918 -2832
rect 912 -2844 918 -2838
rect 912 -2850 918 -2844
rect 912 -2856 918 -2850
rect 912 -2862 918 -2856
rect 912 -2868 918 -2862
rect 912 -2874 918 -2868
rect 912 -2880 918 -2874
rect 912 -2886 918 -2880
rect 912 -2892 918 -2886
rect 912 -2898 918 -2892
rect 912 -2904 918 -2898
rect 912 -2910 918 -2904
rect 912 -2916 918 -2910
rect 912 -2922 918 -2916
rect 912 -2928 918 -2922
rect 912 -2934 918 -2928
rect 912 -2940 918 -2934
rect 912 -2946 918 -2940
rect 912 -2952 918 -2946
rect 912 -2958 918 -2952
rect 912 -2964 918 -2958
rect 912 -2970 918 -2964
rect 912 -2976 918 -2970
rect 912 -2982 918 -2976
rect 912 -2988 918 -2982
rect 912 -2994 918 -2988
rect 912 -3000 918 -2994
rect 912 -3006 918 -3000
rect 912 -3012 918 -3006
rect 912 -3018 918 -3012
rect 912 -3024 918 -3018
rect 912 -3030 918 -3024
rect 912 -3036 918 -3030
rect 912 -3042 918 -3036
rect 912 -3048 918 -3042
rect 912 -3054 918 -3048
rect 912 -3060 918 -3054
rect 912 -3066 918 -3060
rect 912 -3072 918 -3066
rect 912 -3078 918 -3072
rect 912 -3084 918 -3078
rect 912 -3090 918 -3084
rect 912 -3096 918 -3090
rect 912 -3102 918 -3096
rect 912 -3108 918 -3102
rect 912 -3240 918 -3234
rect 912 -3318 918 -3312
rect 912 -3324 918 -3318
rect 912 -3330 918 -3324
rect 912 -3336 918 -3330
rect 912 -3342 918 -3336
rect 912 -3348 918 -3342
rect 912 -3354 918 -3348
rect 912 -3360 918 -3354
rect 912 -3366 918 -3360
rect 912 -3372 918 -3366
rect 912 -3378 918 -3372
rect 912 -3384 918 -3378
rect 912 -3390 918 -3384
rect 912 -3396 918 -3390
rect 912 -3468 918 -3462
rect 912 -3474 918 -3468
rect 912 -3480 918 -3474
rect 918 -1140 924 -1134
rect 918 -1146 924 -1140
rect 918 -1152 924 -1146
rect 918 -1158 924 -1152
rect 918 -1164 924 -1158
rect 918 -1170 924 -1164
rect 918 -1176 924 -1170
rect 918 -1182 924 -1176
rect 918 -1188 924 -1182
rect 918 -1194 924 -1188
rect 918 -1200 924 -1194
rect 918 -1206 924 -1200
rect 918 -1212 924 -1206
rect 918 -1218 924 -1212
rect 918 -1224 924 -1218
rect 918 -1230 924 -1224
rect 918 -1236 924 -1230
rect 918 -1242 924 -1236
rect 918 -1248 924 -1242
rect 918 -1254 924 -1248
rect 918 -1260 924 -1254
rect 918 -1266 924 -1260
rect 918 -1272 924 -1266
rect 918 -1278 924 -1272
rect 918 -1284 924 -1278
rect 918 -1290 924 -1284
rect 918 -1296 924 -1290
rect 918 -1302 924 -1296
rect 918 -1308 924 -1302
rect 918 -1314 924 -1308
rect 918 -1320 924 -1314
rect 918 -1326 924 -1320
rect 918 -1332 924 -1326
rect 918 -1338 924 -1332
rect 918 -1344 924 -1338
rect 918 -1350 924 -1344
rect 918 -2700 924 -2694
rect 918 -2706 924 -2700
rect 918 -2712 924 -2706
rect 918 -2718 924 -2712
rect 918 -2724 924 -2718
rect 918 -2730 924 -2724
rect 918 -2736 924 -2730
rect 918 -2742 924 -2736
rect 918 -2748 924 -2742
rect 918 -2754 924 -2748
rect 918 -2760 924 -2754
rect 918 -2766 924 -2760
rect 918 -2772 924 -2766
rect 918 -2778 924 -2772
rect 918 -2784 924 -2778
rect 918 -2790 924 -2784
rect 918 -2796 924 -2790
rect 918 -2802 924 -2796
rect 918 -2808 924 -2802
rect 918 -2814 924 -2808
rect 918 -2820 924 -2814
rect 918 -2826 924 -2820
rect 918 -2832 924 -2826
rect 918 -2838 924 -2832
rect 918 -2844 924 -2838
rect 918 -2850 924 -2844
rect 918 -2856 924 -2850
rect 918 -2862 924 -2856
rect 918 -2868 924 -2862
rect 918 -2874 924 -2868
rect 918 -2880 924 -2874
rect 918 -2886 924 -2880
rect 918 -2892 924 -2886
rect 918 -2898 924 -2892
rect 918 -2904 924 -2898
rect 918 -2910 924 -2904
rect 918 -2916 924 -2910
rect 918 -2922 924 -2916
rect 918 -2928 924 -2922
rect 918 -2934 924 -2928
rect 918 -2940 924 -2934
rect 918 -2946 924 -2940
rect 918 -2952 924 -2946
rect 918 -2958 924 -2952
rect 918 -2964 924 -2958
rect 918 -2970 924 -2964
rect 918 -2976 924 -2970
rect 918 -2982 924 -2976
rect 918 -2988 924 -2982
rect 918 -2994 924 -2988
rect 918 -3000 924 -2994
rect 918 -3006 924 -3000
rect 918 -3012 924 -3006
rect 918 -3018 924 -3012
rect 918 -3024 924 -3018
rect 918 -3030 924 -3024
rect 918 -3036 924 -3030
rect 918 -3042 924 -3036
rect 918 -3048 924 -3042
rect 918 -3054 924 -3048
rect 918 -3060 924 -3054
rect 918 -3066 924 -3060
rect 918 -3072 924 -3066
rect 918 -3078 924 -3072
rect 918 -3084 924 -3078
rect 918 -3090 924 -3084
rect 918 -3096 924 -3090
rect 918 -3228 924 -3222
rect 918 -3234 924 -3228
rect 918 -3240 924 -3234
rect 918 -3312 924 -3306
rect 918 -3318 924 -3312
rect 918 -3324 924 -3318
rect 918 -3330 924 -3324
rect 918 -3336 924 -3330
rect 918 -3342 924 -3336
rect 918 -3348 924 -3342
rect 918 -3354 924 -3348
rect 918 -3360 924 -3354
rect 918 -3366 924 -3360
rect 918 -3372 924 -3366
rect 918 -3378 924 -3372
rect 918 -3384 924 -3378
rect 918 -3390 924 -3384
rect 918 -3396 924 -3390
rect 918 -3462 924 -3456
rect 918 -3468 924 -3462
rect 918 -3474 924 -3468
rect 918 -3480 924 -3474
rect 918 -3486 924 -3480
rect 924 -1140 930 -1134
rect 924 -1146 930 -1140
rect 924 -1152 930 -1146
rect 924 -1158 930 -1152
rect 924 -1164 930 -1158
rect 924 -1170 930 -1164
rect 924 -1176 930 -1170
rect 924 -1182 930 -1176
rect 924 -1188 930 -1182
rect 924 -1194 930 -1188
rect 924 -1200 930 -1194
rect 924 -1206 930 -1200
rect 924 -1212 930 -1206
rect 924 -1218 930 -1212
rect 924 -1224 930 -1218
rect 924 -1230 930 -1224
rect 924 -1236 930 -1230
rect 924 -1242 930 -1236
rect 924 -1248 930 -1242
rect 924 -1254 930 -1248
rect 924 -1260 930 -1254
rect 924 -1266 930 -1260
rect 924 -1272 930 -1266
rect 924 -1278 930 -1272
rect 924 -1284 930 -1278
rect 924 -1290 930 -1284
rect 924 -1296 930 -1290
rect 924 -1302 930 -1296
rect 924 -1308 930 -1302
rect 924 -1314 930 -1308
rect 924 -1320 930 -1314
rect 924 -1326 930 -1320
rect 924 -1332 930 -1326
rect 924 -1338 930 -1332
rect 924 -1344 930 -1338
rect 924 -1350 930 -1344
rect 924 -2676 930 -2670
rect 924 -2682 930 -2676
rect 924 -2688 930 -2682
rect 924 -2694 930 -2688
rect 924 -2700 930 -2694
rect 924 -2706 930 -2700
rect 924 -2712 930 -2706
rect 924 -2718 930 -2712
rect 924 -2724 930 -2718
rect 924 -2730 930 -2724
rect 924 -2736 930 -2730
rect 924 -2742 930 -2736
rect 924 -2748 930 -2742
rect 924 -2754 930 -2748
rect 924 -2760 930 -2754
rect 924 -2766 930 -2760
rect 924 -2772 930 -2766
rect 924 -2778 930 -2772
rect 924 -2784 930 -2778
rect 924 -2790 930 -2784
rect 924 -2796 930 -2790
rect 924 -2802 930 -2796
rect 924 -2808 930 -2802
rect 924 -2814 930 -2808
rect 924 -2820 930 -2814
rect 924 -2826 930 -2820
rect 924 -2832 930 -2826
rect 924 -2838 930 -2832
rect 924 -2844 930 -2838
rect 924 -2850 930 -2844
rect 924 -2856 930 -2850
rect 924 -2862 930 -2856
rect 924 -2868 930 -2862
rect 924 -2874 930 -2868
rect 924 -2880 930 -2874
rect 924 -2886 930 -2880
rect 924 -2892 930 -2886
rect 924 -2898 930 -2892
rect 924 -2904 930 -2898
rect 924 -2910 930 -2904
rect 924 -2916 930 -2910
rect 924 -2922 930 -2916
rect 924 -2928 930 -2922
rect 924 -2934 930 -2928
rect 924 -2940 930 -2934
rect 924 -2946 930 -2940
rect 924 -2952 930 -2946
rect 924 -2958 930 -2952
rect 924 -2964 930 -2958
rect 924 -2970 930 -2964
rect 924 -2976 930 -2970
rect 924 -2982 930 -2976
rect 924 -2988 930 -2982
rect 924 -2994 930 -2988
rect 924 -3000 930 -2994
rect 924 -3006 930 -3000
rect 924 -3012 930 -3006
rect 924 -3018 930 -3012
rect 924 -3024 930 -3018
rect 924 -3030 930 -3024
rect 924 -3036 930 -3030
rect 924 -3042 930 -3036
rect 924 -3048 930 -3042
rect 924 -3054 930 -3048
rect 924 -3060 930 -3054
rect 924 -3066 930 -3060
rect 924 -3072 930 -3066
rect 924 -3078 930 -3072
rect 924 -3084 930 -3078
rect 924 -3210 930 -3204
rect 924 -3216 930 -3210
rect 924 -3222 930 -3216
rect 924 -3228 930 -3222
rect 924 -3234 930 -3228
rect 924 -3306 930 -3300
rect 924 -3312 930 -3306
rect 924 -3318 930 -3312
rect 924 -3324 930 -3318
rect 924 -3330 930 -3324
rect 924 -3336 930 -3330
rect 924 -3342 930 -3336
rect 924 -3348 930 -3342
rect 924 -3354 930 -3348
rect 924 -3360 930 -3354
rect 924 -3366 930 -3360
rect 924 -3372 930 -3366
rect 924 -3378 930 -3372
rect 924 -3384 930 -3378
rect 924 -3390 930 -3384
rect 924 -3456 930 -3450
rect 924 -3462 930 -3456
rect 924 -3468 930 -3462
rect 924 -3474 930 -3468
rect 924 -3480 930 -3474
rect 924 -3486 930 -3480
rect 930 -1134 936 -1128
rect 930 -1140 936 -1134
rect 930 -1146 936 -1140
rect 930 -1152 936 -1146
rect 930 -1158 936 -1152
rect 930 -1164 936 -1158
rect 930 -1170 936 -1164
rect 930 -1176 936 -1170
rect 930 -1182 936 -1176
rect 930 -1188 936 -1182
rect 930 -1194 936 -1188
rect 930 -1200 936 -1194
rect 930 -1206 936 -1200
rect 930 -1212 936 -1206
rect 930 -1218 936 -1212
rect 930 -1224 936 -1218
rect 930 -1230 936 -1224
rect 930 -1236 936 -1230
rect 930 -1242 936 -1236
rect 930 -1248 936 -1242
rect 930 -1254 936 -1248
rect 930 -1260 936 -1254
rect 930 -1266 936 -1260
rect 930 -1272 936 -1266
rect 930 -1278 936 -1272
rect 930 -1284 936 -1278
rect 930 -1290 936 -1284
rect 930 -1296 936 -1290
rect 930 -1302 936 -1296
rect 930 -1308 936 -1302
rect 930 -1314 936 -1308
rect 930 -1320 936 -1314
rect 930 -1326 936 -1320
rect 930 -1332 936 -1326
rect 930 -1338 936 -1332
rect 930 -1344 936 -1338
rect 930 -2658 936 -2652
rect 930 -2664 936 -2658
rect 930 -2670 936 -2664
rect 930 -2676 936 -2670
rect 930 -2682 936 -2676
rect 930 -2688 936 -2682
rect 930 -2694 936 -2688
rect 930 -2700 936 -2694
rect 930 -2706 936 -2700
rect 930 -2712 936 -2706
rect 930 -2718 936 -2712
rect 930 -2724 936 -2718
rect 930 -2730 936 -2724
rect 930 -2736 936 -2730
rect 930 -2742 936 -2736
rect 930 -2748 936 -2742
rect 930 -2754 936 -2748
rect 930 -2760 936 -2754
rect 930 -2766 936 -2760
rect 930 -2772 936 -2766
rect 930 -2778 936 -2772
rect 930 -2784 936 -2778
rect 930 -2790 936 -2784
rect 930 -2796 936 -2790
rect 930 -2802 936 -2796
rect 930 -2808 936 -2802
rect 930 -2814 936 -2808
rect 930 -2820 936 -2814
rect 930 -2826 936 -2820
rect 930 -2832 936 -2826
rect 930 -2838 936 -2832
rect 930 -2844 936 -2838
rect 930 -2850 936 -2844
rect 930 -2856 936 -2850
rect 930 -2862 936 -2856
rect 930 -2868 936 -2862
rect 930 -2874 936 -2868
rect 930 -2880 936 -2874
rect 930 -2886 936 -2880
rect 930 -2892 936 -2886
rect 930 -2898 936 -2892
rect 930 -2904 936 -2898
rect 930 -2910 936 -2904
rect 930 -2916 936 -2910
rect 930 -2922 936 -2916
rect 930 -2928 936 -2922
rect 930 -2934 936 -2928
rect 930 -2940 936 -2934
rect 930 -2946 936 -2940
rect 930 -2952 936 -2946
rect 930 -2958 936 -2952
rect 930 -2964 936 -2958
rect 930 -2970 936 -2964
rect 930 -2976 936 -2970
rect 930 -2982 936 -2976
rect 930 -2988 936 -2982
rect 930 -2994 936 -2988
rect 930 -3000 936 -2994
rect 930 -3006 936 -3000
rect 930 -3012 936 -3006
rect 930 -3018 936 -3012
rect 930 -3024 936 -3018
rect 930 -3030 936 -3024
rect 930 -3036 936 -3030
rect 930 -3042 936 -3036
rect 930 -3048 936 -3042
rect 930 -3054 936 -3048
rect 930 -3060 936 -3054
rect 930 -3066 936 -3060
rect 930 -3072 936 -3066
rect 930 -3192 936 -3186
rect 930 -3198 936 -3192
rect 930 -3204 936 -3198
rect 930 -3210 936 -3204
rect 930 -3216 936 -3210
rect 930 -3222 936 -3216
rect 930 -3228 936 -3222
rect 930 -3300 936 -3294
rect 930 -3306 936 -3300
rect 930 -3312 936 -3306
rect 930 -3318 936 -3312
rect 930 -3324 936 -3318
rect 930 -3330 936 -3324
rect 930 -3336 936 -3330
rect 930 -3342 936 -3336
rect 930 -3348 936 -3342
rect 930 -3354 936 -3348
rect 930 -3360 936 -3354
rect 930 -3366 936 -3360
rect 930 -3372 936 -3366
rect 930 -3378 936 -3372
rect 930 -3384 936 -3378
rect 930 -3450 936 -3444
rect 930 -3456 936 -3450
rect 930 -3462 936 -3456
rect 930 -3468 936 -3462
rect 930 -3474 936 -3468
rect 930 -3480 936 -3474
rect 930 -3486 936 -3480
rect 936 -1134 942 -1128
rect 936 -1140 942 -1134
rect 936 -1146 942 -1140
rect 936 -1152 942 -1146
rect 936 -1158 942 -1152
rect 936 -1164 942 -1158
rect 936 -1170 942 -1164
rect 936 -1176 942 -1170
rect 936 -1182 942 -1176
rect 936 -1188 942 -1182
rect 936 -1194 942 -1188
rect 936 -1200 942 -1194
rect 936 -1206 942 -1200
rect 936 -1212 942 -1206
rect 936 -1218 942 -1212
rect 936 -1224 942 -1218
rect 936 -1230 942 -1224
rect 936 -1236 942 -1230
rect 936 -1242 942 -1236
rect 936 -1248 942 -1242
rect 936 -1254 942 -1248
rect 936 -1260 942 -1254
rect 936 -1266 942 -1260
rect 936 -1272 942 -1266
rect 936 -1278 942 -1272
rect 936 -1284 942 -1278
rect 936 -1290 942 -1284
rect 936 -1296 942 -1290
rect 936 -1302 942 -1296
rect 936 -1308 942 -1302
rect 936 -1314 942 -1308
rect 936 -1320 942 -1314
rect 936 -1326 942 -1320
rect 936 -1332 942 -1326
rect 936 -1338 942 -1332
rect 936 -1344 942 -1338
rect 936 -2634 942 -2628
rect 936 -2640 942 -2634
rect 936 -2646 942 -2640
rect 936 -2652 942 -2646
rect 936 -2658 942 -2652
rect 936 -2664 942 -2658
rect 936 -2670 942 -2664
rect 936 -2676 942 -2670
rect 936 -2682 942 -2676
rect 936 -2688 942 -2682
rect 936 -2694 942 -2688
rect 936 -2700 942 -2694
rect 936 -2706 942 -2700
rect 936 -2712 942 -2706
rect 936 -2718 942 -2712
rect 936 -2724 942 -2718
rect 936 -2730 942 -2724
rect 936 -2736 942 -2730
rect 936 -2742 942 -2736
rect 936 -2748 942 -2742
rect 936 -2754 942 -2748
rect 936 -2760 942 -2754
rect 936 -2766 942 -2760
rect 936 -2772 942 -2766
rect 936 -2778 942 -2772
rect 936 -2784 942 -2778
rect 936 -2790 942 -2784
rect 936 -2796 942 -2790
rect 936 -2802 942 -2796
rect 936 -2808 942 -2802
rect 936 -2814 942 -2808
rect 936 -2820 942 -2814
rect 936 -2826 942 -2820
rect 936 -2832 942 -2826
rect 936 -2838 942 -2832
rect 936 -2844 942 -2838
rect 936 -2850 942 -2844
rect 936 -2856 942 -2850
rect 936 -2862 942 -2856
rect 936 -2868 942 -2862
rect 936 -2874 942 -2868
rect 936 -2880 942 -2874
rect 936 -2886 942 -2880
rect 936 -2892 942 -2886
rect 936 -2898 942 -2892
rect 936 -2904 942 -2898
rect 936 -2910 942 -2904
rect 936 -2916 942 -2910
rect 936 -2922 942 -2916
rect 936 -2928 942 -2922
rect 936 -2934 942 -2928
rect 936 -2940 942 -2934
rect 936 -2946 942 -2940
rect 936 -2952 942 -2946
rect 936 -2958 942 -2952
rect 936 -2964 942 -2958
rect 936 -2970 942 -2964
rect 936 -2976 942 -2970
rect 936 -2982 942 -2976
rect 936 -2988 942 -2982
rect 936 -2994 942 -2988
rect 936 -3000 942 -2994
rect 936 -3006 942 -3000
rect 936 -3012 942 -3006
rect 936 -3018 942 -3012
rect 936 -3024 942 -3018
rect 936 -3030 942 -3024
rect 936 -3036 942 -3030
rect 936 -3042 942 -3036
rect 936 -3048 942 -3042
rect 936 -3054 942 -3048
rect 936 -3060 942 -3054
rect 936 -3180 942 -3174
rect 936 -3186 942 -3180
rect 936 -3192 942 -3186
rect 936 -3198 942 -3192
rect 936 -3204 942 -3198
rect 936 -3210 942 -3204
rect 936 -3216 942 -3210
rect 936 -3222 942 -3216
rect 936 -3294 942 -3288
rect 936 -3300 942 -3294
rect 936 -3306 942 -3300
rect 936 -3312 942 -3306
rect 936 -3318 942 -3312
rect 936 -3324 942 -3318
rect 936 -3330 942 -3324
rect 936 -3336 942 -3330
rect 936 -3342 942 -3336
rect 936 -3348 942 -3342
rect 936 -3354 942 -3348
rect 936 -3360 942 -3354
rect 936 -3366 942 -3360
rect 936 -3372 942 -3366
rect 936 -3378 942 -3372
rect 936 -3444 942 -3438
rect 936 -3450 942 -3444
rect 936 -3456 942 -3450
rect 936 -3462 942 -3456
rect 936 -3468 942 -3462
rect 936 -3474 942 -3468
rect 936 -3480 942 -3474
rect 936 -3486 942 -3480
rect 942 -1134 948 -1128
rect 942 -1140 948 -1134
rect 942 -1146 948 -1140
rect 942 -1152 948 -1146
rect 942 -1158 948 -1152
rect 942 -1164 948 -1158
rect 942 -1170 948 -1164
rect 942 -1176 948 -1170
rect 942 -1182 948 -1176
rect 942 -1188 948 -1182
rect 942 -1194 948 -1188
rect 942 -1200 948 -1194
rect 942 -1206 948 -1200
rect 942 -1212 948 -1206
rect 942 -1218 948 -1212
rect 942 -1224 948 -1218
rect 942 -1230 948 -1224
rect 942 -1236 948 -1230
rect 942 -1242 948 -1236
rect 942 -1248 948 -1242
rect 942 -1254 948 -1248
rect 942 -1260 948 -1254
rect 942 -1266 948 -1260
rect 942 -1272 948 -1266
rect 942 -1278 948 -1272
rect 942 -1284 948 -1278
rect 942 -1290 948 -1284
rect 942 -1296 948 -1290
rect 942 -1302 948 -1296
rect 942 -1308 948 -1302
rect 942 -1314 948 -1308
rect 942 -1320 948 -1314
rect 942 -1326 948 -1320
rect 942 -1332 948 -1326
rect 942 -1338 948 -1332
rect 942 -1344 948 -1338
rect 942 -2616 948 -2610
rect 942 -2622 948 -2616
rect 942 -2628 948 -2622
rect 942 -2634 948 -2628
rect 942 -2640 948 -2634
rect 942 -2646 948 -2640
rect 942 -2652 948 -2646
rect 942 -2658 948 -2652
rect 942 -2664 948 -2658
rect 942 -2670 948 -2664
rect 942 -2676 948 -2670
rect 942 -2682 948 -2676
rect 942 -2688 948 -2682
rect 942 -2694 948 -2688
rect 942 -2700 948 -2694
rect 942 -2706 948 -2700
rect 942 -2712 948 -2706
rect 942 -2718 948 -2712
rect 942 -2724 948 -2718
rect 942 -2730 948 -2724
rect 942 -2736 948 -2730
rect 942 -2742 948 -2736
rect 942 -2748 948 -2742
rect 942 -2754 948 -2748
rect 942 -2760 948 -2754
rect 942 -2766 948 -2760
rect 942 -2772 948 -2766
rect 942 -2778 948 -2772
rect 942 -2784 948 -2778
rect 942 -2790 948 -2784
rect 942 -2796 948 -2790
rect 942 -2802 948 -2796
rect 942 -2808 948 -2802
rect 942 -2814 948 -2808
rect 942 -2820 948 -2814
rect 942 -2826 948 -2820
rect 942 -2832 948 -2826
rect 942 -2838 948 -2832
rect 942 -2844 948 -2838
rect 942 -2850 948 -2844
rect 942 -2856 948 -2850
rect 942 -2862 948 -2856
rect 942 -2868 948 -2862
rect 942 -2874 948 -2868
rect 942 -2880 948 -2874
rect 942 -2886 948 -2880
rect 942 -2892 948 -2886
rect 942 -2898 948 -2892
rect 942 -2904 948 -2898
rect 942 -2910 948 -2904
rect 942 -2916 948 -2910
rect 942 -2922 948 -2916
rect 942 -2928 948 -2922
rect 942 -2934 948 -2928
rect 942 -2940 948 -2934
rect 942 -2946 948 -2940
rect 942 -2952 948 -2946
rect 942 -2958 948 -2952
rect 942 -2964 948 -2958
rect 942 -2970 948 -2964
rect 942 -2976 948 -2970
rect 942 -2982 948 -2976
rect 942 -2988 948 -2982
rect 942 -2994 948 -2988
rect 942 -3000 948 -2994
rect 942 -3006 948 -3000
rect 942 -3012 948 -3006
rect 942 -3018 948 -3012
rect 942 -3024 948 -3018
rect 942 -3030 948 -3024
rect 942 -3036 948 -3030
rect 942 -3042 948 -3036
rect 942 -3048 948 -3042
rect 942 -3162 948 -3156
rect 942 -3168 948 -3162
rect 942 -3174 948 -3168
rect 942 -3180 948 -3174
rect 942 -3186 948 -3180
rect 942 -3192 948 -3186
rect 942 -3198 948 -3192
rect 942 -3204 948 -3198
rect 942 -3210 948 -3204
rect 942 -3216 948 -3210
rect 942 -3222 948 -3216
rect 942 -3288 948 -3282
rect 942 -3294 948 -3288
rect 942 -3300 948 -3294
rect 942 -3306 948 -3300
rect 942 -3312 948 -3306
rect 942 -3318 948 -3312
rect 942 -3324 948 -3318
rect 942 -3330 948 -3324
rect 942 -3336 948 -3330
rect 942 -3342 948 -3336
rect 942 -3348 948 -3342
rect 942 -3354 948 -3348
rect 942 -3360 948 -3354
rect 942 -3366 948 -3360
rect 942 -3372 948 -3366
rect 942 -3378 948 -3372
rect 942 -3444 948 -3438
rect 942 -3450 948 -3444
rect 942 -3456 948 -3450
rect 942 -3462 948 -3456
rect 942 -3468 948 -3462
rect 942 -3474 948 -3468
rect 942 -3480 948 -3474
rect 942 -3486 948 -3480
rect 948 -1134 954 -1128
rect 948 -1140 954 -1134
rect 948 -1146 954 -1140
rect 948 -1152 954 -1146
rect 948 -1158 954 -1152
rect 948 -1164 954 -1158
rect 948 -1170 954 -1164
rect 948 -1176 954 -1170
rect 948 -1182 954 -1176
rect 948 -1188 954 -1182
rect 948 -1194 954 -1188
rect 948 -1200 954 -1194
rect 948 -1206 954 -1200
rect 948 -1212 954 -1206
rect 948 -1218 954 -1212
rect 948 -1224 954 -1218
rect 948 -1230 954 -1224
rect 948 -1236 954 -1230
rect 948 -1242 954 -1236
rect 948 -1248 954 -1242
rect 948 -1254 954 -1248
rect 948 -1260 954 -1254
rect 948 -1266 954 -1260
rect 948 -1272 954 -1266
rect 948 -1278 954 -1272
rect 948 -1284 954 -1278
rect 948 -1290 954 -1284
rect 948 -1296 954 -1290
rect 948 -1302 954 -1296
rect 948 -1308 954 -1302
rect 948 -1314 954 -1308
rect 948 -1320 954 -1314
rect 948 -1326 954 -1320
rect 948 -1332 954 -1326
rect 948 -1338 954 -1332
rect 948 -1344 954 -1338
rect 948 -2592 954 -2586
rect 948 -2598 954 -2592
rect 948 -2604 954 -2598
rect 948 -2610 954 -2604
rect 948 -2616 954 -2610
rect 948 -2622 954 -2616
rect 948 -2628 954 -2622
rect 948 -2634 954 -2628
rect 948 -2640 954 -2634
rect 948 -2646 954 -2640
rect 948 -2652 954 -2646
rect 948 -2658 954 -2652
rect 948 -2664 954 -2658
rect 948 -2670 954 -2664
rect 948 -2676 954 -2670
rect 948 -2682 954 -2676
rect 948 -2688 954 -2682
rect 948 -2694 954 -2688
rect 948 -2700 954 -2694
rect 948 -2706 954 -2700
rect 948 -2712 954 -2706
rect 948 -2718 954 -2712
rect 948 -2724 954 -2718
rect 948 -2730 954 -2724
rect 948 -2736 954 -2730
rect 948 -2742 954 -2736
rect 948 -2748 954 -2742
rect 948 -2754 954 -2748
rect 948 -2760 954 -2754
rect 948 -2766 954 -2760
rect 948 -2772 954 -2766
rect 948 -2778 954 -2772
rect 948 -2784 954 -2778
rect 948 -2790 954 -2784
rect 948 -2796 954 -2790
rect 948 -2802 954 -2796
rect 948 -2808 954 -2802
rect 948 -2814 954 -2808
rect 948 -2820 954 -2814
rect 948 -2826 954 -2820
rect 948 -2832 954 -2826
rect 948 -2838 954 -2832
rect 948 -2844 954 -2838
rect 948 -2850 954 -2844
rect 948 -2856 954 -2850
rect 948 -2862 954 -2856
rect 948 -2868 954 -2862
rect 948 -2874 954 -2868
rect 948 -2880 954 -2874
rect 948 -2886 954 -2880
rect 948 -2892 954 -2886
rect 948 -2898 954 -2892
rect 948 -2904 954 -2898
rect 948 -2910 954 -2904
rect 948 -2916 954 -2910
rect 948 -2922 954 -2916
rect 948 -2928 954 -2922
rect 948 -2934 954 -2928
rect 948 -2940 954 -2934
rect 948 -2946 954 -2940
rect 948 -2952 954 -2946
rect 948 -2958 954 -2952
rect 948 -2964 954 -2958
rect 948 -2970 954 -2964
rect 948 -2976 954 -2970
rect 948 -2982 954 -2976
rect 948 -2988 954 -2982
rect 948 -2994 954 -2988
rect 948 -3000 954 -2994
rect 948 -3006 954 -3000
rect 948 -3012 954 -3006
rect 948 -3018 954 -3012
rect 948 -3024 954 -3018
rect 948 -3030 954 -3024
rect 948 -3036 954 -3030
rect 948 -3150 954 -3144
rect 948 -3156 954 -3150
rect 948 -3162 954 -3156
rect 948 -3168 954 -3162
rect 948 -3174 954 -3168
rect 948 -3180 954 -3174
rect 948 -3186 954 -3180
rect 948 -3192 954 -3186
rect 948 -3198 954 -3192
rect 948 -3204 954 -3198
rect 948 -3210 954 -3204
rect 948 -3216 954 -3210
rect 948 -3282 954 -3276
rect 948 -3288 954 -3282
rect 948 -3294 954 -3288
rect 948 -3300 954 -3294
rect 948 -3306 954 -3300
rect 948 -3312 954 -3306
rect 948 -3318 954 -3312
rect 948 -3324 954 -3318
rect 948 -3330 954 -3324
rect 948 -3336 954 -3330
rect 948 -3342 954 -3336
rect 948 -3348 954 -3342
rect 948 -3354 954 -3348
rect 948 -3360 954 -3354
rect 948 -3366 954 -3360
rect 948 -3372 954 -3366
rect 948 -3438 954 -3432
rect 948 -3444 954 -3438
rect 948 -3450 954 -3444
rect 948 -3456 954 -3450
rect 948 -3462 954 -3456
rect 948 -3468 954 -3462
rect 948 -3474 954 -3468
rect 948 -3480 954 -3474
rect 948 -3486 954 -3480
rect 954 -1134 960 -1128
rect 954 -1140 960 -1134
rect 954 -1146 960 -1140
rect 954 -1152 960 -1146
rect 954 -1158 960 -1152
rect 954 -1164 960 -1158
rect 954 -1170 960 -1164
rect 954 -1176 960 -1170
rect 954 -1182 960 -1176
rect 954 -1188 960 -1182
rect 954 -1194 960 -1188
rect 954 -1200 960 -1194
rect 954 -1206 960 -1200
rect 954 -1212 960 -1206
rect 954 -1218 960 -1212
rect 954 -1224 960 -1218
rect 954 -1230 960 -1224
rect 954 -1236 960 -1230
rect 954 -1242 960 -1236
rect 954 -1248 960 -1242
rect 954 -1254 960 -1248
rect 954 -1260 960 -1254
rect 954 -1266 960 -1260
rect 954 -1272 960 -1266
rect 954 -1278 960 -1272
rect 954 -1284 960 -1278
rect 954 -1290 960 -1284
rect 954 -1296 960 -1290
rect 954 -1302 960 -1296
rect 954 -1308 960 -1302
rect 954 -1314 960 -1308
rect 954 -1320 960 -1314
rect 954 -1326 960 -1320
rect 954 -1332 960 -1326
rect 954 -1338 960 -1332
rect 954 -2574 960 -2568
rect 954 -2580 960 -2574
rect 954 -2586 960 -2580
rect 954 -2592 960 -2586
rect 954 -2598 960 -2592
rect 954 -2604 960 -2598
rect 954 -2610 960 -2604
rect 954 -2616 960 -2610
rect 954 -2622 960 -2616
rect 954 -2628 960 -2622
rect 954 -2634 960 -2628
rect 954 -2640 960 -2634
rect 954 -2646 960 -2640
rect 954 -2652 960 -2646
rect 954 -2658 960 -2652
rect 954 -2664 960 -2658
rect 954 -2670 960 -2664
rect 954 -2676 960 -2670
rect 954 -2682 960 -2676
rect 954 -2688 960 -2682
rect 954 -2694 960 -2688
rect 954 -2700 960 -2694
rect 954 -2706 960 -2700
rect 954 -2712 960 -2706
rect 954 -2718 960 -2712
rect 954 -2724 960 -2718
rect 954 -2730 960 -2724
rect 954 -2736 960 -2730
rect 954 -2742 960 -2736
rect 954 -2748 960 -2742
rect 954 -2754 960 -2748
rect 954 -2760 960 -2754
rect 954 -2766 960 -2760
rect 954 -2772 960 -2766
rect 954 -2778 960 -2772
rect 954 -2784 960 -2778
rect 954 -2790 960 -2784
rect 954 -2796 960 -2790
rect 954 -2802 960 -2796
rect 954 -2808 960 -2802
rect 954 -2814 960 -2808
rect 954 -2820 960 -2814
rect 954 -2826 960 -2820
rect 954 -2832 960 -2826
rect 954 -2838 960 -2832
rect 954 -2844 960 -2838
rect 954 -2850 960 -2844
rect 954 -2856 960 -2850
rect 954 -2862 960 -2856
rect 954 -2868 960 -2862
rect 954 -2874 960 -2868
rect 954 -2880 960 -2874
rect 954 -2886 960 -2880
rect 954 -2892 960 -2886
rect 954 -2898 960 -2892
rect 954 -2904 960 -2898
rect 954 -2910 960 -2904
rect 954 -2916 960 -2910
rect 954 -2922 960 -2916
rect 954 -2928 960 -2922
rect 954 -2934 960 -2928
rect 954 -2940 960 -2934
rect 954 -2946 960 -2940
rect 954 -2952 960 -2946
rect 954 -2958 960 -2952
rect 954 -2964 960 -2958
rect 954 -2970 960 -2964
rect 954 -2976 960 -2970
rect 954 -2982 960 -2976
rect 954 -2988 960 -2982
rect 954 -2994 960 -2988
rect 954 -3000 960 -2994
rect 954 -3006 960 -3000
rect 954 -3012 960 -3006
rect 954 -3018 960 -3012
rect 954 -3024 960 -3018
rect 954 -3132 960 -3126
rect 954 -3138 960 -3132
rect 954 -3144 960 -3138
rect 954 -3150 960 -3144
rect 954 -3156 960 -3150
rect 954 -3162 960 -3156
rect 954 -3168 960 -3162
rect 954 -3174 960 -3168
rect 954 -3180 960 -3174
rect 954 -3186 960 -3180
rect 954 -3192 960 -3186
rect 954 -3198 960 -3192
rect 954 -3204 960 -3198
rect 954 -3210 960 -3204
rect 954 -3282 960 -3276
rect 954 -3288 960 -3282
rect 954 -3294 960 -3288
rect 954 -3300 960 -3294
rect 954 -3306 960 -3300
rect 954 -3312 960 -3306
rect 954 -3318 960 -3312
rect 954 -3324 960 -3318
rect 954 -3330 960 -3324
rect 954 -3336 960 -3330
rect 954 -3342 960 -3336
rect 954 -3348 960 -3342
rect 954 -3354 960 -3348
rect 954 -3360 960 -3354
rect 954 -3366 960 -3360
rect 954 -3432 960 -3426
rect 954 -3438 960 -3432
rect 954 -3444 960 -3438
rect 954 -3450 960 -3444
rect 954 -3456 960 -3450
rect 954 -3462 960 -3456
rect 954 -3468 960 -3462
rect 954 -3474 960 -3468
rect 954 -3480 960 -3474
rect 954 -3486 960 -3480
rect 954 -3492 960 -3486
rect 960 -1128 966 -1122
rect 960 -1134 966 -1128
rect 960 -1140 966 -1134
rect 960 -1146 966 -1140
rect 960 -1152 966 -1146
rect 960 -1158 966 -1152
rect 960 -1164 966 -1158
rect 960 -1170 966 -1164
rect 960 -1176 966 -1170
rect 960 -1182 966 -1176
rect 960 -1188 966 -1182
rect 960 -1194 966 -1188
rect 960 -1200 966 -1194
rect 960 -1206 966 -1200
rect 960 -1212 966 -1206
rect 960 -1218 966 -1212
rect 960 -1224 966 -1218
rect 960 -1230 966 -1224
rect 960 -1236 966 -1230
rect 960 -1242 966 -1236
rect 960 -1248 966 -1242
rect 960 -1254 966 -1248
rect 960 -1260 966 -1254
rect 960 -1266 966 -1260
rect 960 -1272 966 -1266
rect 960 -1278 966 -1272
rect 960 -1284 966 -1278
rect 960 -1290 966 -1284
rect 960 -1296 966 -1290
rect 960 -1302 966 -1296
rect 960 -1308 966 -1302
rect 960 -1314 966 -1308
rect 960 -1320 966 -1314
rect 960 -1326 966 -1320
rect 960 -1332 966 -1326
rect 960 -1338 966 -1332
rect 960 -2550 966 -2544
rect 960 -2556 966 -2550
rect 960 -2562 966 -2556
rect 960 -2568 966 -2562
rect 960 -2574 966 -2568
rect 960 -2580 966 -2574
rect 960 -2586 966 -2580
rect 960 -2592 966 -2586
rect 960 -2598 966 -2592
rect 960 -2604 966 -2598
rect 960 -2610 966 -2604
rect 960 -2616 966 -2610
rect 960 -2622 966 -2616
rect 960 -2628 966 -2622
rect 960 -2634 966 -2628
rect 960 -2640 966 -2634
rect 960 -2646 966 -2640
rect 960 -2652 966 -2646
rect 960 -2658 966 -2652
rect 960 -2664 966 -2658
rect 960 -2670 966 -2664
rect 960 -2676 966 -2670
rect 960 -2682 966 -2676
rect 960 -2688 966 -2682
rect 960 -2694 966 -2688
rect 960 -2700 966 -2694
rect 960 -2706 966 -2700
rect 960 -2712 966 -2706
rect 960 -2718 966 -2712
rect 960 -2724 966 -2718
rect 960 -2730 966 -2724
rect 960 -2736 966 -2730
rect 960 -2742 966 -2736
rect 960 -2748 966 -2742
rect 960 -2754 966 -2748
rect 960 -2760 966 -2754
rect 960 -2766 966 -2760
rect 960 -2772 966 -2766
rect 960 -2778 966 -2772
rect 960 -2784 966 -2778
rect 960 -2790 966 -2784
rect 960 -2796 966 -2790
rect 960 -2802 966 -2796
rect 960 -2808 966 -2802
rect 960 -2814 966 -2808
rect 960 -2820 966 -2814
rect 960 -2826 966 -2820
rect 960 -2832 966 -2826
rect 960 -2838 966 -2832
rect 960 -2844 966 -2838
rect 960 -2850 966 -2844
rect 960 -2856 966 -2850
rect 960 -2862 966 -2856
rect 960 -2868 966 -2862
rect 960 -2874 966 -2868
rect 960 -2880 966 -2874
rect 960 -2886 966 -2880
rect 960 -2892 966 -2886
rect 960 -2898 966 -2892
rect 960 -2904 966 -2898
rect 960 -2910 966 -2904
rect 960 -2916 966 -2910
rect 960 -2922 966 -2916
rect 960 -2928 966 -2922
rect 960 -2934 966 -2928
rect 960 -2940 966 -2934
rect 960 -2946 966 -2940
rect 960 -2952 966 -2946
rect 960 -2958 966 -2952
rect 960 -2964 966 -2958
rect 960 -2970 966 -2964
rect 960 -2976 966 -2970
rect 960 -2982 966 -2976
rect 960 -2988 966 -2982
rect 960 -2994 966 -2988
rect 960 -3000 966 -2994
rect 960 -3006 966 -3000
rect 960 -3012 966 -3006
rect 960 -3120 966 -3114
rect 960 -3126 966 -3120
rect 960 -3132 966 -3126
rect 960 -3138 966 -3132
rect 960 -3144 966 -3138
rect 960 -3150 966 -3144
rect 960 -3156 966 -3150
rect 960 -3162 966 -3156
rect 960 -3168 966 -3162
rect 960 -3174 966 -3168
rect 960 -3180 966 -3174
rect 960 -3186 966 -3180
rect 960 -3192 966 -3186
rect 960 -3198 966 -3192
rect 960 -3204 966 -3198
rect 960 -3276 966 -3270
rect 960 -3282 966 -3276
rect 960 -3288 966 -3282
rect 960 -3294 966 -3288
rect 960 -3300 966 -3294
rect 960 -3306 966 -3300
rect 960 -3312 966 -3306
rect 960 -3318 966 -3312
rect 960 -3324 966 -3318
rect 960 -3330 966 -3324
rect 960 -3336 966 -3330
rect 960 -3342 966 -3336
rect 960 -3348 966 -3342
rect 960 -3354 966 -3348
rect 960 -3360 966 -3354
rect 960 -3426 966 -3420
rect 960 -3432 966 -3426
rect 960 -3438 966 -3432
rect 960 -3444 966 -3438
rect 960 -3450 966 -3444
rect 960 -3456 966 -3450
rect 960 -3462 966 -3456
rect 960 -3468 966 -3462
rect 960 -3474 966 -3468
rect 960 -3480 966 -3474
rect 960 -3486 966 -3480
rect 960 -3492 966 -3486
rect 966 -1128 972 -1122
rect 966 -1134 972 -1128
rect 966 -1140 972 -1134
rect 966 -1146 972 -1140
rect 966 -1152 972 -1146
rect 966 -1158 972 -1152
rect 966 -1164 972 -1158
rect 966 -1170 972 -1164
rect 966 -1176 972 -1170
rect 966 -1182 972 -1176
rect 966 -1188 972 -1182
rect 966 -1194 972 -1188
rect 966 -1200 972 -1194
rect 966 -1206 972 -1200
rect 966 -1212 972 -1206
rect 966 -1218 972 -1212
rect 966 -1224 972 -1218
rect 966 -1230 972 -1224
rect 966 -1236 972 -1230
rect 966 -1242 972 -1236
rect 966 -1248 972 -1242
rect 966 -1254 972 -1248
rect 966 -1260 972 -1254
rect 966 -1266 972 -1260
rect 966 -1272 972 -1266
rect 966 -1278 972 -1272
rect 966 -1284 972 -1278
rect 966 -1290 972 -1284
rect 966 -1296 972 -1290
rect 966 -1302 972 -1296
rect 966 -1308 972 -1302
rect 966 -1314 972 -1308
rect 966 -1320 972 -1314
rect 966 -1326 972 -1320
rect 966 -1332 972 -1326
rect 966 -1338 972 -1332
rect 966 -2532 972 -2526
rect 966 -2538 972 -2532
rect 966 -2544 972 -2538
rect 966 -2550 972 -2544
rect 966 -2556 972 -2550
rect 966 -2562 972 -2556
rect 966 -2568 972 -2562
rect 966 -2574 972 -2568
rect 966 -2580 972 -2574
rect 966 -2586 972 -2580
rect 966 -2592 972 -2586
rect 966 -2598 972 -2592
rect 966 -2604 972 -2598
rect 966 -2610 972 -2604
rect 966 -2616 972 -2610
rect 966 -2622 972 -2616
rect 966 -2628 972 -2622
rect 966 -2634 972 -2628
rect 966 -2640 972 -2634
rect 966 -2646 972 -2640
rect 966 -2652 972 -2646
rect 966 -2658 972 -2652
rect 966 -2664 972 -2658
rect 966 -2670 972 -2664
rect 966 -2676 972 -2670
rect 966 -2682 972 -2676
rect 966 -2688 972 -2682
rect 966 -2694 972 -2688
rect 966 -2700 972 -2694
rect 966 -2706 972 -2700
rect 966 -2712 972 -2706
rect 966 -2718 972 -2712
rect 966 -2724 972 -2718
rect 966 -2730 972 -2724
rect 966 -2736 972 -2730
rect 966 -2742 972 -2736
rect 966 -2748 972 -2742
rect 966 -2754 972 -2748
rect 966 -2760 972 -2754
rect 966 -2766 972 -2760
rect 966 -2772 972 -2766
rect 966 -2778 972 -2772
rect 966 -2784 972 -2778
rect 966 -2790 972 -2784
rect 966 -2796 972 -2790
rect 966 -2802 972 -2796
rect 966 -2808 972 -2802
rect 966 -2814 972 -2808
rect 966 -2820 972 -2814
rect 966 -2826 972 -2820
rect 966 -2832 972 -2826
rect 966 -2838 972 -2832
rect 966 -2844 972 -2838
rect 966 -2850 972 -2844
rect 966 -2856 972 -2850
rect 966 -2862 972 -2856
rect 966 -2868 972 -2862
rect 966 -2874 972 -2868
rect 966 -2880 972 -2874
rect 966 -2886 972 -2880
rect 966 -2892 972 -2886
rect 966 -2898 972 -2892
rect 966 -2904 972 -2898
rect 966 -2910 972 -2904
rect 966 -2916 972 -2910
rect 966 -2922 972 -2916
rect 966 -2928 972 -2922
rect 966 -2934 972 -2928
rect 966 -2940 972 -2934
rect 966 -2946 972 -2940
rect 966 -2952 972 -2946
rect 966 -2958 972 -2952
rect 966 -2964 972 -2958
rect 966 -2970 972 -2964
rect 966 -2976 972 -2970
rect 966 -2982 972 -2976
rect 966 -2988 972 -2982
rect 966 -2994 972 -2988
rect 966 -3000 972 -2994
rect 966 -3108 972 -3102
rect 966 -3114 972 -3108
rect 966 -3120 972 -3114
rect 966 -3126 972 -3120
rect 966 -3132 972 -3126
rect 966 -3138 972 -3132
rect 966 -3144 972 -3138
rect 966 -3150 972 -3144
rect 966 -3156 972 -3150
rect 966 -3162 972 -3156
rect 966 -3168 972 -3162
rect 966 -3174 972 -3168
rect 966 -3180 972 -3174
rect 966 -3186 972 -3180
rect 966 -3192 972 -3186
rect 966 -3198 972 -3192
rect 966 -3204 972 -3198
rect 966 -3270 972 -3264
rect 966 -3276 972 -3270
rect 966 -3282 972 -3276
rect 966 -3288 972 -3282
rect 966 -3294 972 -3288
rect 966 -3300 972 -3294
rect 966 -3306 972 -3300
rect 966 -3312 972 -3306
rect 966 -3318 972 -3312
rect 966 -3324 972 -3318
rect 966 -3330 972 -3324
rect 966 -3336 972 -3330
rect 966 -3342 972 -3336
rect 966 -3348 972 -3342
rect 966 -3354 972 -3348
rect 966 -3360 972 -3354
rect 966 -3420 972 -3414
rect 966 -3426 972 -3420
rect 966 -3432 972 -3426
rect 966 -3438 972 -3432
rect 966 -3444 972 -3438
rect 966 -3450 972 -3444
rect 966 -3456 972 -3450
rect 966 -3462 972 -3456
rect 966 -3468 972 -3462
rect 966 -3474 972 -3468
rect 966 -3480 972 -3474
rect 966 -3486 972 -3480
rect 966 -3492 972 -3486
rect 972 -1128 978 -1122
rect 972 -1134 978 -1128
rect 972 -1140 978 -1134
rect 972 -1146 978 -1140
rect 972 -1152 978 -1146
rect 972 -1158 978 -1152
rect 972 -1164 978 -1158
rect 972 -1170 978 -1164
rect 972 -1176 978 -1170
rect 972 -1182 978 -1176
rect 972 -1188 978 -1182
rect 972 -1194 978 -1188
rect 972 -1200 978 -1194
rect 972 -1206 978 -1200
rect 972 -1212 978 -1206
rect 972 -1218 978 -1212
rect 972 -1224 978 -1218
rect 972 -1230 978 -1224
rect 972 -1236 978 -1230
rect 972 -1242 978 -1236
rect 972 -1248 978 -1242
rect 972 -1254 978 -1248
rect 972 -1260 978 -1254
rect 972 -1266 978 -1260
rect 972 -1272 978 -1266
rect 972 -1278 978 -1272
rect 972 -1284 978 -1278
rect 972 -1290 978 -1284
rect 972 -1296 978 -1290
rect 972 -1302 978 -1296
rect 972 -1308 978 -1302
rect 972 -1314 978 -1308
rect 972 -1320 978 -1314
rect 972 -1326 978 -1320
rect 972 -1332 978 -1326
rect 972 -1338 978 -1332
rect 972 -2508 978 -2502
rect 972 -2514 978 -2508
rect 972 -2520 978 -2514
rect 972 -2526 978 -2520
rect 972 -2532 978 -2526
rect 972 -2538 978 -2532
rect 972 -2544 978 -2538
rect 972 -2550 978 -2544
rect 972 -2556 978 -2550
rect 972 -2562 978 -2556
rect 972 -2568 978 -2562
rect 972 -2574 978 -2568
rect 972 -2580 978 -2574
rect 972 -2586 978 -2580
rect 972 -2592 978 -2586
rect 972 -2598 978 -2592
rect 972 -2604 978 -2598
rect 972 -2610 978 -2604
rect 972 -2616 978 -2610
rect 972 -2622 978 -2616
rect 972 -2628 978 -2622
rect 972 -2634 978 -2628
rect 972 -2640 978 -2634
rect 972 -2646 978 -2640
rect 972 -2652 978 -2646
rect 972 -2658 978 -2652
rect 972 -2664 978 -2658
rect 972 -2670 978 -2664
rect 972 -2676 978 -2670
rect 972 -2682 978 -2676
rect 972 -2688 978 -2682
rect 972 -2694 978 -2688
rect 972 -2700 978 -2694
rect 972 -2706 978 -2700
rect 972 -2712 978 -2706
rect 972 -2718 978 -2712
rect 972 -2724 978 -2718
rect 972 -2730 978 -2724
rect 972 -2736 978 -2730
rect 972 -2742 978 -2736
rect 972 -2748 978 -2742
rect 972 -2754 978 -2748
rect 972 -2760 978 -2754
rect 972 -2766 978 -2760
rect 972 -2772 978 -2766
rect 972 -2778 978 -2772
rect 972 -2784 978 -2778
rect 972 -2790 978 -2784
rect 972 -2796 978 -2790
rect 972 -2802 978 -2796
rect 972 -2808 978 -2802
rect 972 -2814 978 -2808
rect 972 -2820 978 -2814
rect 972 -2826 978 -2820
rect 972 -2832 978 -2826
rect 972 -2838 978 -2832
rect 972 -2844 978 -2838
rect 972 -2850 978 -2844
rect 972 -2856 978 -2850
rect 972 -2862 978 -2856
rect 972 -2868 978 -2862
rect 972 -2874 978 -2868
rect 972 -2880 978 -2874
rect 972 -2886 978 -2880
rect 972 -2892 978 -2886
rect 972 -2898 978 -2892
rect 972 -2904 978 -2898
rect 972 -2910 978 -2904
rect 972 -2916 978 -2910
rect 972 -2922 978 -2916
rect 972 -2928 978 -2922
rect 972 -2934 978 -2928
rect 972 -2940 978 -2934
rect 972 -2946 978 -2940
rect 972 -2952 978 -2946
rect 972 -2958 978 -2952
rect 972 -2964 978 -2958
rect 972 -2970 978 -2964
rect 972 -2976 978 -2970
rect 972 -2982 978 -2976
rect 972 -2988 978 -2982
rect 972 -3090 978 -3084
rect 972 -3096 978 -3090
rect 972 -3102 978 -3096
rect 972 -3108 978 -3102
rect 972 -3114 978 -3108
rect 972 -3120 978 -3114
rect 972 -3126 978 -3120
rect 972 -3132 978 -3126
rect 972 -3138 978 -3132
rect 972 -3144 978 -3138
rect 972 -3150 978 -3144
rect 972 -3156 978 -3150
rect 972 -3162 978 -3156
rect 972 -3168 978 -3162
rect 972 -3174 978 -3168
rect 972 -3180 978 -3174
rect 972 -3186 978 -3180
rect 972 -3192 978 -3186
rect 972 -3198 978 -3192
rect 972 -3264 978 -3258
rect 972 -3270 978 -3264
rect 972 -3276 978 -3270
rect 972 -3282 978 -3276
rect 972 -3288 978 -3282
rect 972 -3294 978 -3288
rect 972 -3300 978 -3294
rect 972 -3306 978 -3300
rect 972 -3312 978 -3306
rect 972 -3318 978 -3312
rect 972 -3324 978 -3318
rect 972 -3330 978 -3324
rect 972 -3336 978 -3330
rect 972 -3342 978 -3336
rect 972 -3348 978 -3342
rect 972 -3354 978 -3348
rect 972 -3414 978 -3408
rect 972 -3420 978 -3414
rect 972 -3426 978 -3420
rect 972 -3432 978 -3426
rect 972 -3438 978 -3432
rect 972 -3444 978 -3438
rect 972 -3450 978 -3444
rect 972 -3456 978 -3450
rect 972 -3462 978 -3456
rect 972 -3468 978 -3462
rect 972 -3474 978 -3468
rect 972 -3480 978 -3474
rect 972 -3486 978 -3480
rect 972 -3492 978 -3486
rect 978 -1128 984 -1122
rect 978 -1134 984 -1128
rect 978 -1140 984 -1134
rect 978 -1146 984 -1140
rect 978 -1152 984 -1146
rect 978 -1158 984 -1152
rect 978 -1164 984 -1158
rect 978 -1170 984 -1164
rect 978 -1176 984 -1170
rect 978 -1182 984 -1176
rect 978 -1188 984 -1182
rect 978 -1194 984 -1188
rect 978 -1200 984 -1194
rect 978 -1206 984 -1200
rect 978 -1212 984 -1206
rect 978 -1218 984 -1212
rect 978 -1224 984 -1218
rect 978 -1230 984 -1224
rect 978 -1236 984 -1230
rect 978 -1242 984 -1236
rect 978 -1248 984 -1242
rect 978 -1254 984 -1248
rect 978 -1260 984 -1254
rect 978 -1266 984 -1260
rect 978 -1272 984 -1266
rect 978 -1278 984 -1272
rect 978 -1284 984 -1278
rect 978 -1290 984 -1284
rect 978 -1296 984 -1290
rect 978 -1302 984 -1296
rect 978 -1308 984 -1302
rect 978 -1314 984 -1308
rect 978 -1320 984 -1314
rect 978 -1326 984 -1320
rect 978 -1332 984 -1326
rect 978 -2490 984 -2484
rect 978 -2496 984 -2490
rect 978 -2502 984 -2496
rect 978 -2508 984 -2502
rect 978 -2514 984 -2508
rect 978 -2520 984 -2514
rect 978 -2526 984 -2520
rect 978 -2532 984 -2526
rect 978 -2538 984 -2532
rect 978 -2544 984 -2538
rect 978 -2550 984 -2544
rect 978 -2556 984 -2550
rect 978 -2562 984 -2556
rect 978 -2568 984 -2562
rect 978 -2574 984 -2568
rect 978 -2580 984 -2574
rect 978 -2586 984 -2580
rect 978 -2592 984 -2586
rect 978 -2598 984 -2592
rect 978 -2604 984 -2598
rect 978 -2610 984 -2604
rect 978 -2616 984 -2610
rect 978 -2622 984 -2616
rect 978 -2628 984 -2622
rect 978 -2634 984 -2628
rect 978 -2640 984 -2634
rect 978 -2646 984 -2640
rect 978 -2652 984 -2646
rect 978 -2658 984 -2652
rect 978 -2664 984 -2658
rect 978 -2670 984 -2664
rect 978 -2676 984 -2670
rect 978 -2682 984 -2676
rect 978 -2688 984 -2682
rect 978 -2694 984 -2688
rect 978 -2700 984 -2694
rect 978 -2706 984 -2700
rect 978 -2712 984 -2706
rect 978 -2718 984 -2712
rect 978 -2724 984 -2718
rect 978 -2730 984 -2724
rect 978 -2736 984 -2730
rect 978 -2742 984 -2736
rect 978 -2748 984 -2742
rect 978 -2754 984 -2748
rect 978 -2760 984 -2754
rect 978 -2766 984 -2760
rect 978 -2772 984 -2766
rect 978 -2778 984 -2772
rect 978 -2784 984 -2778
rect 978 -2790 984 -2784
rect 978 -2796 984 -2790
rect 978 -2802 984 -2796
rect 978 -2808 984 -2802
rect 978 -2814 984 -2808
rect 978 -2820 984 -2814
rect 978 -2826 984 -2820
rect 978 -2832 984 -2826
rect 978 -2838 984 -2832
rect 978 -2844 984 -2838
rect 978 -2850 984 -2844
rect 978 -2856 984 -2850
rect 978 -2862 984 -2856
rect 978 -2868 984 -2862
rect 978 -2874 984 -2868
rect 978 -2880 984 -2874
rect 978 -2886 984 -2880
rect 978 -2892 984 -2886
rect 978 -2898 984 -2892
rect 978 -2904 984 -2898
rect 978 -2910 984 -2904
rect 978 -2916 984 -2910
rect 978 -2922 984 -2916
rect 978 -2928 984 -2922
rect 978 -2934 984 -2928
rect 978 -2940 984 -2934
rect 978 -2946 984 -2940
rect 978 -2952 984 -2946
rect 978 -2958 984 -2952
rect 978 -2964 984 -2958
rect 978 -2970 984 -2964
rect 978 -2976 984 -2970
rect 978 -3078 984 -3072
rect 978 -3084 984 -3078
rect 978 -3090 984 -3084
rect 978 -3096 984 -3090
rect 978 -3102 984 -3096
rect 978 -3108 984 -3102
rect 978 -3114 984 -3108
rect 978 -3120 984 -3114
rect 978 -3126 984 -3120
rect 978 -3132 984 -3126
rect 978 -3138 984 -3132
rect 978 -3144 984 -3138
rect 978 -3150 984 -3144
rect 978 -3156 984 -3150
rect 978 -3162 984 -3156
rect 978 -3168 984 -3162
rect 978 -3174 984 -3168
rect 978 -3180 984 -3174
rect 978 -3186 984 -3180
rect 978 -3192 984 -3186
rect 978 -3258 984 -3252
rect 978 -3264 984 -3258
rect 978 -3270 984 -3264
rect 978 -3276 984 -3270
rect 978 -3282 984 -3276
rect 978 -3288 984 -3282
rect 978 -3294 984 -3288
rect 978 -3300 984 -3294
rect 978 -3306 984 -3300
rect 978 -3312 984 -3306
rect 978 -3318 984 -3312
rect 978 -3324 984 -3318
rect 978 -3330 984 -3324
rect 978 -3336 984 -3330
rect 978 -3342 984 -3336
rect 978 -3348 984 -3342
rect 978 -3414 984 -3408
rect 978 -3420 984 -3414
rect 978 -3426 984 -3420
rect 978 -3432 984 -3426
rect 978 -3438 984 -3432
rect 978 -3444 984 -3438
rect 978 -3450 984 -3444
rect 978 -3456 984 -3450
rect 978 -3462 984 -3456
rect 978 -3468 984 -3462
rect 978 -3474 984 -3468
rect 978 -3480 984 -3474
rect 978 -3486 984 -3480
rect 978 -3492 984 -3486
rect 984 -1128 990 -1122
rect 984 -1134 990 -1128
rect 984 -1140 990 -1134
rect 984 -1146 990 -1140
rect 984 -1152 990 -1146
rect 984 -1158 990 -1152
rect 984 -1164 990 -1158
rect 984 -1170 990 -1164
rect 984 -1176 990 -1170
rect 984 -1182 990 -1176
rect 984 -1188 990 -1182
rect 984 -1194 990 -1188
rect 984 -1200 990 -1194
rect 984 -1206 990 -1200
rect 984 -1212 990 -1206
rect 984 -1218 990 -1212
rect 984 -1224 990 -1218
rect 984 -1230 990 -1224
rect 984 -1236 990 -1230
rect 984 -1242 990 -1236
rect 984 -1248 990 -1242
rect 984 -1254 990 -1248
rect 984 -1260 990 -1254
rect 984 -1266 990 -1260
rect 984 -1272 990 -1266
rect 984 -1278 990 -1272
rect 984 -1284 990 -1278
rect 984 -1290 990 -1284
rect 984 -1296 990 -1290
rect 984 -1302 990 -1296
rect 984 -1308 990 -1302
rect 984 -1314 990 -1308
rect 984 -1320 990 -1314
rect 984 -1326 990 -1320
rect 984 -1332 990 -1326
rect 984 -2466 990 -2460
rect 984 -2472 990 -2466
rect 984 -2478 990 -2472
rect 984 -2484 990 -2478
rect 984 -2490 990 -2484
rect 984 -2496 990 -2490
rect 984 -2502 990 -2496
rect 984 -2508 990 -2502
rect 984 -2514 990 -2508
rect 984 -2520 990 -2514
rect 984 -2526 990 -2520
rect 984 -2532 990 -2526
rect 984 -2538 990 -2532
rect 984 -2544 990 -2538
rect 984 -2550 990 -2544
rect 984 -2556 990 -2550
rect 984 -2562 990 -2556
rect 984 -2568 990 -2562
rect 984 -2574 990 -2568
rect 984 -2580 990 -2574
rect 984 -2586 990 -2580
rect 984 -2592 990 -2586
rect 984 -2598 990 -2592
rect 984 -2604 990 -2598
rect 984 -2610 990 -2604
rect 984 -2616 990 -2610
rect 984 -2622 990 -2616
rect 984 -2628 990 -2622
rect 984 -2634 990 -2628
rect 984 -2640 990 -2634
rect 984 -2646 990 -2640
rect 984 -2652 990 -2646
rect 984 -2658 990 -2652
rect 984 -2664 990 -2658
rect 984 -2670 990 -2664
rect 984 -2676 990 -2670
rect 984 -2682 990 -2676
rect 984 -2688 990 -2682
rect 984 -2694 990 -2688
rect 984 -2700 990 -2694
rect 984 -2706 990 -2700
rect 984 -2712 990 -2706
rect 984 -2718 990 -2712
rect 984 -2724 990 -2718
rect 984 -2730 990 -2724
rect 984 -2736 990 -2730
rect 984 -2742 990 -2736
rect 984 -2748 990 -2742
rect 984 -2754 990 -2748
rect 984 -2760 990 -2754
rect 984 -2766 990 -2760
rect 984 -2772 990 -2766
rect 984 -2778 990 -2772
rect 984 -2784 990 -2778
rect 984 -2790 990 -2784
rect 984 -2796 990 -2790
rect 984 -2802 990 -2796
rect 984 -2808 990 -2802
rect 984 -2814 990 -2808
rect 984 -2820 990 -2814
rect 984 -2826 990 -2820
rect 984 -2832 990 -2826
rect 984 -2838 990 -2832
rect 984 -2844 990 -2838
rect 984 -2850 990 -2844
rect 984 -2856 990 -2850
rect 984 -2862 990 -2856
rect 984 -2868 990 -2862
rect 984 -2874 990 -2868
rect 984 -2880 990 -2874
rect 984 -2886 990 -2880
rect 984 -2892 990 -2886
rect 984 -2898 990 -2892
rect 984 -2904 990 -2898
rect 984 -2910 990 -2904
rect 984 -2916 990 -2910
rect 984 -2922 990 -2916
rect 984 -2928 990 -2922
rect 984 -2934 990 -2928
rect 984 -2940 990 -2934
rect 984 -2946 990 -2940
rect 984 -2952 990 -2946
rect 984 -2958 990 -2952
rect 984 -2964 990 -2958
rect 984 -3066 990 -3060
rect 984 -3072 990 -3066
rect 984 -3078 990 -3072
rect 984 -3084 990 -3078
rect 984 -3090 990 -3084
rect 984 -3096 990 -3090
rect 984 -3102 990 -3096
rect 984 -3108 990 -3102
rect 984 -3114 990 -3108
rect 984 -3120 990 -3114
rect 984 -3126 990 -3120
rect 984 -3132 990 -3126
rect 984 -3138 990 -3132
rect 984 -3144 990 -3138
rect 984 -3150 990 -3144
rect 984 -3156 990 -3150
rect 984 -3162 990 -3156
rect 984 -3168 990 -3162
rect 984 -3174 990 -3168
rect 984 -3180 990 -3174
rect 984 -3186 990 -3180
rect 984 -3252 990 -3246
rect 984 -3258 990 -3252
rect 984 -3264 990 -3258
rect 984 -3270 990 -3264
rect 984 -3276 990 -3270
rect 984 -3282 990 -3276
rect 984 -3288 990 -3282
rect 984 -3294 990 -3288
rect 984 -3300 990 -3294
rect 984 -3306 990 -3300
rect 984 -3312 990 -3306
rect 984 -3318 990 -3312
rect 984 -3324 990 -3318
rect 984 -3330 990 -3324
rect 984 -3336 990 -3330
rect 984 -3342 990 -3336
rect 984 -3408 990 -3402
rect 984 -3414 990 -3408
rect 984 -3420 990 -3414
rect 984 -3426 990 -3420
rect 984 -3432 990 -3426
rect 984 -3438 990 -3432
rect 984 -3444 990 -3438
rect 984 -3450 990 -3444
rect 984 -3456 990 -3450
rect 984 -3462 990 -3456
rect 984 -3468 990 -3462
rect 984 -3474 990 -3468
rect 984 -3480 990 -3474
rect 984 -3486 990 -3480
rect 984 -3492 990 -3486
rect 990 -1122 996 -1116
rect 990 -1128 996 -1122
rect 990 -1134 996 -1128
rect 990 -1140 996 -1134
rect 990 -1146 996 -1140
rect 990 -1152 996 -1146
rect 990 -1158 996 -1152
rect 990 -1164 996 -1158
rect 990 -1170 996 -1164
rect 990 -1176 996 -1170
rect 990 -1182 996 -1176
rect 990 -1188 996 -1182
rect 990 -1194 996 -1188
rect 990 -1200 996 -1194
rect 990 -1206 996 -1200
rect 990 -1212 996 -1206
rect 990 -1218 996 -1212
rect 990 -1224 996 -1218
rect 990 -1230 996 -1224
rect 990 -1236 996 -1230
rect 990 -1242 996 -1236
rect 990 -1248 996 -1242
rect 990 -1254 996 -1248
rect 990 -1260 996 -1254
rect 990 -1266 996 -1260
rect 990 -1272 996 -1266
rect 990 -1278 996 -1272
rect 990 -1284 996 -1278
rect 990 -1290 996 -1284
rect 990 -1296 996 -1290
rect 990 -1302 996 -1296
rect 990 -1308 996 -1302
rect 990 -1314 996 -1308
rect 990 -1320 996 -1314
rect 990 -1326 996 -1320
rect 990 -1332 996 -1326
rect 990 -2448 996 -2442
rect 990 -2454 996 -2448
rect 990 -2460 996 -2454
rect 990 -2466 996 -2460
rect 990 -2472 996 -2466
rect 990 -2478 996 -2472
rect 990 -2484 996 -2478
rect 990 -2490 996 -2484
rect 990 -2496 996 -2490
rect 990 -2502 996 -2496
rect 990 -2508 996 -2502
rect 990 -2514 996 -2508
rect 990 -2520 996 -2514
rect 990 -2526 996 -2520
rect 990 -2532 996 -2526
rect 990 -2538 996 -2532
rect 990 -2544 996 -2538
rect 990 -2550 996 -2544
rect 990 -2556 996 -2550
rect 990 -2562 996 -2556
rect 990 -2568 996 -2562
rect 990 -2574 996 -2568
rect 990 -2580 996 -2574
rect 990 -2586 996 -2580
rect 990 -2592 996 -2586
rect 990 -2598 996 -2592
rect 990 -2604 996 -2598
rect 990 -2610 996 -2604
rect 990 -2616 996 -2610
rect 990 -2622 996 -2616
rect 990 -2628 996 -2622
rect 990 -2634 996 -2628
rect 990 -2640 996 -2634
rect 990 -2646 996 -2640
rect 990 -2652 996 -2646
rect 990 -2658 996 -2652
rect 990 -2664 996 -2658
rect 990 -2670 996 -2664
rect 990 -2676 996 -2670
rect 990 -2682 996 -2676
rect 990 -2688 996 -2682
rect 990 -2694 996 -2688
rect 990 -2700 996 -2694
rect 990 -2706 996 -2700
rect 990 -2712 996 -2706
rect 990 -2718 996 -2712
rect 990 -2724 996 -2718
rect 990 -2730 996 -2724
rect 990 -2736 996 -2730
rect 990 -2742 996 -2736
rect 990 -2748 996 -2742
rect 990 -2754 996 -2748
rect 990 -2760 996 -2754
rect 990 -2766 996 -2760
rect 990 -2772 996 -2766
rect 990 -2778 996 -2772
rect 990 -2784 996 -2778
rect 990 -2790 996 -2784
rect 990 -2796 996 -2790
rect 990 -2802 996 -2796
rect 990 -2808 996 -2802
rect 990 -2814 996 -2808
rect 990 -2820 996 -2814
rect 990 -2826 996 -2820
rect 990 -2832 996 -2826
rect 990 -2838 996 -2832
rect 990 -2844 996 -2838
rect 990 -2850 996 -2844
rect 990 -2856 996 -2850
rect 990 -2862 996 -2856
rect 990 -2868 996 -2862
rect 990 -2874 996 -2868
rect 990 -2880 996 -2874
rect 990 -2886 996 -2880
rect 990 -2892 996 -2886
rect 990 -2898 996 -2892
rect 990 -2904 996 -2898
rect 990 -2910 996 -2904
rect 990 -2916 996 -2910
rect 990 -2922 996 -2916
rect 990 -2928 996 -2922
rect 990 -2934 996 -2928
rect 990 -2940 996 -2934
rect 990 -2946 996 -2940
rect 990 -2952 996 -2946
rect 990 -3054 996 -3048
rect 990 -3060 996 -3054
rect 990 -3066 996 -3060
rect 990 -3072 996 -3066
rect 990 -3078 996 -3072
rect 990 -3084 996 -3078
rect 990 -3090 996 -3084
rect 990 -3096 996 -3090
rect 990 -3102 996 -3096
rect 990 -3108 996 -3102
rect 990 -3114 996 -3108
rect 990 -3120 996 -3114
rect 990 -3126 996 -3120
rect 990 -3132 996 -3126
rect 990 -3138 996 -3132
rect 990 -3144 996 -3138
rect 990 -3150 996 -3144
rect 990 -3156 996 -3150
rect 990 -3162 996 -3156
rect 990 -3168 996 -3162
rect 990 -3174 996 -3168
rect 990 -3180 996 -3174
rect 990 -3186 996 -3180
rect 990 -3252 996 -3246
rect 990 -3258 996 -3252
rect 990 -3264 996 -3258
rect 990 -3270 996 -3264
rect 990 -3276 996 -3270
rect 990 -3282 996 -3276
rect 990 -3288 996 -3282
rect 990 -3294 996 -3288
rect 990 -3300 996 -3294
rect 990 -3306 996 -3300
rect 990 -3312 996 -3306
rect 990 -3318 996 -3312
rect 990 -3324 996 -3318
rect 990 -3330 996 -3324
rect 990 -3336 996 -3330
rect 990 -3342 996 -3336
rect 990 -3402 996 -3396
rect 990 -3408 996 -3402
rect 990 -3414 996 -3408
rect 990 -3420 996 -3414
rect 990 -3426 996 -3420
rect 990 -3432 996 -3426
rect 990 -3438 996 -3432
rect 990 -3444 996 -3438
rect 990 -3450 996 -3444
rect 990 -3456 996 -3450
rect 990 -3462 996 -3456
rect 990 -3468 996 -3462
rect 990 -3474 996 -3468
rect 990 -3480 996 -3474
rect 990 -3486 996 -3480
rect 990 -3492 996 -3486
rect 996 -1122 1002 -1116
rect 996 -1128 1002 -1122
rect 996 -1134 1002 -1128
rect 996 -1140 1002 -1134
rect 996 -1146 1002 -1140
rect 996 -1152 1002 -1146
rect 996 -1158 1002 -1152
rect 996 -1164 1002 -1158
rect 996 -1170 1002 -1164
rect 996 -1176 1002 -1170
rect 996 -1182 1002 -1176
rect 996 -1188 1002 -1182
rect 996 -1194 1002 -1188
rect 996 -1200 1002 -1194
rect 996 -1206 1002 -1200
rect 996 -1212 1002 -1206
rect 996 -1218 1002 -1212
rect 996 -1224 1002 -1218
rect 996 -1230 1002 -1224
rect 996 -1236 1002 -1230
rect 996 -1242 1002 -1236
rect 996 -1248 1002 -1242
rect 996 -1254 1002 -1248
rect 996 -1260 1002 -1254
rect 996 -1266 1002 -1260
rect 996 -1272 1002 -1266
rect 996 -1278 1002 -1272
rect 996 -1284 1002 -1278
rect 996 -1290 1002 -1284
rect 996 -1296 1002 -1290
rect 996 -1302 1002 -1296
rect 996 -1308 1002 -1302
rect 996 -1314 1002 -1308
rect 996 -1320 1002 -1314
rect 996 -1326 1002 -1320
rect 996 -1332 1002 -1326
rect 996 -2424 1002 -2418
rect 996 -2430 1002 -2424
rect 996 -2436 1002 -2430
rect 996 -2442 1002 -2436
rect 996 -2448 1002 -2442
rect 996 -2454 1002 -2448
rect 996 -2460 1002 -2454
rect 996 -2466 1002 -2460
rect 996 -2472 1002 -2466
rect 996 -2478 1002 -2472
rect 996 -2484 1002 -2478
rect 996 -2490 1002 -2484
rect 996 -2496 1002 -2490
rect 996 -2502 1002 -2496
rect 996 -2508 1002 -2502
rect 996 -2514 1002 -2508
rect 996 -2520 1002 -2514
rect 996 -2526 1002 -2520
rect 996 -2532 1002 -2526
rect 996 -2538 1002 -2532
rect 996 -2544 1002 -2538
rect 996 -2550 1002 -2544
rect 996 -2556 1002 -2550
rect 996 -2562 1002 -2556
rect 996 -2568 1002 -2562
rect 996 -2574 1002 -2568
rect 996 -2580 1002 -2574
rect 996 -2586 1002 -2580
rect 996 -2592 1002 -2586
rect 996 -2598 1002 -2592
rect 996 -2604 1002 -2598
rect 996 -2610 1002 -2604
rect 996 -2616 1002 -2610
rect 996 -2622 1002 -2616
rect 996 -2628 1002 -2622
rect 996 -2634 1002 -2628
rect 996 -2640 1002 -2634
rect 996 -2646 1002 -2640
rect 996 -2652 1002 -2646
rect 996 -2658 1002 -2652
rect 996 -2664 1002 -2658
rect 996 -2670 1002 -2664
rect 996 -2676 1002 -2670
rect 996 -2682 1002 -2676
rect 996 -2688 1002 -2682
rect 996 -2694 1002 -2688
rect 996 -2700 1002 -2694
rect 996 -2706 1002 -2700
rect 996 -2712 1002 -2706
rect 996 -2718 1002 -2712
rect 996 -2724 1002 -2718
rect 996 -2730 1002 -2724
rect 996 -2736 1002 -2730
rect 996 -2742 1002 -2736
rect 996 -2748 1002 -2742
rect 996 -2754 1002 -2748
rect 996 -2760 1002 -2754
rect 996 -2766 1002 -2760
rect 996 -2772 1002 -2766
rect 996 -2778 1002 -2772
rect 996 -2784 1002 -2778
rect 996 -2790 1002 -2784
rect 996 -2796 1002 -2790
rect 996 -2802 1002 -2796
rect 996 -2808 1002 -2802
rect 996 -2814 1002 -2808
rect 996 -2820 1002 -2814
rect 996 -2826 1002 -2820
rect 996 -2832 1002 -2826
rect 996 -2838 1002 -2832
rect 996 -2844 1002 -2838
rect 996 -2850 1002 -2844
rect 996 -2856 1002 -2850
rect 996 -2862 1002 -2856
rect 996 -2868 1002 -2862
rect 996 -2874 1002 -2868
rect 996 -2880 1002 -2874
rect 996 -2886 1002 -2880
rect 996 -2892 1002 -2886
rect 996 -2898 1002 -2892
rect 996 -2904 1002 -2898
rect 996 -2910 1002 -2904
rect 996 -2916 1002 -2910
rect 996 -2922 1002 -2916
rect 996 -2928 1002 -2922
rect 996 -2934 1002 -2928
rect 996 -2940 1002 -2934
rect 996 -3042 1002 -3036
rect 996 -3048 1002 -3042
rect 996 -3054 1002 -3048
rect 996 -3060 1002 -3054
rect 996 -3066 1002 -3060
rect 996 -3072 1002 -3066
rect 996 -3078 1002 -3072
rect 996 -3084 1002 -3078
rect 996 -3090 1002 -3084
rect 996 -3096 1002 -3090
rect 996 -3102 1002 -3096
rect 996 -3108 1002 -3102
rect 996 -3114 1002 -3108
rect 996 -3120 1002 -3114
rect 996 -3126 1002 -3120
rect 996 -3132 1002 -3126
rect 996 -3138 1002 -3132
rect 996 -3144 1002 -3138
rect 996 -3150 1002 -3144
rect 996 -3156 1002 -3150
rect 996 -3162 1002 -3156
rect 996 -3168 1002 -3162
rect 996 -3174 1002 -3168
rect 996 -3180 1002 -3174
rect 996 -3246 1002 -3240
rect 996 -3252 1002 -3246
rect 996 -3258 1002 -3252
rect 996 -3264 1002 -3258
rect 996 -3270 1002 -3264
rect 996 -3276 1002 -3270
rect 996 -3282 1002 -3276
rect 996 -3288 1002 -3282
rect 996 -3294 1002 -3288
rect 996 -3300 1002 -3294
rect 996 -3306 1002 -3300
rect 996 -3312 1002 -3306
rect 996 -3318 1002 -3312
rect 996 -3324 1002 -3318
rect 996 -3330 1002 -3324
rect 996 -3336 1002 -3330
rect 996 -3396 1002 -3390
rect 996 -3402 1002 -3396
rect 996 -3408 1002 -3402
rect 996 -3414 1002 -3408
rect 996 -3420 1002 -3414
rect 996 -3426 1002 -3420
rect 996 -3432 1002 -3426
rect 996 -3438 1002 -3432
rect 996 -3444 1002 -3438
rect 996 -3450 1002 -3444
rect 996 -3456 1002 -3450
rect 996 -3462 1002 -3456
rect 996 -3468 1002 -3462
rect 996 -3474 1002 -3468
rect 996 -3480 1002 -3474
rect 996 -3486 1002 -3480
rect 996 -3492 1002 -3486
rect 996 -3498 1002 -3492
rect 1002 -1122 1008 -1116
rect 1002 -1128 1008 -1122
rect 1002 -1134 1008 -1128
rect 1002 -1140 1008 -1134
rect 1002 -1146 1008 -1140
rect 1002 -1152 1008 -1146
rect 1002 -1158 1008 -1152
rect 1002 -1164 1008 -1158
rect 1002 -1170 1008 -1164
rect 1002 -1176 1008 -1170
rect 1002 -1182 1008 -1176
rect 1002 -1188 1008 -1182
rect 1002 -1194 1008 -1188
rect 1002 -1200 1008 -1194
rect 1002 -1206 1008 -1200
rect 1002 -1212 1008 -1206
rect 1002 -1218 1008 -1212
rect 1002 -1224 1008 -1218
rect 1002 -1230 1008 -1224
rect 1002 -1236 1008 -1230
rect 1002 -1242 1008 -1236
rect 1002 -1248 1008 -1242
rect 1002 -1254 1008 -1248
rect 1002 -1260 1008 -1254
rect 1002 -1266 1008 -1260
rect 1002 -1272 1008 -1266
rect 1002 -1278 1008 -1272
rect 1002 -1284 1008 -1278
rect 1002 -1290 1008 -1284
rect 1002 -1296 1008 -1290
rect 1002 -1302 1008 -1296
rect 1002 -1308 1008 -1302
rect 1002 -1314 1008 -1308
rect 1002 -1320 1008 -1314
rect 1002 -1326 1008 -1320
rect 1002 -2406 1008 -2400
rect 1002 -2412 1008 -2406
rect 1002 -2418 1008 -2412
rect 1002 -2424 1008 -2418
rect 1002 -2430 1008 -2424
rect 1002 -2436 1008 -2430
rect 1002 -2442 1008 -2436
rect 1002 -2448 1008 -2442
rect 1002 -2454 1008 -2448
rect 1002 -2460 1008 -2454
rect 1002 -2466 1008 -2460
rect 1002 -2472 1008 -2466
rect 1002 -2478 1008 -2472
rect 1002 -2484 1008 -2478
rect 1002 -2490 1008 -2484
rect 1002 -2496 1008 -2490
rect 1002 -2502 1008 -2496
rect 1002 -2508 1008 -2502
rect 1002 -2514 1008 -2508
rect 1002 -2520 1008 -2514
rect 1002 -2526 1008 -2520
rect 1002 -2532 1008 -2526
rect 1002 -2538 1008 -2532
rect 1002 -2544 1008 -2538
rect 1002 -2550 1008 -2544
rect 1002 -2556 1008 -2550
rect 1002 -2562 1008 -2556
rect 1002 -2568 1008 -2562
rect 1002 -2574 1008 -2568
rect 1002 -2580 1008 -2574
rect 1002 -2586 1008 -2580
rect 1002 -2592 1008 -2586
rect 1002 -2598 1008 -2592
rect 1002 -2604 1008 -2598
rect 1002 -2610 1008 -2604
rect 1002 -2616 1008 -2610
rect 1002 -2622 1008 -2616
rect 1002 -2628 1008 -2622
rect 1002 -2634 1008 -2628
rect 1002 -2640 1008 -2634
rect 1002 -2646 1008 -2640
rect 1002 -2652 1008 -2646
rect 1002 -2658 1008 -2652
rect 1002 -2664 1008 -2658
rect 1002 -2670 1008 -2664
rect 1002 -2676 1008 -2670
rect 1002 -2682 1008 -2676
rect 1002 -2688 1008 -2682
rect 1002 -2694 1008 -2688
rect 1002 -2700 1008 -2694
rect 1002 -2706 1008 -2700
rect 1002 -2712 1008 -2706
rect 1002 -2718 1008 -2712
rect 1002 -2724 1008 -2718
rect 1002 -2730 1008 -2724
rect 1002 -2736 1008 -2730
rect 1002 -2742 1008 -2736
rect 1002 -2748 1008 -2742
rect 1002 -2754 1008 -2748
rect 1002 -2760 1008 -2754
rect 1002 -2766 1008 -2760
rect 1002 -2772 1008 -2766
rect 1002 -2778 1008 -2772
rect 1002 -2784 1008 -2778
rect 1002 -2790 1008 -2784
rect 1002 -2796 1008 -2790
rect 1002 -2802 1008 -2796
rect 1002 -2808 1008 -2802
rect 1002 -2814 1008 -2808
rect 1002 -2820 1008 -2814
rect 1002 -2826 1008 -2820
rect 1002 -2832 1008 -2826
rect 1002 -2838 1008 -2832
rect 1002 -2844 1008 -2838
rect 1002 -2850 1008 -2844
rect 1002 -2856 1008 -2850
rect 1002 -2862 1008 -2856
rect 1002 -2868 1008 -2862
rect 1002 -2874 1008 -2868
rect 1002 -2880 1008 -2874
rect 1002 -2886 1008 -2880
rect 1002 -2892 1008 -2886
rect 1002 -2898 1008 -2892
rect 1002 -2904 1008 -2898
rect 1002 -2910 1008 -2904
rect 1002 -2916 1008 -2910
rect 1002 -2922 1008 -2916
rect 1002 -2928 1008 -2922
rect 1002 -2934 1008 -2928
rect 1002 -3030 1008 -3024
rect 1002 -3036 1008 -3030
rect 1002 -3042 1008 -3036
rect 1002 -3048 1008 -3042
rect 1002 -3054 1008 -3048
rect 1002 -3060 1008 -3054
rect 1002 -3066 1008 -3060
rect 1002 -3072 1008 -3066
rect 1002 -3078 1008 -3072
rect 1002 -3084 1008 -3078
rect 1002 -3090 1008 -3084
rect 1002 -3096 1008 -3090
rect 1002 -3102 1008 -3096
rect 1002 -3108 1008 -3102
rect 1002 -3114 1008 -3108
rect 1002 -3120 1008 -3114
rect 1002 -3126 1008 -3120
rect 1002 -3132 1008 -3126
rect 1002 -3138 1008 -3132
rect 1002 -3144 1008 -3138
rect 1002 -3150 1008 -3144
rect 1002 -3156 1008 -3150
rect 1002 -3162 1008 -3156
rect 1002 -3168 1008 -3162
rect 1002 -3174 1008 -3168
rect 1002 -3240 1008 -3234
rect 1002 -3246 1008 -3240
rect 1002 -3252 1008 -3246
rect 1002 -3258 1008 -3252
rect 1002 -3264 1008 -3258
rect 1002 -3270 1008 -3264
rect 1002 -3276 1008 -3270
rect 1002 -3282 1008 -3276
rect 1002 -3288 1008 -3282
rect 1002 -3294 1008 -3288
rect 1002 -3300 1008 -3294
rect 1002 -3306 1008 -3300
rect 1002 -3312 1008 -3306
rect 1002 -3318 1008 -3312
rect 1002 -3324 1008 -3318
rect 1002 -3330 1008 -3324
rect 1002 -3390 1008 -3384
rect 1002 -3396 1008 -3390
rect 1002 -3402 1008 -3396
rect 1002 -3408 1008 -3402
rect 1002 -3414 1008 -3408
rect 1002 -3420 1008 -3414
rect 1002 -3426 1008 -3420
rect 1002 -3432 1008 -3426
rect 1002 -3438 1008 -3432
rect 1002 -3444 1008 -3438
rect 1002 -3450 1008 -3444
rect 1002 -3456 1008 -3450
rect 1002 -3462 1008 -3456
rect 1002 -3468 1008 -3462
rect 1002 -3474 1008 -3468
rect 1002 -3480 1008 -3474
rect 1002 -3486 1008 -3480
rect 1002 -3492 1008 -3486
rect 1002 -3498 1008 -3492
rect 1008 -1122 1014 -1116
rect 1008 -1128 1014 -1122
rect 1008 -1134 1014 -1128
rect 1008 -1140 1014 -1134
rect 1008 -1146 1014 -1140
rect 1008 -1152 1014 -1146
rect 1008 -1158 1014 -1152
rect 1008 -1164 1014 -1158
rect 1008 -1170 1014 -1164
rect 1008 -1176 1014 -1170
rect 1008 -1182 1014 -1176
rect 1008 -1188 1014 -1182
rect 1008 -1194 1014 -1188
rect 1008 -1200 1014 -1194
rect 1008 -1206 1014 -1200
rect 1008 -1212 1014 -1206
rect 1008 -1218 1014 -1212
rect 1008 -1224 1014 -1218
rect 1008 -1230 1014 -1224
rect 1008 -1236 1014 -1230
rect 1008 -1242 1014 -1236
rect 1008 -1248 1014 -1242
rect 1008 -1254 1014 -1248
rect 1008 -1260 1014 -1254
rect 1008 -1266 1014 -1260
rect 1008 -1272 1014 -1266
rect 1008 -1278 1014 -1272
rect 1008 -1284 1014 -1278
rect 1008 -1290 1014 -1284
rect 1008 -1296 1014 -1290
rect 1008 -1302 1014 -1296
rect 1008 -1308 1014 -1302
rect 1008 -1314 1014 -1308
rect 1008 -1320 1014 -1314
rect 1008 -1326 1014 -1320
rect 1008 -2388 1014 -2382
rect 1008 -2394 1014 -2388
rect 1008 -2400 1014 -2394
rect 1008 -2406 1014 -2400
rect 1008 -2412 1014 -2406
rect 1008 -2418 1014 -2412
rect 1008 -2424 1014 -2418
rect 1008 -2430 1014 -2424
rect 1008 -2436 1014 -2430
rect 1008 -2442 1014 -2436
rect 1008 -2448 1014 -2442
rect 1008 -2454 1014 -2448
rect 1008 -2460 1014 -2454
rect 1008 -2466 1014 -2460
rect 1008 -2472 1014 -2466
rect 1008 -2478 1014 -2472
rect 1008 -2484 1014 -2478
rect 1008 -2490 1014 -2484
rect 1008 -2496 1014 -2490
rect 1008 -2502 1014 -2496
rect 1008 -2508 1014 -2502
rect 1008 -2514 1014 -2508
rect 1008 -2520 1014 -2514
rect 1008 -2526 1014 -2520
rect 1008 -2532 1014 -2526
rect 1008 -2538 1014 -2532
rect 1008 -2544 1014 -2538
rect 1008 -2550 1014 -2544
rect 1008 -2556 1014 -2550
rect 1008 -2562 1014 -2556
rect 1008 -2568 1014 -2562
rect 1008 -2574 1014 -2568
rect 1008 -2580 1014 -2574
rect 1008 -2586 1014 -2580
rect 1008 -2592 1014 -2586
rect 1008 -2598 1014 -2592
rect 1008 -2604 1014 -2598
rect 1008 -2610 1014 -2604
rect 1008 -2616 1014 -2610
rect 1008 -2622 1014 -2616
rect 1008 -2628 1014 -2622
rect 1008 -2634 1014 -2628
rect 1008 -2640 1014 -2634
rect 1008 -2646 1014 -2640
rect 1008 -2652 1014 -2646
rect 1008 -2658 1014 -2652
rect 1008 -2664 1014 -2658
rect 1008 -2670 1014 -2664
rect 1008 -2676 1014 -2670
rect 1008 -2682 1014 -2676
rect 1008 -2688 1014 -2682
rect 1008 -2694 1014 -2688
rect 1008 -2700 1014 -2694
rect 1008 -2706 1014 -2700
rect 1008 -2712 1014 -2706
rect 1008 -2718 1014 -2712
rect 1008 -2724 1014 -2718
rect 1008 -2730 1014 -2724
rect 1008 -2736 1014 -2730
rect 1008 -2742 1014 -2736
rect 1008 -2748 1014 -2742
rect 1008 -2754 1014 -2748
rect 1008 -2760 1014 -2754
rect 1008 -2766 1014 -2760
rect 1008 -2772 1014 -2766
rect 1008 -2778 1014 -2772
rect 1008 -2784 1014 -2778
rect 1008 -2790 1014 -2784
rect 1008 -2796 1014 -2790
rect 1008 -2802 1014 -2796
rect 1008 -2808 1014 -2802
rect 1008 -2814 1014 -2808
rect 1008 -2820 1014 -2814
rect 1008 -2826 1014 -2820
rect 1008 -2832 1014 -2826
rect 1008 -2838 1014 -2832
rect 1008 -2844 1014 -2838
rect 1008 -2850 1014 -2844
rect 1008 -2856 1014 -2850
rect 1008 -2862 1014 -2856
rect 1008 -2868 1014 -2862
rect 1008 -2874 1014 -2868
rect 1008 -2880 1014 -2874
rect 1008 -2886 1014 -2880
rect 1008 -2892 1014 -2886
rect 1008 -2898 1014 -2892
rect 1008 -2904 1014 -2898
rect 1008 -2910 1014 -2904
rect 1008 -2916 1014 -2910
rect 1008 -2922 1014 -2916
rect 1008 -3018 1014 -3012
rect 1008 -3024 1014 -3018
rect 1008 -3030 1014 -3024
rect 1008 -3036 1014 -3030
rect 1008 -3042 1014 -3036
rect 1008 -3048 1014 -3042
rect 1008 -3054 1014 -3048
rect 1008 -3060 1014 -3054
rect 1008 -3066 1014 -3060
rect 1008 -3072 1014 -3066
rect 1008 -3078 1014 -3072
rect 1008 -3084 1014 -3078
rect 1008 -3090 1014 -3084
rect 1008 -3096 1014 -3090
rect 1008 -3102 1014 -3096
rect 1008 -3108 1014 -3102
rect 1008 -3114 1014 -3108
rect 1008 -3120 1014 -3114
rect 1008 -3126 1014 -3120
rect 1008 -3132 1014 -3126
rect 1008 -3138 1014 -3132
rect 1008 -3144 1014 -3138
rect 1008 -3150 1014 -3144
rect 1008 -3156 1014 -3150
rect 1008 -3162 1014 -3156
rect 1008 -3168 1014 -3162
rect 1008 -3234 1014 -3228
rect 1008 -3240 1014 -3234
rect 1008 -3246 1014 -3240
rect 1008 -3252 1014 -3246
rect 1008 -3258 1014 -3252
rect 1008 -3264 1014 -3258
rect 1008 -3270 1014 -3264
rect 1008 -3276 1014 -3270
rect 1008 -3282 1014 -3276
rect 1008 -3288 1014 -3282
rect 1008 -3294 1014 -3288
rect 1008 -3300 1014 -3294
rect 1008 -3306 1014 -3300
rect 1008 -3312 1014 -3306
rect 1008 -3318 1014 -3312
rect 1008 -3324 1014 -3318
rect 1008 -3330 1014 -3324
rect 1008 -3390 1014 -3384
rect 1008 -3396 1014 -3390
rect 1008 -3402 1014 -3396
rect 1008 -3408 1014 -3402
rect 1008 -3414 1014 -3408
rect 1008 -3420 1014 -3414
rect 1008 -3426 1014 -3420
rect 1008 -3432 1014 -3426
rect 1008 -3438 1014 -3432
rect 1008 -3444 1014 -3438
rect 1008 -3450 1014 -3444
rect 1008 -3456 1014 -3450
rect 1008 -3462 1014 -3456
rect 1008 -3468 1014 -3462
rect 1008 -3474 1014 -3468
rect 1008 -3480 1014 -3474
rect 1008 -3486 1014 -3480
rect 1008 -3492 1014 -3486
rect 1008 -3498 1014 -3492
rect 1014 -1122 1020 -1116
rect 1014 -1128 1020 -1122
rect 1014 -1134 1020 -1128
rect 1014 -1140 1020 -1134
rect 1014 -1146 1020 -1140
rect 1014 -1152 1020 -1146
rect 1014 -1158 1020 -1152
rect 1014 -1164 1020 -1158
rect 1014 -1170 1020 -1164
rect 1014 -1176 1020 -1170
rect 1014 -1182 1020 -1176
rect 1014 -1188 1020 -1182
rect 1014 -1194 1020 -1188
rect 1014 -1200 1020 -1194
rect 1014 -1206 1020 -1200
rect 1014 -1212 1020 -1206
rect 1014 -1218 1020 -1212
rect 1014 -1224 1020 -1218
rect 1014 -1230 1020 -1224
rect 1014 -1236 1020 -1230
rect 1014 -1242 1020 -1236
rect 1014 -1248 1020 -1242
rect 1014 -1254 1020 -1248
rect 1014 -1260 1020 -1254
rect 1014 -1266 1020 -1260
rect 1014 -1272 1020 -1266
rect 1014 -1278 1020 -1272
rect 1014 -1284 1020 -1278
rect 1014 -1290 1020 -1284
rect 1014 -1296 1020 -1290
rect 1014 -1302 1020 -1296
rect 1014 -1308 1020 -1302
rect 1014 -1314 1020 -1308
rect 1014 -1320 1020 -1314
rect 1014 -1326 1020 -1320
rect 1014 -2364 1020 -2358
rect 1014 -2370 1020 -2364
rect 1014 -2376 1020 -2370
rect 1014 -2382 1020 -2376
rect 1014 -2388 1020 -2382
rect 1014 -2394 1020 -2388
rect 1014 -2400 1020 -2394
rect 1014 -2406 1020 -2400
rect 1014 -2412 1020 -2406
rect 1014 -2418 1020 -2412
rect 1014 -2424 1020 -2418
rect 1014 -2430 1020 -2424
rect 1014 -2436 1020 -2430
rect 1014 -2442 1020 -2436
rect 1014 -2448 1020 -2442
rect 1014 -2454 1020 -2448
rect 1014 -2460 1020 -2454
rect 1014 -2466 1020 -2460
rect 1014 -2472 1020 -2466
rect 1014 -2478 1020 -2472
rect 1014 -2484 1020 -2478
rect 1014 -2490 1020 -2484
rect 1014 -2496 1020 -2490
rect 1014 -2502 1020 -2496
rect 1014 -2508 1020 -2502
rect 1014 -2514 1020 -2508
rect 1014 -2520 1020 -2514
rect 1014 -2526 1020 -2520
rect 1014 -2532 1020 -2526
rect 1014 -2538 1020 -2532
rect 1014 -2544 1020 -2538
rect 1014 -2550 1020 -2544
rect 1014 -2556 1020 -2550
rect 1014 -2562 1020 -2556
rect 1014 -2568 1020 -2562
rect 1014 -2574 1020 -2568
rect 1014 -2580 1020 -2574
rect 1014 -2586 1020 -2580
rect 1014 -2592 1020 -2586
rect 1014 -2598 1020 -2592
rect 1014 -2604 1020 -2598
rect 1014 -2610 1020 -2604
rect 1014 -2616 1020 -2610
rect 1014 -2622 1020 -2616
rect 1014 -2628 1020 -2622
rect 1014 -2634 1020 -2628
rect 1014 -2640 1020 -2634
rect 1014 -2646 1020 -2640
rect 1014 -2652 1020 -2646
rect 1014 -2658 1020 -2652
rect 1014 -2664 1020 -2658
rect 1014 -2670 1020 -2664
rect 1014 -2676 1020 -2670
rect 1014 -2682 1020 -2676
rect 1014 -2688 1020 -2682
rect 1014 -2694 1020 -2688
rect 1014 -2700 1020 -2694
rect 1014 -2706 1020 -2700
rect 1014 -2712 1020 -2706
rect 1014 -2718 1020 -2712
rect 1014 -2724 1020 -2718
rect 1014 -2730 1020 -2724
rect 1014 -2736 1020 -2730
rect 1014 -2742 1020 -2736
rect 1014 -2748 1020 -2742
rect 1014 -2754 1020 -2748
rect 1014 -2760 1020 -2754
rect 1014 -2766 1020 -2760
rect 1014 -2772 1020 -2766
rect 1014 -2778 1020 -2772
rect 1014 -2784 1020 -2778
rect 1014 -2790 1020 -2784
rect 1014 -2796 1020 -2790
rect 1014 -2802 1020 -2796
rect 1014 -2808 1020 -2802
rect 1014 -2814 1020 -2808
rect 1014 -2820 1020 -2814
rect 1014 -2826 1020 -2820
rect 1014 -2832 1020 -2826
rect 1014 -2838 1020 -2832
rect 1014 -2844 1020 -2838
rect 1014 -2850 1020 -2844
rect 1014 -2856 1020 -2850
rect 1014 -2862 1020 -2856
rect 1014 -2868 1020 -2862
rect 1014 -2874 1020 -2868
rect 1014 -2880 1020 -2874
rect 1014 -2886 1020 -2880
rect 1014 -2892 1020 -2886
rect 1014 -2898 1020 -2892
rect 1014 -2904 1020 -2898
rect 1014 -2910 1020 -2904
rect 1014 -3012 1020 -3006
rect 1014 -3018 1020 -3012
rect 1014 -3024 1020 -3018
rect 1014 -3030 1020 -3024
rect 1014 -3036 1020 -3030
rect 1014 -3042 1020 -3036
rect 1014 -3048 1020 -3042
rect 1014 -3054 1020 -3048
rect 1014 -3060 1020 -3054
rect 1014 -3066 1020 -3060
rect 1014 -3072 1020 -3066
rect 1014 -3078 1020 -3072
rect 1014 -3084 1020 -3078
rect 1014 -3090 1020 -3084
rect 1014 -3096 1020 -3090
rect 1014 -3102 1020 -3096
rect 1014 -3108 1020 -3102
rect 1014 -3114 1020 -3108
rect 1014 -3120 1020 -3114
rect 1014 -3126 1020 -3120
rect 1014 -3132 1020 -3126
rect 1014 -3138 1020 -3132
rect 1014 -3144 1020 -3138
rect 1014 -3150 1020 -3144
rect 1014 -3156 1020 -3150
rect 1014 -3162 1020 -3156
rect 1014 -3168 1020 -3162
rect 1014 -3234 1020 -3228
rect 1014 -3240 1020 -3234
rect 1014 -3246 1020 -3240
rect 1014 -3252 1020 -3246
rect 1014 -3258 1020 -3252
rect 1014 -3264 1020 -3258
rect 1014 -3270 1020 -3264
rect 1014 -3276 1020 -3270
rect 1014 -3282 1020 -3276
rect 1014 -3288 1020 -3282
rect 1014 -3294 1020 -3288
rect 1014 -3300 1020 -3294
rect 1014 -3306 1020 -3300
rect 1014 -3312 1020 -3306
rect 1014 -3318 1020 -3312
rect 1014 -3324 1020 -3318
rect 1014 -3384 1020 -3378
rect 1014 -3390 1020 -3384
rect 1014 -3396 1020 -3390
rect 1014 -3402 1020 -3396
rect 1014 -3408 1020 -3402
rect 1014 -3414 1020 -3408
rect 1014 -3420 1020 -3414
rect 1014 -3426 1020 -3420
rect 1014 -3432 1020 -3426
rect 1014 -3438 1020 -3432
rect 1014 -3444 1020 -3438
rect 1014 -3450 1020 -3444
rect 1014 -3456 1020 -3450
rect 1014 -3462 1020 -3456
rect 1014 -3468 1020 -3462
rect 1014 -3474 1020 -3468
rect 1014 -3480 1020 -3474
rect 1014 -3486 1020 -3480
rect 1014 -3492 1020 -3486
rect 1014 -3498 1020 -3492
rect 1020 -1116 1026 -1110
rect 1020 -1122 1026 -1116
rect 1020 -1128 1026 -1122
rect 1020 -1134 1026 -1128
rect 1020 -1140 1026 -1134
rect 1020 -1146 1026 -1140
rect 1020 -1152 1026 -1146
rect 1020 -1158 1026 -1152
rect 1020 -1164 1026 -1158
rect 1020 -1170 1026 -1164
rect 1020 -1176 1026 -1170
rect 1020 -1182 1026 -1176
rect 1020 -1188 1026 -1182
rect 1020 -1194 1026 -1188
rect 1020 -1200 1026 -1194
rect 1020 -1206 1026 -1200
rect 1020 -1212 1026 -1206
rect 1020 -1218 1026 -1212
rect 1020 -1224 1026 -1218
rect 1020 -1230 1026 -1224
rect 1020 -1236 1026 -1230
rect 1020 -1242 1026 -1236
rect 1020 -1248 1026 -1242
rect 1020 -1254 1026 -1248
rect 1020 -1260 1026 -1254
rect 1020 -1266 1026 -1260
rect 1020 -1272 1026 -1266
rect 1020 -1278 1026 -1272
rect 1020 -1284 1026 -1278
rect 1020 -1290 1026 -1284
rect 1020 -1296 1026 -1290
rect 1020 -1302 1026 -1296
rect 1020 -1308 1026 -1302
rect 1020 -1314 1026 -1308
rect 1020 -1320 1026 -1314
rect 1020 -1326 1026 -1320
rect 1020 -2346 1026 -2340
rect 1020 -2352 1026 -2346
rect 1020 -2358 1026 -2352
rect 1020 -2364 1026 -2358
rect 1020 -2370 1026 -2364
rect 1020 -2376 1026 -2370
rect 1020 -2382 1026 -2376
rect 1020 -2388 1026 -2382
rect 1020 -2394 1026 -2388
rect 1020 -2400 1026 -2394
rect 1020 -2406 1026 -2400
rect 1020 -2412 1026 -2406
rect 1020 -2418 1026 -2412
rect 1020 -2424 1026 -2418
rect 1020 -2430 1026 -2424
rect 1020 -2436 1026 -2430
rect 1020 -2442 1026 -2436
rect 1020 -2448 1026 -2442
rect 1020 -2454 1026 -2448
rect 1020 -2460 1026 -2454
rect 1020 -2466 1026 -2460
rect 1020 -2472 1026 -2466
rect 1020 -2478 1026 -2472
rect 1020 -2484 1026 -2478
rect 1020 -2490 1026 -2484
rect 1020 -2496 1026 -2490
rect 1020 -2502 1026 -2496
rect 1020 -2508 1026 -2502
rect 1020 -2514 1026 -2508
rect 1020 -2520 1026 -2514
rect 1020 -2526 1026 -2520
rect 1020 -2532 1026 -2526
rect 1020 -2538 1026 -2532
rect 1020 -2544 1026 -2538
rect 1020 -2550 1026 -2544
rect 1020 -2556 1026 -2550
rect 1020 -2562 1026 -2556
rect 1020 -2568 1026 -2562
rect 1020 -2574 1026 -2568
rect 1020 -2580 1026 -2574
rect 1020 -2586 1026 -2580
rect 1020 -2592 1026 -2586
rect 1020 -2598 1026 -2592
rect 1020 -2604 1026 -2598
rect 1020 -2610 1026 -2604
rect 1020 -2616 1026 -2610
rect 1020 -2622 1026 -2616
rect 1020 -2628 1026 -2622
rect 1020 -2634 1026 -2628
rect 1020 -2640 1026 -2634
rect 1020 -2646 1026 -2640
rect 1020 -2652 1026 -2646
rect 1020 -2658 1026 -2652
rect 1020 -2664 1026 -2658
rect 1020 -2670 1026 -2664
rect 1020 -2676 1026 -2670
rect 1020 -2682 1026 -2676
rect 1020 -2688 1026 -2682
rect 1020 -2694 1026 -2688
rect 1020 -2700 1026 -2694
rect 1020 -2706 1026 -2700
rect 1020 -2712 1026 -2706
rect 1020 -2718 1026 -2712
rect 1020 -2724 1026 -2718
rect 1020 -2730 1026 -2724
rect 1020 -2736 1026 -2730
rect 1020 -2742 1026 -2736
rect 1020 -2748 1026 -2742
rect 1020 -2754 1026 -2748
rect 1020 -2760 1026 -2754
rect 1020 -2766 1026 -2760
rect 1020 -2772 1026 -2766
rect 1020 -2778 1026 -2772
rect 1020 -2784 1026 -2778
rect 1020 -2790 1026 -2784
rect 1020 -2796 1026 -2790
rect 1020 -2802 1026 -2796
rect 1020 -2808 1026 -2802
rect 1020 -2814 1026 -2808
rect 1020 -2820 1026 -2814
rect 1020 -2826 1026 -2820
rect 1020 -2832 1026 -2826
rect 1020 -2838 1026 -2832
rect 1020 -2844 1026 -2838
rect 1020 -2850 1026 -2844
rect 1020 -2856 1026 -2850
rect 1020 -2862 1026 -2856
rect 1020 -2868 1026 -2862
rect 1020 -2874 1026 -2868
rect 1020 -2880 1026 -2874
rect 1020 -2886 1026 -2880
rect 1020 -2892 1026 -2886
rect 1020 -2898 1026 -2892
rect 1020 -3000 1026 -2994
rect 1020 -3006 1026 -3000
rect 1020 -3012 1026 -3006
rect 1020 -3018 1026 -3012
rect 1020 -3024 1026 -3018
rect 1020 -3030 1026 -3024
rect 1020 -3036 1026 -3030
rect 1020 -3042 1026 -3036
rect 1020 -3048 1026 -3042
rect 1020 -3054 1026 -3048
rect 1020 -3060 1026 -3054
rect 1020 -3066 1026 -3060
rect 1020 -3072 1026 -3066
rect 1020 -3078 1026 -3072
rect 1020 -3084 1026 -3078
rect 1020 -3090 1026 -3084
rect 1020 -3096 1026 -3090
rect 1020 -3102 1026 -3096
rect 1020 -3108 1026 -3102
rect 1020 -3114 1026 -3108
rect 1020 -3120 1026 -3114
rect 1020 -3126 1026 -3120
rect 1020 -3132 1026 -3126
rect 1020 -3138 1026 -3132
rect 1020 -3144 1026 -3138
rect 1020 -3150 1026 -3144
rect 1020 -3156 1026 -3150
rect 1020 -3162 1026 -3156
rect 1020 -3228 1026 -3222
rect 1020 -3234 1026 -3228
rect 1020 -3240 1026 -3234
rect 1020 -3246 1026 -3240
rect 1020 -3252 1026 -3246
rect 1020 -3258 1026 -3252
rect 1020 -3264 1026 -3258
rect 1020 -3270 1026 -3264
rect 1020 -3276 1026 -3270
rect 1020 -3282 1026 -3276
rect 1020 -3288 1026 -3282
rect 1020 -3294 1026 -3288
rect 1020 -3300 1026 -3294
rect 1020 -3306 1026 -3300
rect 1020 -3312 1026 -3306
rect 1020 -3318 1026 -3312
rect 1020 -3378 1026 -3372
rect 1020 -3384 1026 -3378
rect 1020 -3390 1026 -3384
rect 1020 -3396 1026 -3390
rect 1020 -3402 1026 -3396
rect 1020 -3408 1026 -3402
rect 1020 -3414 1026 -3408
rect 1020 -3420 1026 -3414
rect 1020 -3426 1026 -3420
rect 1020 -3432 1026 -3426
rect 1020 -3438 1026 -3432
rect 1020 -3444 1026 -3438
rect 1020 -3450 1026 -3444
rect 1020 -3456 1026 -3450
rect 1020 -3462 1026 -3456
rect 1020 -3468 1026 -3462
rect 1020 -3474 1026 -3468
rect 1020 -3480 1026 -3474
rect 1020 -3486 1026 -3480
rect 1020 -3492 1026 -3486
rect 1020 -3498 1026 -3492
rect 1026 -1116 1032 -1110
rect 1026 -1122 1032 -1116
rect 1026 -1128 1032 -1122
rect 1026 -1134 1032 -1128
rect 1026 -1140 1032 -1134
rect 1026 -1146 1032 -1140
rect 1026 -1152 1032 -1146
rect 1026 -1158 1032 -1152
rect 1026 -1164 1032 -1158
rect 1026 -1170 1032 -1164
rect 1026 -1176 1032 -1170
rect 1026 -1182 1032 -1176
rect 1026 -1188 1032 -1182
rect 1026 -1194 1032 -1188
rect 1026 -1200 1032 -1194
rect 1026 -1206 1032 -1200
rect 1026 -1212 1032 -1206
rect 1026 -1218 1032 -1212
rect 1026 -1224 1032 -1218
rect 1026 -1230 1032 -1224
rect 1026 -1236 1032 -1230
rect 1026 -1242 1032 -1236
rect 1026 -1248 1032 -1242
rect 1026 -1254 1032 -1248
rect 1026 -1260 1032 -1254
rect 1026 -1266 1032 -1260
rect 1026 -1272 1032 -1266
rect 1026 -1278 1032 -1272
rect 1026 -1284 1032 -1278
rect 1026 -1290 1032 -1284
rect 1026 -1296 1032 -1290
rect 1026 -1302 1032 -1296
rect 1026 -1308 1032 -1302
rect 1026 -1314 1032 -1308
rect 1026 -1320 1032 -1314
rect 1026 -1326 1032 -1320
rect 1026 -2322 1032 -2316
rect 1026 -2328 1032 -2322
rect 1026 -2334 1032 -2328
rect 1026 -2340 1032 -2334
rect 1026 -2346 1032 -2340
rect 1026 -2352 1032 -2346
rect 1026 -2358 1032 -2352
rect 1026 -2364 1032 -2358
rect 1026 -2370 1032 -2364
rect 1026 -2376 1032 -2370
rect 1026 -2382 1032 -2376
rect 1026 -2388 1032 -2382
rect 1026 -2394 1032 -2388
rect 1026 -2400 1032 -2394
rect 1026 -2406 1032 -2400
rect 1026 -2412 1032 -2406
rect 1026 -2418 1032 -2412
rect 1026 -2424 1032 -2418
rect 1026 -2430 1032 -2424
rect 1026 -2436 1032 -2430
rect 1026 -2442 1032 -2436
rect 1026 -2448 1032 -2442
rect 1026 -2454 1032 -2448
rect 1026 -2460 1032 -2454
rect 1026 -2466 1032 -2460
rect 1026 -2472 1032 -2466
rect 1026 -2478 1032 -2472
rect 1026 -2484 1032 -2478
rect 1026 -2490 1032 -2484
rect 1026 -2496 1032 -2490
rect 1026 -2502 1032 -2496
rect 1026 -2508 1032 -2502
rect 1026 -2514 1032 -2508
rect 1026 -2520 1032 -2514
rect 1026 -2526 1032 -2520
rect 1026 -2532 1032 -2526
rect 1026 -2538 1032 -2532
rect 1026 -2544 1032 -2538
rect 1026 -2550 1032 -2544
rect 1026 -2556 1032 -2550
rect 1026 -2562 1032 -2556
rect 1026 -2568 1032 -2562
rect 1026 -2574 1032 -2568
rect 1026 -2580 1032 -2574
rect 1026 -2586 1032 -2580
rect 1026 -2592 1032 -2586
rect 1026 -2598 1032 -2592
rect 1026 -2604 1032 -2598
rect 1026 -2610 1032 -2604
rect 1026 -2616 1032 -2610
rect 1026 -2622 1032 -2616
rect 1026 -2628 1032 -2622
rect 1026 -2634 1032 -2628
rect 1026 -2640 1032 -2634
rect 1026 -2646 1032 -2640
rect 1026 -2652 1032 -2646
rect 1026 -2658 1032 -2652
rect 1026 -2664 1032 -2658
rect 1026 -2670 1032 -2664
rect 1026 -2676 1032 -2670
rect 1026 -2682 1032 -2676
rect 1026 -2688 1032 -2682
rect 1026 -2694 1032 -2688
rect 1026 -2700 1032 -2694
rect 1026 -2706 1032 -2700
rect 1026 -2712 1032 -2706
rect 1026 -2718 1032 -2712
rect 1026 -2724 1032 -2718
rect 1026 -2730 1032 -2724
rect 1026 -2736 1032 -2730
rect 1026 -2742 1032 -2736
rect 1026 -2748 1032 -2742
rect 1026 -2754 1032 -2748
rect 1026 -2760 1032 -2754
rect 1026 -2766 1032 -2760
rect 1026 -2772 1032 -2766
rect 1026 -2778 1032 -2772
rect 1026 -2784 1032 -2778
rect 1026 -2790 1032 -2784
rect 1026 -2796 1032 -2790
rect 1026 -2802 1032 -2796
rect 1026 -2808 1032 -2802
rect 1026 -2814 1032 -2808
rect 1026 -2820 1032 -2814
rect 1026 -2826 1032 -2820
rect 1026 -2832 1032 -2826
rect 1026 -2838 1032 -2832
rect 1026 -2844 1032 -2838
rect 1026 -2850 1032 -2844
rect 1026 -2856 1032 -2850
rect 1026 -2862 1032 -2856
rect 1026 -2868 1032 -2862
rect 1026 -2874 1032 -2868
rect 1026 -2880 1032 -2874
rect 1026 -2886 1032 -2880
rect 1026 -2988 1032 -2982
rect 1026 -2994 1032 -2988
rect 1026 -3000 1032 -2994
rect 1026 -3006 1032 -3000
rect 1026 -3012 1032 -3006
rect 1026 -3018 1032 -3012
rect 1026 -3024 1032 -3018
rect 1026 -3030 1032 -3024
rect 1026 -3036 1032 -3030
rect 1026 -3042 1032 -3036
rect 1026 -3048 1032 -3042
rect 1026 -3054 1032 -3048
rect 1026 -3060 1032 -3054
rect 1026 -3066 1032 -3060
rect 1026 -3072 1032 -3066
rect 1026 -3078 1032 -3072
rect 1026 -3084 1032 -3078
rect 1026 -3090 1032 -3084
rect 1026 -3096 1032 -3090
rect 1026 -3102 1032 -3096
rect 1026 -3108 1032 -3102
rect 1026 -3114 1032 -3108
rect 1026 -3120 1032 -3114
rect 1026 -3126 1032 -3120
rect 1026 -3132 1032 -3126
rect 1026 -3138 1032 -3132
rect 1026 -3144 1032 -3138
rect 1026 -3150 1032 -3144
rect 1026 -3156 1032 -3150
rect 1026 -3222 1032 -3216
rect 1026 -3228 1032 -3222
rect 1026 -3234 1032 -3228
rect 1026 -3240 1032 -3234
rect 1026 -3246 1032 -3240
rect 1026 -3252 1032 -3246
rect 1026 -3258 1032 -3252
rect 1026 -3264 1032 -3258
rect 1026 -3270 1032 -3264
rect 1026 -3276 1032 -3270
rect 1026 -3282 1032 -3276
rect 1026 -3288 1032 -3282
rect 1026 -3294 1032 -3288
rect 1026 -3300 1032 -3294
rect 1026 -3306 1032 -3300
rect 1026 -3312 1032 -3306
rect 1026 -3318 1032 -3312
rect 1026 -3372 1032 -3366
rect 1026 -3378 1032 -3372
rect 1026 -3384 1032 -3378
rect 1026 -3390 1032 -3384
rect 1026 -3396 1032 -3390
rect 1026 -3402 1032 -3396
rect 1026 -3408 1032 -3402
rect 1026 -3414 1032 -3408
rect 1026 -3420 1032 -3414
rect 1026 -3426 1032 -3420
rect 1026 -3432 1032 -3426
rect 1026 -3438 1032 -3432
rect 1026 -3444 1032 -3438
rect 1026 -3450 1032 -3444
rect 1026 -3456 1032 -3450
rect 1026 -3462 1032 -3456
rect 1026 -3468 1032 -3462
rect 1026 -3474 1032 -3468
rect 1026 -3480 1032 -3474
rect 1026 -3486 1032 -3480
rect 1026 -3492 1032 -3486
rect 1026 -3498 1032 -3492
rect 1032 -1116 1038 -1110
rect 1032 -1122 1038 -1116
rect 1032 -1128 1038 -1122
rect 1032 -1134 1038 -1128
rect 1032 -1140 1038 -1134
rect 1032 -1146 1038 -1140
rect 1032 -1152 1038 -1146
rect 1032 -1158 1038 -1152
rect 1032 -1164 1038 -1158
rect 1032 -1170 1038 -1164
rect 1032 -1176 1038 -1170
rect 1032 -1182 1038 -1176
rect 1032 -1188 1038 -1182
rect 1032 -1194 1038 -1188
rect 1032 -1200 1038 -1194
rect 1032 -1206 1038 -1200
rect 1032 -1212 1038 -1206
rect 1032 -1218 1038 -1212
rect 1032 -1224 1038 -1218
rect 1032 -1230 1038 -1224
rect 1032 -1236 1038 -1230
rect 1032 -1242 1038 -1236
rect 1032 -1248 1038 -1242
rect 1032 -1254 1038 -1248
rect 1032 -1260 1038 -1254
rect 1032 -1266 1038 -1260
rect 1032 -1272 1038 -1266
rect 1032 -1278 1038 -1272
rect 1032 -1284 1038 -1278
rect 1032 -1290 1038 -1284
rect 1032 -1296 1038 -1290
rect 1032 -1302 1038 -1296
rect 1032 -1308 1038 -1302
rect 1032 -1314 1038 -1308
rect 1032 -1320 1038 -1314
rect 1032 -2304 1038 -2298
rect 1032 -2310 1038 -2304
rect 1032 -2316 1038 -2310
rect 1032 -2322 1038 -2316
rect 1032 -2328 1038 -2322
rect 1032 -2334 1038 -2328
rect 1032 -2340 1038 -2334
rect 1032 -2346 1038 -2340
rect 1032 -2352 1038 -2346
rect 1032 -2358 1038 -2352
rect 1032 -2364 1038 -2358
rect 1032 -2370 1038 -2364
rect 1032 -2376 1038 -2370
rect 1032 -2382 1038 -2376
rect 1032 -2388 1038 -2382
rect 1032 -2394 1038 -2388
rect 1032 -2400 1038 -2394
rect 1032 -2406 1038 -2400
rect 1032 -2412 1038 -2406
rect 1032 -2418 1038 -2412
rect 1032 -2424 1038 -2418
rect 1032 -2430 1038 -2424
rect 1032 -2436 1038 -2430
rect 1032 -2442 1038 -2436
rect 1032 -2448 1038 -2442
rect 1032 -2454 1038 -2448
rect 1032 -2460 1038 -2454
rect 1032 -2466 1038 -2460
rect 1032 -2472 1038 -2466
rect 1032 -2478 1038 -2472
rect 1032 -2484 1038 -2478
rect 1032 -2490 1038 -2484
rect 1032 -2496 1038 -2490
rect 1032 -2502 1038 -2496
rect 1032 -2508 1038 -2502
rect 1032 -2514 1038 -2508
rect 1032 -2520 1038 -2514
rect 1032 -2526 1038 -2520
rect 1032 -2532 1038 -2526
rect 1032 -2538 1038 -2532
rect 1032 -2544 1038 -2538
rect 1032 -2550 1038 -2544
rect 1032 -2556 1038 -2550
rect 1032 -2562 1038 -2556
rect 1032 -2568 1038 -2562
rect 1032 -2574 1038 -2568
rect 1032 -2580 1038 -2574
rect 1032 -2586 1038 -2580
rect 1032 -2592 1038 -2586
rect 1032 -2598 1038 -2592
rect 1032 -2604 1038 -2598
rect 1032 -2610 1038 -2604
rect 1032 -2616 1038 -2610
rect 1032 -2622 1038 -2616
rect 1032 -2628 1038 -2622
rect 1032 -2634 1038 -2628
rect 1032 -2640 1038 -2634
rect 1032 -2646 1038 -2640
rect 1032 -2652 1038 -2646
rect 1032 -2658 1038 -2652
rect 1032 -2664 1038 -2658
rect 1032 -2670 1038 -2664
rect 1032 -2676 1038 -2670
rect 1032 -2682 1038 -2676
rect 1032 -2688 1038 -2682
rect 1032 -2694 1038 -2688
rect 1032 -2700 1038 -2694
rect 1032 -2706 1038 -2700
rect 1032 -2712 1038 -2706
rect 1032 -2718 1038 -2712
rect 1032 -2724 1038 -2718
rect 1032 -2730 1038 -2724
rect 1032 -2736 1038 -2730
rect 1032 -2742 1038 -2736
rect 1032 -2748 1038 -2742
rect 1032 -2754 1038 -2748
rect 1032 -2760 1038 -2754
rect 1032 -2766 1038 -2760
rect 1032 -2772 1038 -2766
rect 1032 -2778 1038 -2772
rect 1032 -2784 1038 -2778
rect 1032 -2790 1038 -2784
rect 1032 -2796 1038 -2790
rect 1032 -2802 1038 -2796
rect 1032 -2808 1038 -2802
rect 1032 -2814 1038 -2808
rect 1032 -2820 1038 -2814
rect 1032 -2826 1038 -2820
rect 1032 -2832 1038 -2826
rect 1032 -2838 1038 -2832
rect 1032 -2844 1038 -2838
rect 1032 -2850 1038 -2844
rect 1032 -2856 1038 -2850
rect 1032 -2862 1038 -2856
rect 1032 -2868 1038 -2862
rect 1032 -2874 1038 -2868
rect 1032 -2976 1038 -2970
rect 1032 -2982 1038 -2976
rect 1032 -2988 1038 -2982
rect 1032 -2994 1038 -2988
rect 1032 -3000 1038 -2994
rect 1032 -3006 1038 -3000
rect 1032 -3012 1038 -3006
rect 1032 -3018 1038 -3012
rect 1032 -3024 1038 -3018
rect 1032 -3030 1038 -3024
rect 1032 -3036 1038 -3030
rect 1032 -3042 1038 -3036
rect 1032 -3048 1038 -3042
rect 1032 -3054 1038 -3048
rect 1032 -3060 1038 -3054
rect 1032 -3066 1038 -3060
rect 1032 -3072 1038 -3066
rect 1032 -3078 1038 -3072
rect 1032 -3084 1038 -3078
rect 1032 -3090 1038 -3084
rect 1032 -3096 1038 -3090
rect 1032 -3102 1038 -3096
rect 1032 -3108 1038 -3102
rect 1032 -3114 1038 -3108
rect 1032 -3120 1038 -3114
rect 1032 -3126 1038 -3120
rect 1032 -3132 1038 -3126
rect 1032 -3138 1038 -3132
rect 1032 -3144 1038 -3138
rect 1032 -3150 1038 -3144
rect 1032 -3216 1038 -3210
rect 1032 -3222 1038 -3216
rect 1032 -3228 1038 -3222
rect 1032 -3234 1038 -3228
rect 1032 -3240 1038 -3234
rect 1032 -3246 1038 -3240
rect 1032 -3252 1038 -3246
rect 1032 -3258 1038 -3252
rect 1032 -3264 1038 -3258
rect 1032 -3270 1038 -3264
rect 1032 -3276 1038 -3270
rect 1032 -3282 1038 -3276
rect 1032 -3288 1038 -3282
rect 1032 -3294 1038 -3288
rect 1032 -3300 1038 -3294
rect 1032 -3306 1038 -3300
rect 1032 -3312 1038 -3306
rect 1032 -3366 1038 -3360
rect 1032 -3372 1038 -3366
rect 1032 -3378 1038 -3372
rect 1032 -3384 1038 -3378
rect 1032 -3390 1038 -3384
rect 1032 -3396 1038 -3390
rect 1032 -3402 1038 -3396
rect 1032 -3408 1038 -3402
rect 1032 -3414 1038 -3408
rect 1032 -3420 1038 -3414
rect 1032 -3426 1038 -3420
rect 1032 -3432 1038 -3426
rect 1032 -3438 1038 -3432
rect 1032 -3444 1038 -3438
rect 1032 -3450 1038 -3444
rect 1032 -3456 1038 -3450
rect 1032 -3462 1038 -3456
rect 1032 -3468 1038 -3462
rect 1032 -3474 1038 -3468
rect 1032 -3480 1038 -3474
rect 1032 -3486 1038 -3480
rect 1032 -3492 1038 -3486
rect 1032 -3498 1038 -3492
rect 1032 -3504 1038 -3498
rect 1038 -1116 1044 -1110
rect 1038 -1122 1044 -1116
rect 1038 -1128 1044 -1122
rect 1038 -1134 1044 -1128
rect 1038 -1140 1044 -1134
rect 1038 -1146 1044 -1140
rect 1038 -1152 1044 -1146
rect 1038 -1158 1044 -1152
rect 1038 -1164 1044 -1158
rect 1038 -1170 1044 -1164
rect 1038 -1176 1044 -1170
rect 1038 -1182 1044 -1176
rect 1038 -1188 1044 -1182
rect 1038 -1194 1044 -1188
rect 1038 -1200 1044 -1194
rect 1038 -1206 1044 -1200
rect 1038 -1212 1044 -1206
rect 1038 -1218 1044 -1212
rect 1038 -1224 1044 -1218
rect 1038 -1230 1044 -1224
rect 1038 -1236 1044 -1230
rect 1038 -1242 1044 -1236
rect 1038 -1248 1044 -1242
rect 1038 -1254 1044 -1248
rect 1038 -1260 1044 -1254
rect 1038 -1266 1044 -1260
rect 1038 -1272 1044 -1266
rect 1038 -1278 1044 -1272
rect 1038 -1284 1044 -1278
rect 1038 -1290 1044 -1284
rect 1038 -1296 1044 -1290
rect 1038 -1302 1044 -1296
rect 1038 -1308 1044 -1302
rect 1038 -1314 1044 -1308
rect 1038 -1320 1044 -1314
rect 1038 -2286 1044 -2280
rect 1038 -2292 1044 -2286
rect 1038 -2298 1044 -2292
rect 1038 -2304 1044 -2298
rect 1038 -2310 1044 -2304
rect 1038 -2316 1044 -2310
rect 1038 -2322 1044 -2316
rect 1038 -2328 1044 -2322
rect 1038 -2334 1044 -2328
rect 1038 -2340 1044 -2334
rect 1038 -2346 1044 -2340
rect 1038 -2352 1044 -2346
rect 1038 -2358 1044 -2352
rect 1038 -2364 1044 -2358
rect 1038 -2370 1044 -2364
rect 1038 -2376 1044 -2370
rect 1038 -2382 1044 -2376
rect 1038 -2388 1044 -2382
rect 1038 -2394 1044 -2388
rect 1038 -2400 1044 -2394
rect 1038 -2406 1044 -2400
rect 1038 -2412 1044 -2406
rect 1038 -2418 1044 -2412
rect 1038 -2424 1044 -2418
rect 1038 -2430 1044 -2424
rect 1038 -2436 1044 -2430
rect 1038 -2442 1044 -2436
rect 1038 -2448 1044 -2442
rect 1038 -2454 1044 -2448
rect 1038 -2460 1044 -2454
rect 1038 -2466 1044 -2460
rect 1038 -2472 1044 -2466
rect 1038 -2478 1044 -2472
rect 1038 -2484 1044 -2478
rect 1038 -2490 1044 -2484
rect 1038 -2496 1044 -2490
rect 1038 -2502 1044 -2496
rect 1038 -2508 1044 -2502
rect 1038 -2514 1044 -2508
rect 1038 -2520 1044 -2514
rect 1038 -2526 1044 -2520
rect 1038 -2532 1044 -2526
rect 1038 -2538 1044 -2532
rect 1038 -2544 1044 -2538
rect 1038 -2550 1044 -2544
rect 1038 -2556 1044 -2550
rect 1038 -2562 1044 -2556
rect 1038 -2568 1044 -2562
rect 1038 -2574 1044 -2568
rect 1038 -2580 1044 -2574
rect 1038 -2586 1044 -2580
rect 1038 -2592 1044 -2586
rect 1038 -2598 1044 -2592
rect 1038 -2604 1044 -2598
rect 1038 -2610 1044 -2604
rect 1038 -2616 1044 -2610
rect 1038 -2622 1044 -2616
rect 1038 -2628 1044 -2622
rect 1038 -2634 1044 -2628
rect 1038 -2640 1044 -2634
rect 1038 -2646 1044 -2640
rect 1038 -2652 1044 -2646
rect 1038 -2658 1044 -2652
rect 1038 -2664 1044 -2658
rect 1038 -2670 1044 -2664
rect 1038 -2676 1044 -2670
rect 1038 -2682 1044 -2676
rect 1038 -2688 1044 -2682
rect 1038 -2694 1044 -2688
rect 1038 -2700 1044 -2694
rect 1038 -2706 1044 -2700
rect 1038 -2712 1044 -2706
rect 1038 -2718 1044 -2712
rect 1038 -2724 1044 -2718
rect 1038 -2730 1044 -2724
rect 1038 -2736 1044 -2730
rect 1038 -2742 1044 -2736
rect 1038 -2748 1044 -2742
rect 1038 -2754 1044 -2748
rect 1038 -2760 1044 -2754
rect 1038 -2766 1044 -2760
rect 1038 -2772 1044 -2766
rect 1038 -2778 1044 -2772
rect 1038 -2784 1044 -2778
rect 1038 -2790 1044 -2784
rect 1038 -2796 1044 -2790
rect 1038 -2802 1044 -2796
rect 1038 -2808 1044 -2802
rect 1038 -2814 1044 -2808
rect 1038 -2820 1044 -2814
rect 1038 -2826 1044 -2820
rect 1038 -2832 1044 -2826
rect 1038 -2838 1044 -2832
rect 1038 -2844 1044 -2838
rect 1038 -2850 1044 -2844
rect 1038 -2856 1044 -2850
rect 1038 -2862 1044 -2856
rect 1038 -2868 1044 -2862
rect 1038 -2964 1044 -2958
rect 1038 -2970 1044 -2964
rect 1038 -2976 1044 -2970
rect 1038 -2982 1044 -2976
rect 1038 -2988 1044 -2982
rect 1038 -2994 1044 -2988
rect 1038 -3000 1044 -2994
rect 1038 -3006 1044 -3000
rect 1038 -3012 1044 -3006
rect 1038 -3018 1044 -3012
rect 1038 -3024 1044 -3018
rect 1038 -3030 1044 -3024
rect 1038 -3036 1044 -3030
rect 1038 -3042 1044 -3036
rect 1038 -3048 1044 -3042
rect 1038 -3054 1044 -3048
rect 1038 -3060 1044 -3054
rect 1038 -3066 1044 -3060
rect 1038 -3072 1044 -3066
rect 1038 -3078 1044 -3072
rect 1038 -3084 1044 -3078
rect 1038 -3090 1044 -3084
rect 1038 -3096 1044 -3090
rect 1038 -3102 1044 -3096
rect 1038 -3108 1044 -3102
rect 1038 -3114 1044 -3108
rect 1038 -3120 1044 -3114
rect 1038 -3126 1044 -3120
rect 1038 -3132 1044 -3126
rect 1038 -3138 1044 -3132
rect 1038 -3144 1044 -3138
rect 1038 -3216 1044 -3210
rect 1038 -3222 1044 -3216
rect 1038 -3228 1044 -3222
rect 1038 -3234 1044 -3228
rect 1038 -3240 1044 -3234
rect 1038 -3246 1044 -3240
rect 1038 -3252 1044 -3246
rect 1038 -3258 1044 -3252
rect 1038 -3264 1044 -3258
rect 1038 -3270 1044 -3264
rect 1038 -3276 1044 -3270
rect 1038 -3282 1044 -3276
rect 1038 -3288 1044 -3282
rect 1038 -3294 1044 -3288
rect 1038 -3300 1044 -3294
rect 1038 -3306 1044 -3300
rect 1038 -3366 1044 -3360
rect 1038 -3372 1044 -3366
rect 1038 -3378 1044 -3372
rect 1038 -3384 1044 -3378
rect 1038 -3390 1044 -3384
rect 1038 -3396 1044 -3390
rect 1038 -3402 1044 -3396
rect 1038 -3408 1044 -3402
rect 1038 -3414 1044 -3408
rect 1038 -3420 1044 -3414
rect 1038 -3426 1044 -3420
rect 1038 -3432 1044 -3426
rect 1038 -3438 1044 -3432
rect 1038 -3444 1044 -3438
rect 1038 -3450 1044 -3444
rect 1038 -3456 1044 -3450
rect 1038 -3462 1044 -3456
rect 1038 -3468 1044 -3462
rect 1038 -3474 1044 -3468
rect 1038 -3480 1044 -3474
rect 1038 -3486 1044 -3480
rect 1038 -3492 1044 -3486
rect 1038 -3498 1044 -3492
rect 1038 -3504 1044 -3498
rect 1044 -1116 1050 -1110
rect 1044 -1122 1050 -1116
rect 1044 -1128 1050 -1122
rect 1044 -1134 1050 -1128
rect 1044 -1140 1050 -1134
rect 1044 -1146 1050 -1140
rect 1044 -1152 1050 -1146
rect 1044 -1158 1050 -1152
rect 1044 -1164 1050 -1158
rect 1044 -1170 1050 -1164
rect 1044 -1176 1050 -1170
rect 1044 -1182 1050 -1176
rect 1044 -1188 1050 -1182
rect 1044 -1194 1050 -1188
rect 1044 -1200 1050 -1194
rect 1044 -1206 1050 -1200
rect 1044 -1212 1050 -1206
rect 1044 -1218 1050 -1212
rect 1044 -1224 1050 -1218
rect 1044 -1230 1050 -1224
rect 1044 -1236 1050 -1230
rect 1044 -1242 1050 -1236
rect 1044 -1248 1050 -1242
rect 1044 -1254 1050 -1248
rect 1044 -1260 1050 -1254
rect 1044 -1266 1050 -1260
rect 1044 -1272 1050 -1266
rect 1044 -1278 1050 -1272
rect 1044 -1284 1050 -1278
rect 1044 -1290 1050 -1284
rect 1044 -1296 1050 -1290
rect 1044 -1302 1050 -1296
rect 1044 -1308 1050 -1302
rect 1044 -1314 1050 -1308
rect 1044 -1320 1050 -1314
rect 1044 -2262 1050 -2256
rect 1044 -2268 1050 -2262
rect 1044 -2274 1050 -2268
rect 1044 -2280 1050 -2274
rect 1044 -2286 1050 -2280
rect 1044 -2292 1050 -2286
rect 1044 -2298 1050 -2292
rect 1044 -2304 1050 -2298
rect 1044 -2310 1050 -2304
rect 1044 -2316 1050 -2310
rect 1044 -2322 1050 -2316
rect 1044 -2328 1050 -2322
rect 1044 -2334 1050 -2328
rect 1044 -2340 1050 -2334
rect 1044 -2346 1050 -2340
rect 1044 -2352 1050 -2346
rect 1044 -2358 1050 -2352
rect 1044 -2364 1050 -2358
rect 1044 -2370 1050 -2364
rect 1044 -2376 1050 -2370
rect 1044 -2382 1050 -2376
rect 1044 -2388 1050 -2382
rect 1044 -2394 1050 -2388
rect 1044 -2400 1050 -2394
rect 1044 -2406 1050 -2400
rect 1044 -2412 1050 -2406
rect 1044 -2418 1050 -2412
rect 1044 -2424 1050 -2418
rect 1044 -2430 1050 -2424
rect 1044 -2436 1050 -2430
rect 1044 -2442 1050 -2436
rect 1044 -2448 1050 -2442
rect 1044 -2454 1050 -2448
rect 1044 -2460 1050 -2454
rect 1044 -2466 1050 -2460
rect 1044 -2472 1050 -2466
rect 1044 -2478 1050 -2472
rect 1044 -2484 1050 -2478
rect 1044 -2490 1050 -2484
rect 1044 -2496 1050 -2490
rect 1044 -2502 1050 -2496
rect 1044 -2508 1050 -2502
rect 1044 -2514 1050 -2508
rect 1044 -2520 1050 -2514
rect 1044 -2526 1050 -2520
rect 1044 -2532 1050 -2526
rect 1044 -2538 1050 -2532
rect 1044 -2544 1050 -2538
rect 1044 -2550 1050 -2544
rect 1044 -2556 1050 -2550
rect 1044 -2562 1050 -2556
rect 1044 -2568 1050 -2562
rect 1044 -2574 1050 -2568
rect 1044 -2580 1050 -2574
rect 1044 -2586 1050 -2580
rect 1044 -2592 1050 -2586
rect 1044 -2598 1050 -2592
rect 1044 -2604 1050 -2598
rect 1044 -2610 1050 -2604
rect 1044 -2616 1050 -2610
rect 1044 -2622 1050 -2616
rect 1044 -2628 1050 -2622
rect 1044 -2634 1050 -2628
rect 1044 -2640 1050 -2634
rect 1044 -2646 1050 -2640
rect 1044 -2652 1050 -2646
rect 1044 -2658 1050 -2652
rect 1044 -2664 1050 -2658
rect 1044 -2670 1050 -2664
rect 1044 -2676 1050 -2670
rect 1044 -2682 1050 -2676
rect 1044 -2688 1050 -2682
rect 1044 -2694 1050 -2688
rect 1044 -2700 1050 -2694
rect 1044 -2706 1050 -2700
rect 1044 -2712 1050 -2706
rect 1044 -2718 1050 -2712
rect 1044 -2724 1050 -2718
rect 1044 -2730 1050 -2724
rect 1044 -2736 1050 -2730
rect 1044 -2742 1050 -2736
rect 1044 -2748 1050 -2742
rect 1044 -2754 1050 -2748
rect 1044 -2760 1050 -2754
rect 1044 -2766 1050 -2760
rect 1044 -2772 1050 -2766
rect 1044 -2778 1050 -2772
rect 1044 -2784 1050 -2778
rect 1044 -2790 1050 -2784
rect 1044 -2796 1050 -2790
rect 1044 -2802 1050 -2796
rect 1044 -2808 1050 -2802
rect 1044 -2814 1050 -2808
rect 1044 -2820 1050 -2814
rect 1044 -2826 1050 -2820
rect 1044 -2832 1050 -2826
rect 1044 -2838 1050 -2832
rect 1044 -2844 1050 -2838
rect 1044 -2850 1050 -2844
rect 1044 -2856 1050 -2850
rect 1044 -2952 1050 -2946
rect 1044 -2958 1050 -2952
rect 1044 -2964 1050 -2958
rect 1044 -2970 1050 -2964
rect 1044 -2976 1050 -2970
rect 1044 -2982 1050 -2976
rect 1044 -2988 1050 -2982
rect 1044 -2994 1050 -2988
rect 1044 -3000 1050 -2994
rect 1044 -3006 1050 -3000
rect 1044 -3012 1050 -3006
rect 1044 -3018 1050 -3012
rect 1044 -3024 1050 -3018
rect 1044 -3030 1050 -3024
rect 1044 -3036 1050 -3030
rect 1044 -3042 1050 -3036
rect 1044 -3048 1050 -3042
rect 1044 -3054 1050 -3048
rect 1044 -3060 1050 -3054
rect 1044 -3066 1050 -3060
rect 1044 -3072 1050 -3066
rect 1044 -3078 1050 -3072
rect 1044 -3084 1050 -3078
rect 1044 -3090 1050 -3084
rect 1044 -3096 1050 -3090
rect 1044 -3102 1050 -3096
rect 1044 -3108 1050 -3102
rect 1044 -3114 1050 -3108
rect 1044 -3120 1050 -3114
rect 1044 -3126 1050 -3120
rect 1044 -3132 1050 -3126
rect 1044 -3138 1050 -3132
rect 1044 -3144 1050 -3138
rect 1044 -3210 1050 -3204
rect 1044 -3216 1050 -3210
rect 1044 -3222 1050 -3216
rect 1044 -3228 1050 -3222
rect 1044 -3234 1050 -3228
rect 1044 -3240 1050 -3234
rect 1044 -3246 1050 -3240
rect 1044 -3252 1050 -3246
rect 1044 -3258 1050 -3252
rect 1044 -3264 1050 -3258
rect 1044 -3270 1050 -3264
rect 1044 -3276 1050 -3270
rect 1044 -3282 1050 -3276
rect 1044 -3288 1050 -3282
rect 1044 -3294 1050 -3288
rect 1044 -3300 1050 -3294
rect 1044 -3306 1050 -3300
rect 1044 -3360 1050 -3354
rect 1044 -3366 1050 -3360
rect 1044 -3372 1050 -3366
rect 1044 -3378 1050 -3372
rect 1044 -3384 1050 -3378
rect 1044 -3390 1050 -3384
rect 1044 -3396 1050 -3390
rect 1044 -3402 1050 -3396
rect 1044 -3408 1050 -3402
rect 1044 -3414 1050 -3408
rect 1044 -3420 1050 -3414
rect 1044 -3426 1050 -3420
rect 1044 -3432 1050 -3426
rect 1044 -3438 1050 -3432
rect 1044 -3444 1050 -3438
rect 1044 -3450 1050 -3444
rect 1044 -3456 1050 -3450
rect 1044 -3462 1050 -3456
rect 1044 -3468 1050 -3462
rect 1044 -3474 1050 -3468
rect 1044 -3480 1050 -3474
rect 1044 -3486 1050 -3480
rect 1044 -3492 1050 -3486
rect 1044 -3498 1050 -3492
rect 1044 -3504 1050 -3498
rect 1050 -1116 1056 -1110
rect 1050 -1122 1056 -1116
rect 1050 -1128 1056 -1122
rect 1050 -1134 1056 -1128
rect 1050 -1140 1056 -1134
rect 1050 -1146 1056 -1140
rect 1050 -1152 1056 -1146
rect 1050 -1158 1056 -1152
rect 1050 -1164 1056 -1158
rect 1050 -1170 1056 -1164
rect 1050 -1176 1056 -1170
rect 1050 -1182 1056 -1176
rect 1050 -1188 1056 -1182
rect 1050 -1194 1056 -1188
rect 1050 -1200 1056 -1194
rect 1050 -1206 1056 -1200
rect 1050 -1212 1056 -1206
rect 1050 -1218 1056 -1212
rect 1050 -1224 1056 -1218
rect 1050 -1230 1056 -1224
rect 1050 -1236 1056 -1230
rect 1050 -1242 1056 -1236
rect 1050 -1248 1056 -1242
rect 1050 -1254 1056 -1248
rect 1050 -1260 1056 -1254
rect 1050 -1266 1056 -1260
rect 1050 -1272 1056 -1266
rect 1050 -1278 1056 -1272
rect 1050 -1284 1056 -1278
rect 1050 -1290 1056 -1284
rect 1050 -1296 1056 -1290
rect 1050 -1302 1056 -1296
rect 1050 -1308 1056 -1302
rect 1050 -1314 1056 -1308
rect 1050 -1320 1056 -1314
rect 1050 -2244 1056 -2238
rect 1050 -2250 1056 -2244
rect 1050 -2256 1056 -2250
rect 1050 -2262 1056 -2256
rect 1050 -2268 1056 -2262
rect 1050 -2274 1056 -2268
rect 1050 -2280 1056 -2274
rect 1050 -2286 1056 -2280
rect 1050 -2292 1056 -2286
rect 1050 -2298 1056 -2292
rect 1050 -2304 1056 -2298
rect 1050 -2310 1056 -2304
rect 1050 -2316 1056 -2310
rect 1050 -2322 1056 -2316
rect 1050 -2328 1056 -2322
rect 1050 -2334 1056 -2328
rect 1050 -2340 1056 -2334
rect 1050 -2346 1056 -2340
rect 1050 -2352 1056 -2346
rect 1050 -2358 1056 -2352
rect 1050 -2364 1056 -2358
rect 1050 -2370 1056 -2364
rect 1050 -2376 1056 -2370
rect 1050 -2382 1056 -2376
rect 1050 -2388 1056 -2382
rect 1050 -2394 1056 -2388
rect 1050 -2400 1056 -2394
rect 1050 -2406 1056 -2400
rect 1050 -2412 1056 -2406
rect 1050 -2418 1056 -2412
rect 1050 -2424 1056 -2418
rect 1050 -2430 1056 -2424
rect 1050 -2436 1056 -2430
rect 1050 -2442 1056 -2436
rect 1050 -2448 1056 -2442
rect 1050 -2454 1056 -2448
rect 1050 -2460 1056 -2454
rect 1050 -2466 1056 -2460
rect 1050 -2472 1056 -2466
rect 1050 -2478 1056 -2472
rect 1050 -2484 1056 -2478
rect 1050 -2490 1056 -2484
rect 1050 -2496 1056 -2490
rect 1050 -2502 1056 -2496
rect 1050 -2508 1056 -2502
rect 1050 -2514 1056 -2508
rect 1050 -2520 1056 -2514
rect 1050 -2526 1056 -2520
rect 1050 -2532 1056 -2526
rect 1050 -2538 1056 -2532
rect 1050 -2544 1056 -2538
rect 1050 -2550 1056 -2544
rect 1050 -2556 1056 -2550
rect 1050 -2562 1056 -2556
rect 1050 -2568 1056 -2562
rect 1050 -2574 1056 -2568
rect 1050 -2580 1056 -2574
rect 1050 -2586 1056 -2580
rect 1050 -2592 1056 -2586
rect 1050 -2598 1056 -2592
rect 1050 -2604 1056 -2598
rect 1050 -2610 1056 -2604
rect 1050 -2616 1056 -2610
rect 1050 -2622 1056 -2616
rect 1050 -2628 1056 -2622
rect 1050 -2634 1056 -2628
rect 1050 -2640 1056 -2634
rect 1050 -2646 1056 -2640
rect 1050 -2652 1056 -2646
rect 1050 -2658 1056 -2652
rect 1050 -2664 1056 -2658
rect 1050 -2670 1056 -2664
rect 1050 -2676 1056 -2670
rect 1050 -2682 1056 -2676
rect 1050 -2688 1056 -2682
rect 1050 -2694 1056 -2688
rect 1050 -2700 1056 -2694
rect 1050 -2706 1056 -2700
rect 1050 -2712 1056 -2706
rect 1050 -2718 1056 -2712
rect 1050 -2724 1056 -2718
rect 1050 -2730 1056 -2724
rect 1050 -2736 1056 -2730
rect 1050 -2742 1056 -2736
rect 1050 -2748 1056 -2742
rect 1050 -2754 1056 -2748
rect 1050 -2760 1056 -2754
rect 1050 -2766 1056 -2760
rect 1050 -2772 1056 -2766
rect 1050 -2778 1056 -2772
rect 1050 -2784 1056 -2778
rect 1050 -2790 1056 -2784
rect 1050 -2796 1056 -2790
rect 1050 -2802 1056 -2796
rect 1050 -2808 1056 -2802
rect 1050 -2814 1056 -2808
rect 1050 -2820 1056 -2814
rect 1050 -2826 1056 -2820
rect 1050 -2832 1056 -2826
rect 1050 -2838 1056 -2832
rect 1050 -2844 1056 -2838
rect 1050 -2946 1056 -2940
rect 1050 -2952 1056 -2946
rect 1050 -2958 1056 -2952
rect 1050 -2964 1056 -2958
rect 1050 -2970 1056 -2964
rect 1050 -2976 1056 -2970
rect 1050 -2982 1056 -2976
rect 1050 -2988 1056 -2982
rect 1050 -2994 1056 -2988
rect 1050 -3000 1056 -2994
rect 1050 -3006 1056 -3000
rect 1050 -3012 1056 -3006
rect 1050 -3018 1056 -3012
rect 1050 -3024 1056 -3018
rect 1050 -3030 1056 -3024
rect 1050 -3036 1056 -3030
rect 1050 -3042 1056 -3036
rect 1050 -3048 1056 -3042
rect 1050 -3054 1056 -3048
rect 1050 -3060 1056 -3054
rect 1050 -3066 1056 -3060
rect 1050 -3072 1056 -3066
rect 1050 -3078 1056 -3072
rect 1050 -3084 1056 -3078
rect 1050 -3090 1056 -3084
rect 1050 -3096 1056 -3090
rect 1050 -3102 1056 -3096
rect 1050 -3108 1056 -3102
rect 1050 -3114 1056 -3108
rect 1050 -3120 1056 -3114
rect 1050 -3126 1056 -3120
rect 1050 -3132 1056 -3126
rect 1050 -3138 1056 -3132
rect 1050 -3204 1056 -3198
rect 1050 -3210 1056 -3204
rect 1050 -3216 1056 -3210
rect 1050 -3222 1056 -3216
rect 1050 -3228 1056 -3222
rect 1050 -3234 1056 -3228
rect 1050 -3240 1056 -3234
rect 1050 -3246 1056 -3240
rect 1050 -3252 1056 -3246
rect 1050 -3258 1056 -3252
rect 1050 -3264 1056 -3258
rect 1050 -3270 1056 -3264
rect 1050 -3276 1056 -3270
rect 1050 -3282 1056 -3276
rect 1050 -3288 1056 -3282
rect 1050 -3294 1056 -3288
rect 1050 -3300 1056 -3294
rect 1050 -3354 1056 -3348
rect 1050 -3360 1056 -3354
rect 1050 -3366 1056 -3360
rect 1050 -3372 1056 -3366
rect 1050 -3378 1056 -3372
rect 1050 -3384 1056 -3378
rect 1050 -3390 1056 -3384
rect 1050 -3396 1056 -3390
rect 1050 -3402 1056 -3396
rect 1050 -3408 1056 -3402
rect 1050 -3414 1056 -3408
rect 1050 -3420 1056 -3414
rect 1050 -3426 1056 -3420
rect 1050 -3432 1056 -3426
rect 1050 -3438 1056 -3432
rect 1050 -3444 1056 -3438
rect 1050 -3450 1056 -3444
rect 1050 -3456 1056 -3450
rect 1050 -3462 1056 -3456
rect 1050 -3468 1056 -3462
rect 1050 -3474 1056 -3468
rect 1050 -3480 1056 -3474
rect 1050 -3486 1056 -3480
rect 1050 -3492 1056 -3486
rect 1050 -3498 1056 -3492
rect 1050 -3504 1056 -3498
rect 1056 -1116 1062 -1110
rect 1056 -1122 1062 -1116
rect 1056 -1128 1062 -1122
rect 1056 -1134 1062 -1128
rect 1056 -1140 1062 -1134
rect 1056 -1146 1062 -1140
rect 1056 -1152 1062 -1146
rect 1056 -1158 1062 -1152
rect 1056 -1164 1062 -1158
rect 1056 -1170 1062 -1164
rect 1056 -1176 1062 -1170
rect 1056 -1182 1062 -1176
rect 1056 -1188 1062 -1182
rect 1056 -1194 1062 -1188
rect 1056 -1200 1062 -1194
rect 1056 -1206 1062 -1200
rect 1056 -1212 1062 -1206
rect 1056 -1218 1062 -1212
rect 1056 -1224 1062 -1218
rect 1056 -1230 1062 -1224
rect 1056 -1236 1062 -1230
rect 1056 -1242 1062 -1236
rect 1056 -1248 1062 -1242
rect 1056 -1254 1062 -1248
rect 1056 -1260 1062 -1254
rect 1056 -1266 1062 -1260
rect 1056 -1272 1062 -1266
rect 1056 -1278 1062 -1272
rect 1056 -1284 1062 -1278
rect 1056 -1290 1062 -1284
rect 1056 -1296 1062 -1290
rect 1056 -1302 1062 -1296
rect 1056 -1308 1062 -1302
rect 1056 -1314 1062 -1308
rect 1056 -1320 1062 -1314
rect 1056 -2226 1062 -2220
rect 1056 -2232 1062 -2226
rect 1056 -2238 1062 -2232
rect 1056 -2244 1062 -2238
rect 1056 -2250 1062 -2244
rect 1056 -2256 1062 -2250
rect 1056 -2262 1062 -2256
rect 1056 -2268 1062 -2262
rect 1056 -2274 1062 -2268
rect 1056 -2280 1062 -2274
rect 1056 -2286 1062 -2280
rect 1056 -2292 1062 -2286
rect 1056 -2298 1062 -2292
rect 1056 -2304 1062 -2298
rect 1056 -2310 1062 -2304
rect 1056 -2316 1062 -2310
rect 1056 -2322 1062 -2316
rect 1056 -2328 1062 -2322
rect 1056 -2334 1062 -2328
rect 1056 -2340 1062 -2334
rect 1056 -2346 1062 -2340
rect 1056 -2352 1062 -2346
rect 1056 -2358 1062 -2352
rect 1056 -2364 1062 -2358
rect 1056 -2370 1062 -2364
rect 1056 -2376 1062 -2370
rect 1056 -2382 1062 -2376
rect 1056 -2388 1062 -2382
rect 1056 -2394 1062 -2388
rect 1056 -2400 1062 -2394
rect 1056 -2406 1062 -2400
rect 1056 -2412 1062 -2406
rect 1056 -2418 1062 -2412
rect 1056 -2424 1062 -2418
rect 1056 -2430 1062 -2424
rect 1056 -2436 1062 -2430
rect 1056 -2442 1062 -2436
rect 1056 -2448 1062 -2442
rect 1056 -2454 1062 -2448
rect 1056 -2460 1062 -2454
rect 1056 -2466 1062 -2460
rect 1056 -2472 1062 -2466
rect 1056 -2478 1062 -2472
rect 1056 -2484 1062 -2478
rect 1056 -2490 1062 -2484
rect 1056 -2496 1062 -2490
rect 1056 -2502 1062 -2496
rect 1056 -2508 1062 -2502
rect 1056 -2514 1062 -2508
rect 1056 -2520 1062 -2514
rect 1056 -2526 1062 -2520
rect 1056 -2532 1062 -2526
rect 1056 -2538 1062 -2532
rect 1056 -2544 1062 -2538
rect 1056 -2550 1062 -2544
rect 1056 -2556 1062 -2550
rect 1056 -2562 1062 -2556
rect 1056 -2568 1062 -2562
rect 1056 -2574 1062 -2568
rect 1056 -2580 1062 -2574
rect 1056 -2586 1062 -2580
rect 1056 -2592 1062 -2586
rect 1056 -2598 1062 -2592
rect 1056 -2604 1062 -2598
rect 1056 -2610 1062 -2604
rect 1056 -2616 1062 -2610
rect 1056 -2622 1062 -2616
rect 1056 -2628 1062 -2622
rect 1056 -2634 1062 -2628
rect 1056 -2640 1062 -2634
rect 1056 -2646 1062 -2640
rect 1056 -2652 1062 -2646
rect 1056 -2658 1062 -2652
rect 1056 -2664 1062 -2658
rect 1056 -2670 1062 -2664
rect 1056 -2676 1062 -2670
rect 1056 -2682 1062 -2676
rect 1056 -2688 1062 -2682
rect 1056 -2694 1062 -2688
rect 1056 -2700 1062 -2694
rect 1056 -2706 1062 -2700
rect 1056 -2712 1062 -2706
rect 1056 -2718 1062 -2712
rect 1056 -2724 1062 -2718
rect 1056 -2730 1062 -2724
rect 1056 -2736 1062 -2730
rect 1056 -2742 1062 -2736
rect 1056 -2748 1062 -2742
rect 1056 -2754 1062 -2748
rect 1056 -2760 1062 -2754
rect 1056 -2766 1062 -2760
rect 1056 -2772 1062 -2766
rect 1056 -2778 1062 -2772
rect 1056 -2784 1062 -2778
rect 1056 -2790 1062 -2784
rect 1056 -2796 1062 -2790
rect 1056 -2802 1062 -2796
rect 1056 -2808 1062 -2802
rect 1056 -2814 1062 -2808
rect 1056 -2820 1062 -2814
rect 1056 -2826 1062 -2820
rect 1056 -2832 1062 -2826
rect 1056 -2934 1062 -2928
rect 1056 -2940 1062 -2934
rect 1056 -2946 1062 -2940
rect 1056 -2952 1062 -2946
rect 1056 -2958 1062 -2952
rect 1056 -2964 1062 -2958
rect 1056 -2970 1062 -2964
rect 1056 -2976 1062 -2970
rect 1056 -2982 1062 -2976
rect 1056 -2988 1062 -2982
rect 1056 -2994 1062 -2988
rect 1056 -3000 1062 -2994
rect 1056 -3006 1062 -3000
rect 1056 -3012 1062 -3006
rect 1056 -3018 1062 -3012
rect 1056 -3024 1062 -3018
rect 1056 -3030 1062 -3024
rect 1056 -3036 1062 -3030
rect 1056 -3042 1062 -3036
rect 1056 -3048 1062 -3042
rect 1056 -3054 1062 -3048
rect 1056 -3060 1062 -3054
rect 1056 -3066 1062 -3060
rect 1056 -3072 1062 -3066
rect 1056 -3078 1062 -3072
rect 1056 -3084 1062 -3078
rect 1056 -3090 1062 -3084
rect 1056 -3096 1062 -3090
rect 1056 -3102 1062 -3096
rect 1056 -3108 1062 -3102
rect 1056 -3114 1062 -3108
rect 1056 -3120 1062 -3114
rect 1056 -3126 1062 -3120
rect 1056 -3132 1062 -3126
rect 1056 -3198 1062 -3192
rect 1056 -3204 1062 -3198
rect 1056 -3210 1062 -3204
rect 1056 -3216 1062 -3210
rect 1056 -3222 1062 -3216
rect 1056 -3228 1062 -3222
rect 1056 -3234 1062 -3228
rect 1056 -3240 1062 -3234
rect 1056 -3246 1062 -3240
rect 1056 -3252 1062 -3246
rect 1056 -3258 1062 -3252
rect 1056 -3264 1062 -3258
rect 1056 -3270 1062 -3264
rect 1056 -3276 1062 -3270
rect 1056 -3282 1062 -3276
rect 1056 -3288 1062 -3282
rect 1056 -3294 1062 -3288
rect 1056 -3300 1062 -3294
rect 1056 -3348 1062 -3342
rect 1056 -3354 1062 -3348
rect 1056 -3360 1062 -3354
rect 1056 -3366 1062 -3360
rect 1056 -3372 1062 -3366
rect 1056 -3378 1062 -3372
rect 1056 -3384 1062 -3378
rect 1056 -3390 1062 -3384
rect 1056 -3396 1062 -3390
rect 1056 -3402 1062 -3396
rect 1056 -3408 1062 -3402
rect 1056 -3414 1062 -3408
rect 1056 -3420 1062 -3414
rect 1056 -3426 1062 -3420
rect 1056 -3432 1062 -3426
rect 1056 -3438 1062 -3432
rect 1056 -3444 1062 -3438
rect 1056 -3450 1062 -3444
rect 1056 -3456 1062 -3450
rect 1056 -3462 1062 -3456
rect 1056 -3468 1062 -3462
rect 1056 -3474 1062 -3468
rect 1056 -3480 1062 -3474
rect 1056 -3486 1062 -3480
rect 1056 -3492 1062 -3486
rect 1056 -3498 1062 -3492
rect 1056 -3504 1062 -3498
rect 1062 -1116 1068 -1110
rect 1062 -1122 1068 -1116
rect 1062 -1128 1068 -1122
rect 1062 -1134 1068 -1128
rect 1062 -1140 1068 -1134
rect 1062 -1146 1068 -1140
rect 1062 -1152 1068 -1146
rect 1062 -1158 1068 -1152
rect 1062 -1164 1068 -1158
rect 1062 -1170 1068 -1164
rect 1062 -1176 1068 -1170
rect 1062 -1182 1068 -1176
rect 1062 -1188 1068 -1182
rect 1062 -1194 1068 -1188
rect 1062 -1200 1068 -1194
rect 1062 -1206 1068 -1200
rect 1062 -1212 1068 -1206
rect 1062 -1218 1068 -1212
rect 1062 -1224 1068 -1218
rect 1062 -1230 1068 -1224
rect 1062 -1236 1068 -1230
rect 1062 -1242 1068 -1236
rect 1062 -1248 1068 -1242
rect 1062 -1254 1068 -1248
rect 1062 -1260 1068 -1254
rect 1062 -1266 1068 -1260
rect 1062 -1272 1068 -1266
rect 1062 -1278 1068 -1272
rect 1062 -1284 1068 -1278
rect 1062 -1290 1068 -1284
rect 1062 -1296 1068 -1290
rect 1062 -1302 1068 -1296
rect 1062 -1308 1068 -1302
rect 1062 -1314 1068 -1308
rect 1062 -1320 1068 -1314
rect 1062 -2208 1068 -2202
rect 1062 -2214 1068 -2208
rect 1062 -2220 1068 -2214
rect 1062 -2226 1068 -2220
rect 1062 -2232 1068 -2226
rect 1062 -2238 1068 -2232
rect 1062 -2244 1068 -2238
rect 1062 -2250 1068 -2244
rect 1062 -2256 1068 -2250
rect 1062 -2262 1068 -2256
rect 1062 -2268 1068 -2262
rect 1062 -2274 1068 -2268
rect 1062 -2280 1068 -2274
rect 1062 -2286 1068 -2280
rect 1062 -2292 1068 -2286
rect 1062 -2298 1068 -2292
rect 1062 -2304 1068 -2298
rect 1062 -2310 1068 -2304
rect 1062 -2316 1068 -2310
rect 1062 -2322 1068 -2316
rect 1062 -2328 1068 -2322
rect 1062 -2334 1068 -2328
rect 1062 -2340 1068 -2334
rect 1062 -2346 1068 -2340
rect 1062 -2352 1068 -2346
rect 1062 -2358 1068 -2352
rect 1062 -2364 1068 -2358
rect 1062 -2370 1068 -2364
rect 1062 -2376 1068 -2370
rect 1062 -2382 1068 -2376
rect 1062 -2388 1068 -2382
rect 1062 -2394 1068 -2388
rect 1062 -2400 1068 -2394
rect 1062 -2406 1068 -2400
rect 1062 -2412 1068 -2406
rect 1062 -2418 1068 -2412
rect 1062 -2424 1068 -2418
rect 1062 -2430 1068 -2424
rect 1062 -2436 1068 -2430
rect 1062 -2442 1068 -2436
rect 1062 -2448 1068 -2442
rect 1062 -2454 1068 -2448
rect 1062 -2460 1068 -2454
rect 1062 -2466 1068 -2460
rect 1062 -2472 1068 -2466
rect 1062 -2478 1068 -2472
rect 1062 -2484 1068 -2478
rect 1062 -2490 1068 -2484
rect 1062 -2496 1068 -2490
rect 1062 -2502 1068 -2496
rect 1062 -2508 1068 -2502
rect 1062 -2514 1068 -2508
rect 1062 -2520 1068 -2514
rect 1062 -2526 1068 -2520
rect 1062 -2532 1068 -2526
rect 1062 -2538 1068 -2532
rect 1062 -2544 1068 -2538
rect 1062 -2550 1068 -2544
rect 1062 -2556 1068 -2550
rect 1062 -2562 1068 -2556
rect 1062 -2568 1068 -2562
rect 1062 -2574 1068 -2568
rect 1062 -2580 1068 -2574
rect 1062 -2586 1068 -2580
rect 1062 -2592 1068 -2586
rect 1062 -2598 1068 -2592
rect 1062 -2604 1068 -2598
rect 1062 -2610 1068 -2604
rect 1062 -2616 1068 -2610
rect 1062 -2622 1068 -2616
rect 1062 -2628 1068 -2622
rect 1062 -2634 1068 -2628
rect 1062 -2640 1068 -2634
rect 1062 -2646 1068 -2640
rect 1062 -2652 1068 -2646
rect 1062 -2658 1068 -2652
rect 1062 -2664 1068 -2658
rect 1062 -2670 1068 -2664
rect 1062 -2676 1068 -2670
rect 1062 -2682 1068 -2676
rect 1062 -2688 1068 -2682
rect 1062 -2694 1068 -2688
rect 1062 -2700 1068 -2694
rect 1062 -2706 1068 -2700
rect 1062 -2712 1068 -2706
rect 1062 -2718 1068 -2712
rect 1062 -2724 1068 -2718
rect 1062 -2730 1068 -2724
rect 1062 -2736 1068 -2730
rect 1062 -2742 1068 -2736
rect 1062 -2748 1068 -2742
rect 1062 -2754 1068 -2748
rect 1062 -2760 1068 -2754
rect 1062 -2766 1068 -2760
rect 1062 -2772 1068 -2766
rect 1062 -2778 1068 -2772
rect 1062 -2784 1068 -2778
rect 1062 -2790 1068 -2784
rect 1062 -2796 1068 -2790
rect 1062 -2802 1068 -2796
rect 1062 -2808 1068 -2802
rect 1062 -2814 1068 -2808
rect 1062 -2820 1068 -2814
rect 1062 -2826 1068 -2820
rect 1062 -2922 1068 -2916
rect 1062 -2928 1068 -2922
rect 1062 -2934 1068 -2928
rect 1062 -2940 1068 -2934
rect 1062 -2946 1068 -2940
rect 1062 -2952 1068 -2946
rect 1062 -2958 1068 -2952
rect 1062 -2964 1068 -2958
rect 1062 -2970 1068 -2964
rect 1062 -2976 1068 -2970
rect 1062 -2982 1068 -2976
rect 1062 -2988 1068 -2982
rect 1062 -2994 1068 -2988
rect 1062 -3000 1068 -2994
rect 1062 -3006 1068 -3000
rect 1062 -3012 1068 -3006
rect 1062 -3018 1068 -3012
rect 1062 -3024 1068 -3018
rect 1062 -3030 1068 -3024
rect 1062 -3036 1068 -3030
rect 1062 -3042 1068 -3036
rect 1062 -3048 1068 -3042
rect 1062 -3054 1068 -3048
rect 1062 -3060 1068 -3054
rect 1062 -3066 1068 -3060
rect 1062 -3072 1068 -3066
rect 1062 -3078 1068 -3072
rect 1062 -3084 1068 -3078
rect 1062 -3090 1068 -3084
rect 1062 -3096 1068 -3090
rect 1062 -3102 1068 -3096
rect 1062 -3108 1068 -3102
rect 1062 -3114 1068 -3108
rect 1062 -3120 1068 -3114
rect 1062 -3126 1068 -3120
rect 1062 -3198 1068 -3192
rect 1062 -3204 1068 -3198
rect 1062 -3210 1068 -3204
rect 1062 -3216 1068 -3210
rect 1062 -3222 1068 -3216
rect 1062 -3228 1068 -3222
rect 1062 -3234 1068 -3228
rect 1062 -3240 1068 -3234
rect 1062 -3246 1068 -3240
rect 1062 -3252 1068 -3246
rect 1062 -3258 1068 -3252
rect 1062 -3264 1068 -3258
rect 1062 -3270 1068 -3264
rect 1062 -3276 1068 -3270
rect 1062 -3282 1068 -3276
rect 1062 -3288 1068 -3282
rect 1062 -3294 1068 -3288
rect 1062 -3342 1068 -3336
rect 1062 -3348 1068 -3342
rect 1062 -3354 1068 -3348
rect 1062 -3360 1068 -3354
rect 1062 -3366 1068 -3360
rect 1062 -3372 1068 -3366
rect 1062 -3378 1068 -3372
rect 1062 -3384 1068 -3378
rect 1062 -3390 1068 -3384
rect 1062 -3396 1068 -3390
rect 1062 -3402 1068 -3396
rect 1062 -3408 1068 -3402
rect 1062 -3414 1068 -3408
rect 1062 -3420 1068 -3414
rect 1062 -3426 1068 -3420
rect 1062 -3432 1068 -3426
rect 1062 -3438 1068 -3432
rect 1062 -3444 1068 -3438
rect 1062 -3450 1068 -3444
rect 1062 -3456 1068 -3450
rect 1062 -3462 1068 -3456
rect 1062 -3468 1068 -3462
rect 1062 -3474 1068 -3468
rect 1062 -3480 1068 -3474
rect 1062 -3486 1068 -3480
rect 1062 -3492 1068 -3486
rect 1062 -3498 1068 -3492
rect 1062 -3504 1068 -3498
rect 1068 -1110 1074 -1104
rect 1068 -1116 1074 -1110
rect 1068 -1122 1074 -1116
rect 1068 -1128 1074 -1122
rect 1068 -1134 1074 -1128
rect 1068 -1140 1074 -1134
rect 1068 -1146 1074 -1140
rect 1068 -1152 1074 -1146
rect 1068 -1158 1074 -1152
rect 1068 -1164 1074 -1158
rect 1068 -1170 1074 -1164
rect 1068 -1176 1074 -1170
rect 1068 -1182 1074 -1176
rect 1068 -1188 1074 -1182
rect 1068 -1194 1074 -1188
rect 1068 -1200 1074 -1194
rect 1068 -1206 1074 -1200
rect 1068 -1212 1074 -1206
rect 1068 -1218 1074 -1212
rect 1068 -1224 1074 -1218
rect 1068 -1230 1074 -1224
rect 1068 -1236 1074 -1230
rect 1068 -1242 1074 -1236
rect 1068 -1248 1074 -1242
rect 1068 -1254 1074 -1248
rect 1068 -1260 1074 -1254
rect 1068 -1266 1074 -1260
rect 1068 -1272 1074 -1266
rect 1068 -1278 1074 -1272
rect 1068 -1284 1074 -1278
rect 1068 -1290 1074 -1284
rect 1068 -1296 1074 -1290
rect 1068 -1302 1074 -1296
rect 1068 -1308 1074 -1302
rect 1068 -1314 1074 -1308
rect 1068 -2190 1074 -2184
rect 1068 -2196 1074 -2190
rect 1068 -2202 1074 -2196
rect 1068 -2208 1074 -2202
rect 1068 -2214 1074 -2208
rect 1068 -2220 1074 -2214
rect 1068 -2226 1074 -2220
rect 1068 -2232 1074 -2226
rect 1068 -2238 1074 -2232
rect 1068 -2244 1074 -2238
rect 1068 -2250 1074 -2244
rect 1068 -2256 1074 -2250
rect 1068 -2262 1074 -2256
rect 1068 -2268 1074 -2262
rect 1068 -2274 1074 -2268
rect 1068 -2280 1074 -2274
rect 1068 -2286 1074 -2280
rect 1068 -2292 1074 -2286
rect 1068 -2298 1074 -2292
rect 1068 -2304 1074 -2298
rect 1068 -2310 1074 -2304
rect 1068 -2316 1074 -2310
rect 1068 -2322 1074 -2316
rect 1068 -2328 1074 -2322
rect 1068 -2334 1074 -2328
rect 1068 -2340 1074 -2334
rect 1068 -2346 1074 -2340
rect 1068 -2352 1074 -2346
rect 1068 -2358 1074 -2352
rect 1068 -2364 1074 -2358
rect 1068 -2370 1074 -2364
rect 1068 -2376 1074 -2370
rect 1068 -2382 1074 -2376
rect 1068 -2388 1074 -2382
rect 1068 -2394 1074 -2388
rect 1068 -2400 1074 -2394
rect 1068 -2406 1074 -2400
rect 1068 -2412 1074 -2406
rect 1068 -2418 1074 -2412
rect 1068 -2424 1074 -2418
rect 1068 -2430 1074 -2424
rect 1068 -2436 1074 -2430
rect 1068 -2442 1074 -2436
rect 1068 -2448 1074 -2442
rect 1068 -2454 1074 -2448
rect 1068 -2460 1074 -2454
rect 1068 -2466 1074 -2460
rect 1068 -2472 1074 -2466
rect 1068 -2478 1074 -2472
rect 1068 -2484 1074 -2478
rect 1068 -2490 1074 -2484
rect 1068 -2496 1074 -2490
rect 1068 -2502 1074 -2496
rect 1068 -2508 1074 -2502
rect 1068 -2514 1074 -2508
rect 1068 -2520 1074 -2514
rect 1068 -2526 1074 -2520
rect 1068 -2532 1074 -2526
rect 1068 -2538 1074 -2532
rect 1068 -2544 1074 -2538
rect 1068 -2550 1074 -2544
rect 1068 -2556 1074 -2550
rect 1068 -2562 1074 -2556
rect 1068 -2568 1074 -2562
rect 1068 -2574 1074 -2568
rect 1068 -2580 1074 -2574
rect 1068 -2586 1074 -2580
rect 1068 -2592 1074 -2586
rect 1068 -2598 1074 -2592
rect 1068 -2604 1074 -2598
rect 1068 -2610 1074 -2604
rect 1068 -2616 1074 -2610
rect 1068 -2622 1074 -2616
rect 1068 -2628 1074 -2622
rect 1068 -2634 1074 -2628
rect 1068 -2640 1074 -2634
rect 1068 -2646 1074 -2640
rect 1068 -2652 1074 -2646
rect 1068 -2658 1074 -2652
rect 1068 -2664 1074 -2658
rect 1068 -2670 1074 -2664
rect 1068 -2676 1074 -2670
rect 1068 -2682 1074 -2676
rect 1068 -2688 1074 -2682
rect 1068 -2694 1074 -2688
rect 1068 -2700 1074 -2694
rect 1068 -2706 1074 -2700
rect 1068 -2712 1074 -2706
rect 1068 -2718 1074 -2712
rect 1068 -2724 1074 -2718
rect 1068 -2730 1074 -2724
rect 1068 -2736 1074 -2730
rect 1068 -2742 1074 -2736
rect 1068 -2748 1074 -2742
rect 1068 -2754 1074 -2748
rect 1068 -2760 1074 -2754
rect 1068 -2766 1074 -2760
rect 1068 -2772 1074 -2766
rect 1068 -2778 1074 -2772
rect 1068 -2784 1074 -2778
rect 1068 -2790 1074 -2784
rect 1068 -2796 1074 -2790
rect 1068 -2802 1074 -2796
rect 1068 -2808 1074 -2802
rect 1068 -2814 1074 -2808
rect 1068 -2916 1074 -2910
rect 1068 -2922 1074 -2916
rect 1068 -2928 1074 -2922
rect 1068 -2934 1074 -2928
rect 1068 -2940 1074 -2934
rect 1068 -2946 1074 -2940
rect 1068 -2952 1074 -2946
rect 1068 -2958 1074 -2952
rect 1068 -2964 1074 -2958
rect 1068 -2970 1074 -2964
rect 1068 -2976 1074 -2970
rect 1068 -2982 1074 -2976
rect 1068 -2988 1074 -2982
rect 1068 -2994 1074 -2988
rect 1068 -3000 1074 -2994
rect 1068 -3006 1074 -3000
rect 1068 -3012 1074 -3006
rect 1068 -3018 1074 -3012
rect 1068 -3024 1074 -3018
rect 1068 -3030 1074 -3024
rect 1068 -3036 1074 -3030
rect 1068 -3042 1074 -3036
rect 1068 -3048 1074 -3042
rect 1068 -3054 1074 -3048
rect 1068 -3060 1074 -3054
rect 1068 -3066 1074 -3060
rect 1068 -3072 1074 -3066
rect 1068 -3078 1074 -3072
rect 1068 -3084 1074 -3078
rect 1068 -3090 1074 -3084
rect 1068 -3096 1074 -3090
rect 1068 -3102 1074 -3096
rect 1068 -3108 1074 -3102
rect 1068 -3114 1074 -3108
rect 1068 -3120 1074 -3114
rect 1068 -3126 1074 -3120
rect 1068 -3192 1074 -3186
rect 1068 -3198 1074 -3192
rect 1068 -3204 1074 -3198
rect 1068 -3210 1074 -3204
rect 1068 -3216 1074 -3210
rect 1068 -3222 1074 -3216
rect 1068 -3228 1074 -3222
rect 1068 -3234 1074 -3228
rect 1068 -3240 1074 -3234
rect 1068 -3246 1074 -3240
rect 1068 -3252 1074 -3246
rect 1068 -3258 1074 -3252
rect 1068 -3264 1074 -3258
rect 1068 -3270 1074 -3264
rect 1068 -3276 1074 -3270
rect 1068 -3282 1074 -3276
rect 1068 -3288 1074 -3282
rect 1068 -3294 1074 -3288
rect 1068 -3336 1074 -3330
rect 1068 -3342 1074 -3336
rect 1068 -3348 1074 -3342
rect 1068 -3354 1074 -3348
rect 1068 -3360 1074 -3354
rect 1068 -3366 1074 -3360
rect 1068 -3372 1074 -3366
rect 1068 -3378 1074 -3372
rect 1068 -3384 1074 -3378
rect 1068 -3390 1074 -3384
rect 1068 -3396 1074 -3390
rect 1068 -3402 1074 -3396
rect 1068 -3408 1074 -3402
rect 1068 -3414 1074 -3408
rect 1068 -3420 1074 -3414
rect 1068 -3426 1074 -3420
rect 1068 -3432 1074 -3426
rect 1068 -3438 1074 -3432
rect 1068 -3444 1074 -3438
rect 1068 -3450 1074 -3444
rect 1068 -3456 1074 -3450
rect 1068 -3462 1074 -3456
rect 1068 -3468 1074 -3462
rect 1068 -3474 1074 -3468
rect 1068 -3480 1074 -3474
rect 1068 -3486 1074 -3480
rect 1068 -3492 1074 -3486
rect 1068 -3498 1074 -3492
rect 1068 -3504 1074 -3498
rect 1074 -1110 1080 -1104
rect 1074 -1116 1080 -1110
rect 1074 -1122 1080 -1116
rect 1074 -1128 1080 -1122
rect 1074 -1134 1080 -1128
rect 1074 -1140 1080 -1134
rect 1074 -1146 1080 -1140
rect 1074 -1152 1080 -1146
rect 1074 -1158 1080 -1152
rect 1074 -1164 1080 -1158
rect 1074 -1170 1080 -1164
rect 1074 -1176 1080 -1170
rect 1074 -1182 1080 -1176
rect 1074 -1188 1080 -1182
rect 1074 -1194 1080 -1188
rect 1074 -1200 1080 -1194
rect 1074 -1206 1080 -1200
rect 1074 -1212 1080 -1206
rect 1074 -1218 1080 -1212
rect 1074 -1224 1080 -1218
rect 1074 -1230 1080 -1224
rect 1074 -1236 1080 -1230
rect 1074 -1242 1080 -1236
rect 1074 -1248 1080 -1242
rect 1074 -1254 1080 -1248
rect 1074 -1260 1080 -1254
rect 1074 -1266 1080 -1260
rect 1074 -1272 1080 -1266
rect 1074 -1278 1080 -1272
rect 1074 -1284 1080 -1278
rect 1074 -1290 1080 -1284
rect 1074 -1296 1080 -1290
rect 1074 -1302 1080 -1296
rect 1074 -1308 1080 -1302
rect 1074 -1314 1080 -1308
rect 1074 -2166 1080 -2160
rect 1074 -2172 1080 -2166
rect 1074 -2178 1080 -2172
rect 1074 -2184 1080 -2178
rect 1074 -2190 1080 -2184
rect 1074 -2196 1080 -2190
rect 1074 -2202 1080 -2196
rect 1074 -2208 1080 -2202
rect 1074 -2214 1080 -2208
rect 1074 -2220 1080 -2214
rect 1074 -2226 1080 -2220
rect 1074 -2232 1080 -2226
rect 1074 -2238 1080 -2232
rect 1074 -2244 1080 -2238
rect 1074 -2250 1080 -2244
rect 1074 -2256 1080 -2250
rect 1074 -2262 1080 -2256
rect 1074 -2268 1080 -2262
rect 1074 -2274 1080 -2268
rect 1074 -2280 1080 -2274
rect 1074 -2286 1080 -2280
rect 1074 -2292 1080 -2286
rect 1074 -2298 1080 -2292
rect 1074 -2304 1080 -2298
rect 1074 -2310 1080 -2304
rect 1074 -2316 1080 -2310
rect 1074 -2322 1080 -2316
rect 1074 -2328 1080 -2322
rect 1074 -2334 1080 -2328
rect 1074 -2340 1080 -2334
rect 1074 -2346 1080 -2340
rect 1074 -2352 1080 -2346
rect 1074 -2358 1080 -2352
rect 1074 -2364 1080 -2358
rect 1074 -2370 1080 -2364
rect 1074 -2376 1080 -2370
rect 1074 -2382 1080 -2376
rect 1074 -2388 1080 -2382
rect 1074 -2394 1080 -2388
rect 1074 -2400 1080 -2394
rect 1074 -2406 1080 -2400
rect 1074 -2412 1080 -2406
rect 1074 -2418 1080 -2412
rect 1074 -2424 1080 -2418
rect 1074 -2430 1080 -2424
rect 1074 -2436 1080 -2430
rect 1074 -2442 1080 -2436
rect 1074 -2448 1080 -2442
rect 1074 -2454 1080 -2448
rect 1074 -2460 1080 -2454
rect 1074 -2466 1080 -2460
rect 1074 -2472 1080 -2466
rect 1074 -2478 1080 -2472
rect 1074 -2484 1080 -2478
rect 1074 -2490 1080 -2484
rect 1074 -2496 1080 -2490
rect 1074 -2502 1080 -2496
rect 1074 -2508 1080 -2502
rect 1074 -2514 1080 -2508
rect 1074 -2520 1080 -2514
rect 1074 -2526 1080 -2520
rect 1074 -2532 1080 -2526
rect 1074 -2538 1080 -2532
rect 1074 -2544 1080 -2538
rect 1074 -2550 1080 -2544
rect 1074 -2556 1080 -2550
rect 1074 -2562 1080 -2556
rect 1074 -2568 1080 -2562
rect 1074 -2574 1080 -2568
rect 1074 -2580 1080 -2574
rect 1074 -2586 1080 -2580
rect 1074 -2592 1080 -2586
rect 1074 -2598 1080 -2592
rect 1074 -2604 1080 -2598
rect 1074 -2610 1080 -2604
rect 1074 -2616 1080 -2610
rect 1074 -2622 1080 -2616
rect 1074 -2628 1080 -2622
rect 1074 -2634 1080 -2628
rect 1074 -2640 1080 -2634
rect 1074 -2646 1080 -2640
rect 1074 -2652 1080 -2646
rect 1074 -2658 1080 -2652
rect 1074 -2664 1080 -2658
rect 1074 -2670 1080 -2664
rect 1074 -2676 1080 -2670
rect 1074 -2682 1080 -2676
rect 1074 -2688 1080 -2682
rect 1074 -2694 1080 -2688
rect 1074 -2700 1080 -2694
rect 1074 -2706 1080 -2700
rect 1074 -2712 1080 -2706
rect 1074 -2718 1080 -2712
rect 1074 -2724 1080 -2718
rect 1074 -2730 1080 -2724
rect 1074 -2736 1080 -2730
rect 1074 -2742 1080 -2736
rect 1074 -2748 1080 -2742
rect 1074 -2754 1080 -2748
rect 1074 -2760 1080 -2754
rect 1074 -2766 1080 -2760
rect 1074 -2772 1080 -2766
rect 1074 -2778 1080 -2772
rect 1074 -2784 1080 -2778
rect 1074 -2790 1080 -2784
rect 1074 -2796 1080 -2790
rect 1074 -2802 1080 -2796
rect 1074 -2904 1080 -2898
rect 1074 -2910 1080 -2904
rect 1074 -2916 1080 -2910
rect 1074 -2922 1080 -2916
rect 1074 -2928 1080 -2922
rect 1074 -2934 1080 -2928
rect 1074 -2940 1080 -2934
rect 1074 -2946 1080 -2940
rect 1074 -2952 1080 -2946
rect 1074 -2958 1080 -2952
rect 1074 -2964 1080 -2958
rect 1074 -2970 1080 -2964
rect 1074 -2976 1080 -2970
rect 1074 -2982 1080 -2976
rect 1074 -2988 1080 -2982
rect 1074 -2994 1080 -2988
rect 1074 -3000 1080 -2994
rect 1074 -3006 1080 -3000
rect 1074 -3012 1080 -3006
rect 1074 -3018 1080 -3012
rect 1074 -3024 1080 -3018
rect 1074 -3030 1080 -3024
rect 1074 -3036 1080 -3030
rect 1074 -3042 1080 -3036
rect 1074 -3048 1080 -3042
rect 1074 -3054 1080 -3048
rect 1074 -3060 1080 -3054
rect 1074 -3066 1080 -3060
rect 1074 -3072 1080 -3066
rect 1074 -3078 1080 -3072
rect 1074 -3084 1080 -3078
rect 1074 -3090 1080 -3084
rect 1074 -3096 1080 -3090
rect 1074 -3102 1080 -3096
rect 1074 -3108 1080 -3102
rect 1074 -3114 1080 -3108
rect 1074 -3120 1080 -3114
rect 1074 -3186 1080 -3180
rect 1074 -3192 1080 -3186
rect 1074 -3198 1080 -3192
rect 1074 -3204 1080 -3198
rect 1074 -3210 1080 -3204
rect 1074 -3216 1080 -3210
rect 1074 -3222 1080 -3216
rect 1074 -3228 1080 -3222
rect 1074 -3234 1080 -3228
rect 1074 -3240 1080 -3234
rect 1074 -3246 1080 -3240
rect 1074 -3252 1080 -3246
rect 1074 -3258 1080 -3252
rect 1074 -3264 1080 -3258
rect 1074 -3270 1080 -3264
rect 1074 -3276 1080 -3270
rect 1074 -3282 1080 -3276
rect 1074 -3288 1080 -3282
rect 1074 -3336 1080 -3330
rect 1074 -3342 1080 -3336
rect 1074 -3348 1080 -3342
rect 1074 -3354 1080 -3348
rect 1074 -3360 1080 -3354
rect 1074 -3366 1080 -3360
rect 1074 -3372 1080 -3366
rect 1074 -3378 1080 -3372
rect 1074 -3384 1080 -3378
rect 1074 -3390 1080 -3384
rect 1074 -3396 1080 -3390
rect 1074 -3402 1080 -3396
rect 1074 -3408 1080 -3402
rect 1074 -3414 1080 -3408
rect 1074 -3420 1080 -3414
rect 1074 -3426 1080 -3420
rect 1074 -3432 1080 -3426
rect 1074 -3438 1080 -3432
rect 1074 -3444 1080 -3438
rect 1074 -3450 1080 -3444
rect 1074 -3456 1080 -3450
rect 1074 -3462 1080 -3456
rect 1074 -3468 1080 -3462
rect 1074 -3474 1080 -3468
rect 1074 -3480 1080 -3474
rect 1074 -3486 1080 -3480
rect 1074 -3492 1080 -3486
rect 1074 -3498 1080 -3492
rect 1074 -3504 1080 -3498
rect 1080 -1110 1086 -1104
rect 1080 -1116 1086 -1110
rect 1080 -1122 1086 -1116
rect 1080 -1128 1086 -1122
rect 1080 -1134 1086 -1128
rect 1080 -1140 1086 -1134
rect 1080 -1146 1086 -1140
rect 1080 -1152 1086 -1146
rect 1080 -1158 1086 -1152
rect 1080 -1164 1086 -1158
rect 1080 -1170 1086 -1164
rect 1080 -1176 1086 -1170
rect 1080 -1182 1086 -1176
rect 1080 -1188 1086 -1182
rect 1080 -1194 1086 -1188
rect 1080 -1200 1086 -1194
rect 1080 -1206 1086 -1200
rect 1080 -1212 1086 -1206
rect 1080 -1218 1086 -1212
rect 1080 -1224 1086 -1218
rect 1080 -1230 1086 -1224
rect 1080 -1236 1086 -1230
rect 1080 -1242 1086 -1236
rect 1080 -1248 1086 -1242
rect 1080 -1254 1086 -1248
rect 1080 -1260 1086 -1254
rect 1080 -1266 1086 -1260
rect 1080 -1272 1086 -1266
rect 1080 -1278 1086 -1272
rect 1080 -1284 1086 -1278
rect 1080 -1290 1086 -1284
rect 1080 -1296 1086 -1290
rect 1080 -1302 1086 -1296
rect 1080 -1308 1086 -1302
rect 1080 -1314 1086 -1308
rect 1080 -2148 1086 -2142
rect 1080 -2154 1086 -2148
rect 1080 -2160 1086 -2154
rect 1080 -2166 1086 -2160
rect 1080 -2172 1086 -2166
rect 1080 -2178 1086 -2172
rect 1080 -2184 1086 -2178
rect 1080 -2190 1086 -2184
rect 1080 -2196 1086 -2190
rect 1080 -2202 1086 -2196
rect 1080 -2208 1086 -2202
rect 1080 -2214 1086 -2208
rect 1080 -2220 1086 -2214
rect 1080 -2226 1086 -2220
rect 1080 -2232 1086 -2226
rect 1080 -2238 1086 -2232
rect 1080 -2244 1086 -2238
rect 1080 -2250 1086 -2244
rect 1080 -2256 1086 -2250
rect 1080 -2262 1086 -2256
rect 1080 -2268 1086 -2262
rect 1080 -2274 1086 -2268
rect 1080 -2280 1086 -2274
rect 1080 -2286 1086 -2280
rect 1080 -2292 1086 -2286
rect 1080 -2298 1086 -2292
rect 1080 -2304 1086 -2298
rect 1080 -2310 1086 -2304
rect 1080 -2316 1086 -2310
rect 1080 -2322 1086 -2316
rect 1080 -2328 1086 -2322
rect 1080 -2334 1086 -2328
rect 1080 -2340 1086 -2334
rect 1080 -2346 1086 -2340
rect 1080 -2352 1086 -2346
rect 1080 -2358 1086 -2352
rect 1080 -2364 1086 -2358
rect 1080 -2370 1086 -2364
rect 1080 -2376 1086 -2370
rect 1080 -2382 1086 -2376
rect 1080 -2388 1086 -2382
rect 1080 -2394 1086 -2388
rect 1080 -2400 1086 -2394
rect 1080 -2406 1086 -2400
rect 1080 -2412 1086 -2406
rect 1080 -2418 1086 -2412
rect 1080 -2424 1086 -2418
rect 1080 -2430 1086 -2424
rect 1080 -2436 1086 -2430
rect 1080 -2442 1086 -2436
rect 1080 -2448 1086 -2442
rect 1080 -2454 1086 -2448
rect 1080 -2460 1086 -2454
rect 1080 -2466 1086 -2460
rect 1080 -2472 1086 -2466
rect 1080 -2478 1086 -2472
rect 1080 -2484 1086 -2478
rect 1080 -2490 1086 -2484
rect 1080 -2496 1086 -2490
rect 1080 -2502 1086 -2496
rect 1080 -2508 1086 -2502
rect 1080 -2514 1086 -2508
rect 1080 -2520 1086 -2514
rect 1080 -2526 1086 -2520
rect 1080 -2532 1086 -2526
rect 1080 -2538 1086 -2532
rect 1080 -2544 1086 -2538
rect 1080 -2550 1086 -2544
rect 1080 -2556 1086 -2550
rect 1080 -2562 1086 -2556
rect 1080 -2568 1086 -2562
rect 1080 -2574 1086 -2568
rect 1080 -2580 1086 -2574
rect 1080 -2586 1086 -2580
rect 1080 -2592 1086 -2586
rect 1080 -2598 1086 -2592
rect 1080 -2604 1086 -2598
rect 1080 -2610 1086 -2604
rect 1080 -2616 1086 -2610
rect 1080 -2622 1086 -2616
rect 1080 -2628 1086 -2622
rect 1080 -2634 1086 -2628
rect 1080 -2640 1086 -2634
rect 1080 -2646 1086 -2640
rect 1080 -2652 1086 -2646
rect 1080 -2658 1086 -2652
rect 1080 -2664 1086 -2658
rect 1080 -2670 1086 -2664
rect 1080 -2676 1086 -2670
rect 1080 -2682 1086 -2676
rect 1080 -2688 1086 -2682
rect 1080 -2694 1086 -2688
rect 1080 -2700 1086 -2694
rect 1080 -2706 1086 -2700
rect 1080 -2712 1086 -2706
rect 1080 -2718 1086 -2712
rect 1080 -2724 1086 -2718
rect 1080 -2730 1086 -2724
rect 1080 -2736 1086 -2730
rect 1080 -2742 1086 -2736
rect 1080 -2748 1086 -2742
rect 1080 -2754 1086 -2748
rect 1080 -2760 1086 -2754
rect 1080 -2766 1086 -2760
rect 1080 -2772 1086 -2766
rect 1080 -2778 1086 -2772
rect 1080 -2784 1086 -2778
rect 1080 -2790 1086 -2784
rect 1080 -2892 1086 -2886
rect 1080 -2898 1086 -2892
rect 1080 -2904 1086 -2898
rect 1080 -2910 1086 -2904
rect 1080 -2916 1086 -2910
rect 1080 -2922 1086 -2916
rect 1080 -2928 1086 -2922
rect 1080 -2934 1086 -2928
rect 1080 -2940 1086 -2934
rect 1080 -2946 1086 -2940
rect 1080 -2952 1086 -2946
rect 1080 -2958 1086 -2952
rect 1080 -2964 1086 -2958
rect 1080 -2970 1086 -2964
rect 1080 -2976 1086 -2970
rect 1080 -2982 1086 -2976
rect 1080 -2988 1086 -2982
rect 1080 -2994 1086 -2988
rect 1080 -3000 1086 -2994
rect 1080 -3006 1086 -3000
rect 1080 -3012 1086 -3006
rect 1080 -3018 1086 -3012
rect 1080 -3024 1086 -3018
rect 1080 -3030 1086 -3024
rect 1080 -3036 1086 -3030
rect 1080 -3042 1086 -3036
rect 1080 -3048 1086 -3042
rect 1080 -3054 1086 -3048
rect 1080 -3060 1086 -3054
rect 1080 -3066 1086 -3060
rect 1080 -3072 1086 -3066
rect 1080 -3078 1086 -3072
rect 1080 -3084 1086 -3078
rect 1080 -3090 1086 -3084
rect 1080 -3096 1086 -3090
rect 1080 -3102 1086 -3096
rect 1080 -3108 1086 -3102
rect 1080 -3114 1086 -3108
rect 1080 -3180 1086 -3174
rect 1080 -3186 1086 -3180
rect 1080 -3192 1086 -3186
rect 1080 -3198 1086 -3192
rect 1080 -3204 1086 -3198
rect 1080 -3210 1086 -3204
rect 1080 -3216 1086 -3210
rect 1080 -3222 1086 -3216
rect 1080 -3228 1086 -3222
rect 1080 -3234 1086 -3228
rect 1080 -3240 1086 -3234
rect 1080 -3246 1086 -3240
rect 1080 -3252 1086 -3246
rect 1080 -3258 1086 -3252
rect 1080 -3264 1086 -3258
rect 1080 -3270 1086 -3264
rect 1080 -3276 1086 -3270
rect 1080 -3282 1086 -3276
rect 1080 -3330 1086 -3324
rect 1080 -3336 1086 -3330
rect 1080 -3342 1086 -3336
rect 1080 -3348 1086 -3342
rect 1080 -3354 1086 -3348
rect 1080 -3360 1086 -3354
rect 1080 -3366 1086 -3360
rect 1080 -3372 1086 -3366
rect 1080 -3378 1086 -3372
rect 1080 -3384 1086 -3378
rect 1080 -3390 1086 -3384
rect 1080 -3396 1086 -3390
rect 1080 -3402 1086 -3396
rect 1080 -3408 1086 -3402
rect 1080 -3414 1086 -3408
rect 1080 -3420 1086 -3414
rect 1080 -3426 1086 -3420
rect 1080 -3432 1086 -3426
rect 1080 -3438 1086 -3432
rect 1080 -3444 1086 -3438
rect 1080 -3450 1086 -3444
rect 1080 -3456 1086 -3450
rect 1080 -3462 1086 -3456
rect 1080 -3468 1086 -3462
rect 1080 -3474 1086 -3468
rect 1080 -3480 1086 -3474
rect 1080 -3486 1086 -3480
rect 1080 -3492 1086 -3486
rect 1080 -3498 1086 -3492
rect 1080 -3504 1086 -3498
rect 1080 -3510 1086 -3504
rect 1086 -1110 1092 -1104
rect 1086 -1116 1092 -1110
rect 1086 -1122 1092 -1116
rect 1086 -1128 1092 -1122
rect 1086 -1134 1092 -1128
rect 1086 -1140 1092 -1134
rect 1086 -1146 1092 -1140
rect 1086 -1152 1092 -1146
rect 1086 -1158 1092 -1152
rect 1086 -1164 1092 -1158
rect 1086 -1170 1092 -1164
rect 1086 -1176 1092 -1170
rect 1086 -1182 1092 -1176
rect 1086 -1188 1092 -1182
rect 1086 -1194 1092 -1188
rect 1086 -1200 1092 -1194
rect 1086 -1206 1092 -1200
rect 1086 -1212 1092 -1206
rect 1086 -1218 1092 -1212
rect 1086 -1224 1092 -1218
rect 1086 -1230 1092 -1224
rect 1086 -1236 1092 -1230
rect 1086 -1242 1092 -1236
rect 1086 -1248 1092 -1242
rect 1086 -1254 1092 -1248
rect 1086 -1260 1092 -1254
rect 1086 -1266 1092 -1260
rect 1086 -1272 1092 -1266
rect 1086 -1278 1092 -1272
rect 1086 -1284 1092 -1278
rect 1086 -1290 1092 -1284
rect 1086 -1296 1092 -1290
rect 1086 -1302 1092 -1296
rect 1086 -1308 1092 -1302
rect 1086 -1314 1092 -1308
rect 1086 -2130 1092 -2124
rect 1086 -2136 1092 -2130
rect 1086 -2142 1092 -2136
rect 1086 -2148 1092 -2142
rect 1086 -2154 1092 -2148
rect 1086 -2160 1092 -2154
rect 1086 -2166 1092 -2160
rect 1086 -2172 1092 -2166
rect 1086 -2178 1092 -2172
rect 1086 -2184 1092 -2178
rect 1086 -2190 1092 -2184
rect 1086 -2196 1092 -2190
rect 1086 -2202 1092 -2196
rect 1086 -2208 1092 -2202
rect 1086 -2214 1092 -2208
rect 1086 -2220 1092 -2214
rect 1086 -2226 1092 -2220
rect 1086 -2232 1092 -2226
rect 1086 -2238 1092 -2232
rect 1086 -2244 1092 -2238
rect 1086 -2250 1092 -2244
rect 1086 -2256 1092 -2250
rect 1086 -2262 1092 -2256
rect 1086 -2268 1092 -2262
rect 1086 -2274 1092 -2268
rect 1086 -2280 1092 -2274
rect 1086 -2286 1092 -2280
rect 1086 -2292 1092 -2286
rect 1086 -2298 1092 -2292
rect 1086 -2304 1092 -2298
rect 1086 -2310 1092 -2304
rect 1086 -2316 1092 -2310
rect 1086 -2322 1092 -2316
rect 1086 -2328 1092 -2322
rect 1086 -2334 1092 -2328
rect 1086 -2340 1092 -2334
rect 1086 -2346 1092 -2340
rect 1086 -2352 1092 -2346
rect 1086 -2358 1092 -2352
rect 1086 -2364 1092 -2358
rect 1086 -2370 1092 -2364
rect 1086 -2376 1092 -2370
rect 1086 -2382 1092 -2376
rect 1086 -2388 1092 -2382
rect 1086 -2394 1092 -2388
rect 1086 -2400 1092 -2394
rect 1086 -2406 1092 -2400
rect 1086 -2412 1092 -2406
rect 1086 -2418 1092 -2412
rect 1086 -2424 1092 -2418
rect 1086 -2430 1092 -2424
rect 1086 -2436 1092 -2430
rect 1086 -2442 1092 -2436
rect 1086 -2448 1092 -2442
rect 1086 -2454 1092 -2448
rect 1086 -2460 1092 -2454
rect 1086 -2466 1092 -2460
rect 1086 -2472 1092 -2466
rect 1086 -2478 1092 -2472
rect 1086 -2484 1092 -2478
rect 1086 -2490 1092 -2484
rect 1086 -2496 1092 -2490
rect 1086 -2502 1092 -2496
rect 1086 -2508 1092 -2502
rect 1086 -2514 1092 -2508
rect 1086 -2520 1092 -2514
rect 1086 -2526 1092 -2520
rect 1086 -2532 1092 -2526
rect 1086 -2538 1092 -2532
rect 1086 -2544 1092 -2538
rect 1086 -2550 1092 -2544
rect 1086 -2556 1092 -2550
rect 1086 -2562 1092 -2556
rect 1086 -2568 1092 -2562
rect 1086 -2574 1092 -2568
rect 1086 -2580 1092 -2574
rect 1086 -2586 1092 -2580
rect 1086 -2592 1092 -2586
rect 1086 -2598 1092 -2592
rect 1086 -2604 1092 -2598
rect 1086 -2610 1092 -2604
rect 1086 -2616 1092 -2610
rect 1086 -2622 1092 -2616
rect 1086 -2628 1092 -2622
rect 1086 -2634 1092 -2628
rect 1086 -2640 1092 -2634
rect 1086 -2646 1092 -2640
rect 1086 -2652 1092 -2646
rect 1086 -2658 1092 -2652
rect 1086 -2664 1092 -2658
rect 1086 -2670 1092 -2664
rect 1086 -2676 1092 -2670
rect 1086 -2682 1092 -2676
rect 1086 -2688 1092 -2682
rect 1086 -2694 1092 -2688
rect 1086 -2700 1092 -2694
rect 1086 -2706 1092 -2700
rect 1086 -2712 1092 -2706
rect 1086 -2718 1092 -2712
rect 1086 -2724 1092 -2718
rect 1086 -2730 1092 -2724
rect 1086 -2736 1092 -2730
rect 1086 -2742 1092 -2736
rect 1086 -2748 1092 -2742
rect 1086 -2754 1092 -2748
rect 1086 -2760 1092 -2754
rect 1086 -2766 1092 -2760
rect 1086 -2772 1092 -2766
rect 1086 -2778 1092 -2772
rect 1086 -2784 1092 -2778
rect 1086 -2880 1092 -2874
rect 1086 -2886 1092 -2880
rect 1086 -2892 1092 -2886
rect 1086 -2898 1092 -2892
rect 1086 -2904 1092 -2898
rect 1086 -2910 1092 -2904
rect 1086 -2916 1092 -2910
rect 1086 -2922 1092 -2916
rect 1086 -2928 1092 -2922
rect 1086 -2934 1092 -2928
rect 1086 -2940 1092 -2934
rect 1086 -2946 1092 -2940
rect 1086 -2952 1092 -2946
rect 1086 -2958 1092 -2952
rect 1086 -2964 1092 -2958
rect 1086 -2970 1092 -2964
rect 1086 -2976 1092 -2970
rect 1086 -2982 1092 -2976
rect 1086 -2988 1092 -2982
rect 1086 -2994 1092 -2988
rect 1086 -3000 1092 -2994
rect 1086 -3006 1092 -3000
rect 1086 -3012 1092 -3006
rect 1086 -3018 1092 -3012
rect 1086 -3024 1092 -3018
rect 1086 -3030 1092 -3024
rect 1086 -3036 1092 -3030
rect 1086 -3042 1092 -3036
rect 1086 -3048 1092 -3042
rect 1086 -3054 1092 -3048
rect 1086 -3060 1092 -3054
rect 1086 -3066 1092 -3060
rect 1086 -3072 1092 -3066
rect 1086 -3078 1092 -3072
rect 1086 -3084 1092 -3078
rect 1086 -3090 1092 -3084
rect 1086 -3096 1092 -3090
rect 1086 -3102 1092 -3096
rect 1086 -3108 1092 -3102
rect 1086 -3180 1092 -3174
rect 1086 -3186 1092 -3180
rect 1086 -3192 1092 -3186
rect 1086 -3198 1092 -3192
rect 1086 -3204 1092 -3198
rect 1086 -3210 1092 -3204
rect 1086 -3216 1092 -3210
rect 1086 -3222 1092 -3216
rect 1086 -3228 1092 -3222
rect 1086 -3234 1092 -3228
rect 1086 -3240 1092 -3234
rect 1086 -3246 1092 -3240
rect 1086 -3252 1092 -3246
rect 1086 -3258 1092 -3252
rect 1086 -3264 1092 -3258
rect 1086 -3270 1092 -3264
rect 1086 -3276 1092 -3270
rect 1086 -3282 1092 -3276
rect 1086 -3324 1092 -3318
rect 1086 -3330 1092 -3324
rect 1086 -3336 1092 -3330
rect 1086 -3342 1092 -3336
rect 1086 -3348 1092 -3342
rect 1086 -3354 1092 -3348
rect 1086 -3360 1092 -3354
rect 1086 -3366 1092 -3360
rect 1086 -3372 1092 -3366
rect 1086 -3378 1092 -3372
rect 1086 -3384 1092 -3378
rect 1086 -3390 1092 -3384
rect 1086 -3396 1092 -3390
rect 1086 -3402 1092 -3396
rect 1086 -3408 1092 -3402
rect 1086 -3414 1092 -3408
rect 1086 -3420 1092 -3414
rect 1086 -3426 1092 -3420
rect 1086 -3432 1092 -3426
rect 1086 -3438 1092 -3432
rect 1086 -3444 1092 -3438
rect 1086 -3450 1092 -3444
rect 1086 -3456 1092 -3450
rect 1086 -3462 1092 -3456
rect 1086 -3468 1092 -3462
rect 1086 -3474 1092 -3468
rect 1086 -3480 1092 -3474
rect 1086 -3486 1092 -3480
rect 1086 -3492 1092 -3486
rect 1086 -3498 1092 -3492
rect 1086 -3504 1092 -3498
rect 1086 -3510 1092 -3504
rect 1092 -1110 1098 -1104
rect 1092 -1116 1098 -1110
rect 1092 -1122 1098 -1116
rect 1092 -1128 1098 -1122
rect 1092 -1134 1098 -1128
rect 1092 -1140 1098 -1134
rect 1092 -1146 1098 -1140
rect 1092 -1152 1098 -1146
rect 1092 -1158 1098 -1152
rect 1092 -1164 1098 -1158
rect 1092 -1170 1098 -1164
rect 1092 -1176 1098 -1170
rect 1092 -1182 1098 -1176
rect 1092 -1188 1098 -1182
rect 1092 -1194 1098 -1188
rect 1092 -1200 1098 -1194
rect 1092 -1206 1098 -1200
rect 1092 -1212 1098 -1206
rect 1092 -1218 1098 -1212
rect 1092 -1224 1098 -1218
rect 1092 -1230 1098 -1224
rect 1092 -1236 1098 -1230
rect 1092 -1242 1098 -1236
rect 1092 -1248 1098 -1242
rect 1092 -1254 1098 -1248
rect 1092 -1260 1098 -1254
rect 1092 -1266 1098 -1260
rect 1092 -1272 1098 -1266
rect 1092 -1278 1098 -1272
rect 1092 -1284 1098 -1278
rect 1092 -1290 1098 -1284
rect 1092 -1296 1098 -1290
rect 1092 -1302 1098 -1296
rect 1092 -1308 1098 -1302
rect 1092 -1314 1098 -1308
rect 1092 -2112 1098 -2106
rect 1092 -2118 1098 -2112
rect 1092 -2124 1098 -2118
rect 1092 -2130 1098 -2124
rect 1092 -2136 1098 -2130
rect 1092 -2142 1098 -2136
rect 1092 -2148 1098 -2142
rect 1092 -2154 1098 -2148
rect 1092 -2160 1098 -2154
rect 1092 -2166 1098 -2160
rect 1092 -2172 1098 -2166
rect 1092 -2178 1098 -2172
rect 1092 -2184 1098 -2178
rect 1092 -2190 1098 -2184
rect 1092 -2196 1098 -2190
rect 1092 -2202 1098 -2196
rect 1092 -2208 1098 -2202
rect 1092 -2214 1098 -2208
rect 1092 -2220 1098 -2214
rect 1092 -2226 1098 -2220
rect 1092 -2232 1098 -2226
rect 1092 -2238 1098 -2232
rect 1092 -2244 1098 -2238
rect 1092 -2250 1098 -2244
rect 1092 -2256 1098 -2250
rect 1092 -2262 1098 -2256
rect 1092 -2268 1098 -2262
rect 1092 -2274 1098 -2268
rect 1092 -2280 1098 -2274
rect 1092 -2286 1098 -2280
rect 1092 -2292 1098 -2286
rect 1092 -2298 1098 -2292
rect 1092 -2304 1098 -2298
rect 1092 -2310 1098 -2304
rect 1092 -2316 1098 -2310
rect 1092 -2322 1098 -2316
rect 1092 -2328 1098 -2322
rect 1092 -2334 1098 -2328
rect 1092 -2340 1098 -2334
rect 1092 -2346 1098 -2340
rect 1092 -2352 1098 -2346
rect 1092 -2358 1098 -2352
rect 1092 -2364 1098 -2358
rect 1092 -2370 1098 -2364
rect 1092 -2376 1098 -2370
rect 1092 -2382 1098 -2376
rect 1092 -2388 1098 -2382
rect 1092 -2394 1098 -2388
rect 1092 -2400 1098 -2394
rect 1092 -2406 1098 -2400
rect 1092 -2412 1098 -2406
rect 1092 -2418 1098 -2412
rect 1092 -2424 1098 -2418
rect 1092 -2430 1098 -2424
rect 1092 -2436 1098 -2430
rect 1092 -2442 1098 -2436
rect 1092 -2448 1098 -2442
rect 1092 -2454 1098 -2448
rect 1092 -2460 1098 -2454
rect 1092 -2466 1098 -2460
rect 1092 -2472 1098 -2466
rect 1092 -2478 1098 -2472
rect 1092 -2484 1098 -2478
rect 1092 -2490 1098 -2484
rect 1092 -2496 1098 -2490
rect 1092 -2502 1098 -2496
rect 1092 -2508 1098 -2502
rect 1092 -2514 1098 -2508
rect 1092 -2520 1098 -2514
rect 1092 -2526 1098 -2520
rect 1092 -2532 1098 -2526
rect 1092 -2538 1098 -2532
rect 1092 -2544 1098 -2538
rect 1092 -2550 1098 -2544
rect 1092 -2556 1098 -2550
rect 1092 -2562 1098 -2556
rect 1092 -2568 1098 -2562
rect 1092 -2574 1098 -2568
rect 1092 -2580 1098 -2574
rect 1092 -2586 1098 -2580
rect 1092 -2592 1098 -2586
rect 1092 -2598 1098 -2592
rect 1092 -2604 1098 -2598
rect 1092 -2610 1098 -2604
rect 1092 -2616 1098 -2610
rect 1092 -2622 1098 -2616
rect 1092 -2628 1098 -2622
rect 1092 -2634 1098 -2628
rect 1092 -2640 1098 -2634
rect 1092 -2646 1098 -2640
rect 1092 -2652 1098 -2646
rect 1092 -2658 1098 -2652
rect 1092 -2664 1098 -2658
rect 1092 -2670 1098 -2664
rect 1092 -2676 1098 -2670
rect 1092 -2682 1098 -2676
rect 1092 -2688 1098 -2682
rect 1092 -2694 1098 -2688
rect 1092 -2700 1098 -2694
rect 1092 -2706 1098 -2700
rect 1092 -2712 1098 -2706
rect 1092 -2718 1098 -2712
rect 1092 -2724 1098 -2718
rect 1092 -2730 1098 -2724
rect 1092 -2736 1098 -2730
rect 1092 -2742 1098 -2736
rect 1092 -2748 1098 -2742
rect 1092 -2754 1098 -2748
rect 1092 -2760 1098 -2754
rect 1092 -2766 1098 -2760
rect 1092 -2772 1098 -2766
rect 1092 -2874 1098 -2868
rect 1092 -2880 1098 -2874
rect 1092 -2886 1098 -2880
rect 1092 -2892 1098 -2886
rect 1092 -2898 1098 -2892
rect 1092 -2904 1098 -2898
rect 1092 -2910 1098 -2904
rect 1092 -2916 1098 -2910
rect 1092 -2922 1098 -2916
rect 1092 -2928 1098 -2922
rect 1092 -2934 1098 -2928
rect 1092 -2940 1098 -2934
rect 1092 -2946 1098 -2940
rect 1092 -2952 1098 -2946
rect 1092 -2958 1098 -2952
rect 1092 -2964 1098 -2958
rect 1092 -2970 1098 -2964
rect 1092 -2976 1098 -2970
rect 1092 -2982 1098 -2976
rect 1092 -2988 1098 -2982
rect 1092 -2994 1098 -2988
rect 1092 -3000 1098 -2994
rect 1092 -3006 1098 -3000
rect 1092 -3012 1098 -3006
rect 1092 -3018 1098 -3012
rect 1092 -3024 1098 -3018
rect 1092 -3030 1098 -3024
rect 1092 -3036 1098 -3030
rect 1092 -3042 1098 -3036
rect 1092 -3048 1098 -3042
rect 1092 -3054 1098 -3048
rect 1092 -3060 1098 -3054
rect 1092 -3066 1098 -3060
rect 1092 -3072 1098 -3066
rect 1092 -3078 1098 -3072
rect 1092 -3084 1098 -3078
rect 1092 -3090 1098 -3084
rect 1092 -3096 1098 -3090
rect 1092 -3102 1098 -3096
rect 1092 -3174 1098 -3168
rect 1092 -3180 1098 -3174
rect 1092 -3186 1098 -3180
rect 1092 -3192 1098 -3186
rect 1092 -3198 1098 -3192
rect 1092 -3204 1098 -3198
rect 1092 -3210 1098 -3204
rect 1092 -3216 1098 -3210
rect 1092 -3222 1098 -3216
rect 1092 -3228 1098 -3222
rect 1092 -3234 1098 -3228
rect 1092 -3240 1098 -3234
rect 1092 -3246 1098 -3240
rect 1092 -3252 1098 -3246
rect 1092 -3258 1098 -3252
rect 1092 -3264 1098 -3258
rect 1092 -3270 1098 -3264
rect 1092 -3276 1098 -3270
rect 1092 -3282 1098 -3276
rect 1092 -3318 1098 -3312
rect 1092 -3324 1098 -3318
rect 1092 -3330 1098 -3324
rect 1092 -3336 1098 -3330
rect 1092 -3342 1098 -3336
rect 1092 -3348 1098 -3342
rect 1092 -3354 1098 -3348
rect 1092 -3360 1098 -3354
rect 1092 -3366 1098 -3360
rect 1092 -3372 1098 -3366
rect 1092 -3378 1098 -3372
rect 1092 -3384 1098 -3378
rect 1092 -3390 1098 -3384
rect 1092 -3396 1098 -3390
rect 1092 -3402 1098 -3396
rect 1092 -3408 1098 -3402
rect 1092 -3414 1098 -3408
rect 1092 -3420 1098 -3414
rect 1092 -3426 1098 -3420
rect 1092 -3432 1098 -3426
rect 1092 -3438 1098 -3432
rect 1092 -3444 1098 -3438
rect 1092 -3450 1098 -3444
rect 1092 -3456 1098 -3450
rect 1092 -3462 1098 -3456
rect 1092 -3468 1098 -3462
rect 1092 -3474 1098 -3468
rect 1092 -3480 1098 -3474
rect 1092 -3486 1098 -3480
rect 1092 -3492 1098 -3486
rect 1092 -3498 1098 -3492
rect 1092 -3504 1098 -3498
rect 1092 -3510 1098 -3504
rect 1098 -1110 1104 -1104
rect 1098 -1116 1104 -1110
rect 1098 -1122 1104 -1116
rect 1098 -1128 1104 -1122
rect 1098 -1134 1104 -1128
rect 1098 -1140 1104 -1134
rect 1098 -1146 1104 -1140
rect 1098 -1152 1104 -1146
rect 1098 -1158 1104 -1152
rect 1098 -1164 1104 -1158
rect 1098 -1170 1104 -1164
rect 1098 -1176 1104 -1170
rect 1098 -1182 1104 -1176
rect 1098 -1188 1104 -1182
rect 1098 -1194 1104 -1188
rect 1098 -1200 1104 -1194
rect 1098 -1206 1104 -1200
rect 1098 -1212 1104 -1206
rect 1098 -1218 1104 -1212
rect 1098 -1224 1104 -1218
rect 1098 -1230 1104 -1224
rect 1098 -1236 1104 -1230
rect 1098 -1242 1104 -1236
rect 1098 -1248 1104 -1242
rect 1098 -1254 1104 -1248
rect 1098 -1260 1104 -1254
rect 1098 -1266 1104 -1260
rect 1098 -1272 1104 -1266
rect 1098 -1278 1104 -1272
rect 1098 -1284 1104 -1278
rect 1098 -1290 1104 -1284
rect 1098 -1296 1104 -1290
rect 1098 -1302 1104 -1296
rect 1098 -1308 1104 -1302
rect 1098 -1314 1104 -1308
rect 1098 -2094 1104 -2088
rect 1098 -2100 1104 -2094
rect 1098 -2106 1104 -2100
rect 1098 -2112 1104 -2106
rect 1098 -2118 1104 -2112
rect 1098 -2124 1104 -2118
rect 1098 -2130 1104 -2124
rect 1098 -2136 1104 -2130
rect 1098 -2142 1104 -2136
rect 1098 -2148 1104 -2142
rect 1098 -2154 1104 -2148
rect 1098 -2160 1104 -2154
rect 1098 -2166 1104 -2160
rect 1098 -2172 1104 -2166
rect 1098 -2178 1104 -2172
rect 1098 -2184 1104 -2178
rect 1098 -2190 1104 -2184
rect 1098 -2196 1104 -2190
rect 1098 -2202 1104 -2196
rect 1098 -2208 1104 -2202
rect 1098 -2214 1104 -2208
rect 1098 -2220 1104 -2214
rect 1098 -2226 1104 -2220
rect 1098 -2232 1104 -2226
rect 1098 -2238 1104 -2232
rect 1098 -2244 1104 -2238
rect 1098 -2250 1104 -2244
rect 1098 -2256 1104 -2250
rect 1098 -2262 1104 -2256
rect 1098 -2268 1104 -2262
rect 1098 -2274 1104 -2268
rect 1098 -2280 1104 -2274
rect 1098 -2286 1104 -2280
rect 1098 -2292 1104 -2286
rect 1098 -2298 1104 -2292
rect 1098 -2304 1104 -2298
rect 1098 -2310 1104 -2304
rect 1098 -2316 1104 -2310
rect 1098 -2322 1104 -2316
rect 1098 -2328 1104 -2322
rect 1098 -2334 1104 -2328
rect 1098 -2340 1104 -2334
rect 1098 -2346 1104 -2340
rect 1098 -2352 1104 -2346
rect 1098 -2358 1104 -2352
rect 1098 -2364 1104 -2358
rect 1098 -2370 1104 -2364
rect 1098 -2376 1104 -2370
rect 1098 -2382 1104 -2376
rect 1098 -2388 1104 -2382
rect 1098 -2394 1104 -2388
rect 1098 -2400 1104 -2394
rect 1098 -2406 1104 -2400
rect 1098 -2412 1104 -2406
rect 1098 -2418 1104 -2412
rect 1098 -2424 1104 -2418
rect 1098 -2430 1104 -2424
rect 1098 -2436 1104 -2430
rect 1098 -2442 1104 -2436
rect 1098 -2448 1104 -2442
rect 1098 -2454 1104 -2448
rect 1098 -2460 1104 -2454
rect 1098 -2466 1104 -2460
rect 1098 -2472 1104 -2466
rect 1098 -2478 1104 -2472
rect 1098 -2484 1104 -2478
rect 1098 -2490 1104 -2484
rect 1098 -2496 1104 -2490
rect 1098 -2502 1104 -2496
rect 1098 -2508 1104 -2502
rect 1098 -2514 1104 -2508
rect 1098 -2520 1104 -2514
rect 1098 -2526 1104 -2520
rect 1098 -2532 1104 -2526
rect 1098 -2538 1104 -2532
rect 1098 -2544 1104 -2538
rect 1098 -2550 1104 -2544
rect 1098 -2556 1104 -2550
rect 1098 -2562 1104 -2556
rect 1098 -2568 1104 -2562
rect 1098 -2574 1104 -2568
rect 1098 -2580 1104 -2574
rect 1098 -2586 1104 -2580
rect 1098 -2592 1104 -2586
rect 1098 -2598 1104 -2592
rect 1098 -2604 1104 -2598
rect 1098 -2610 1104 -2604
rect 1098 -2616 1104 -2610
rect 1098 -2622 1104 -2616
rect 1098 -2628 1104 -2622
rect 1098 -2634 1104 -2628
rect 1098 -2640 1104 -2634
rect 1098 -2646 1104 -2640
rect 1098 -2652 1104 -2646
rect 1098 -2658 1104 -2652
rect 1098 -2664 1104 -2658
rect 1098 -2670 1104 -2664
rect 1098 -2676 1104 -2670
rect 1098 -2682 1104 -2676
rect 1098 -2688 1104 -2682
rect 1098 -2694 1104 -2688
rect 1098 -2700 1104 -2694
rect 1098 -2706 1104 -2700
rect 1098 -2712 1104 -2706
rect 1098 -2718 1104 -2712
rect 1098 -2724 1104 -2718
rect 1098 -2730 1104 -2724
rect 1098 -2736 1104 -2730
rect 1098 -2742 1104 -2736
rect 1098 -2748 1104 -2742
rect 1098 -2754 1104 -2748
rect 1098 -2760 1104 -2754
rect 1098 -2766 1104 -2760
rect 1098 -2862 1104 -2856
rect 1098 -2868 1104 -2862
rect 1098 -2874 1104 -2868
rect 1098 -2880 1104 -2874
rect 1098 -2886 1104 -2880
rect 1098 -2892 1104 -2886
rect 1098 -2898 1104 -2892
rect 1098 -2904 1104 -2898
rect 1098 -2910 1104 -2904
rect 1098 -2916 1104 -2910
rect 1098 -2922 1104 -2916
rect 1098 -2928 1104 -2922
rect 1098 -2934 1104 -2928
rect 1098 -2940 1104 -2934
rect 1098 -2946 1104 -2940
rect 1098 -2952 1104 -2946
rect 1098 -2958 1104 -2952
rect 1098 -2964 1104 -2958
rect 1098 -2970 1104 -2964
rect 1098 -2976 1104 -2970
rect 1098 -2982 1104 -2976
rect 1098 -2988 1104 -2982
rect 1098 -2994 1104 -2988
rect 1098 -3000 1104 -2994
rect 1098 -3006 1104 -3000
rect 1098 -3012 1104 -3006
rect 1098 -3018 1104 -3012
rect 1098 -3024 1104 -3018
rect 1098 -3030 1104 -3024
rect 1098 -3036 1104 -3030
rect 1098 -3042 1104 -3036
rect 1098 -3048 1104 -3042
rect 1098 -3054 1104 -3048
rect 1098 -3060 1104 -3054
rect 1098 -3066 1104 -3060
rect 1098 -3072 1104 -3066
rect 1098 -3078 1104 -3072
rect 1098 -3084 1104 -3078
rect 1098 -3090 1104 -3084
rect 1098 -3096 1104 -3090
rect 1098 -3102 1104 -3096
rect 1098 -3168 1104 -3162
rect 1098 -3174 1104 -3168
rect 1098 -3180 1104 -3174
rect 1098 -3186 1104 -3180
rect 1098 -3192 1104 -3186
rect 1098 -3198 1104 -3192
rect 1098 -3204 1104 -3198
rect 1098 -3210 1104 -3204
rect 1098 -3216 1104 -3210
rect 1098 -3222 1104 -3216
rect 1098 -3228 1104 -3222
rect 1098 -3234 1104 -3228
rect 1098 -3240 1104 -3234
rect 1098 -3246 1104 -3240
rect 1098 -3252 1104 -3246
rect 1098 -3258 1104 -3252
rect 1098 -3264 1104 -3258
rect 1098 -3270 1104 -3264
rect 1098 -3276 1104 -3270
rect 1098 -3318 1104 -3312
rect 1098 -3324 1104 -3318
rect 1098 -3330 1104 -3324
rect 1098 -3336 1104 -3330
rect 1098 -3342 1104 -3336
rect 1098 -3348 1104 -3342
rect 1098 -3354 1104 -3348
rect 1098 -3360 1104 -3354
rect 1098 -3366 1104 -3360
rect 1098 -3372 1104 -3366
rect 1098 -3378 1104 -3372
rect 1098 -3384 1104 -3378
rect 1098 -3390 1104 -3384
rect 1098 -3396 1104 -3390
rect 1098 -3402 1104 -3396
rect 1098 -3408 1104 -3402
rect 1098 -3414 1104 -3408
rect 1098 -3420 1104 -3414
rect 1098 -3426 1104 -3420
rect 1098 -3432 1104 -3426
rect 1098 -3438 1104 -3432
rect 1098 -3444 1104 -3438
rect 1098 -3450 1104 -3444
rect 1098 -3456 1104 -3450
rect 1098 -3462 1104 -3456
rect 1098 -3468 1104 -3462
rect 1098 -3474 1104 -3468
rect 1098 -3480 1104 -3474
rect 1098 -3486 1104 -3480
rect 1098 -3492 1104 -3486
rect 1098 -3498 1104 -3492
rect 1098 -3504 1104 -3498
rect 1098 -3510 1104 -3504
rect 1104 -1110 1110 -1104
rect 1104 -1116 1110 -1110
rect 1104 -1122 1110 -1116
rect 1104 -1128 1110 -1122
rect 1104 -1134 1110 -1128
rect 1104 -1140 1110 -1134
rect 1104 -1146 1110 -1140
rect 1104 -1152 1110 -1146
rect 1104 -1158 1110 -1152
rect 1104 -1164 1110 -1158
rect 1104 -1170 1110 -1164
rect 1104 -1176 1110 -1170
rect 1104 -1182 1110 -1176
rect 1104 -1188 1110 -1182
rect 1104 -1194 1110 -1188
rect 1104 -1200 1110 -1194
rect 1104 -1206 1110 -1200
rect 1104 -1212 1110 -1206
rect 1104 -1218 1110 -1212
rect 1104 -1224 1110 -1218
rect 1104 -1230 1110 -1224
rect 1104 -1236 1110 -1230
rect 1104 -1242 1110 -1236
rect 1104 -1248 1110 -1242
rect 1104 -1254 1110 -1248
rect 1104 -1260 1110 -1254
rect 1104 -1266 1110 -1260
rect 1104 -1272 1110 -1266
rect 1104 -1278 1110 -1272
rect 1104 -1284 1110 -1278
rect 1104 -1290 1110 -1284
rect 1104 -1296 1110 -1290
rect 1104 -1302 1110 -1296
rect 1104 -1308 1110 -1302
rect 1104 -1314 1110 -1308
rect 1104 -2076 1110 -2070
rect 1104 -2082 1110 -2076
rect 1104 -2088 1110 -2082
rect 1104 -2094 1110 -2088
rect 1104 -2100 1110 -2094
rect 1104 -2106 1110 -2100
rect 1104 -2112 1110 -2106
rect 1104 -2118 1110 -2112
rect 1104 -2124 1110 -2118
rect 1104 -2130 1110 -2124
rect 1104 -2136 1110 -2130
rect 1104 -2142 1110 -2136
rect 1104 -2148 1110 -2142
rect 1104 -2154 1110 -2148
rect 1104 -2160 1110 -2154
rect 1104 -2166 1110 -2160
rect 1104 -2172 1110 -2166
rect 1104 -2178 1110 -2172
rect 1104 -2184 1110 -2178
rect 1104 -2190 1110 -2184
rect 1104 -2196 1110 -2190
rect 1104 -2202 1110 -2196
rect 1104 -2208 1110 -2202
rect 1104 -2214 1110 -2208
rect 1104 -2220 1110 -2214
rect 1104 -2226 1110 -2220
rect 1104 -2232 1110 -2226
rect 1104 -2238 1110 -2232
rect 1104 -2244 1110 -2238
rect 1104 -2250 1110 -2244
rect 1104 -2256 1110 -2250
rect 1104 -2262 1110 -2256
rect 1104 -2268 1110 -2262
rect 1104 -2274 1110 -2268
rect 1104 -2280 1110 -2274
rect 1104 -2286 1110 -2280
rect 1104 -2292 1110 -2286
rect 1104 -2298 1110 -2292
rect 1104 -2304 1110 -2298
rect 1104 -2310 1110 -2304
rect 1104 -2316 1110 -2310
rect 1104 -2322 1110 -2316
rect 1104 -2328 1110 -2322
rect 1104 -2334 1110 -2328
rect 1104 -2340 1110 -2334
rect 1104 -2346 1110 -2340
rect 1104 -2352 1110 -2346
rect 1104 -2358 1110 -2352
rect 1104 -2364 1110 -2358
rect 1104 -2370 1110 -2364
rect 1104 -2376 1110 -2370
rect 1104 -2382 1110 -2376
rect 1104 -2388 1110 -2382
rect 1104 -2394 1110 -2388
rect 1104 -2400 1110 -2394
rect 1104 -2406 1110 -2400
rect 1104 -2412 1110 -2406
rect 1104 -2418 1110 -2412
rect 1104 -2424 1110 -2418
rect 1104 -2430 1110 -2424
rect 1104 -2436 1110 -2430
rect 1104 -2442 1110 -2436
rect 1104 -2448 1110 -2442
rect 1104 -2454 1110 -2448
rect 1104 -2460 1110 -2454
rect 1104 -2466 1110 -2460
rect 1104 -2472 1110 -2466
rect 1104 -2478 1110 -2472
rect 1104 -2484 1110 -2478
rect 1104 -2490 1110 -2484
rect 1104 -2496 1110 -2490
rect 1104 -2502 1110 -2496
rect 1104 -2508 1110 -2502
rect 1104 -2514 1110 -2508
rect 1104 -2520 1110 -2514
rect 1104 -2526 1110 -2520
rect 1104 -2532 1110 -2526
rect 1104 -2538 1110 -2532
rect 1104 -2544 1110 -2538
rect 1104 -2550 1110 -2544
rect 1104 -2556 1110 -2550
rect 1104 -2562 1110 -2556
rect 1104 -2568 1110 -2562
rect 1104 -2574 1110 -2568
rect 1104 -2580 1110 -2574
rect 1104 -2586 1110 -2580
rect 1104 -2592 1110 -2586
rect 1104 -2598 1110 -2592
rect 1104 -2604 1110 -2598
rect 1104 -2610 1110 -2604
rect 1104 -2616 1110 -2610
rect 1104 -2622 1110 -2616
rect 1104 -2628 1110 -2622
rect 1104 -2634 1110 -2628
rect 1104 -2640 1110 -2634
rect 1104 -2646 1110 -2640
rect 1104 -2652 1110 -2646
rect 1104 -2658 1110 -2652
rect 1104 -2664 1110 -2658
rect 1104 -2670 1110 -2664
rect 1104 -2676 1110 -2670
rect 1104 -2682 1110 -2676
rect 1104 -2688 1110 -2682
rect 1104 -2694 1110 -2688
rect 1104 -2700 1110 -2694
rect 1104 -2706 1110 -2700
rect 1104 -2712 1110 -2706
rect 1104 -2718 1110 -2712
rect 1104 -2724 1110 -2718
rect 1104 -2730 1110 -2724
rect 1104 -2736 1110 -2730
rect 1104 -2742 1110 -2736
rect 1104 -2748 1110 -2742
rect 1104 -2754 1110 -2748
rect 1104 -2850 1110 -2844
rect 1104 -2856 1110 -2850
rect 1104 -2862 1110 -2856
rect 1104 -2868 1110 -2862
rect 1104 -2874 1110 -2868
rect 1104 -2880 1110 -2874
rect 1104 -2886 1110 -2880
rect 1104 -2892 1110 -2886
rect 1104 -2898 1110 -2892
rect 1104 -2904 1110 -2898
rect 1104 -2910 1110 -2904
rect 1104 -2916 1110 -2910
rect 1104 -2922 1110 -2916
rect 1104 -2928 1110 -2922
rect 1104 -2934 1110 -2928
rect 1104 -2940 1110 -2934
rect 1104 -2946 1110 -2940
rect 1104 -2952 1110 -2946
rect 1104 -2958 1110 -2952
rect 1104 -2964 1110 -2958
rect 1104 -2970 1110 -2964
rect 1104 -2976 1110 -2970
rect 1104 -2982 1110 -2976
rect 1104 -2988 1110 -2982
rect 1104 -2994 1110 -2988
rect 1104 -3000 1110 -2994
rect 1104 -3006 1110 -3000
rect 1104 -3012 1110 -3006
rect 1104 -3018 1110 -3012
rect 1104 -3024 1110 -3018
rect 1104 -3030 1110 -3024
rect 1104 -3036 1110 -3030
rect 1104 -3042 1110 -3036
rect 1104 -3048 1110 -3042
rect 1104 -3054 1110 -3048
rect 1104 -3060 1110 -3054
rect 1104 -3066 1110 -3060
rect 1104 -3072 1110 -3066
rect 1104 -3078 1110 -3072
rect 1104 -3084 1110 -3078
rect 1104 -3090 1110 -3084
rect 1104 -3096 1110 -3090
rect 1104 -3168 1110 -3162
rect 1104 -3174 1110 -3168
rect 1104 -3180 1110 -3174
rect 1104 -3186 1110 -3180
rect 1104 -3192 1110 -3186
rect 1104 -3198 1110 -3192
rect 1104 -3204 1110 -3198
rect 1104 -3210 1110 -3204
rect 1104 -3216 1110 -3210
rect 1104 -3222 1110 -3216
rect 1104 -3228 1110 -3222
rect 1104 -3234 1110 -3228
rect 1104 -3240 1110 -3234
rect 1104 -3246 1110 -3240
rect 1104 -3252 1110 -3246
rect 1104 -3258 1110 -3252
rect 1104 -3264 1110 -3258
rect 1104 -3270 1110 -3264
rect 1104 -3276 1110 -3270
rect 1104 -3318 1110 -3312
rect 1104 -3324 1110 -3318
rect 1104 -3330 1110 -3324
rect 1104 -3336 1110 -3330
rect 1104 -3342 1110 -3336
rect 1104 -3348 1110 -3342
rect 1104 -3354 1110 -3348
rect 1104 -3360 1110 -3354
rect 1104 -3366 1110 -3360
rect 1104 -3372 1110 -3366
rect 1104 -3378 1110 -3372
rect 1104 -3384 1110 -3378
rect 1104 -3390 1110 -3384
rect 1104 -3396 1110 -3390
rect 1104 -3402 1110 -3396
rect 1104 -3408 1110 -3402
rect 1104 -3414 1110 -3408
rect 1104 -3420 1110 -3414
rect 1104 -3426 1110 -3420
rect 1104 -3432 1110 -3426
rect 1104 -3438 1110 -3432
rect 1104 -3444 1110 -3438
rect 1104 -3450 1110 -3444
rect 1104 -3456 1110 -3450
rect 1104 -3462 1110 -3456
rect 1104 -3468 1110 -3462
rect 1104 -3474 1110 -3468
rect 1104 -3480 1110 -3474
rect 1104 -3486 1110 -3480
rect 1104 -3492 1110 -3486
rect 1104 -3498 1110 -3492
rect 1104 -3504 1110 -3498
rect 1104 -3510 1110 -3504
rect 1110 -1110 1116 -1104
rect 1110 -1116 1116 -1110
rect 1110 -1122 1116 -1116
rect 1110 -1128 1116 -1122
rect 1110 -1134 1116 -1128
rect 1110 -1140 1116 -1134
rect 1110 -1146 1116 -1140
rect 1110 -1152 1116 -1146
rect 1110 -1158 1116 -1152
rect 1110 -1164 1116 -1158
rect 1110 -1170 1116 -1164
rect 1110 -1176 1116 -1170
rect 1110 -1182 1116 -1176
rect 1110 -1188 1116 -1182
rect 1110 -1194 1116 -1188
rect 1110 -1200 1116 -1194
rect 1110 -1206 1116 -1200
rect 1110 -1212 1116 -1206
rect 1110 -1218 1116 -1212
rect 1110 -1224 1116 -1218
rect 1110 -1230 1116 -1224
rect 1110 -1236 1116 -1230
rect 1110 -1242 1116 -1236
rect 1110 -1248 1116 -1242
rect 1110 -1254 1116 -1248
rect 1110 -1260 1116 -1254
rect 1110 -1266 1116 -1260
rect 1110 -1272 1116 -1266
rect 1110 -1278 1116 -1272
rect 1110 -1284 1116 -1278
rect 1110 -1290 1116 -1284
rect 1110 -1296 1116 -1290
rect 1110 -1302 1116 -1296
rect 1110 -1308 1116 -1302
rect 1110 -1314 1116 -1308
rect 1110 -2058 1116 -2052
rect 1110 -2064 1116 -2058
rect 1110 -2070 1116 -2064
rect 1110 -2076 1116 -2070
rect 1110 -2082 1116 -2076
rect 1110 -2088 1116 -2082
rect 1110 -2094 1116 -2088
rect 1110 -2100 1116 -2094
rect 1110 -2106 1116 -2100
rect 1110 -2112 1116 -2106
rect 1110 -2118 1116 -2112
rect 1110 -2124 1116 -2118
rect 1110 -2130 1116 -2124
rect 1110 -2136 1116 -2130
rect 1110 -2142 1116 -2136
rect 1110 -2148 1116 -2142
rect 1110 -2154 1116 -2148
rect 1110 -2160 1116 -2154
rect 1110 -2166 1116 -2160
rect 1110 -2172 1116 -2166
rect 1110 -2178 1116 -2172
rect 1110 -2184 1116 -2178
rect 1110 -2190 1116 -2184
rect 1110 -2196 1116 -2190
rect 1110 -2202 1116 -2196
rect 1110 -2208 1116 -2202
rect 1110 -2214 1116 -2208
rect 1110 -2220 1116 -2214
rect 1110 -2226 1116 -2220
rect 1110 -2232 1116 -2226
rect 1110 -2238 1116 -2232
rect 1110 -2244 1116 -2238
rect 1110 -2250 1116 -2244
rect 1110 -2256 1116 -2250
rect 1110 -2262 1116 -2256
rect 1110 -2268 1116 -2262
rect 1110 -2274 1116 -2268
rect 1110 -2280 1116 -2274
rect 1110 -2286 1116 -2280
rect 1110 -2292 1116 -2286
rect 1110 -2298 1116 -2292
rect 1110 -2304 1116 -2298
rect 1110 -2310 1116 -2304
rect 1110 -2316 1116 -2310
rect 1110 -2322 1116 -2316
rect 1110 -2328 1116 -2322
rect 1110 -2334 1116 -2328
rect 1110 -2340 1116 -2334
rect 1110 -2346 1116 -2340
rect 1110 -2352 1116 -2346
rect 1110 -2358 1116 -2352
rect 1110 -2364 1116 -2358
rect 1110 -2370 1116 -2364
rect 1110 -2376 1116 -2370
rect 1110 -2382 1116 -2376
rect 1110 -2388 1116 -2382
rect 1110 -2394 1116 -2388
rect 1110 -2400 1116 -2394
rect 1110 -2406 1116 -2400
rect 1110 -2412 1116 -2406
rect 1110 -2418 1116 -2412
rect 1110 -2424 1116 -2418
rect 1110 -2430 1116 -2424
rect 1110 -2436 1116 -2430
rect 1110 -2442 1116 -2436
rect 1110 -2448 1116 -2442
rect 1110 -2454 1116 -2448
rect 1110 -2460 1116 -2454
rect 1110 -2466 1116 -2460
rect 1110 -2472 1116 -2466
rect 1110 -2478 1116 -2472
rect 1110 -2484 1116 -2478
rect 1110 -2490 1116 -2484
rect 1110 -2496 1116 -2490
rect 1110 -2502 1116 -2496
rect 1110 -2508 1116 -2502
rect 1110 -2514 1116 -2508
rect 1110 -2520 1116 -2514
rect 1110 -2526 1116 -2520
rect 1110 -2532 1116 -2526
rect 1110 -2538 1116 -2532
rect 1110 -2544 1116 -2538
rect 1110 -2550 1116 -2544
rect 1110 -2556 1116 -2550
rect 1110 -2562 1116 -2556
rect 1110 -2568 1116 -2562
rect 1110 -2574 1116 -2568
rect 1110 -2580 1116 -2574
rect 1110 -2586 1116 -2580
rect 1110 -2592 1116 -2586
rect 1110 -2598 1116 -2592
rect 1110 -2604 1116 -2598
rect 1110 -2610 1116 -2604
rect 1110 -2616 1116 -2610
rect 1110 -2622 1116 -2616
rect 1110 -2628 1116 -2622
rect 1110 -2634 1116 -2628
rect 1110 -2640 1116 -2634
rect 1110 -2646 1116 -2640
rect 1110 -2652 1116 -2646
rect 1110 -2658 1116 -2652
rect 1110 -2664 1116 -2658
rect 1110 -2670 1116 -2664
rect 1110 -2676 1116 -2670
rect 1110 -2682 1116 -2676
rect 1110 -2688 1116 -2682
rect 1110 -2694 1116 -2688
rect 1110 -2700 1116 -2694
rect 1110 -2706 1116 -2700
rect 1110 -2712 1116 -2706
rect 1110 -2718 1116 -2712
rect 1110 -2724 1116 -2718
rect 1110 -2730 1116 -2724
rect 1110 -2736 1116 -2730
rect 1110 -2742 1116 -2736
rect 1110 -2844 1116 -2838
rect 1110 -2850 1116 -2844
rect 1110 -2856 1116 -2850
rect 1110 -2862 1116 -2856
rect 1110 -2868 1116 -2862
rect 1110 -2874 1116 -2868
rect 1110 -2880 1116 -2874
rect 1110 -2886 1116 -2880
rect 1110 -2892 1116 -2886
rect 1110 -2898 1116 -2892
rect 1110 -2904 1116 -2898
rect 1110 -2910 1116 -2904
rect 1110 -2916 1116 -2910
rect 1110 -2922 1116 -2916
rect 1110 -2928 1116 -2922
rect 1110 -2934 1116 -2928
rect 1110 -2940 1116 -2934
rect 1110 -2946 1116 -2940
rect 1110 -2952 1116 -2946
rect 1110 -2958 1116 -2952
rect 1110 -2964 1116 -2958
rect 1110 -2970 1116 -2964
rect 1110 -2976 1116 -2970
rect 1110 -2982 1116 -2976
rect 1110 -2988 1116 -2982
rect 1110 -2994 1116 -2988
rect 1110 -3000 1116 -2994
rect 1110 -3006 1116 -3000
rect 1110 -3012 1116 -3006
rect 1110 -3018 1116 -3012
rect 1110 -3024 1116 -3018
rect 1110 -3030 1116 -3024
rect 1110 -3036 1116 -3030
rect 1110 -3042 1116 -3036
rect 1110 -3048 1116 -3042
rect 1110 -3054 1116 -3048
rect 1110 -3060 1116 -3054
rect 1110 -3066 1116 -3060
rect 1110 -3072 1116 -3066
rect 1110 -3078 1116 -3072
rect 1110 -3084 1116 -3078
rect 1110 -3090 1116 -3084
rect 1110 -3162 1116 -3156
rect 1110 -3168 1116 -3162
rect 1110 -3174 1116 -3168
rect 1110 -3180 1116 -3174
rect 1110 -3186 1116 -3180
rect 1110 -3192 1116 -3186
rect 1110 -3198 1116 -3192
rect 1110 -3204 1116 -3198
rect 1110 -3210 1116 -3204
rect 1110 -3216 1116 -3210
rect 1110 -3222 1116 -3216
rect 1110 -3228 1116 -3222
rect 1110 -3234 1116 -3228
rect 1110 -3240 1116 -3234
rect 1110 -3246 1116 -3240
rect 1110 -3252 1116 -3246
rect 1110 -3258 1116 -3252
rect 1110 -3264 1116 -3258
rect 1110 -3270 1116 -3264
rect 1110 -3318 1116 -3312
rect 1110 -3324 1116 -3318
rect 1110 -3330 1116 -3324
rect 1110 -3336 1116 -3330
rect 1110 -3342 1116 -3336
rect 1110 -3348 1116 -3342
rect 1110 -3354 1116 -3348
rect 1110 -3360 1116 -3354
rect 1110 -3366 1116 -3360
rect 1110 -3372 1116 -3366
rect 1110 -3378 1116 -3372
rect 1110 -3384 1116 -3378
rect 1110 -3390 1116 -3384
rect 1110 -3396 1116 -3390
rect 1110 -3402 1116 -3396
rect 1110 -3408 1116 -3402
rect 1110 -3414 1116 -3408
rect 1110 -3420 1116 -3414
rect 1110 -3426 1116 -3420
rect 1110 -3432 1116 -3426
rect 1110 -3438 1116 -3432
rect 1110 -3444 1116 -3438
rect 1110 -3450 1116 -3444
rect 1110 -3456 1116 -3450
rect 1110 -3462 1116 -3456
rect 1110 -3468 1116 -3462
rect 1110 -3474 1116 -3468
rect 1110 -3480 1116 -3474
rect 1110 -3486 1116 -3480
rect 1110 -3492 1116 -3486
rect 1110 -3498 1116 -3492
rect 1110 -3504 1116 -3498
rect 1110 -3510 1116 -3504
rect 1116 -1110 1122 -1104
rect 1116 -1116 1122 -1110
rect 1116 -1122 1122 -1116
rect 1116 -1128 1122 -1122
rect 1116 -1134 1122 -1128
rect 1116 -1140 1122 -1134
rect 1116 -1146 1122 -1140
rect 1116 -1152 1122 -1146
rect 1116 -1158 1122 -1152
rect 1116 -1164 1122 -1158
rect 1116 -1170 1122 -1164
rect 1116 -1176 1122 -1170
rect 1116 -1182 1122 -1176
rect 1116 -1188 1122 -1182
rect 1116 -1194 1122 -1188
rect 1116 -1200 1122 -1194
rect 1116 -1206 1122 -1200
rect 1116 -1212 1122 -1206
rect 1116 -1218 1122 -1212
rect 1116 -1224 1122 -1218
rect 1116 -1230 1122 -1224
rect 1116 -1236 1122 -1230
rect 1116 -1242 1122 -1236
rect 1116 -1248 1122 -1242
rect 1116 -1254 1122 -1248
rect 1116 -1260 1122 -1254
rect 1116 -1266 1122 -1260
rect 1116 -1272 1122 -1266
rect 1116 -1278 1122 -1272
rect 1116 -1284 1122 -1278
rect 1116 -1290 1122 -1284
rect 1116 -1296 1122 -1290
rect 1116 -1302 1122 -1296
rect 1116 -1308 1122 -1302
rect 1116 -2040 1122 -2034
rect 1116 -2046 1122 -2040
rect 1116 -2052 1122 -2046
rect 1116 -2058 1122 -2052
rect 1116 -2064 1122 -2058
rect 1116 -2070 1122 -2064
rect 1116 -2076 1122 -2070
rect 1116 -2082 1122 -2076
rect 1116 -2088 1122 -2082
rect 1116 -2094 1122 -2088
rect 1116 -2100 1122 -2094
rect 1116 -2106 1122 -2100
rect 1116 -2112 1122 -2106
rect 1116 -2118 1122 -2112
rect 1116 -2124 1122 -2118
rect 1116 -2130 1122 -2124
rect 1116 -2136 1122 -2130
rect 1116 -2142 1122 -2136
rect 1116 -2148 1122 -2142
rect 1116 -2154 1122 -2148
rect 1116 -2160 1122 -2154
rect 1116 -2166 1122 -2160
rect 1116 -2172 1122 -2166
rect 1116 -2178 1122 -2172
rect 1116 -2184 1122 -2178
rect 1116 -2190 1122 -2184
rect 1116 -2196 1122 -2190
rect 1116 -2202 1122 -2196
rect 1116 -2208 1122 -2202
rect 1116 -2214 1122 -2208
rect 1116 -2220 1122 -2214
rect 1116 -2226 1122 -2220
rect 1116 -2232 1122 -2226
rect 1116 -2238 1122 -2232
rect 1116 -2244 1122 -2238
rect 1116 -2250 1122 -2244
rect 1116 -2256 1122 -2250
rect 1116 -2262 1122 -2256
rect 1116 -2268 1122 -2262
rect 1116 -2274 1122 -2268
rect 1116 -2280 1122 -2274
rect 1116 -2286 1122 -2280
rect 1116 -2292 1122 -2286
rect 1116 -2298 1122 -2292
rect 1116 -2304 1122 -2298
rect 1116 -2310 1122 -2304
rect 1116 -2316 1122 -2310
rect 1116 -2322 1122 -2316
rect 1116 -2328 1122 -2322
rect 1116 -2334 1122 -2328
rect 1116 -2340 1122 -2334
rect 1116 -2346 1122 -2340
rect 1116 -2352 1122 -2346
rect 1116 -2358 1122 -2352
rect 1116 -2364 1122 -2358
rect 1116 -2370 1122 -2364
rect 1116 -2376 1122 -2370
rect 1116 -2382 1122 -2376
rect 1116 -2388 1122 -2382
rect 1116 -2394 1122 -2388
rect 1116 -2400 1122 -2394
rect 1116 -2406 1122 -2400
rect 1116 -2412 1122 -2406
rect 1116 -2418 1122 -2412
rect 1116 -2424 1122 -2418
rect 1116 -2430 1122 -2424
rect 1116 -2436 1122 -2430
rect 1116 -2442 1122 -2436
rect 1116 -2448 1122 -2442
rect 1116 -2454 1122 -2448
rect 1116 -2460 1122 -2454
rect 1116 -2466 1122 -2460
rect 1116 -2472 1122 -2466
rect 1116 -2478 1122 -2472
rect 1116 -2484 1122 -2478
rect 1116 -2490 1122 -2484
rect 1116 -2496 1122 -2490
rect 1116 -2502 1122 -2496
rect 1116 -2508 1122 -2502
rect 1116 -2514 1122 -2508
rect 1116 -2520 1122 -2514
rect 1116 -2526 1122 -2520
rect 1116 -2532 1122 -2526
rect 1116 -2538 1122 -2532
rect 1116 -2544 1122 -2538
rect 1116 -2550 1122 -2544
rect 1116 -2556 1122 -2550
rect 1116 -2562 1122 -2556
rect 1116 -2568 1122 -2562
rect 1116 -2574 1122 -2568
rect 1116 -2580 1122 -2574
rect 1116 -2586 1122 -2580
rect 1116 -2592 1122 -2586
rect 1116 -2598 1122 -2592
rect 1116 -2604 1122 -2598
rect 1116 -2610 1122 -2604
rect 1116 -2616 1122 -2610
rect 1116 -2622 1122 -2616
rect 1116 -2628 1122 -2622
rect 1116 -2634 1122 -2628
rect 1116 -2640 1122 -2634
rect 1116 -2646 1122 -2640
rect 1116 -2652 1122 -2646
rect 1116 -2658 1122 -2652
rect 1116 -2664 1122 -2658
rect 1116 -2670 1122 -2664
rect 1116 -2676 1122 -2670
rect 1116 -2682 1122 -2676
rect 1116 -2688 1122 -2682
rect 1116 -2694 1122 -2688
rect 1116 -2700 1122 -2694
rect 1116 -2706 1122 -2700
rect 1116 -2712 1122 -2706
rect 1116 -2718 1122 -2712
rect 1116 -2724 1122 -2718
rect 1116 -2730 1122 -2724
rect 1116 -2736 1122 -2730
rect 1116 -2832 1122 -2826
rect 1116 -2838 1122 -2832
rect 1116 -2844 1122 -2838
rect 1116 -2850 1122 -2844
rect 1116 -2856 1122 -2850
rect 1116 -2862 1122 -2856
rect 1116 -2868 1122 -2862
rect 1116 -2874 1122 -2868
rect 1116 -2880 1122 -2874
rect 1116 -2886 1122 -2880
rect 1116 -2892 1122 -2886
rect 1116 -2898 1122 -2892
rect 1116 -2904 1122 -2898
rect 1116 -2910 1122 -2904
rect 1116 -2916 1122 -2910
rect 1116 -2922 1122 -2916
rect 1116 -2928 1122 -2922
rect 1116 -2934 1122 -2928
rect 1116 -2940 1122 -2934
rect 1116 -2946 1122 -2940
rect 1116 -2952 1122 -2946
rect 1116 -2958 1122 -2952
rect 1116 -2964 1122 -2958
rect 1116 -2970 1122 -2964
rect 1116 -2976 1122 -2970
rect 1116 -2982 1122 -2976
rect 1116 -2988 1122 -2982
rect 1116 -2994 1122 -2988
rect 1116 -3000 1122 -2994
rect 1116 -3006 1122 -3000
rect 1116 -3012 1122 -3006
rect 1116 -3018 1122 -3012
rect 1116 -3024 1122 -3018
rect 1116 -3030 1122 -3024
rect 1116 -3036 1122 -3030
rect 1116 -3042 1122 -3036
rect 1116 -3048 1122 -3042
rect 1116 -3054 1122 -3048
rect 1116 -3060 1122 -3054
rect 1116 -3066 1122 -3060
rect 1116 -3072 1122 -3066
rect 1116 -3078 1122 -3072
rect 1116 -3084 1122 -3078
rect 1116 -3156 1122 -3150
rect 1116 -3162 1122 -3156
rect 1116 -3168 1122 -3162
rect 1116 -3174 1122 -3168
rect 1116 -3180 1122 -3174
rect 1116 -3186 1122 -3180
rect 1116 -3192 1122 -3186
rect 1116 -3198 1122 -3192
rect 1116 -3204 1122 -3198
rect 1116 -3210 1122 -3204
rect 1116 -3216 1122 -3210
rect 1116 -3222 1122 -3216
rect 1116 -3228 1122 -3222
rect 1116 -3234 1122 -3228
rect 1116 -3240 1122 -3234
rect 1116 -3246 1122 -3240
rect 1116 -3252 1122 -3246
rect 1116 -3258 1122 -3252
rect 1116 -3264 1122 -3258
rect 1116 -3270 1122 -3264
rect 1116 -3318 1122 -3312
rect 1116 -3324 1122 -3318
rect 1116 -3330 1122 -3324
rect 1116 -3336 1122 -3330
rect 1116 -3342 1122 -3336
rect 1116 -3348 1122 -3342
rect 1116 -3354 1122 -3348
rect 1116 -3360 1122 -3354
rect 1116 -3366 1122 -3360
rect 1116 -3372 1122 -3366
rect 1116 -3378 1122 -3372
rect 1116 -3384 1122 -3378
rect 1116 -3390 1122 -3384
rect 1116 -3396 1122 -3390
rect 1116 -3402 1122 -3396
rect 1116 -3408 1122 -3402
rect 1116 -3414 1122 -3408
rect 1116 -3420 1122 -3414
rect 1116 -3426 1122 -3420
rect 1116 -3432 1122 -3426
rect 1116 -3438 1122 -3432
rect 1116 -3444 1122 -3438
rect 1116 -3450 1122 -3444
rect 1116 -3456 1122 -3450
rect 1116 -3462 1122 -3456
rect 1116 -3468 1122 -3462
rect 1116 -3474 1122 -3468
rect 1116 -3480 1122 -3474
rect 1116 -3486 1122 -3480
rect 1116 -3492 1122 -3486
rect 1116 -3498 1122 -3492
rect 1116 -3504 1122 -3498
rect 1116 -3510 1122 -3504
rect 1122 -1110 1128 -1104
rect 1122 -1116 1128 -1110
rect 1122 -1122 1128 -1116
rect 1122 -1128 1128 -1122
rect 1122 -1134 1128 -1128
rect 1122 -1140 1128 -1134
rect 1122 -1146 1128 -1140
rect 1122 -1152 1128 -1146
rect 1122 -1158 1128 -1152
rect 1122 -1164 1128 -1158
rect 1122 -1170 1128 -1164
rect 1122 -1176 1128 -1170
rect 1122 -1182 1128 -1176
rect 1122 -1188 1128 -1182
rect 1122 -1194 1128 -1188
rect 1122 -1200 1128 -1194
rect 1122 -1206 1128 -1200
rect 1122 -1212 1128 -1206
rect 1122 -1218 1128 -1212
rect 1122 -1224 1128 -1218
rect 1122 -1230 1128 -1224
rect 1122 -1236 1128 -1230
rect 1122 -1242 1128 -1236
rect 1122 -1248 1128 -1242
rect 1122 -1254 1128 -1248
rect 1122 -1260 1128 -1254
rect 1122 -1266 1128 -1260
rect 1122 -1272 1128 -1266
rect 1122 -1278 1128 -1272
rect 1122 -1284 1128 -1278
rect 1122 -1290 1128 -1284
rect 1122 -1296 1128 -1290
rect 1122 -1302 1128 -1296
rect 1122 -1308 1128 -1302
rect 1122 -2022 1128 -2016
rect 1122 -2028 1128 -2022
rect 1122 -2034 1128 -2028
rect 1122 -2040 1128 -2034
rect 1122 -2046 1128 -2040
rect 1122 -2052 1128 -2046
rect 1122 -2058 1128 -2052
rect 1122 -2064 1128 -2058
rect 1122 -2070 1128 -2064
rect 1122 -2076 1128 -2070
rect 1122 -2082 1128 -2076
rect 1122 -2088 1128 -2082
rect 1122 -2094 1128 -2088
rect 1122 -2100 1128 -2094
rect 1122 -2106 1128 -2100
rect 1122 -2112 1128 -2106
rect 1122 -2118 1128 -2112
rect 1122 -2124 1128 -2118
rect 1122 -2130 1128 -2124
rect 1122 -2136 1128 -2130
rect 1122 -2142 1128 -2136
rect 1122 -2148 1128 -2142
rect 1122 -2154 1128 -2148
rect 1122 -2160 1128 -2154
rect 1122 -2166 1128 -2160
rect 1122 -2172 1128 -2166
rect 1122 -2178 1128 -2172
rect 1122 -2184 1128 -2178
rect 1122 -2190 1128 -2184
rect 1122 -2196 1128 -2190
rect 1122 -2202 1128 -2196
rect 1122 -2208 1128 -2202
rect 1122 -2214 1128 -2208
rect 1122 -2220 1128 -2214
rect 1122 -2226 1128 -2220
rect 1122 -2232 1128 -2226
rect 1122 -2238 1128 -2232
rect 1122 -2244 1128 -2238
rect 1122 -2250 1128 -2244
rect 1122 -2256 1128 -2250
rect 1122 -2262 1128 -2256
rect 1122 -2268 1128 -2262
rect 1122 -2274 1128 -2268
rect 1122 -2280 1128 -2274
rect 1122 -2286 1128 -2280
rect 1122 -2292 1128 -2286
rect 1122 -2298 1128 -2292
rect 1122 -2304 1128 -2298
rect 1122 -2310 1128 -2304
rect 1122 -2316 1128 -2310
rect 1122 -2322 1128 -2316
rect 1122 -2328 1128 -2322
rect 1122 -2334 1128 -2328
rect 1122 -2340 1128 -2334
rect 1122 -2346 1128 -2340
rect 1122 -2352 1128 -2346
rect 1122 -2358 1128 -2352
rect 1122 -2364 1128 -2358
rect 1122 -2370 1128 -2364
rect 1122 -2376 1128 -2370
rect 1122 -2382 1128 -2376
rect 1122 -2388 1128 -2382
rect 1122 -2394 1128 -2388
rect 1122 -2400 1128 -2394
rect 1122 -2406 1128 -2400
rect 1122 -2412 1128 -2406
rect 1122 -2418 1128 -2412
rect 1122 -2424 1128 -2418
rect 1122 -2430 1128 -2424
rect 1122 -2436 1128 -2430
rect 1122 -2442 1128 -2436
rect 1122 -2448 1128 -2442
rect 1122 -2454 1128 -2448
rect 1122 -2460 1128 -2454
rect 1122 -2466 1128 -2460
rect 1122 -2472 1128 -2466
rect 1122 -2478 1128 -2472
rect 1122 -2484 1128 -2478
rect 1122 -2490 1128 -2484
rect 1122 -2496 1128 -2490
rect 1122 -2502 1128 -2496
rect 1122 -2508 1128 -2502
rect 1122 -2514 1128 -2508
rect 1122 -2520 1128 -2514
rect 1122 -2526 1128 -2520
rect 1122 -2532 1128 -2526
rect 1122 -2538 1128 -2532
rect 1122 -2544 1128 -2538
rect 1122 -2550 1128 -2544
rect 1122 -2556 1128 -2550
rect 1122 -2562 1128 -2556
rect 1122 -2568 1128 -2562
rect 1122 -2574 1128 -2568
rect 1122 -2580 1128 -2574
rect 1122 -2586 1128 -2580
rect 1122 -2592 1128 -2586
rect 1122 -2598 1128 -2592
rect 1122 -2604 1128 -2598
rect 1122 -2610 1128 -2604
rect 1122 -2616 1128 -2610
rect 1122 -2622 1128 -2616
rect 1122 -2628 1128 -2622
rect 1122 -2634 1128 -2628
rect 1122 -2640 1128 -2634
rect 1122 -2646 1128 -2640
rect 1122 -2652 1128 -2646
rect 1122 -2658 1128 -2652
rect 1122 -2664 1128 -2658
rect 1122 -2670 1128 -2664
rect 1122 -2676 1128 -2670
rect 1122 -2682 1128 -2676
rect 1122 -2688 1128 -2682
rect 1122 -2694 1128 -2688
rect 1122 -2700 1128 -2694
rect 1122 -2706 1128 -2700
rect 1122 -2712 1128 -2706
rect 1122 -2718 1128 -2712
rect 1122 -2724 1128 -2718
rect 1122 -2826 1128 -2820
rect 1122 -2832 1128 -2826
rect 1122 -2838 1128 -2832
rect 1122 -2844 1128 -2838
rect 1122 -2850 1128 -2844
rect 1122 -2856 1128 -2850
rect 1122 -2862 1128 -2856
rect 1122 -2868 1128 -2862
rect 1122 -2874 1128 -2868
rect 1122 -2880 1128 -2874
rect 1122 -2886 1128 -2880
rect 1122 -2892 1128 -2886
rect 1122 -2898 1128 -2892
rect 1122 -2904 1128 -2898
rect 1122 -2910 1128 -2904
rect 1122 -2916 1128 -2910
rect 1122 -2922 1128 -2916
rect 1122 -2928 1128 -2922
rect 1122 -2934 1128 -2928
rect 1122 -2940 1128 -2934
rect 1122 -2946 1128 -2940
rect 1122 -2952 1128 -2946
rect 1122 -2958 1128 -2952
rect 1122 -2964 1128 -2958
rect 1122 -2970 1128 -2964
rect 1122 -2976 1128 -2970
rect 1122 -2982 1128 -2976
rect 1122 -2988 1128 -2982
rect 1122 -2994 1128 -2988
rect 1122 -3000 1128 -2994
rect 1122 -3006 1128 -3000
rect 1122 -3012 1128 -3006
rect 1122 -3018 1128 -3012
rect 1122 -3024 1128 -3018
rect 1122 -3030 1128 -3024
rect 1122 -3036 1128 -3030
rect 1122 -3042 1128 -3036
rect 1122 -3048 1128 -3042
rect 1122 -3054 1128 -3048
rect 1122 -3060 1128 -3054
rect 1122 -3066 1128 -3060
rect 1122 -3072 1128 -3066
rect 1122 -3078 1128 -3072
rect 1122 -3150 1128 -3144
rect 1122 -3156 1128 -3150
rect 1122 -3162 1128 -3156
rect 1122 -3168 1128 -3162
rect 1122 -3174 1128 -3168
rect 1122 -3180 1128 -3174
rect 1122 -3186 1128 -3180
rect 1122 -3192 1128 -3186
rect 1122 -3198 1128 -3192
rect 1122 -3204 1128 -3198
rect 1122 -3210 1128 -3204
rect 1122 -3216 1128 -3210
rect 1122 -3222 1128 -3216
rect 1122 -3228 1128 -3222
rect 1122 -3234 1128 -3228
rect 1122 -3240 1128 -3234
rect 1122 -3246 1128 -3240
rect 1122 -3252 1128 -3246
rect 1122 -3258 1128 -3252
rect 1122 -3264 1128 -3258
rect 1122 -3318 1128 -3312
rect 1122 -3324 1128 -3318
rect 1122 -3330 1128 -3324
rect 1122 -3336 1128 -3330
rect 1122 -3342 1128 -3336
rect 1122 -3348 1128 -3342
rect 1122 -3354 1128 -3348
rect 1122 -3360 1128 -3354
rect 1122 -3366 1128 -3360
rect 1122 -3372 1128 -3366
rect 1122 -3378 1128 -3372
rect 1122 -3384 1128 -3378
rect 1122 -3390 1128 -3384
rect 1122 -3396 1128 -3390
rect 1122 -3402 1128 -3396
rect 1122 -3408 1128 -3402
rect 1122 -3414 1128 -3408
rect 1122 -3420 1128 -3414
rect 1122 -3426 1128 -3420
rect 1122 -3432 1128 -3426
rect 1122 -3438 1128 -3432
rect 1122 -3444 1128 -3438
rect 1122 -3450 1128 -3444
rect 1122 -3456 1128 -3450
rect 1122 -3462 1128 -3456
rect 1122 -3468 1128 -3462
rect 1122 -3474 1128 -3468
rect 1122 -3480 1128 -3474
rect 1122 -3486 1128 -3480
rect 1122 -3492 1128 -3486
rect 1122 -3498 1128 -3492
rect 1122 -3504 1128 -3498
rect 1122 -3510 1128 -3504
rect 1128 -1104 1134 -1098
rect 1128 -1110 1134 -1104
rect 1128 -1116 1134 -1110
rect 1128 -1122 1134 -1116
rect 1128 -1128 1134 -1122
rect 1128 -1134 1134 -1128
rect 1128 -1140 1134 -1134
rect 1128 -1146 1134 -1140
rect 1128 -1152 1134 -1146
rect 1128 -1158 1134 -1152
rect 1128 -1164 1134 -1158
rect 1128 -1170 1134 -1164
rect 1128 -1176 1134 -1170
rect 1128 -1182 1134 -1176
rect 1128 -1188 1134 -1182
rect 1128 -1194 1134 -1188
rect 1128 -1200 1134 -1194
rect 1128 -1206 1134 -1200
rect 1128 -1212 1134 -1206
rect 1128 -1218 1134 -1212
rect 1128 -1224 1134 -1218
rect 1128 -1230 1134 -1224
rect 1128 -1236 1134 -1230
rect 1128 -1242 1134 -1236
rect 1128 -1248 1134 -1242
rect 1128 -1254 1134 -1248
rect 1128 -1260 1134 -1254
rect 1128 -1266 1134 -1260
rect 1128 -1272 1134 -1266
rect 1128 -1278 1134 -1272
rect 1128 -1284 1134 -1278
rect 1128 -1290 1134 -1284
rect 1128 -1296 1134 -1290
rect 1128 -1302 1134 -1296
rect 1128 -1308 1134 -1302
rect 1128 -2004 1134 -1998
rect 1128 -2010 1134 -2004
rect 1128 -2016 1134 -2010
rect 1128 -2022 1134 -2016
rect 1128 -2028 1134 -2022
rect 1128 -2034 1134 -2028
rect 1128 -2040 1134 -2034
rect 1128 -2046 1134 -2040
rect 1128 -2052 1134 -2046
rect 1128 -2058 1134 -2052
rect 1128 -2064 1134 -2058
rect 1128 -2070 1134 -2064
rect 1128 -2076 1134 -2070
rect 1128 -2082 1134 -2076
rect 1128 -2088 1134 -2082
rect 1128 -2094 1134 -2088
rect 1128 -2100 1134 -2094
rect 1128 -2106 1134 -2100
rect 1128 -2112 1134 -2106
rect 1128 -2118 1134 -2112
rect 1128 -2124 1134 -2118
rect 1128 -2130 1134 -2124
rect 1128 -2136 1134 -2130
rect 1128 -2142 1134 -2136
rect 1128 -2148 1134 -2142
rect 1128 -2154 1134 -2148
rect 1128 -2160 1134 -2154
rect 1128 -2166 1134 -2160
rect 1128 -2172 1134 -2166
rect 1128 -2178 1134 -2172
rect 1128 -2184 1134 -2178
rect 1128 -2190 1134 -2184
rect 1128 -2196 1134 -2190
rect 1128 -2202 1134 -2196
rect 1128 -2208 1134 -2202
rect 1128 -2214 1134 -2208
rect 1128 -2220 1134 -2214
rect 1128 -2226 1134 -2220
rect 1128 -2232 1134 -2226
rect 1128 -2238 1134 -2232
rect 1128 -2244 1134 -2238
rect 1128 -2250 1134 -2244
rect 1128 -2256 1134 -2250
rect 1128 -2262 1134 -2256
rect 1128 -2268 1134 -2262
rect 1128 -2274 1134 -2268
rect 1128 -2280 1134 -2274
rect 1128 -2286 1134 -2280
rect 1128 -2292 1134 -2286
rect 1128 -2298 1134 -2292
rect 1128 -2304 1134 -2298
rect 1128 -2310 1134 -2304
rect 1128 -2316 1134 -2310
rect 1128 -2322 1134 -2316
rect 1128 -2328 1134 -2322
rect 1128 -2334 1134 -2328
rect 1128 -2340 1134 -2334
rect 1128 -2346 1134 -2340
rect 1128 -2352 1134 -2346
rect 1128 -2358 1134 -2352
rect 1128 -2364 1134 -2358
rect 1128 -2370 1134 -2364
rect 1128 -2376 1134 -2370
rect 1128 -2382 1134 -2376
rect 1128 -2388 1134 -2382
rect 1128 -2394 1134 -2388
rect 1128 -2400 1134 -2394
rect 1128 -2406 1134 -2400
rect 1128 -2412 1134 -2406
rect 1128 -2418 1134 -2412
rect 1128 -2424 1134 -2418
rect 1128 -2430 1134 -2424
rect 1128 -2436 1134 -2430
rect 1128 -2442 1134 -2436
rect 1128 -2448 1134 -2442
rect 1128 -2454 1134 -2448
rect 1128 -2460 1134 -2454
rect 1128 -2466 1134 -2460
rect 1128 -2472 1134 -2466
rect 1128 -2478 1134 -2472
rect 1128 -2484 1134 -2478
rect 1128 -2490 1134 -2484
rect 1128 -2496 1134 -2490
rect 1128 -2502 1134 -2496
rect 1128 -2508 1134 -2502
rect 1128 -2514 1134 -2508
rect 1128 -2520 1134 -2514
rect 1128 -2526 1134 -2520
rect 1128 -2532 1134 -2526
rect 1128 -2538 1134 -2532
rect 1128 -2544 1134 -2538
rect 1128 -2550 1134 -2544
rect 1128 -2556 1134 -2550
rect 1128 -2562 1134 -2556
rect 1128 -2568 1134 -2562
rect 1128 -2574 1134 -2568
rect 1128 -2580 1134 -2574
rect 1128 -2586 1134 -2580
rect 1128 -2592 1134 -2586
rect 1128 -2598 1134 -2592
rect 1128 -2604 1134 -2598
rect 1128 -2610 1134 -2604
rect 1128 -2616 1134 -2610
rect 1128 -2622 1134 -2616
rect 1128 -2628 1134 -2622
rect 1128 -2634 1134 -2628
rect 1128 -2640 1134 -2634
rect 1128 -2646 1134 -2640
rect 1128 -2652 1134 -2646
rect 1128 -2658 1134 -2652
rect 1128 -2664 1134 -2658
rect 1128 -2670 1134 -2664
rect 1128 -2676 1134 -2670
rect 1128 -2682 1134 -2676
rect 1128 -2688 1134 -2682
rect 1128 -2694 1134 -2688
rect 1128 -2700 1134 -2694
rect 1128 -2706 1134 -2700
rect 1128 -2712 1134 -2706
rect 1128 -2814 1134 -2808
rect 1128 -2820 1134 -2814
rect 1128 -2826 1134 -2820
rect 1128 -2832 1134 -2826
rect 1128 -2838 1134 -2832
rect 1128 -2844 1134 -2838
rect 1128 -2850 1134 -2844
rect 1128 -2856 1134 -2850
rect 1128 -2862 1134 -2856
rect 1128 -2868 1134 -2862
rect 1128 -2874 1134 -2868
rect 1128 -2880 1134 -2874
rect 1128 -2886 1134 -2880
rect 1128 -2892 1134 -2886
rect 1128 -2898 1134 -2892
rect 1128 -2904 1134 -2898
rect 1128 -2910 1134 -2904
rect 1128 -2916 1134 -2910
rect 1128 -2922 1134 -2916
rect 1128 -2928 1134 -2922
rect 1128 -2934 1134 -2928
rect 1128 -2940 1134 -2934
rect 1128 -2946 1134 -2940
rect 1128 -2952 1134 -2946
rect 1128 -2958 1134 -2952
rect 1128 -2964 1134 -2958
rect 1128 -2970 1134 -2964
rect 1128 -2976 1134 -2970
rect 1128 -2982 1134 -2976
rect 1128 -2988 1134 -2982
rect 1128 -2994 1134 -2988
rect 1128 -3000 1134 -2994
rect 1128 -3006 1134 -3000
rect 1128 -3012 1134 -3006
rect 1128 -3018 1134 -3012
rect 1128 -3024 1134 -3018
rect 1128 -3030 1134 -3024
rect 1128 -3036 1134 -3030
rect 1128 -3042 1134 -3036
rect 1128 -3048 1134 -3042
rect 1128 -3054 1134 -3048
rect 1128 -3060 1134 -3054
rect 1128 -3066 1134 -3060
rect 1128 -3072 1134 -3066
rect 1128 -3078 1134 -3072
rect 1128 -3150 1134 -3144
rect 1128 -3156 1134 -3150
rect 1128 -3162 1134 -3156
rect 1128 -3168 1134 -3162
rect 1128 -3174 1134 -3168
rect 1128 -3180 1134 -3174
rect 1128 -3186 1134 -3180
rect 1128 -3192 1134 -3186
rect 1128 -3198 1134 -3192
rect 1128 -3204 1134 -3198
rect 1128 -3210 1134 -3204
rect 1128 -3216 1134 -3210
rect 1128 -3222 1134 -3216
rect 1128 -3228 1134 -3222
rect 1128 -3234 1134 -3228
rect 1128 -3240 1134 -3234
rect 1128 -3246 1134 -3240
rect 1128 -3252 1134 -3246
rect 1128 -3258 1134 -3252
rect 1128 -3264 1134 -3258
rect 1128 -3318 1134 -3312
rect 1128 -3324 1134 -3318
rect 1128 -3330 1134 -3324
rect 1128 -3336 1134 -3330
rect 1128 -3342 1134 -3336
rect 1128 -3348 1134 -3342
rect 1128 -3354 1134 -3348
rect 1128 -3360 1134 -3354
rect 1128 -3366 1134 -3360
rect 1128 -3372 1134 -3366
rect 1128 -3378 1134 -3372
rect 1128 -3384 1134 -3378
rect 1128 -3390 1134 -3384
rect 1128 -3396 1134 -3390
rect 1128 -3402 1134 -3396
rect 1128 -3408 1134 -3402
rect 1128 -3414 1134 -3408
rect 1128 -3420 1134 -3414
rect 1128 -3426 1134 -3420
rect 1128 -3432 1134 -3426
rect 1128 -3438 1134 -3432
rect 1128 -3444 1134 -3438
rect 1128 -3450 1134 -3444
rect 1128 -3456 1134 -3450
rect 1128 -3462 1134 -3456
rect 1128 -3468 1134 -3462
rect 1128 -3474 1134 -3468
rect 1128 -3480 1134 -3474
rect 1128 -3486 1134 -3480
rect 1128 -3492 1134 -3486
rect 1128 -3498 1134 -3492
rect 1128 -3504 1134 -3498
rect 1128 -3510 1134 -3504
rect 1128 -3516 1134 -3510
rect 1134 -1104 1140 -1098
rect 1134 -1110 1140 -1104
rect 1134 -1116 1140 -1110
rect 1134 -1122 1140 -1116
rect 1134 -1128 1140 -1122
rect 1134 -1134 1140 -1128
rect 1134 -1140 1140 -1134
rect 1134 -1146 1140 -1140
rect 1134 -1152 1140 -1146
rect 1134 -1158 1140 -1152
rect 1134 -1164 1140 -1158
rect 1134 -1170 1140 -1164
rect 1134 -1176 1140 -1170
rect 1134 -1182 1140 -1176
rect 1134 -1188 1140 -1182
rect 1134 -1194 1140 -1188
rect 1134 -1200 1140 -1194
rect 1134 -1206 1140 -1200
rect 1134 -1212 1140 -1206
rect 1134 -1218 1140 -1212
rect 1134 -1224 1140 -1218
rect 1134 -1230 1140 -1224
rect 1134 -1236 1140 -1230
rect 1134 -1242 1140 -1236
rect 1134 -1248 1140 -1242
rect 1134 -1254 1140 -1248
rect 1134 -1260 1140 -1254
rect 1134 -1266 1140 -1260
rect 1134 -1272 1140 -1266
rect 1134 -1278 1140 -1272
rect 1134 -1284 1140 -1278
rect 1134 -1290 1140 -1284
rect 1134 -1296 1140 -1290
rect 1134 -1302 1140 -1296
rect 1134 -1308 1140 -1302
rect 1134 -1986 1140 -1980
rect 1134 -1992 1140 -1986
rect 1134 -1998 1140 -1992
rect 1134 -2004 1140 -1998
rect 1134 -2010 1140 -2004
rect 1134 -2016 1140 -2010
rect 1134 -2022 1140 -2016
rect 1134 -2028 1140 -2022
rect 1134 -2034 1140 -2028
rect 1134 -2040 1140 -2034
rect 1134 -2046 1140 -2040
rect 1134 -2052 1140 -2046
rect 1134 -2058 1140 -2052
rect 1134 -2064 1140 -2058
rect 1134 -2070 1140 -2064
rect 1134 -2076 1140 -2070
rect 1134 -2082 1140 -2076
rect 1134 -2088 1140 -2082
rect 1134 -2094 1140 -2088
rect 1134 -2100 1140 -2094
rect 1134 -2106 1140 -2100
rect 1134 -2112 1140 -2106
rect 1134 -2118 1140 -2112
rect 1134 -2124 1140 -2118
rect 1134 -2130 1140 -2124
rect 1134 -2136 1140 -2130
rect 1134 -2142 1140 -2136
rect 1134 -2148 1140 -2142
rect 1134 -2154 1140 -2148
rect 1134 -2160 1140 -2154
rect 1134 -2166 1140 -2160
rect 1134 -2172 1140 -2166
rect 1134 -2178 1140 -2172
rect 1134 -2184 1140 -2178
rect 1134 -2190 1140 -2184
rect 1134 -2196 1140 -2190
rect 1134 -2202 1140 -2196
rect 1134 -2208 1140 -2202
rect 1134 -2214 1140 -2208
rect 1134 -2220 1140 -2214
rect 1134 -2226 1140 -2220
rect 1134 -2232 1140 -2226
rect 1134 -2238 1140 -2232
rect 1134 -2244 1140 -2238
rect 1134 -2250 1140 -2244
rect 1134 -2256 1140 -2250
rect 1134 -2262 1140 -2256
rect 1134 -2268 1140 -2262
rect 1134 -2274 1140 -2268
rect 1134 -2280 1140 -2274
rect 1134 -2286 1140 -2280
rect 1134 -2292 1140 -2286
rect 1134 -2298 1140 -2292
rect 1134 -2304 1140 -2298
rect 1134 -2310 1140 -2304
rect 1134 -2316 1140 -2310
rect 1134 -2322 1140 -2316
rect 1134 -2328 1140 -2322
rect 1134 -2334 1140 -2328
rect 1134 -2340 1140 -2334
rect 1134 -2346 1140 -2340
rect 1134 -2352 1140 -2346
rect 1134 -2358 1140 -2352
rect 1134 -2364 1140 -2358
rect 1134 -2370 1140 -2364
rect 1134 -2376 1140 -2370
rect 1134 -2382 1140 -2376
rect 1134 -2388 1140 -2382
rect 1134 -2394 1140 -2388
rect 1134 -2400 1140 -2394
rect 1134 -2406 1140 -2400
rect 1134 -2412 1140 -2406
rect 1134 -2418 1140 -2412
rect 1134 -2424 1140 -2418
rect 1134 -2430 1140 -2424
rect 1134 -2436 1140 -2430
rect 1134 -2442 1140 -2436
rect 1134 -2448 1140 -2442
rect 1134 -2454 1140 -2448
rect 1134 -2460 1140 -2454
rect 1134 -2466 1140 -2460
rect 1134 -2472 1140 -2466
rect 1134 -2478 1140 -2472
rect 1134 -2484 1140 -2478
rect 1134 -2490 1140 -2484
rect 1134 -2496 1140 -2490
rect 1134 -2502 1140 -2496
rect 1134 -2508 1140 -2502
rect 1134 -2514 1140 -2508
rect 1134 -2520 1140 -2514
rect 1134 -2526 1140 -2520
rect 1134 -2532 1140 -2526
rect 1134 -2538 1140 -2532
rect 1134 -2544 1140 -2538
rect 1134 -2550 1140 -2544
rect 1134 -2556 1140 -2550
rect 1134 -2562 1140 -2556
rect 1134 -2568 1140 -2562
rect 1134 -2574 1140 -2568
rect 1134 -2580 1140 -2574
rect 1134 -2586 1140 -2580
rect 1134 -2592 1140 -2586
rect 1134 -2598 1140 -2592
rect 1134 -2604 1140 -2598
rect 1134 -2610 1140 -2604
rect 1134 -2616 1140 -2610
rect 1134 -2622 1140 -2616
rect 1134 -2628 1140 -2622
rect 1134 -2634 1140 -2628
rect 1134 -2640 1140 -2634
rect 1134 -2646 1140 -2640
rect 1134 -2652 1140 -2646
rect 1134 -2658 1140 -2652
rect 1134 -2664 1140 -2658
rect 1134 -2670 1140 -2664
rect 1134 -2676 1140 -2670
rect 1134 -2682 1140 -2676
rect 1134 -2688 1140 -2682
rect 1134 -2694 1140 -2688
rect 1134 -2700 1140 -2694
rect 1134 -2706 1140 -2700
rect 1134 -2802 1140 -2796
rect 1134 -2808 1140 -2802
rect 1134 -2814 1140 -2808
rect 1134 -2820 1140 -2814
rect 1134 -2826 1140 -2820
rect 1134 -2832 1140 -2826
rect 1134 -2838 1140 -2832
rect 1134 -2844 1140 -2838
rect 1134 -2850 1140 -2844
rect 1134 -2856 1140 -2850
rect 1134 -2862 1140 -2856
rect 1134 -2868 1140 -2862
rect 1134 -2874 1140 -2868
rect 1134 -2880 1140 -2874
rect 1134 -2886 1140 -2880
rect 1134 -2892 1140 -2886
rect 1134 -2898 1140 -2892
rect 1134 -2904 1140 -2898
rect 1134 -2910 1140 -2904
rect 1134 -2916 1140 -2910
rect 1134 -2922 1140 -2916
rect 1134 -2928 1140 -2922
rect 1134 -2934 1140 -2928
rect 1134 -2940 1140 -2934
rect 1134 -2946 1140 -2940
rect 1134 -2952 1140 -2946
rect 1134 -2958 1140 -2952
rect 1134 -2964 1140 -2958
rect 1134 -2970 1140 -2964
rect 1134 -2976 1140 -2970
rect 1134 -2982 1140 -2976
rect 1134 -2988 1140 -2982
rect 1134 -2994 1140 -2988
rect 1134 -3000 1140 -2994
rect 1134 -3006 1140 -3000
rect 1134 -3012 1140 -3006
rect 1134 -3018 1140 -3012
rect 1134 -3024 1140 -3018
rect 1134 -3030 1140 -3024
rect 1134 -3036 1140 -3030
rect 1134 -3042 1140 -3036
rect 1134 -3048 1140 -3042
rect 1134 -3054 1140 -3048
rect 1134 -3060 1140 -3054
rect 1134 -3066 1140 -3060
rect 1134 -3072 1140 -3066
rect 1134 -3144 1140 -3138
rect 1134 -3150 1140 -3144
rect 1134 -3156 1140 -3150
rect 1134 -3162 1140 -3156
rect 1134 -3168 1140 -3162
rect 1134 -3174 1140 -3168
rect 1134 -3180 1140 -3174
rect 1134 -3186 1140 -3180
rect 1134 -3192 1140 -3186
rect 1134 -3198 1140 -3192
rect 1134 -3204 1140 -3198
rect 1134 -3210 1140 -3204
rect 1134 -3216 1140 -3210
rect 1134 -3222 1140 -3216
rect 1134 -3228 1140 -3222
rect 1134 -3234 1140 -3228
rect 1134 -3240 1140 -3234
rect 1134 -3246 1140 -3240
rect 1134 -3252 1140 -3246
rect 1134 -3258 1140 -3252
rect 1134 -3264 1140 -3258
rect 1134 -3318 1140 -3312
rect 1134 -3324 1140 -3318
rect 1134 -3330 1140 -3324
rect 1134 -3336 1140 -3330
rect 1134 -3342 1140 -3336
rect 1134 -3348 1140 -3342
rect 1134 -3354 1140 -3348
rect 1134 -3360 1140 -3354
rect 1134 -3366 1140 -3360
rect 1134 -3372 1140 -3366
rect 1134 -3378 1140 -3372
rect 1134 -3384 1140 -3378
rect 1134 -3390 1140 -3384
rect 1134 -3396 1140 -3390
rect 1134 -3402 1140 -3396
rect 1134 -3408 1140 -3402
rect 1134 -3414 1140 -3408
rect 1134 -3420 1140 -3414
rect 1134 -3426 1140 -3420
rect 1134 -3432 1140 -3426
rect 1134 -3438 1140 -3432
rect 1134 -3444 1140 -3438
rect 1134 -3450 1140 -3444
rect 1134 -3456 1140 -3450
rect 1134 -3462 1140 -3456
rect 1134 -3468 1140 -3462
rect 1134 -3474 1140 -3468
rect 1134 -3480 1140 -3474
rect 1134 -3486 1140 -3480
rect 1134 -3492 1140 -3486
rect 1134 -3498 1140 -3492
rect 1134 -3504 1140 -3498
rect 1134 -3510 1140 -3504
rect 1134 -3516 1140 -3510
rect 1140 -1104 1146 -1098
rect 1140 -1110 1146 -1104
rect 1140 -1116 1146 -1110
rect 1140 -1122 1146 -1116
rect 1140 -1128 1146 -1122
rect 1140 -1134 1146 -1128
rect 1140 -1140 1146 -1134
rect 1140 -1146 1146 -1140
rect 1140 -1152 1146 -1146
rect 1140 -1158 1146 -1152
rect 1140 -1164 1146 -1158
rect 1140 -1170 1146 -1164
rect 1140 -1176 1146 -1170
rect 1140 -1182 1146 -1176
rect 1140 -1188 1146 -1182
rect 1140 -1194 1146 -1188
rect 1140 -1200 1146 -1194
rect 1140 -1206 1146 -1200
rect 1140 -1212 1146 -1206
rect 1140 -1218 1146 -1212
rect 1140 -1224 1146 -1218
rect 1140 -1230 1146 -1224
rect 1140 -1236 1146 -1230
rect 1140 -1242 1146 -1236
rect 1140 -1248 1146 -1242
rect 1140 -1254 1146 -1248
rect 1140 -1260 1146 -1254
rect 1140 -1266 1146 -1260
rect 1140 -1272 1146 -1266
rect 1140 -1278 1146 -1272
rect 1140 -1284 1146 -1278
rect 1140 -1290 1146 -1284
rect 1140 -1296 1146 -1290
rect 1140 -1302 1146 -1296
rect 1140 -1308 1146 -1302
rect 1140 -1974 1146 -1968
rect 1140 -1980 1146 -1974
rect 1140 -1986 1146 -1980
rect 1140 -1992 1146 -1986
rect 1140 -1998 1146 -1992
rect 1140 -2004 1146 -1998
rect 1140 -2010 1146 -2004
rect 1140 -2016 1146 -2010
rect 1140 -2022 1146 -2016
rect 1140 -2028 1146 -2022
rect 1140 -2034 1146 -2028
rect 1140 -2040 1146 -2034
rect 1140 -2046 1146 -2040
rect 1140 -2052 1146 -2046
rect 1140 -2058 1146 -2052
rect 1140 -2064 1146 -2058
rect 1140 -2070 1146 -2064
rect 1140 -2076 1146 -2070
rect 1140 -2082 1146 -2076
rect 1140 -2088 1146 -2082
rect 1140 -2094 1146 -2088
rect 1140 -2100 1146 -2094
rect 1140 -2106 1146 -2100
rect 1140 -2112 1146 -2106
rect 1140 -2118 1146 -2112
rect 1140 -2124 1146 -2118
rect 1140 -2130 1146 -2124
rect 1140 -2136 1146 -2130
rect 1140 -2142 1146 -2136
rect 1140 -2148 1146 -2142
rect 1140 -2154 1146 -2148
rect 1140 -2160 1146 -2154
rect 1140 -2166 1146 -2160
rect 1140 -2172 1146 -2166
rect 1140 -2178 1146 -2172
rect 1140 -2184 1146 -2178
rect 1140 -2190 1146 -2184
rect 1140 -2196 1146 -2190
rect 1140 -2202 1146 -2196
rect 1140 -2208 1146 -2202
rect 1140 -2214 1146 -2208
rect 1140 -2220 1146 -2214
rect 1140 -2226 1146 -2220
rect 1140 -2232 1146 -2226
rect 1140 -2238 1146 -2232
rect 1140 -2244 1146 -2238
rect 1140 -2250 1146 -2244
rect 1140 -2256 1146 -2250
rect 1140 -2262 1146 -2256
rect 1140 -2268 1146 -2262
rect 1140 -2274 1146 -2268
rect 1140 -2280 1146 -2274
rect 1140 -2286 1146 -2280
rect 1140 -2292 1146 -2286
rect 1140 -2298 1146 -2292
rect 1140 -2304 1146 -2298
rect 1140 -2310 1146 -2304
rect 1140 -2316 1146 -2310
rect 1140 -2322 1146 -2316
rect 1140 -2328 1146 -2322
rect 1140 -2334 1146 -2328
rect 1140 -2340 1146 -2334
rect 1140 -2346 1146 -2340
rect 1140 -2352 1146 -2346
rect 1140 -2358 1146 -2352
rect 1140 -2364 1146 -2358
rect 1140 -2370 1146 -2364
rect 1140 -2376 1146 -2370
rect 1140 -2382 1146 -2376
rect 1140 -2388 1146 -2382
rect 1140 -2394 1146 -2388
rect 1140 -2400 1146 -2394
rect 1140 -2406 1146 -2400
rect 1140 -2412 1146 -2406
rect 1140 -2418 1146 -2412
rect 1140 -2424 1146 -2418
rect 1140 -2430 1146 -2424
rect 1140 -2436 1146 -2430
rect 1140 -2442 1146 -2436
rect 1140 -2448 1146 -2442
rect 1140 -2454 1146 -2448
rect 1140 -2460 1146 -2454
rect 1140 -2466 1146 -2460
rect 1140 -2472 1146 -2466
rect 1140 -2478 1146 -2472
rect 1140 -2484 1146 -2478
rect 1140 -2490 1146 -2484
rect 1140 -2496 1146 -2490
rect 1140 -2502 1146 -2496
rect 1140 -2508 1146 -2502
rect 1140 -2514 1146 -2508
rect 1140 -2520 1146 -2514
rect 1140 -2526 1146 -2520
rect 1140 -2532 1146 -2526
rect 1140 -2538 1146 -2532
rect 1140 -2544 1146 -2538
rect 1140 -2550 1146 -2544
rect 1140 -2556 1146 -2550
rect 1140 -2562 1146 -2556
rect 1140 -2568 1146 -2562
rect 1140 -2574 1146 -2568
rect 1140 -2580 1146 -2574
rect 1140 -2586 1146 -2580
rect 1140 -2592 1146 -2586
rect 1140 -2598 1146 -2592
rect 1140 -2604 1146 -2598
rect 1140 -2610 1146 -2604
rect 1140 -2616 1146 -2610
rect 1140 -2622 1146 -2616
rect 1140 -2628 1146 -2622
rect 1140 -2634 1146 -2628
rect 1140 -2640 1146 -2634
rect 1140 -2646 1146 -2640
rect 1140 -2652 1146 -2646
rect 1140 -2658 1146 -2652
rect 1140 -2664 1146 -2658
rect 1140 -2670 1146 -2664
rect 1140 -2676 1146 -2670
rect 1140 -2682 1146 -2676
rect 1140 -2688 1146 -2682
rect 1140 -2694 1146 -2688
rect 1140 -2796 1146 -2790
rect 1140 -2802 1146 -2796
rect 1140 -2808 1146 -2802
rect 1140 -2814 1146 -2808
rect 1140 -2820 1146 -2814
rect 1140 -2826 1146 -2820
rect 1140 -2832 1146 -2826
rect 1140 -2838 1146 -2832
rect 1140 -2844 1146 -2838
rect 1140 -2850 1146 -2844
rect 1140 -2856 1146 -2850
rect 1140 -2862 1146 -2856
rect 1140 -2868 1146 -2862
rect 1140 -2874 1146 -2868
rect 1140 -2880 1146 -2874
rect 1140 -2886 1146 -2880
rect 1140 -2892 1146 -2886
rect 1140 -2898 1146 -2892
rect 1140 -2904 1146 -2898
rect 1140 -2910 1146 -2904
rect 1140 -2916 1146 -2910
rect 1140 -2922 1146 -2916
rect 1140 -2928 1146 -2922
rect 1140 -2934 1146 -2928
rect 1140 -2940 1146 -2934
rect 1140 -2946 1146 -2940
rect 1140 -2952 1146 -2946
rect 1140 -2958 1146 -2952
rect 1140 -2964 1146 -2958
rect 1140 -2970 1146 -2964
rect 1140 -2976 1146 -2970
rect 1140 -2982 1146 -2976
rect 1140 -2988 1146 -2982
rect 1140 -2994 1146 -2988
rect 1140 -3000 1146 -2994
rect 1140 -3006 1146 -3000
rect 1140 -3012 1146 -3006
rect 1140 -3018 1146 -3012
rect 1140 -3024 1146 -3018
rect 1140 -3030 1146 -3024
rect 1140 -3036 1146 -3030
rect 1140 -3042 1146 -3036
rect 1140 -3048 1146 -3042
rect 1140 -3054 1146 -3048
rect 1140 -3060 1146 -3054
rect 1140 -3066 1146 -3060
rect 1140 -3138 1146 -3132
rect 1140 -3144 1146 -3138
rect 1140 -3150 1146 -3144
rect 1140 -3156 1146 -3150
rect 1140 -3162 1146 -3156
rect 1140 -3168 1146 -3162
rect 1140 -3174 1146 -3168
rect 1140 -3180 1146 -3174
rect 1140 -3186 1146 -3180
rect 1140 -3192 1146 -3186
rect 1140 -3198 1146 -3192
rect 1140 -3204 1146 -3198
rect 1140 -3210 1146 -3204
rect 1140 -3216 1146 -3210
rect 1140 -3222 1146 -3216
rect 1140 -3228 1146 -3222
rect 1140 -3234 1146 -3228
rect 1140 -3240 1146 -3234
rect 1140 -3246 1146 -3240
rect 1140 -3252 1146 -3246
rect 1140 -3258 1146 -3252
rect 1140 -3318 1146 -3312
rect 1140 -3324 1146 -3318
rect 1140 -3330 1146 -3324
rect 1140 -3336 1146 -3330
rect 1140 -3342 1146 -3336
rect 1140 -3348 1146 -3342
rect 1140 -3354 1146 -3348
rect 1140 -3360 1146 -3354
rect 1140 -3366 1146 -3360
rect 1140 -3372 1146 -3366
rect 1140 -3378 1146 -3372
rect 1140 -3384 1146 -3378
rect 1140 -3390 1146 -3384
rect 1140 -3396 1146 -3390
rect 1140 -3402 1146 -3396
rect 1140 -3408 1146 -3402
rect 1140 -3414 1146 -3408
rect 1140 -3420 1146 -3414
rect 1140 -3426 1146 -3420
rect 1140 -3432 1146 -3426
rect 1140 -3438 1146 -3432
rect 1140 -3444 1146 -3438
rect 1140 -3450 1146 -3444
rect 1140 -3456 1146 -3450
rect 1140 -3462 1146 -3456
rect 1140 -3468 1146 -3462
rect 1140 -3474 1146 -3468
rect 1140 -3480 1146 -3474
rect 1140 -3486 1146 -3480
rect 1140 -3492 1146 -3486
rect 1140 -3498 1146 -3492
rect 1140 -3504 1146 -3498
rect 1140 -3510 1146 -3504
rect 1140 -3516 1146 -3510
rect 1146 -1104 1152 -1098
rect 1146 -1110 1152 -1104
rect 1146 -1116 1152 -1110
rect 1146 -1122 1152 -1116
rect 1146 -1128 1152 -1122
rect 1146 -1134 1152 -1128
rect 1146 -1140 1152 -1134
rect 1146 -1146 1152 -1140
rect 1146 -1152 1152 -1146
rect 1146 -1158 1152 -1152
rect 1146 -1164 1152 -1158
rect 1146 -1170 1152 -1164
rect 1146 -1176 1152 -1170
rect 1146 -1182 1152 -1176
rect 1146 -1188 1152 -1182
rect 1146 -1194 1152 -1188
rect 1146 -1200 1152 -1194
rect 1146 -1206 1152 -1200
rect 1146 -1212 1152 -1206
rect 1146 -1218 1152 -1212
rect 1146 -1224 1152 -1218
rect 1146 -1230 1152 -1224
rect 1146 -1236 1152 -1230
rect 1146 -1242 1152 -1236
rect 1146 -1248 1152 -1242
rect 1146 -1254 1152 -1248
rect 1146 -1260 1152 -1254
rect 1146 -1266 1152 -1260
rect 1146 -1272 1152 -1266
rect 1146 -1278 1152 -1272
rect 1146 -1284 1152 -1278
rect 1146 -1290 1152 -1284
rect 1146 -1296 1152 -1290
rect 1146 -1302 1152 -1296
rect 1146 -1308 1152 -1302
rect 1146 -1956 1152 -1950
rect 1146 -1962 1152 -1956
rect 1146 -1968 1152 -1962
rect 1146 -1974 1152 -1968
rect 1146 -1980 1152 -1974
rect 1146 -1986 1152 -1980
rect 1146 -1992 1152 -1986
rect 1146 -1998 1152 -1992
rect 1146 -2004 1152 -1998
rect 1146 -2010 1152 -2004
rect 1146 -2016 1152 -2010
rect 1146 -2022 1152 -2016
rect 1146 -2028 1152 -2022
rect 1146 -2034 1152 -2028
rect 1146 -2040 1152 -2034
rect 1146 -2046 1152 -2040
rect 1146 -2052 1152 -2046
rect 1146 -2058 1152 -2052
rect 1146 -2064 1152 -2058
rect 1146 -2070 1152 -2064
rect 1146 -2076 1152 -2070
rect 1146 -2082 1152 -2076
rect 1146 -2088 1152 -2082
rect 1146 -2094 1152 -2088
rect 1146 -2100 1152 -2094
rect 1146 -2106 1152 -2100
rect 1146 -2112 1152 -2106
rect 1146 -2118 1152 -2112
rect 1146 -2124 1152 -2118
rect 1146 -2130 1152 -2124
rect 1146 -2136 1152 -2130
rect 1146 -2142 1152 -2136
rect 1146 -2148 1152 -2142
rect 1146 -2154 1152 -2148
rect 1146 -2160 1152 -2154
rect 1146 -2166 1152 -2160
rect 1146 -2172 1152 -2166
rect 1146 -2178 1152 -2172
rect 1146 -2184 1152 -2178
rect 1146 -2190 1152 -2184
rect 1146 -2196 1152 -2190
rect 1146 -2202 1152 -2196
rect 1146 -2208 1152 -2202
rect 1146 -2214 1152 -2208
rect 1146 -2220 1152 -2214
rect 1146 -2226 1152 -2220
rect 1146 -2232 1152 -2226
rect 1146 -2238 1152 -2232
rect 1146 -2244 1152 -2238
rect 1146 -2250 1152 -2244
rect 1146 -2256 1152 -2250
rect 1146 -2262 1152 -2256
rect 1146 -2268 1152 -2262
rect 1146 -2274 1152 -2268
rect 1146 -2280 1152 -2274
rect 1146 -2286 1152 -2280
rect 1146 -2292 1152 -2286
rect 1146 -2298 1152 -2292
rect 1146 -2304 1152 -2298
rect 1146 -2310 1152 -2304
rect 1146 -2316 1152 -2310
rect 1146 -2322 1152 -2316
rect 1146 -2328 1152 -2322
rect 1146 -2334 1152 -2328
rect 1146 -2340 1152 -2334
rect 1146 -2346 1152 -2340
rect 1146 -2352 1152 -2346
rect 1146 -2358 1152 -2352
rect 1146 -2364 1152 -2358
rect 1146 -2370 1152 -2364
rect 1146 -2376 1152 -2370
rect 1146 -2382 1152 -2376
rect 1146 -2388 1152 -2382
rect 1146 -2394 1152 -2388
rect 1146 -2400 1152 -2394
rect 1146 -2406 1152 -2400
rect 1146 -2412 1152 -2406
rect 1146 -2418 1152 -2412
rect 1146 -2424 1152 -2418
rect 1146 -2430 1152 -2424
rect 1146 -2436 1152 -2430
rect 1146 -2442 1152 -2436
rect 1146 -2448 1152 -2442
rect 1146 -2454 1152 -2448
rect 1146 -2460 1152 -2454
rect 1146 -2466 1152 -2460
rect 1146 -2472 1152 -2466
rect 1146 -2478 1152 -2472
rect 1146 -2484 1152 -2478
rect 1146 -2490 1152 -2484
rect 1146 -2496 1152 -2490
rect 1146 -2502 1152 -2496
rect 1146 -2508 1152 -2502
rect 1146 -2514 1152 -2508
rect 1146 -2520 1152 -2514
rect 1146 -2526 1152 -2520
rect 1146 -2532 1152 -2526
rect 1146 -2538 1152 -2532
rect 1146 -2544 1152 -2538
rect 1146 -2550 1152 -2544
rect 1146 -2556 1152 -2550
rect 1146 -2562 1152 -2556
rect 1146 -2568 1152 -2562
rect 1146 -2574 1152 -2568
rect 1146 -2580 1152 -2574
rect 1146 -2586 1152 -2580
rect 1146 -2592 1152 -2586
rect 1146 -2598 1152 -2592
rect 1146 -2604 1152 -2598
rect 1146 -2610 1152 -2604
rect 1146 -2616 1152 -2610
rect 1146 -2622 1152 -2616
rect 1146 -2628 1152 -2622
rect 1146 -2634 1152 -2628
rect 1146 -2640 1152 -2634
rect 1146 -2646 1152 -2640
rect 1146 -2652 1152 -2646
rect 1146 -2658 1152 -2652
rect 1146 -2664 1152 -2658
rect 1146 -2670 1152 -2664
rect 1146 -2676 1152 -2670
rect 1146 -2682 1152 -2676
rect 1146 -2688 1152 -2682
rect 1146 -2784 1152 -2778
rect 1146 -2790 1152 -2784
rect 1146 -2796 1152 -2790
rect 1146 -2802 1152 -2796
rect 1146 -2808 1152 -2802
rect 1146 -2814 1152 -2808
rect 1146 -2820 1152 -2814
rect 1146 -2826 1152 -2820
rect 1146 -2832 1152 -2826
rect 1146 -2838 1152 -2832
rect 1146 -2844 1152 -2838
rect 1146 -2850 1152 -2844
rect 1146 -2856 1152 -2850
rect 1146 -2862 1152 -2856
rect 1146 -2868 1152 -2862
rect 1146 -2874 1152 -2868
rect 1146 -2880 1152 -2874
rect 1146 -2886 1152 -2880
rect 1146 -2892 1152 -2886
rect 1146 -2898 1152 -2892
rect 1146 -2904 1152 -2898
rect 1146 -2910 1152 -2904
rect 1146 -2916 1152 -2910
rect 1146 -2922 1152 -2916
rect 1146 -2928 1152 -2922
rect 1146 -2934 1152 -2928
rect 1146 -2940 1152 -2934
rect 1146 -2946 1152 -2940
rect 1146 -2952 1152 -2946
rect 1146 -2958 1152 -2952
rect 1146 -2964 1152 -2958
rect 1146 -2970 1152 -2964
rect 1146 -2976 1152 -2970
rect 1146 -2982 1152 -2976
rect 1146 -2988 1152 -2982
rect 1146 -2994 1152 -2988
rect 1146 -3000 1152 -2994
rect 1146 -3006 1152 -3000
rect 1146 -3012 1152 -3006
rect 1146 -3018 1152 -3012
rect 1146 -3024 1152 -3018
rect 1146 -3030 1152 -3024
rect 1146 -3036 1152 -3030
rect 1146 -3042 1152 -3036
rect 1146 -3048 1152 -3042
rect 1146 -3054 1152 -3048
rect 1146 -3060 1152 -3054
rect 1146 -3132 1152 -3126
rect 1146 -3138 1152 -3132
rect 1146 -3144 1152 -3138
rect 1146 -3150 1152 -3144
rect 1146 -3156 1152 -3150
rect 1146 -3162 1152 -3156
rect 1146 -3168 1152 -3162
rect 1146 -3174 1152 -3168
rect 1146 -3180 1152 -3174
rect 1146 -3186 1152 -3180
rect 1146 -3192 1152 -3186
rect 1146 -3198 1152 -3192
rect 1146 -3204 1152 -3198
rect 1146 -3210 1152 -3204
rect 1146 -3216 1152 -3210
rect 1146 -3222 1152 -3216
rect 1146 -3228 1152 -3222
rect 1146 -3234 1152 -3228
rect 1146 -3240 1152 -3234
rect 1146 -3246 1152 -3240
rect 1146 -3252 1152 -3246
rect 1146 -3258 1152 -3252
rect 1146 -3318 1152 -3312
rect 1146 -3324 1152 -3318
rect 1146 -3330 1152 -3324
rect 1146 -3336 1152 -3330
rect 1146 -3342 1152 -3336
rect 1146 -3348 1152 -3342
rect 1146 -3354 1152 -3348
rect 1146 -3360 1152 -3354
rect 1146 -3366 1152 -3360
rect 1146 -3372 1152 -3366
rect 1146 -3378 1152 -3372
rect 1146 -3384 1152 -3378
rect 1146 -3390 1152 -3384
rect 1146 -3396 1152 -3390
rect 1146 -3402 1152 -3396
rect 1146 -3408 1152 -3402
rect 1146 -3414 1152 -3408
rect 1146 -3420 1152 -3414
rect 1146 -3426 1152 -3420
rect 1146 -3432 1152 -3426
rect 1146 -3438 1152 -3432
rect 1146 -3444 1152 -3438
rect 1146 -3450 1152 -3444
rect 1146 -3456 1152 -3450
rect 1146 -3462 1152 -3456
rect 1146 -3468 1152 -3462
rect 1146 -3474 1152 -3468
rect 1146 -3480 1152 -3474
rect 1146 -3486 1152 -3480
rect 1146 -3492 1152 -3486
rect 1146 -3498 1152 -3492
rect 1146 -3504 1152 -3498
rect 1146 -3510 1152 -3504
rect 1146 -3516 1152 -3510
rect 1152 -1104 1158 -1098
rect 1152 -1110 1158 -1104
rect 1152 -1116 1158 -1110
rect 1152 -1122 1158 -1116
rect 1152 -1128 1158 -1122
rect 1152 -1134 1158 -1128
rect 1152 -1140 1158 -1134
rect 1152 -1146 1158 -1140
rect 1152 -1152 1158 -1146
rect 1152 -1158 1158 -1152
rect 1152 -1164 1158 -1158
rect 1152 -1170 1158 -1164
rect 1152 -1176 1158 -1170
rect 1152 -1182 1158 -1176
rect 1152 -1188 1158 -1182
rect 1152 -1194 1158 -1188
rect 1152 -1200 1158 -1194
rect 1152 -1206 1158 -1200
rect 1152 -1212 1158 -1206
rect 1152 -1218 1158 -1212
rect 1152 -1224 1158 -1218
rect 1152 -1230 1158 -1224
rect 1152 -1236 1158 -1230
rect 1152 -1242 1158 -1236
rect 1152 -1248 1158 -1242
rect 1152 -1254 1158 -1248
rect 1152 -1260 1158 -1254
rect 1152 -1266 1158 -1260
rect 1152 -1272 1158 -1266
rect 1152 -1278 1158 -1272
rect 1152 -1284 1158 -1278
rect 1152 -1290 1158 -1284
rect 1152 -1296 1158 -1290
rect 1152 -1302 1158 -1296
rect 1152 -1308 1158 -1302
rect 1152 -1938 1158 -1932
rect 1152 -1944 1158 -1938
rect 1152 -1950 1158 -1944
rect 1152 -1956 1158 -1950
rect 1152 -1962 1158 -1956
rect 1152 -1968 1158 -1962
rect 1152 -1974 1158 -1968
rect 1152 -1980 1158 -1974
rect 1152 -1986 1158 -1980
rect 1152 -1992 1158 -1986
rect 1152 -1998 1158 -1992
rect 1152 -2004 1158 -1998
rect 1152 -2010 1158 -2004
rect 1152 -2016 1158 -2010
rect 1152 -2022 1158 -2016
rect 1152 -2028 1158 -2022
rect 1152 -2034 1158 -2028
rect 1152 -2040 1158 -2034
rect 1152 -2046 1158 -2040
rect 1152 -2052 1158 -2046
rect 1152 -2058 1158 -2052
rect 1152 -2064 1158 -2058
rect 1152 -2070 1158 -2064
rect 1152 -2076 1158 -2070
rect 1152 -2082 1158 -2076
rect 1152 -2088 1158 -2082
rect 1152 -2094 1158 -2088
rect 1152 -2100 1158 -2094
rect 1152 -2106 1158 -2100
rect 1152 -2112 1158 -2106
rect 1152 -2118 1158 -2112
rect 1152 -2124 1158 -2118
rect 1152 -2130 1158 -2124
rect 1152 -2136 1158 -2130
rect 1152 -2142 1158 -2136
rect 1152 -2148 1158 -2142
rect 1152 -2154 1158 -2148
rect 1152 -2160 1158 -2154
rect 1152 -2166 1158 -2160
rect 1152 -2172 1158 -2166
rect 1152 -2178 1158 -2172
rect 1152 -2184 1158 -2178
rect 1152 -2190 1158 -2184
rect 1152 -2196 1158 -2190
rect 1152 -2202 1158 -2196
rect 1152 -2208 1158 -2202
rect 1152 -2214 1158 -2208
rect 1152 -2220 1158 -2214
rect 1152 -2226 1158 -2220
rect 1152 -2232 1158 -2226
rect 1152 -2238 1158 -2232
rect 1152 -2244 1158 -2238
rect 1152 -2250 1158 -2244
rect 1152 -2256 1158 -2250
rect 1152 -2262 1158 -2256
rect 1152 -2268 1158 -2262
rect 1152 -2274 1158 -2268
rect 1152 -2280 1158 -2274
rect 1152 -2286 1158 -2280
rect 1152 -2292 1158 -2286
rect 1152 -2298 1158 -2292
rect 1152 -2304 1158 -2298
rect 1152 -2310 1158 -2304
rect 1152 -2316 1158 -2310
rect 1152 -2322 1158 -2316
rect 1152 -2328 1158 -2322
rect 1152 -2334 1158 -2328
rect 1152 -2340 1158 -2334
rect 1152 -2346 1158 -2340
rect 1152 -2352 1158 -2346
rect 1152 -2358 1158 -2352
rect 1152 -2364 1158 -2358
rect 1152 -2370 1158 -2364
rect 1152 -2376 1158 -2370
rect 1152 -2382 1158 -2376
rect 1152 -2388 1158 -2382
rect 1152 -2394 1158 -2388
rect 1152 -2400 1158 -2394
rect 1152 -2406 1158 -2400
rect 1152 -2412 1158 -2406
rect 1152 -2418 1158 -2412
rect 1152 -2424 1158 -2418
rect 1152 -2430 1158 -2424
rect 1152 -2436 1158 -2430
rect 1152 -2442 1158 -2436
rect 1152 -2448 1158 -2442
rect 1152 -2454 1158 -2448
rect 1152 -2460 1158 -2454
rect 1152 -2466 1158 -2460
rect 1152 -2472 1158 -2466
rect 1152 -2478 1158 -2472
rect 1152 -2484 1158 -2478
rect 1152 -2490 1158 -2484
rect 1152 -2496 1158 -2490
rect 1152 -2502 1158 -2496
rect 1152 -2508 1158 -2502
rect 1152 -2514 1158 -2508
rect 1152 -2520 1158 -2514
rect 1152 -2526 1158 -2520
rect 1152 -2532 1158 -2526
rect 1152 -2538 1158 -2532
rect 1152 -2544 1158 -2538
rect 1152 -2550 1158 -2544
rect 1152 -2556 1158 -2550
rect 1152 -2562 1158 -2556
rect 1152 -2568 1158 -2562
rect 1152 -2574 1158 -2568
rect 1152 -2580 1158 -2574
rect 1152 -2586 1158 -2580
rect 1152 -2592 1158 -2586
rect 1152 -2598 1158 -2592
rect 1152 -2604 1158 -2598
rect 1152 -2610 1158 -2604
rect 1152 -2616 1158 -2610
rect 1152 -2622 1158 -2616
rect 1152 -2628 1158 -2622
rect 1152 -2634 1158 -2628
rect 1152 -2640 1158 -2634
rect 1152 -2646 1158 -2640
rect 1152 -2652 1158 -2646
rect 1152 -2658 1158 -2652
rect 1152 -2664 1158 -2658
rect 1152 -2670 1158 -2664
rect 1152 -2676 1158 -2670
rect 1152 -2772 1158 -2766
rect 1152 -2778 1158 -2772
rect 1152 -2784 1158 -2778
rect 1152 -2790 1158 -2784
rect 1152 -2796 1158 -2790
rect 1152 -2802 1158 -2796
rect 1152 -2808 1158 -2802
rect 1152 -2814 1158 -2808
rect 1152 -2820 1158 -2814
rect 1152 -2826 1158 -2820
rect 1152 -2832 1158 -2826
rect 1152 -2838 1158 -2832
rect 1152 -2844 1158 -2838
rect 1152 -2850 1158 -2844
rect 1152 -2856 1158 -2850
rect 1152 -2862 1158 -2856
rect 1152 -2868 1158 -2862
rect 1152 -2874 1158 -2868
rect 1152 -2880 1158 -2874
rect 1152 -2886 1158 -2880
rect 1152 -2892 1158 -2886
rect 1152 -2898 1158 -2892
rect 1152 -2904 1158 -2898
rect 1152 -2910 1158 -2904
rect 1152 -2916 1158 -2910
rect 1152 -2922 1158 -2916
rect 1152 -2928 1158 -2922
rect 1152 -2934 1158 -2928
rect 1152 -2940 1158 -2934
rect 1152 -2946 1158 -2940
rect 1152 -2952 1158 -2946
rect 1152 -2958 1158 -2952
rect 1152 -2964 1158 -2958
rect 1152 -2970 1158 -2964
rect 1152 -2976 1158 -2970
rect 1152 -2982 1158 -2976
rect 1152 -2988 1158 -2982
rect 1152 -2994 1158 -2988
rect 1152 -3000 1158 -2994
rect 1152 -3006 1158 -3000
rect 1152 -3012 1158 -3006
rect 1152 -3018 1158 -3012
rect 1152 -3024 1158 -3018
rect 1152 -3030 1158 -3024
rect 1152 -3036 1158 -3030
rect 1152 -3042 1158 -3036
rect 1152 -3048 1158 -3042
rect 1152 -3054 1158 -3048
rect 1152 -3132 1158 -3126
rect 1152 -3138 1158 -3132
rect 1152 -3144 1158 -3138
rect 1152 -3150 1158 -3144
rect 1152 -3156 1158 -3150
rect 1152 -3162 1158 -3156
rect 1152 -3168 1158 -3162
rect 1152 -3174 1158 -3168
rect 1152 -3180 1158 -3174
rect 1152 -3186 1158 -3180
rect 1152 -3192 1158 -3186
rect 1152 -3198 1158 -3192
rect 1152 -3204 1158 -3198
rect 1152 -3210 1158 -3204
rect 1152 -3216 1158 -3210
rect 1152 -3222 1158 -3216
rect 1152 -3228 1158 -3222
rect 1152 -3234 1158 -3228
rect 1152 -3240 1158 -3234
rect 1152 -3246 1158 -3240
rect 1152 -3252 1158 -3246
rect 1152 -3318 1158 -3312
rect 1152 -3324 1158 -3318
rect 1152 -3330 1158 -3324
rect 1152 -3336 1158 -3330
rect 1152 -3342 1158 -3336
rect 1152 -3348 1158 -3342
rect 1152 -3354 1158 -3348
rect 1152 -3360 1158 -3354
rect 1152 -3366 1158 -3360
rect 1152 -3372 1158 -3366
rect 1152 -3378 1158 -3372
rect 1152 -3384 1158 -3378
rect 1152 -3390 1158 -3384
rect 1152 -3396 1158 -3390
rect 1152 -3402 1158 -3396
rect 1152 -3408 1158 -3402
rect 1152 -3414 1158 -3408
rect 1152 -3420 1158 -3414
rect 1152 -3426 1158 -3420
rect 1152 -3432 1158 -3426
rect 1152 -3438 1158 -3432
rect 1152 -3444 1158 -3438
rect 1152 -3450 1158 -3444
rect 1152 -3456 1158 -3450
rect 1152 -3462 1158 -3456
rect 1152 -3468 1158 -3462
rect 1152 -3474 1158 -3468
rect 1152 -3480 1158 -3474
rect 1152 -3486 1158 -3480
rect 1152 -3492 1158 -3486
rect 1152 -3498 1158 -3492
rect 1152 -3504 1158 -3498
rect 1152 -3510 1158 -3504
rect 1152 -3516 1158 -3510
rect 1158 -1104 1164 -1098
rect 1158 -1110 1164 -1104
rect 1158 -1116 1164 -1110
rect 1158 -1122 1164 -1116
rect 1158 -1128 1164 -1122
rect 1158 -1134 1164 -1128
rect 1158 -1140 1164 -1134
rect 1158 -1146 1164 -1140
rect 1158 -1152 1164 -1146
rect 1158 -1158 1164 -1152
rect 1158 -1164 1164 -1158
rect 1158 -1170 1164 -1164
rect 1158 -1176 1164 -1170
rect 1158 -1182 1164 -1176
rect 1158 -1188 1164 -1182
rect 1158 -1194 1164 -1188
rect 1158 -1200 1164 -1194
rect 1158 -1206 1164 -1200
rect 1158 -1212 1164 -1206
rect 1158 -1218 1164 -1212
rect 1158 -1224 1164 -1218
rect 1158 -1230 1164 -1224
rect 1158 -1236 1164 -1230
rect 1158 -1242 1164 -1236
rect 1158 -1248 1164 -1242
rect 1158 -1254 1164 -1248
rect 1158 -1260 1164 -1254
rect 1158 -1266 1164 -1260
rect 1158 -1272 1164 -1266
rect 1158 -1278 1164 -1272
rect 1158 -1284 1164 -1278
rect 1158 -1290 1164 -1284
rect 1158 -1296 1164 -1290
rect 1158 -1302 1164 -1296
rect 1158 -1308 1164 -1302
rect 1158 -1920 1164 -1914
rect 1158 -1926 1164 -1920
rect 1158 -1932 1164 -1926
rect 1158 -1938 1164 -1932
rect 1158 -1944 1164 -1938
rect 1158 -1950 1164 -1944
rect 1158 -1956 1164 -1950
rect 1158 -1962 1164 -1956
rect 1158 -1968 1164 -1962
rect 1158 -1974 1164 -1968
rect 1158 -1980 1164 -1974
rect 1158 -1986 1164 -1980
rect 1158 -1992 1164 -1986
rect 1158 -1998 1164 -1992
rect 1158 -2004 1164 -1998
rect 1158 -2010 1164 -2004
rect 1158 -2016 1164 -2010
rect 1158 -2022 1164 -2016
rect 1158 -2028 1164 -2022
rect 1158 -2034 1164 -2028
rect 1158 -2040 1164 -2034
rect 1158 -2046 1164 -2040
rect 1158 -2052 1164 -2046
rect 1158 -2058 1164 -2052
rect 1158 -2064 1164 -2058
rect 1158 -2070 1164 -2064
rect 1158 -2076 1164 -2070
rect 1158 -2082 1164 -2076
rect 1158 -2088 1164 -2082
rect 1158 -2094 1164 -2088
rect 1158 -2100 1164 -2094
rect 1158 -2106 1164 -2100
rect 1158 -2112 1164 -2106
rect 1158 -2118 1164 -2112
rect 1158 -2124 1164 -2118
rect 1158 -2130 1164 -2124
rect 1158 -2136 1164 -2130
rect 1158 -2142 1164 -2136
rect 1158 -2148 1164 -2142
rect 1158 -2154 1164 -2148
rect 1158 -2160 1164 -2154
rect 1158 -2166 1164 -2160
rect 1158 -2172 1164 -2166
rect 1158 -2178 1164 -2172
rect 1158 -2184 1164 -2178
rect 1158 -2190 1164 -2184
rect 1158 -2196 1164 -2190
rect 1158 -2202 1164 -2196
rect 1158 -2208 1164 -2202
rect 1158 -2214 1164 -2208
rect 1158 -2220 1164 -2214
rect 1158 -2226 1164 -2220
rect 1158 -2232 1164 -2226
rect 1158 -2238 1164 -2232
rect 1158 -2244 1164 -2238
rect 1158 -2250 1164 -2244
rect 1158 -2256 1164 -2250
rect 1158 -2262 1164 -2256
rect 1158 -2268 1164 -2262
rect 1158 -2274 1164 -2268
rect 1158 -2280 1164 -2274
rect 1158 -2286 1164 -2280
rect 1158 -2292 1164 -2286
rect 1158 -2298 1164 -2292
rect 1158 -2304 1164 -2298
rect 1158 -2310 1164 -2304
rect 1158 -2316 1164 -2310
rect 1158 -2322 1164 -2316
rect 1158 -2328 1164 -2322
rect 1158 -2334 1164 -2328
rect 1158 -2340 1164 -2334
rect 1158 -2346 1164 -2340
rect 1158 -2352 1164 -2346
rect 1158 -2358 1164 -2352
rect 1158 -2364 1164 -2358
rect 1158 -2370 1164 -2364
rect 1158 -2376 1164 -2370
rect 1158 -2382 1164 -2376
rect 1158 -2388 1164 -2382
rect 1158 -2394 1164 -2388
rect 1158 -2400 1164 -2394
rect 1158 -2406 1164 -2400
rect 1158 -2412 1164 -2406
rect 1158 -2418 1164 -2412
rect 1158 -2424 1164 -2418
rect 1158 -2430 1164 -2424
rect 1158 -2436 1164 -2430
rect 1158 -2442 1164 -2436
rect 1158 -2448 1164 -2442
rect 1158 -2454 1164 -2448
rect 1158 -2460 1164 -2454
rect 1158 -2466 1164 -2460
rect 1158 -2472 1164 -2466
rect 1158 -2478 1164 -2472
rect 1158 -2484 1164 -2478
rect 1158 -2490 1164 -2484
rect 1158 -2496 1164 -2490
rect 1158 -2502 1164 -2496
rect 1158 -2508 1164 -2502
rect 1158 -2514 1164 -2508
rect 1158 -2520 1164 -2514
rect 1158 -2526 1164 -2520
rect 1158 -2532 1164 -2526
rect 1158 -2538 1164 -2532
rect 1158 -2544 1164 -2538
rect 1158 -2550 1164 -2544
rect 1158 -2556 1164 -2550
rect 1158 -2562 1164 -2556
rect 1158 -2568 1164 -2562
rect 1158 -2574 1164 -2568
rect 1158 -2580 1164 -2574
rect 1158 -2586 1164 -2580
rect 1158 -2592 1164 -2586
rect 1158 -2598 1164 -2592
rect 1158 -2604 1164 -2598
rect 1158 -2610 1164 -2604
rect 1158 -2616 1164 -2610
rect 1158 -2622 1164 -2616
rect 1158 -2628 1164 -2622
rect 1158 -2634 1164 -2628
rect 1158 -2640 1164 -2634
rect 1158 -2646 1164 -2640
rect 1158 -2652 1164 -2646
rect 1158 -2658 1164 -2652
rect 1158 -2664 1164 -2658
rect 1158 -2670 1164 -2664
rect 1158 -2766 1164 -2760
rect 1158 -2772 1164 -2766
rect 1158 -2778 1164 -2772
rect 1158 -2784 1164 -2778
rect 1158 -2790 1164 -2784
rect 1158 -2796 1164 -2790
rect 1158 -2802 1164 -2796
rect 1158 -2808 1164 -2802
rect 1158 -2814 1164 -2808
rect 1158 -2820 1164 -2814
rect 1158 -2826 1164 -2820
rect 1158 -2832 1164 -2826
rect 1158 -2838 1164 -2832
rect 1158 -2844 1164 -2838
rect 1158 -2850 1164 -2844
rect 1158 -2856 1164 -2850
rect 1158 -2862 1164 -2856
rect 1158 -2868 1164 -2862
rect 1158 -2874 1164 -2868
rect 1158 -2880 1164 -2874
rect 1158 -2886 1164 -2880
rect 1158 -2892 1164 -2886
rect 1158 -2898 1164 -2892
rect 1158 -2904 1164 -2898
rect 1158 -2910 1164 -2904
rect 1158 -2916 1164 -2910
rect 1158 -2922 1164 -2916
rect 1158 -2928 1164 -2922
rect 1158 -2934 1164 -2928
rect 1158 -2940 1164 -2934
rect 1158 -2946 1164 -2940
rect 1158 -2952 1164 -2946
rect 1158 -2958 1164 -2952
rect 1158 -2964 1164 -2958
rect 1158 -2970 1164 -2964
rect 1158 -2976 1164 -2970
rect 1158 -2982 1164 -2976
rect 1158 -2988 1164 -2982
rect 1158 -2994 1164 -2988
rect 1158 -3000 1164 -2994
rect 1158 -3006 1164 -3000
rect 1158 -3012 1164 -3006
rect 1158 -3018 1164 -3012
rect 1158 -3024 1164 -3018
rect 1158 -3030 1164 -3024
rect 1158 -3036 1164 -3030
rect 1158 -3042 1164 -3036
rect 1158 -3048 1164 -3042
rect 1158 -3054 1164 -3048
rect 1158 -3126 1164 -3120
rect 1158 -3132 1164 -3126
rect 1158 -3138 1164 -3132
rect 1158 -3144 1164 -3138
rect 1158 -3150 1164 -3144
rect 1158 -3156 1164 -3150
rect 1158 -3162 1164 -3156
rect 1158 -3168 1164 -3162
rect 1158 -3174 1164 -3168
rect 1158 -3180 1164 -3174
rect 1158 -3186 1164 -3180
rect 1158 -3192 1164 -3186
rect 1158 -3198 1164 -3192
rect 1158 -3204 1164 -3198
rect 1158 -3210 1164 -3204
rect 1158 -3216 1164 -3210
rect 1158 -3222 1164 -3216
rect 1158 -3228 1164 -3222
rect 1158 -3234 1164 -3228
rect 1158 -3240 1164 -3234
rect 1158 -3246 1164 -3240
rect 1158 -3252 1164 -3246
rect 1158 -3318 1164 -3312
rect 1158 -3324 1164 -3318
rect 1158 -3330 1164 -3324
rect 1158 -3336 1164 -3330
rect 1158 -3342 1164 -3336
rect 1158 -3348 1164 -3342
rect 1158 -3354 1164 -3348
rect 1158 -3360 1164 -3354
rect 1158 -3366 1164 -3360
rect 1158 -3372 1164 -3366
rect 1158 -3378 1164 -3372
rect 1158 -3384 1164 -3378
rect 1158 -3390 1164 -3384
rect 1158 -3396 1164 -3390
rect 1158 -3402 1164 -3396
rect 1158 -3408 1164 -3402
rect 1158 -3414 1164 -3408
rect 1158 -3420 1164 -3414
rect 1158 -3426 1164 -3420
rect 1158 -3432 1164 -3426
rect 1158 -3438 1164 -3432
rect 1158 -3444 1164 -3438
rect 1158 -3450 1164 -3444
rect 1158 -3456 1164 -3450
rect 1158 -3462 1164 -3456
rect 1158 -3468 1164 -3462
rect 1158 -3474 1164 -3468
rect 1158 -3480 1164 -3474
rect 1158 -3486 1164 -3480
rect 1158 -3492 1164 -3486
rect 1158 -3498 1164 -3492
rect 1158 -3504 1164 -3498
rect 1158 -3510 1164 -3504
rect 1158 -3516 1164 -3510
rect 1164 -1104 1170 -1098
rect 1164 -1110 1170 -1104
rect 1164 -1116 1170 -1110
rect 1164 -1122 1170 -1116
rect 1164 -1128 1170 -1122
rect 1164 -1134 1170 -1128
rect 1164 -1140 1170 -1134
rect 1164 -1146 1170 -1140
rect 1164 -1152 1170 -1146
rect 1164 -1158 1170 -1152
rect 1164 -1164 1170 -1158
rect 1164 -1170 1170 -1164
rect 1164 -1176 1170 -1170
rect 1164 -1182 1170 -1176
rect 1164 -1188 1170 -1182
rect 1164 -1194 1170 -1188
rect 1164 -1200 1170 -1194
rect 1164 -1206 1170 -1200
rect 1164 -1212 1170 -1206
rect 1164 -1218 1170 -1212
rect 1164 -1224 1170 -1218
rect 1164 -1230 1170 -1224
rect 1164 -1236 1170 -1230
rect 1164 -1242 1170 -1236
rect 1164 -1248 1170 -1242
rect 1164 -1254 1170 -1248
rect 1164 -1260 1170 -1254
rect 1164 -1266 1170 -1260
rect 1164 -1272 1170 -1266
rect 1164 -1278 1170 -1272
rect 1164 -1284 1170 -1278
rect 1164 -1290 1170 -1284
rect 1164 -1296 1170 -1290
rect 1164 -1302 1170 -1296
rect 1164 -1308 1170 -1302
rect 1164 -1908 1170 -1902
rect 1164 -1914 1170 -1908
rect 1164 -1920 1170 -1914
rect 1164 -1926 1170 -1920
rect 1164 -1932 1170 -1926
rect 1164 -1938 1170 -1932
rect 1164 -1944 1170 -1938
rect 1164 -1950 1170 -1944
rect 1164 -1956 1170 -1950
rect 1164 -1962 1170 -1956
rect 1164 -1968 1170 -1962
rect 1164 -1974 1170 -1968
rect 1164 -1980 1170 -1974
rect 1164 -1986 1170 -1980
rect 1164 -1992 1170 -1986
rect 1164 -1998 1170 -1992
rect 1164 -2004 1170 -1998
rect 1164 -2010 1170 -2004
rect 1164 -2016 1170 -2010
rect 1164 -2022 1170 -2016
rect 1164 -2028 1170 -2022
rect 1164 -2034 1170 -2028
rect 1164 -2040 1170 -2034
rect 1164 -2046 1170 -2040
rect 1164 -2052 1170 -2046
rect 1164 -2058 1170 -2052
rect 1164 -2064 1170 -2058
rect 1164 -2070 1170 -2064
rect 1164 -2076 1170 -2070
rect 1164 -2082 1170 -2076
rect 1164 -2088 1170 -2082
rect 1164 -2094 1170 -2088
rect 1164 -2100 1170 -2094
rect 1164 -2106 1170 -2100
rect 1164 -2112 1170 -2106
rect 1164 -2118 1170 -2112
rect 1164 -2124 1170 -2118
rect 1164 -2130 1170 -2124
rect 1164 -2136 1170 -2130
rect 1164 -2142 1170 -2136
rect 1164 -2148 1170 -2142
rect 1164 -2154 1170 -2148
rect 1164 -2160 1170 -2154
rect 1164 -2166 1170 -2160
rect 1164 -2172 1170 -2166
rect 1164 -2178 1170 -2172
rect 1164 -2184 1170 -2178
rect 1164 -2190 1170 -2184
rect 1164 -2196 1170 -2190
rect 1164 -2202 1170 -2196
rect 1164 -2208 1170 -2202
rect 1164 -2214 1170 -2208
rect 1164 -2220 1170 -2214
rect 1164 -2226 1170 -2220
rect 1164 -2232 1170 -2226
rect 1164 -2238 1170 -2232
rect 1164 -2244 1170 -2238
rect 1164 -2250 1170 -2244
rect 1164 -2256 1170 -2250
rect 1164 -2262 1170 -2256
rect 1164 -2268 1170 -2262
rect 1164 -2274 1170 -2268
rect 1164 -2280 1170 -2274
rect 1164 -2286 1170 -2280
rect 1164 -2292 1170 -2286
rect 1164 -2298 1170 -2292
rect 1164 -2304 1170 -2298
rect 1164 -2310 1170 -2304
rect 1164 -2316 1170 -2310
rect 1164 -2322 1170 -2316
rect 1164 -2328 1170 -2322
rect 1164 -2334 1170 -2328
rect 1164 -2340 1170 -2334
rect 1164 -2346 1170 -2340
rect 1164 -2352 1170 -2346
rect 1164 -2358 1170 -2352
rect 1164 -2364 1170 -2358
rect 1164 -2370 1170 -2364
rect 1164 -2376 1170 -2370
rect 1164 -2382 1170 -2376
rect 1164 -2388 1170 -2382
rect 1164 -2394 1170 -2388
rect 1164 -2400 1170 -2394
rect 1164 -2406 1170 -2400
rect 1164 -2412 1170 -2406
rect 1164 -2418 1170 -2412
rect 1164 -2424 1170 -2418
rect 1164 -2430 1170 -2424
rect 1164 -2436 1170 -2430
rect 1164 -2442 1170 -2436
rect 1164 -2448 1170 -2442
rect 1164 -2454 1170 -2448
rect 1164 -2460 1170 -2454
rect 1164 -2466 1170 -2460
rect 1164 -2472 1170 -2466
rect 1164 -2478 1170 -2472
rect 1164 -2484 1170 -2478
rect 1164 -2490 1170 -2484
rect 1164 -2496 1170 -2490
rect 1164 -2502 1170 -2496
rect 1164 -2508 1170 -2502
rect 1164 -2514 1170 -2508
rect 1164 -2520 1170 -2514
rect 1164 -2526 1170 -2520
rect 1164 -2532 1170 -2526
rect 1164 -2538 1170 -2532
rect 1164 -2544 1170 -2538
rect 1164 -2550 1170 -2544
rect 1164 -2556 1170 -2550
rect 1164 -2562 1170 -2556
rect 1164 -2568 1170 -2562
rect 1164 -2574 1170 -2568
rect 1164 -2580 1170 -2574
rect 1164 -2586 1170 -2580
rect 1164 -2592 1170 -2586
rect 1164 -2598 1170 -2592
rect 1164 -2604 1170 -2598
rect 1164 -2610 1170 -2604
rect 1164 -2616 1170 -2610
rect 1164 -2622 1170 -2616
rect 1164 -2628 1170 -2622
rect 1164 -2634 1170 -2628
rect 1164 -2640 1170 -2634
rect 1164 -2646 1170 -2640
rect 1164 -2652 1170 -2646
rect 1164 -2658 1170 -2652
rect 1164 -2754 1170 -2748
rect 1164 -2760 1170 -2754
rect 1164 -2766 1170 -2760
rect 1164 -2772 1170 -2766
rect 1164 -2778 1170 -2772
rect 1164 -2784 1170 -2778
rect 1164 -2790 1170 -2784
rect 1164 -2796 1170 -2790
rect 1164 -2802 1170 -2796
rect 1164 -2808 1170 -2802
rect 1164 -2814 1170 -2808
rect 1164 -2820 1170 -2814
rect 1164 -2826 1170 -2820
rect 1164 -2832 1170 -2826
rect 1164 -2838 1170 -2832
rect 1164 -2844 1170 -2838
rect 1164 -2850 1170 -2844
rect 1164 -2856 1170 -2850
rect 1164 -2862 1170 -2856
rect 1164 -2868 1170 -2862
rect 1164 -2874 1170 -2868
rect 1164 -2880 1170 -2874
rect 1164 -2886 1170 -2880
rect 1164 -2892 1170 -2886
rect 1164 -2898 1170 -2892
rect 1164 -2904 1170 -2898
rect 1164 -2910 1170 -2904
rect 1164 -2916 1170 -2910
rect 1164 -2922 1170 -2916
rect 1164 -2928 1170 -2922
rect 1164 -2934 1170 -2928
rect 1164 -2940 1170 -2934
rect 1164 -2946 1170 -2940
rect 1164 -2952 1170 -2946
rect 1164 -2958 1170 -2952
rect 1164 -2964 1170 -2958
rect 1164 -2970 1170 -2964
rect 1164 -2976 1170 -2970
rect 1164 -2982 1170 -2976
rect 1164 -2988 1170 -2982
rect 1164 -2994 1170 -2988
rect 1164 -3000 1170 -2994
rect 1164 -3006 1170 -3000
rect 1164 -3012 1170 -3006
rect 1164 -3018 1170 -3012
rect 1164 -3024 1170 -3018
rect 1164 -3030 1170 -3024
rect 1164 -3036 1170 -3030
rect 1164 -3042 1170 -3036
rect 1164 -3048 1170 -3042
rect 1164 -3120 1170 -3114
rect 1164 -3126 1170 -3120
rect 1164 -3132 1170 -3126
rect 1164 -3138 1170 -3132
rect 1164 -3144 1170 -3138
rect 1164 -3150 1170 -3144
rect 1164 -3156 1170 -3150
rect 1164 -3162 1170 -3156
rect 1164 -3168 1170 -3162
rect 1164 -3174 1170 -3168
rect 1164 -3180 1170 -3174
rect 1164 -3186 1170 -3180
rect 1164 -3192 1170 -3186
rect 1164 -3198 1170 -3192
rect 1164 -3204 1170 -3198
rect 1164 -3210 1170 -3204
rect 1164 -3216 1170 -3210
rect 1164 -3222 1170 -3216
rect 1164 -3228 1170 -3222
rect 1164 -3234 1170 -3228
rect 1164 -3240 1170 -3234
rect 1164 -3246 1170 -3240
rect 1164 -3252 1170 -3246
rect 1164 -3318 1170 -3312
rect 1164 -3324 1170 -3318
rect 1164 -3330 1170 -3324
rect 1164 -3336 1170 -3330
rect 1164 -3342 1170 -3336
rect 1164 -3348 1170 -3342
rect 1164 -3354 1170 -3348
rect 1164 -3360 1170 -3354
rect 1164 -3366 1170 -3360
rect 1164 -3372 1170 -3366
rect 1164 -3378 1170 -3372
rect 1164 -3384 1170 -3378
rect 1164 -3390 1170 -3384
rect 1164 -3396 1170 -3390
rect 1164 -3402 1170 -3396
rect 1164 -3408 1170 -3402
rect 1164 -3414 1170 -3408
rect 1164 -3420 1170 -3414
rect 1164 -3426 1170 -3420
rect 1164 -3432 1170 -3426
rect 1164 -3438 1170 -3432
rect 1164 -3444 1170 -3438
rect 1164 -3450 1170 -3444
rect 1164 -3456 1170 -3450
rect 1164 -3462 1170 -3456
rect 1164 -3468 1170 -3462
rect 1164 -3474 1170 -3468
rect 1164 -3480 1170 -3474
rect 1164 -3486 1170 -3480
rect 1164 -3492 1170 -3486
rect 1164 -3498 1170 -3492
rect 1164 -3504 1170 -3498
rect 1164 -3510 1170 -3504
rect 1164 -3516 1170 -3510
rect 1170 -1104 1176 -1098
rect 1170 -1110 1176 -1104
rect 1170 -1116 1176 -1110
rect 1170 -1122 1176 -1116
rect 1170 -1128 1176 -1122
rect 1170 -1134 1176 -1128
rect 1170 -1140 1176 -1134
rect 1170 -1146 1176 -1140
rect 1170 -1152 1176 -1146
rect 1170 -1158 1176 -1152
rect 1170 -1164 1176 -1158
rect 1170 -1170 1176 -1164
rect 1170 -1176 1176 -1170
rect 1170 -1182 1176 -1176
rect 1170 -1188 1176 -1182
rect 1170 -1194 1176 -1188
rect 1170 -1200 1176 -1194
rect 1170 -1206 1176 -1200
rect 1170 -1212 1176 -1206
rect 1170 -1218 1176 -1212
rect 1170 -1224 1176 -1218
rect 1170 -1230 1176 -1224
rect 1170 -1236 1176 -1230
rect 1170 -1242 1176 -1236
rect 1170 -1248 1176 -1242
rect 1170 -1254 1176 -1248
rect 1170 -1260 1176 -1254
rect 1170 -1266 1176 -1260
rect 1170 -1272 1176 -1266
rect 1170 -1278 1176 -1272
rect 1170 -1284 1176 -1278
rect 1170 -1290 1176 -1284
rect 1170 -1296 1176 -1290
rect 1170 -1302 1176 -1296
rect 1170 -1308 1176 -1302
rect 1170 -1890 1176 -1884
rect 1170 -1896 1176 -1890
rect 1170 -1902 1176 -1896
rect 1170 -1908 1176 -1902
rect 1170 -1914 1176 -1908
rect 1170 -1920 1176 -1914
rect 1170 -1926 1176 -1920
rect 1170 -1932 1176 -1926
rect 1170 -1938 1176 -1932
rect 1170 -1944 1176 -1938
rect 1170 -1950 1176 -1944
rect 1170 -1956 1176 -1950
rect 1170 -1962 1176 -1956
rect 1170 -1968 1176 -1962
rect 1170 -1974 1176 -1968
rect 1170 -1980 1176 -1974
rect 1170 -1986 1176 -1980
rect 1170 -1992 1176 -1986
rect 1170 -1998 1176 -1992
rect 1170 -2004 1176 -1998
rect 1170 -2010 1176 -2004
rect 1170 -2016 1176 -2010
rect 1170 -2022 1176 -2016
rect 1170 -2028 1176 -2022
rect 1170 -2034 1176 -2028
rect 1170 -2040 1176 -2034
rect 1170 -2046 1176 -2040
rect 1170 -2052 1176 -2046
rect 1170 -2058 1176 -2052
rect 1170 -2064 1176 -2058
rect 1170 -2070 1176 -2064
rect 1170 -2076 1176 -2070
rect 1170 -2082 1176 -2076
rect 1170 -2088 1176 -2082
rect 1170 -2094 1176 -2088
rect 1170 -2100 1176 -2094
rect 1170 -2106 1176 -2100
rect 1170 -2112 1176 -2106
rect 1170 -2118 1176 -2112
rect 1170 -2124 1176 -2118
rect 1170 -2130 1176 -2124
rect 1170 -2136 1176 -2130
rect 1170 -2142 1176 -2136
rect 1170 -2148 1176 -2142
rect 1170 -2154 1176 -2148
rect 1170 -2160 1176 -2154
rect 1170 -2166 1176 -2160
rect 1170 -2172 1176 -2166
rect 1170 -2178 1176 -2172
rect 1170 -2184 1176 -2178
rect 1170 -2190 1176 -2184
rect 1170 -2196 1176 -2190
rect 1170 -2202 1176 -2196
rect 1170 -2208 1176 -2202
rect 1170 -2214 1176 -2208
rect 1170 -2220 1176 -2214
rect 1170 -2226 1176 -2220
rect 1170 -2232 1176 -2226
rect 1170 -2238 1176 -2232
rect 1170 -2244 1176 -2238
rect 1170 -2250 1176 -2244
rect 1170 -2256 1176 -2250
rect 1170 -2262 1176 -2256
rect 1170 -2268 1176 -2262
rect 1170 -2274 1176 -2268
rect 1170 -2280 1176 -2274
rect 1170 -2286 1176 -2280
rect 1170 -2292 1176 -2286
rect 1170 -2298 1176 -2292
rect 1170 -2304 1176 -2298
rect 1170 -2310 1176 -2304
rect 1170 -2316 1176 -2310
rect 1170 -2322 1176 -2316
rect 1170 -2328 1176 -2322
rect 1170 -2334 1176 -2328
rect 1170 -2340 1176 -2334
rect 1170 -2346 1176 -2340
rect 1170 -2352 1176 -2346
rect 1170 -2358 1176 -2352
rect 1170 -2364 1176 -2358
rect 1170 -2370 1176 -2364
rect 1170 -2376 1176 -2370
rect 1170 -2382 1176 -2376
rect 1170 -2388 1176 -2382
rect 1170 -2394 1176 -2388
rect 1170 -2400 1176 -2394
rect 1170 -2406 1176 -2400
rect 1170 -2412 1176 -2406
rect 1170 -2418 1176 -2412
rect 1170 -2424 1176 -2418
rect 1170 -2430 1176 -2424
rect 1170 -2436 1176 -2430
rect 1170 -2442 1176 -2436
rect 1170 -2448 1176 -2442
rect 1170 -2454 1176 -2448
rect 1170 -2460 1176 -2454
rect 1170 -2466 1176 -2460
rect 1170 -2472 1176 -2466
rect 1170 -2478 1176 -2472
rect 1170 -2484 1176 -2478
rect 1170 -2490 1176 -2484
rect 1170 -2496 1176 -2490
rect 1170 -2502 1176 -2496
rect 1170 -2508 1176 -2502
rect 1170 -2514 1176 -2508
rect 1170 -2520 1176 -2514
rect 1170 -2526 1176 -2520
rect 1170 -2532 1176 -2526
rect 1170 -2538 1176 -2532
rect 1170 -2544 1176 -2538
rect 1170 -2550 1176 -2544
rect 1170 -2556 1176 -2550
rect 1170 -2562 1176 -2556
rect 1170 -2568 1176 -2562
rect 1170 -2574 1176 -2568
rect 1170 -2580 1176 -2574
rect 1170 -2586 1176 -2580
rect 1170 -2592 1176 -2586
rect 1170 -2598 1176 -2592
rect 1170 -2604 1176 -2598
rect 1170 -2610 1176 -2604
rect 1170 -2616 1176 -2610
rect 1170 -2622 1176 -2616
rect 1170 -2628 1176 -2622
rect 1170 -2634 1176 -2628
rect 1170 -2640 1176 -2634
rect 1170 -2646 1176 -2640
rect 1170 -2652 1176 -2646
rect 1170 -2748 1176 -2742
rect 1170 -2754 1176 -2748
rect 1170 -2760 1176 -2754
rect 1170 -2766 1176 -2760
rect 1170 -2772 1176 -2766
rect 1170 -2778 1176 -2772
rect 1170 -2784 1176 -2778
rect 1170 -2790 1176 -2784
rect 1170 -2796 1176 -2790
rect 1170 -2802 1176 -2796
rect 1170 -2808 1176 -2802
rect 1170 -2814 1176 -2808
rect 1170 -2820 1176 -2814
rect 1170 -2826 1176 -2820
rect 1170 -2832 1176 -2826
rect 1170 -2838 1176 -2832
rect 1170 -2844 1176 -2838
rect 1170 -2850 1176 -2844
rect 1170 -2856 1176 -2850
rect 1170 -2862 1176 -2856
rect 1170 -2868 1176 -2862
rect 1170 -2874 1176 -2868
rect 1170 -2880 1176 -2874
rect 1170 -2886 1176 -2880
rect 1170 -2892 1176 -2886
rect 1170 -2898 1176 -2892
rect 1170 -2904 1176 -2898
rect 1170 -2910 1176 -2904
rect 1170 -2916 1176 -2910
rect 1170 -2922 1176 -2916
rect 1170 -2928 1176 -2922
rect 1170 -2934 1176 -2928
rect 1170 -2940 1176 -2934
rect 1170 -2946 1176 -2940
rect 1170 -2952 1176 -2946
rect 1170 -2958 1176 -2952
rect 1170 -2964 1176 -2958
rect 1170 -2970 1176 -2964
rect 1170 -2976 1176 -2970
rect 1170 -2982 1176 -2976
rect 1170 -2988 1176 -2982
rect 1170 -2994 1176 -2988
rect 1170 -3000 1176 -2994
rect 1170 -3006 1176 -3000
rect 1170 -3012 1176 -3006
rect 1170 -3018 1176 -3012
rect 1170 -3024 1176 -3018
rect 1170 -3030 1176 -3024
rect 1170 -3036 1176 -3030
rect 1170 -3042 1176 -3036
rect 1170 -3120 1176 -3114
rect 1170 -3126 1176 -3120
rect 1170 -3132 1176 -3126
rect 1170 -3138 1176 -3132
rect 1170 -3144 1176 -3138
rect 1170 -3150 1176 -3144
rect 1170 -3156 1176 -3150
rect 1170 -3162 1176 -3156
rect 1170 -3168 1176 -3162
rect 1170 -3174 1176 -3168
rect 1170 -3180 1176 -3174
rect 1170 -3186 1176 -3180
rect 1170 -3192 1176 -3186
rect 1170 -3198 1176 -3192
rect 1170 -3204 1176 -3198
rect 1170 -3210 1176 -3204
rect 1170 -3216 1176 -3210
rect 1170 -3222 1176 -3216
rect 1170 -3228 1176 -3222
rect 1170 -3234 1176 -3228
rect 1170 -3240 1176 -3234
rect 1170 -3246 1176 -3240
rect 1170 -3252 1176 -3246
rect 1170 -3324 1176 -3318
rect 1170 -3330 1176 -3324
rect 1170 -3336 1176 -3330
rect 1170 -3342 1176 -3336
rect 1170 -3348 1176 -3342
rect 1170 -3354 1176 -3348
rect 1170 -3360 1176 -3354
rect 1170 -3366 1176 -3360
rect 1170 -3372 1176 -3366
rect 1170 -3378 1176 -3372
rect 1170 -3384 1176 -3378
rect 1170 -3390 1176 -3384
rect 1170 -3396 1176 -3390
rect 1170 -3402 1176 -3396
rect 1170 -3408 1176 -3402
rect 1170 -3414 1176 -3408
rect 1170 -3420 1176 -3414
rect 1170 -3426 1176 -3420
rect 1170 -3432 1176 -3426
rect 1170 -3438 1176 -3432
rect 1170 -3444 1176 -3438
rect 1170 -3450 1176 -3444
rect 1170 -3456 1176 -3450
rect 1170 -3462 1176 -3456
rect 1170 -3468 1176 -3462
rect 1170 -3474 1176 -3468
rect 1170 -3480 1176 -3474
rect 1170 -3486 1176 -3480
rect 1170 -3492 1176 -3486
rect 1170 -3498 1176 -3492
rect 1170 -3504 1176 -3498
rect 1170 -3510 1176 -3504
rect 1170 -3516 1176 -3510
rect 1176 -1104 1182 -1098
rect 1176 -1110 1182 -1104
rect 1176 -1116 1182 -1110
rect 1176 -1122 1182 -1116
rect 1176 -1128 1182 -1122
rect 1176 -1134 1182 -1128
rect 1176 -1140 1182 -1134
rect 1176 -1146 1182 -1140
rect 1176 -1152 1182 -1146
rect 1176 -1158 1182 -1152
rect 1176 -1164 1182 -1158
rect 1176 -1170 1182 -1164
rect 1176 -1176 1182 -1170
rect 1176 -1182 1182 -1176
rect 1176 -1188 1182 -1182
rect 1176 -1194 1182 -1188
rect 1176 -1200 1182 -1194
rect 1176 -1206 1182 -1200
rect 1176 -1212 1182 -1206
rect 1176 -1218 1182 -1212
rect 1176 -1224 1182 -1218
rect 1176 -1230 1182 -1224
rect 1176 -1236 1182 -1230
rect 1176 -1242 1182 -1236
rect 1176 -1248 1182 -1242
rect 1176 -1254 1182 -1248
rect 1176 -1260 1182 -1254
rect 1176 -1266 1182 -1260
rect 1176 -1272 1182 -1266
rect 1176 -1278 1182 -1272
rect 1176 -1284 1182 -1278
rect 1176 -1290 1182 -1284
rect 1176 -1296 1182 -1290
rect 1176 -1302 1182 -1296
rect 1176 -1308 1182 -1302
rect 1176 -1872 1182 -1866
rect 1176 -1878 1182 -1872
rect 1176 -1884 1182 -1878
rect 1176 -1890 1182 -1884
rect 1176 -1896 1182 -1890
rect 1176 -1902 1182 -1896
rect 1176 -1908 1182 -1902
rect 1176 -1914 1182 -1908
rect 1176 -1920 1182 -1914
rect 1176 -1926 1182 -1920
rect 1176 -1932 1182 -1926
rect 1176 -1938 1182 -1932
rect 1176 -1944 1182 -1938
rect 1176 -1950 1182 -1944
rect 1176 -1956 1182 -1950
rect 1176 -1962 1182 -1956
rect 1176 -1968 1182 -1962
rect 1176 -1974 1182 -1968
rect 1176 -1980 1182 -1974
rect 1176 -1986 1182 -1980
rect 1176 -1992 1182 -1986
rect 1176 -1998 1182 -1992
rect 1176 -2004 1182 -1998
rect 1176 -2010 1182 -2004
rect 1176 -2016 1182 -2010
rect 1176 -2022 1182 -2016
rect 1176 -2028 1182 -2022
rect 1176 -2034 1182 -2028
rect 1176 -2040 1182 -2034
rect 1176 -2046 1182 -2040
rect 1176 -2052 1182 -2046
rect 1176 -2058 1182 -2052
rect 1176 -2064 1182 -2058
rect 1176 -2070 1182 -2064
rect 1176 -2076 1182 -2070
rect 1176 -2082 1182 -2076
rect 1176 -2088 1182 -2082
rect 1176 -2094 1182 -2088
rect 1176 -2100 1182 -2094
rect 1176 -2106 1182 -2100
rect 1176 -2112 1182 -2106
rect 1176 -2118 1182 -2112
rect 1176 -2124 1182 -2118
rect 1176 -2130 1182 -2124
rect 1176 -2136 1182 -2130
rect 1176 -2142 1182 -2136
rect 1176 -2148 1182 -2142
rect 1176 -2154 1182 -2148
rect 1176 -2160 1182 -2154
rect 1176 -2166 1182 -2160
rect 1176 -2172 1182 -2166
rect 1176 -2178 1182 -2172
rect 1176 -2184 1182 -2178
rect 1176 -2190 1182 -2184
rect 1176 -2196 1182 -2190
rect 1176 -2202 1182 -2196
rect 1176 -2208 1182 -2202
rect 1176 -2214 1182 -2208
rect 1176 -2220 1182 -2214
rect 1176 -2226 1182 -2220
rect 1176 -2232 1182 -2226
rect 1176 -2238 1182 -2232
rect 1176 -2244 1182 -2238
rect 1176 -2250 1182 -2244
rect 1176 -2256 1182 -2250
rect 1176 -2262 1182 -2256
rect 1176 -2268 1182 -2262
rect 1176 -2274 1182 -2268
rect 1176 -2280 1182 -2274
rect 1176 -2286 1182 -2280
rect 1176 -2292 1182 -2286
rect 1176 -2298 1182 -2292
rect 1176 -2304 1182 -2298
rect 1176 -2310 1182 -2304
rect 1176 -2316 1182 -2310
rect 1176 -2322 1182 -2316
rect 1176 -2328 1182 -2322
rect 1176 -2334 1182 -2328
rect 1176 -2340 1182 -2334
rect 1176 -2346 1182 -2340
rect 1176 -2352 1182 -2346
rect 1176 -2358 1182 -2352
rect 1176 -2364 1182 -2358
rect 1176 -2370 1182 -2364
rect 1176 -2376 1182 -2370
rect 1176 -2382 1182 -2376
rect 1176 -2388 1182 -2382
rect 1176 -2394 1182 -2388
rect 1176 -2400 1182 -2394
rect 1176 -2406 1182 -2400
rect 1176 -2412 1182 -2406
rect 1176 -2418 1182 -2412
rect 1176 -2424 1182 -2418
rect 1176 -2430 1182 -2424
rect 1176 -2436 1182 -2430
rect 1176 -2442 1182 -2436
rect 1176 -2448 1182 -2442
rect 1176 -2454 1182 -2448
rect 1176 -2460 1182 -2454
rect 1176 -2466 1182 -2460
rect 1176 -2472 1182 -2466
rect 1176 -2478 1182 -2472
rect 1176 -2484 1182 -2478
rect 1176 -2490 1182 -2484
rect 1176 -2496 1182 -2490
rect 1176 -2502 1182 -2496
rect 1176 -2508 1182 -2502
rect 1176 -2514 1182 -2508
rect 1176 -2520 1182 -2514
rect 1176 -2526 1182 -2520
rect 1176 -2532 1182 -2526
rect 1176 -2538 1182 -2532
rect 1176 -2544 1182 -2538
rect 1176 -2550 1182 -2544
rect 1176 -2556 1182 -2550
rect 1176 -2562 1182 -2556
rect 1176 -2568 1182 -2562
rect 1176 -2574 1182 -2568
rect 1176 -2580 1182 -2574
rect 1176 -2586 1182 -2580
rect 1176 -2592 1182 -2586
rect 1176 -2598 1182 -2592
rect 1176 -2604 1182 -2598
rect 1176 -2610 1182 -2604
rect 1176 -2616 1182 -2610
rect 1176 -2622 1182 -2616
rect 1176 -2628 1182 -2622
rect 1176 -2634 1182 -2628
rect 1176 -2640 1182 -2634
rect 1176 -2736 1182 -2730
rect 1176 -2742 1182 -2736
rect 1176 -2748 1182 -2742
rect 1176 -2754 1182 -2748
rect 1176 -2760 1182 -2754
rect 1176 -2766 1182 -2760
rect 1176 -2772 1182 -2766
rect 1176 -2778 1182 -2772
rect 1176 -2784 1182 -2778
rect 1176 -2790 1182 -2784
rect 1176 -2796 1182 -2790
rect 1176 -2802 1182 -2796
rect 1176 -2808 1182 -2802
rect 1176 -2814 1182 -2808
rect 1176 -2820 1182 -2814
rect 1176 -2826 1182 -2820
rect 1176 -2832 1182 -2826
rect 1176 -2838 1182 -2832
rect 1176 -2844 1182 -2838
rect 1176 -2850 1182 -2844
rect 1176 -2856 1182 -2850
rect 1176 -2862 1182 -2856
rect 1176 -2868 1182 -2862
rect 1176 -2874 1182 -2868
rect 1176 -2880 1182 -2874
rect 1176 -2886 1182 -2880
rect 1176 -2892 1182 -2886
rect 1176 -2898 1182 -2892
rect 1176 -2904 1182 -2898
rect 1176 -2910 1182 -2904
rect 1176 -2916 1182 -2910
rect 1176 -2922 1182 -2916
rect 1176 -2928 1182 -2922
rect 1176 -2934 1182 -2928
rect 1176 -2940 1182 -2934
rect 1176 -2946 1182 -2940
rect 1176 -2952 1182 -2946
rect 1176 -2958 1182 -2952
rect 1176 -2964 1182 -2958
rect 1176 -2970 1182 -2964
rect 1176 -2976 1182 -2970
rect 1176 -2982 1182 -2976
rect 1176 -2988 1182 -2982
rect 1176 -2994 1182 -2988
rect 1176 -3000 1182 -2994
rect 1176 -3006 1182 -3000
rect 1176 -3012 1182 -3006
rect 1176 -3018 1182 -3012
rect 1176 -3024 1182 -3018
rect 1176 -3030 1182 -3024
rect 1176 -3036 1182 -3030
rect 1176 -3114 1182 -3108
rect 1176 -3120 1182 -3114
rect 1176 -3126 1182 -3120
rect 1176 -3132 1182 -3126
rect 1176 -3138 1182 -3132
rect 1176 -3144 1182 -3138
rect 1176 -3150 1182 -3144
rect 1176 -3156 1182 -3150
rect 1176 -3162 1182 -3156
rect 1176 -3168 1182 -3162
rect 1176 -3174 1182 -3168
rect 1176 -3180 1182 -3174
rect 1176 -3186 1182 -3180
rect 1176 -3192 1182 -3186
rect 1176 -3198 1182 -3192
rect 1176 -3204 1182 -3198
rect 1176 -3210 1182 -3204
rect 1176 -3216 1182 -3210
rect 1176 -3222 1182 -3216
rect 1176 -3228 1182 -3222
rect 1176 -3234 1182 -3228
rect 1176 -3240 1182 -3234
rect 1176 -3246 1182 -3240
rect 1176 -3324 1182 -3318
rect 1176 -3330 1182 -3324
rect 1176 -3336 1182 -3330
rect 1176 -3342 1182 -3336
rect 1176 -3348 1182 -3342
rect 1176 -3354 1182 -3348
rect 1176 -3360 1182 -3354
rect 1176 -3366 1182 -3360
rect 1176 -3372 1182 -3366
rect 1176 -3378 1182 -3372
rect 1176 -3384 1182 -3378
rect 1176 -3390 1182 -3384
rect 1176 -3396 1182 -3390
rect 1176 -3402 1182 -3396
rect 1176 -3408 1182 -3402
rect 1176 -3414 1182 -3408
rect 1176 -3420 1182 -3414
rect 1176 -3426 1182 -3420
rect 1176 -3432 1182 -3426
rect 1176 -3438 1182 -3432
rect 1176 -3444 1182 -3438
rect 1176 -3450 1182 -3444
rect 1176 -3456 1182 -3450
rect 1176 -3462 1182 -3456
rect 1176 -3468 1182 -3462
rect 1176 -3474 1182 -3468
rect 1176 -3480 1182 -3474
rect 1176 -3486 1182 -3480
rect 1176 -3492 1182 -3486
rect 1176 -3498 1182 -3492
rect 1176 -3504 1182 -3498
rect 1176 -3510 1182 -3504
rect 1176 -3516 1182 -3510
rect 1182 -1104 1188 -1098
rect 1182 -1110 1188 -1104
rect 1182 -1116 1188 -1110
rect 1182 -1122 1188 -1116
rect 1182 -1128 1188 -1122
rect 1182 -1134 1188 -1128
rect 1182 -1140 1188 -1134
rect 1182 -1146 1188 -1140
rect 1182 -1152 1188 -1146
rect 1182 -1158 1188 -1152
rect 1182 -1164 1188 -1158
rect 1182 -1170 1188 -1164
rect 1182 -1176 1188 -1170
rect 1182 -1182 1188 -1176
rect 1182 -1188 1188 -1182
rect 1182 -1194 1188 -1188
rect 1182 -1200 1188 -1194
rect 1182 -1206 1188 -1200
rect 1182 -1212 1188 -1206
rect 1182 -1218 1188 -1212
rect 1182 -1224 1188 -1218
rect 1182 -1230 1188 -1224
rect 1182 -1236 1188 -1230
rect 1182 -1242 1188 -1236
rect 1182 -1248 1188 -1242
rect 1182 -1254 1188 -1248
rect 1182 -1260 1188 -1254
rect 1182 -1266 1188 -1260
rect 1182 -1272 1188 -1266
rect 1182 -1278 1188 -1272
rect 1182 -1284 1188 -1278
rect 1182 -1290 1188 -1284
rect 1182 -1296 1188 -1290
rect 1182 -1302 1188 -1296
rect 1182 -1308 1188 -1302
rect 1182 -1860 1188 -1854
rect 1182 -1866 1188 -1860
rect 1182 -1872 1188 -1866
rect 1182 -1878 1188 -1872
rect 1182 -1884 1188 -1878
rect 1182 -1890 1188 -1884
rect 1182 -1896 1188 -1890
rect 1182 -1902 1188 -1896
rect 1182 -1908 1188 -1902
rect 1182 -1914 1188 -1908
rect 1182 -1920 1188 -1914
rect 1182 -1926 1188 -1920
rect 1182 -1932 1188 -1926
rect 1182 -1938 1188 -1932
rect 1182 -1944 1188 -1938
rect 1182 -1950 1188 -1944
rect 1182 -1956 1188 -1950
rect 1182 -1962 1188 -1956
rect 1182 -1968 1188 -1962
rect 1182 -1974 1188 -1968
rect 1182 -1980 1188 -1974
rect 1182 -1986 1188 -1980
rect 1182 -1992 1188 -1986
rect 1182 -1998 1188 -1992
rect 1182 -2004 1188 -1998
rect 1182 -2010 1188 -2004
rect 1182 -2016 1188 -2010
rect 1182 -2022 1188 -2016
rect 1182 -2028 1188 -2022
rect 1182 -2034 1188 -2028
rect 1182 -2040 1188 -2034
rect 1182 -2046 1188 -2040
rect 1182 -2052 1188 -2046
rect 1182 -2058 1188 -2052
rect 1182 -2064 1188 -2058
rect 1182 -2070 1188 -2064
rect 1182 -2076 1188 -2070
rect 1182 -2082 1188 -2076
rect 1182 -2088 1188 -2082
rect 1182 -2094 1188 -2088
rect 1182 -2100 1188 -2094
rect 1182 -2106 1188 -2100
rect 1182 -2112 1188 -2106
rect 1182 -2118 1188 -2112
rect 1182 -2124 1188 -2118
rect 1182 -2130 1188 -2124
rect 1182 -2136 1188 -2130
rect 1182 -2142 1188 -2136
rect 1182 -2148 1188 -2142
rect 1182 -2154 1188 -2148
rect 1182 -2160 1188 -2154
rect 1182 -2166 1188 -2160
rect 1182 -2172 1188 -2166
rect 1182 -2178 1188 -2172
rect 1182 -2184 1188 -2178
rect 1182 -2190 1188 -2184
rect 1182 -2196 1188 -2190
rect 1182 -2202 1188 -2196
rect 1182 -2208 1188 -2202
rect 1182 -2214 1188 -2208
rect 1182 -2220 1188 -2214
rect 1182 -2226 1188 -2220
rect 1182 -2232 1188 -2226
rect 1182 -2238 1188 -2232
rect 1182 -2244 1188 -2238
rect 1182 -2250 1188 -2244
rect 1182 -2256 1188 -2250
rect 1182 -2262 1188 -2256
rect 1182 -2268 1188 -2262
rect 1182 -2274 1188 -2268
rect 1182 -2280 1188 -2274
rect 1182 -2286 1188 -2280
rect 1182 -2292 1188 -2286
rect 1182 -2298 1188 -2292
rect 1182 -2304 1188 -2298
rect 1182 -2310 1188 -2304
rect 1182 -2316 1188 -2310
rect 1182 -2322 1188 -2316
rect 1182 -2328 1188 -2322
rect 1182 -2334 1188 -2328
rect 1182 -2340 1188 -2334
rect 1182 -2346 1188 -2340
rect 1182 -2352 1188 -2346
rect 1182 -2358 1188 -2352
rect 1182 -2364 1188 -2358
rect 1182 -2370 1188 -2364
rect 1182 -2376 1188 -2370
rect 1182 -2382 1188 -2376
rect 1182 -2388 1188 -2382
rect 1182 -2394 1188 -2388
rect 1182 -2400 1188 -2394
rect 1182 -2406 1188 -2400
rect 1182 -2412 1188 -2406
rect 1182 -2418 1188 -2412
rect 1182 -2424 1188 -2418
rect 1182 -2430 1188 -2424
rect 1182 -2436 1188 -2430
rect 1182 -2442 1188 -2436
rect 1182 -2448 1188 -2442
rect 1182 -2454 1188 -2448
rect 1182 -2460 1188 -2454
rect 1182 -2466 1188 -2460
rect 1182 -2472 1188 -2466
rect 1182 -2478 1188 -2472
rect 1182 -2484 1188 -2478
rect 1182 -2490 1188 -2484
rect 1182 -2496 1188 -2490
rect 1182 -2502 1188 -2496
rect 1182 -2508 1188 -2502
rect 1182 -2514 1188 -2508
rect 1182 -2520 1188 -2514
rect 1182 -2526 1188 -2520
rect 1182 -2532 1188 -2526
rect 1182 -2538 1188 -2532
rect 1182 -2544 1188 -2538
rect 1182 -2550 1188 -2544
rect 1182 -2556 1188 -2550
rect 1182 -2562 1188 -2556
rect 1182 -2568 1188 -2562
rect 1182 -2574 1188 -2568
rect 1182 -2580 1188 -2574
rect 1182 -2586 1188 -2580
rect 1182 -2592 1188 -2586
rect 1182 -2598 1188 -2592
rect 1182 -2604 1188 -2598
rect 1182 -2610 1188 -2604
rect 1182 -2616 1188 -2610
rect 1182 -2622 1188 -2616
rect 1182 -2628 1188 -2622
rect 1182 -2634 1188 -2628
rect 1182 -2724 1188 -2718
rect 1182 -2730 1188 -2724
rect 1182 -2736 1188 -2730
rect 1182 -2742 1188 -2736
rect 1182 -2748 1188 -2742
rect 1182 -2754 1188 -2748
rect 1182 -2760 1188 -2754
rect 1182 -2766 1188 -2760
rect 1182 -2772 1188 -2766
rect 1182 -2778 1188 -2772
rect 1182 -2784 1188 -2778
rect 1182 -2790 1188 -2784
rect 1182 -2796 1188 -2790
rect 1182 -2802 1188 -2796
rect 1182 -2808 1188 -2802
rect 1182 -2814 1188 -2808
rect 1182 -2820 1188 -2814
rect 1182 -2826 1188 -2820
rect 1182 -2832 1188 -2826
rect 1182 -2838 1188 -2832
rect 1182 -2844 1188 -2838
rect 1182 -2850 1188 -2844
rect 1182 -2856 1188 -2850
rect 1182 -2862 1188 -2856
rect 1182 -2868 1188 -2862
rect 1182 -2874 1188 -2868
rect 1182 -2880 1188 -2874
rect 1182 -2886 1188 -2880
rect 1182 -2892 1188 -2886
rect 1182 -2898 1188 -2892
rect 1182 -2904 1188 -2898
rect 1182 -2910 1188 -2904
rect 1182 -2916 1188 -2910
rect 1182 -2922 1188 -2916
rect 1182 -2928 1188 -2922
rect 1182 -2934 1188 -2928
rect 1182 -2940 1188 -2934
rect 1182 -2946 1188 -2940
rect 1182 -2952 1188 -2946
rect 1182 -2958 1188 -2952
rect 1182 -2964 1188 -2958
rect 1182 -2970 1188 -2964
rect 1182 -2976 1188 -2970
rect 1182 -2982 1188 -2976
rect 1182 -2988 1188 -2982
rect 1182 -2994 1188 -2988
rect 1182 -3000 1188 -2994
rect 1182 -3006 1188 -3000
rect 1182 -3012 1188 -3006
rect 1182 -3018 1188 -3012
rect 1182 -3024 1188 -3018
rect 1182 -3030 1188 -3024
rect 1182 -3036 1188 -3030
rect 1182 -3108 1188 -3102
rect 1182 -3114 1188 -3108
rect 1182 -3120 1188 -3114
rect 1182 -3126 1188 -3120
rect 1182 -3132 1188 -3126
rect 1182 -3138 1188 -3132
rect 1182 -3144 1188 -3138
rect 1182 -3150 1188 -3144
rect 1182 -3156 1188 -3150
rect 1182 -3162 1188 -3156
rect 1182 -3168 1188 -3162
rect 1182 -3174 1188 -3168
rect 1182 -3180 1188 -3174
rect 1182 -3186 1188 -3180
rect 1182 -3192 1188 -3186
rect 1182 -3198 1188 -3192
rect 1182 -3204 1188 -3198
rect 1182 -3210 1188 -3204
rect 1182 -3216 1188 -3210
rect 1182 -3222 1188 -3216
rect 1182 -3228 1188 -3222
rect 1182 -3234 1188 -3228
rect 1182 -3240 1188 -3234
rect 1182 -3246 1188 -3240
rect 1182 -3324 1188 -3318
rect 1182 -3330 1188 -3324
rect 1182 -3336 1188 -3330
rect 1182 -3342 1188 -3336
rect 1182 -3348 1188 -3342
rect 1182 -3354 1188 -3348
rect 1182 -3360 1188 -3354
rect 1182 -3366 1188 -3360
rect 1182 -3372 1188 -3366
rect 1182 -3378 1188 -3372
rect 1182 -3384 1188 -3378
rect 1182 -3390 1188 -3384
rect 1182 -3396 1188 -3390
rect 1182 -3402 1188 -3396
rect 1182 -3408 1188 -3402
rect 1182 -3414 1188 -3408
rect 1182 -3420 1188 -3414
rect 1182 -3426 1188 -3420
rect 1182 -3432 1188 -3426
rect 1182 -3438 1188 -3432
rect 1182 -3444 1188 -3438
rect 1182 -3450 1188 -3444
rect 1182 -3456 1188 -3450
rect 1182 -3462 1188 -3456
rect 1182 -3468 1188 -3462
rect 1182 -3474 1188 -3468
rect 1182 -3480 1188 -3474
rect 1182 -3486 1188 -3480
rect 1182 -3492 1188 -3486
rect 1182 -3498 1188 -3492
rect 1182 -3504 1188 -3498
rect 1182 -3510 1188 -3504
rect 1182 -3516 1188 -3510
rect 1188 -1104 1194 -1098
rect 1188 -1110 1194 -1104
rect 1188 -1116 1194 -1110
rect 1188 -1122 1194 -1116
rect 1188 -1128 1194 -1122
rect 1188 -1134 1194 -1128
rect 1188 -1140 1194 -1134
rect 1188 -1146 1194 -1140
rect 1188 -1152 1194 -1146
rect 1188 -1158 1194 -1152
rect 1188 -1164 1194 -1158
rect 1188 -1170 1194 -1164
rect 1188 -1176 1194 -1170
rect 1188 -1182 1194 -1176
rect 1188 -1188 1194 -1182
rect 1188 -1194 1194 -1188
rect 1188 -1200 1194 -1194
rect 1188 -1206 1194 -1200
rect 1188 -1212 1194 -1206
rect 1188 -1218 1194 -1212
rect 1188 -1224 1194 -1218
rect 1188 -1230 1194 -1224
rect 1188 -1236 1194 -1230
rect 1188 -1242 1194 -1236
rect 1188 -1248 1194 -1242
rect 1188 -1254 1194 -1248
rect 1188 -1260 1194 -1254
rect 1188 -1266 1194 -1260
rect 1188 -1272 1194 -1266
rect 1188 -1278 1194 -1272
rect 1188 -1284 1194 -1278
rect 1188 -1290 1194 -1284
rect 1188 -1296 1194 -1290
rect 1188 -1302 1194 -1296
rect 1188 -1308 1194 -1302
rect 1188 -1842 1194 -1836
rect 1188 -1848 1194 -1842
rect 1188 -1854 1194 -1848
rect 1188 -1860 1194 -1854
rect 1188 -1866 1194 -1860
rect 1188 -1872 1194 -1866
rect 1188 -1878 1194 -1872
rect 1188 -1884 1194 -1878
rect 1188 -1890 1194 -1884
rect 1188 -1896 1194 -1890
rect 1188 -1902 1194 -1896
rect 1188 -1908 1194 -1902
rect 1188 -1914 1194 -1908
rect 1188 -1920 1194 -1914
rect 1188 -1926 1194 -1920
rect 1188 -1932 1194 -1926
rect 1188 -1938 1194 -1932
rect 1188 -1944 1194 -1938
rect 1188 -1950 1194 -1944
rect 1188 -1956 1194 -1950
rect 1188 -1962 1194 -1956
rect 1188 -1968 1194 -1962
rect 1188 -1974 1194 -1968
rect 1188 -1980 1194 -1974
rect 1188 -1986 1194 -1980
rect 1188 -1992 1194 -1986
rect 1188 -1998 1194 -1992
rect 1188 -2004 1194 -1998
rect 1188 -2010 1194 -2004
rect 1188 -2016 1194 -2010
rect 1188 -2022 1194 -2016
rect 1188 -2028 1194 -2022
rect 1188 -2034 1194 -2028
rect 1188 -2040 1194 -2034
rect 1188 -2046 1194 -2040
rect 1188 -2052 1194 -2046
rect 1188 -2058 1194 -2052
rect 1188 -2064 1194 -2058
rect 1188 -2070 1194 -2064
rect 1188 -2076 1194 -2070
rect 1188 -2082 1194 -2076
rect 1188 -2088 1194 -2082
rect 1188 -2094 1194 -2088
rect 1188 -2100 1194 -2094
rect 1188 -2106 1194 -2100
rect 1188 -2112 1194 -2106
rect 1188 -2118 1194 -2112
rect 1188 -2124 1194 -2118
rect 1188 -2130 1194 -2124
rect 1188 -2136 1194 -2130
rect 1188 -2142 1194 -2136
rect 1188 -2148 1194 -2142
rect 1188 -2154 1194 -2148
rect 1188 -2160 1194 -2154
rect 1188 -2166 1194 -2160
rect 1188 -2172 1194 -2166
rect 1188 -2178 1194 -2172
rect 1188 -2184 1194 -2178
rect 1188 -2190 1194 -2184
rect 1188 -2196 1194 -2190
rect 1188 -2202 1194 -2196
rect 1188 -2208 1194 -2202
rect 1188 -2214 1194 -2208
rect 1188 -2220 1194 -2214
rect 1188 -2226 1194 -2220
rect 1188 -2232 1194 -2226
rect 1188 -2238 1194 -2232
rect 1188 -2244 1194 -2238
rect 1188 -2250 1194 -2244
rect 1188 -2256 1194 -2250
rect 1188 -2262 1194 -2256
rect 1188 -2268 1194 -2262
rect 1188 -2274 1194 -2268
rect 1188 -2280 1194 -2274
rect 1188 -2286 1194 -2280
rect 1188 -2292 1194 -2286
rect 1188 -2298 1194 -2292
rect 1188 -2304 1194 -2298
rect 1188 -2310 1194 -2304
rect 1188 -2316 1194 -2310
rect 1188 -2322 1194 -2316
rect 1188 -2328 1194 -2322
rect 1188 -2334 1194 -2328
rect 1188 -2340 1194 -2334
rect 1188 -2346 1194 -2340
rect 1188 -2352 1194 -2346
rect 1188 -2358 1194 -2352
rect 1188 -2364 1194 -2358
rect 1188 -2370 1194 -2364
rect 1188 -2376 1194 -2370
rect 1188 -2382 1194 -2376
rect 1188 -2388 1194 -2382
rect 1188 -2394 1194 -2388
rect 1188 -2400 1194 -2394
rect 1188 -2406 1194 -2400
rect 1188 -2412 1194 -2406
rect 1188 -2418 1194 -2412
rect 1188 -2424 1194 -2418
rect 1188 -2430 1194 -2424
rect 1188 -2436 1194 -2430
rect 1188 -2442 1194 -2436
rect 1188 -2448 1194 -2442
rect 1188 -2454 1194 -2448
rect 1188 -2460 1194 -2454
rect 1188 -2466 1194 -2460
rect 1188 -2472 1194 -2466
rect 1188 -2478 1194 -2472
rect 1188 -2484 1194 -2478
rect 1188 -2490 1194 -2484
rect 1188 -2496 1194 -2490
rect 1188 -2502 1194 -2496
rect 1188 -2508 1194 -2502
rect 1188 -2514 1194 -2508
rect 1188 -2520 1194 -2514
rect 1188 -2526 1194 -2520
rect 1188 -2532 1194 -2526
rect 1188 -2538 1194 -2532
rect 1188 -2544 1194 -2538
rect 1188 -2550 1194 -2544
rect 1188 -2556 1194 -2550
rect 1188 -2562 1194 -2556
rect 1188 -2568 1194 -2562
rect 1188 -2574 1194 -2568
rect 1188 -2580 1194 -2574
rect 1188 -2586 1194 -2580
rect 1188 -2592 1194 -2586
rect 1188 -2598 1194 -2592
rect 1188 -2604 1194 -2598
rect 1188 -2610 1194 -2604
rect 1188 -2616 1194 -2610
rect 1188 -2622 1194 -2616
rect 1188 -2718 1194 -2712
rect 1188 -2724 1194 -2718
rect 1188 -2730 1194 -2724
rect 1188 -2736 1194 -2730
rect 1188 -2742 1194 -2736
rect 1188 -2748 1194 -2742
rect 1188 -2754 1194 -2748
rect 1188 -2760 1194 -2754
rect 1188 -2766 1194 -2760
rect 1188 -2772 1194 -2766
rect 1188 -2778 1194 -2772
rect 1188 -2784 1194 -2778
rect 1188 -2790 1194 -2784
rect 1188 -2796 1194 -2790
rect 1188 -2802 1194 -2796
rect 1188 -2808 1194 -2802
rect 1188 -2814 1194 -2808
rect 1188 -2820 1194 -2814
rect 1188 -2826 1194 -2820
rect 1188 -2832 1194 -2826
rect 1188 -2838 1194 -2832
rect 1188 -2844 1194 -2838
rect 1188 -2850 1194 -2844
rect 1188 -2856 1194 -2850
rect 1188 -2862 1194 -2856
rect 1188 -2868 1194 -2862
rect 1188 -2874 1194 -2868
rect 1188 -2880 1194 -2874
rect 1188 -2886 1194 -2880
rect 1188 -2892 1194 -2886
rect 1188 -2898 1194 -2892
rect 1188 -2904 1194 -2898
rect 1188 -2910 1194 -2904
rect 1188 -2916 1194 -2910
rect 1188 -2922 1194 -2916
rect 1188 -2928 1194 -2922
rect 1188 -2934 1194 -2928
rect 1188 -2940 1194 -2934
rect 1188 -2946 1194 -2940
rect 1188 -2952 1194 -2946
rect 1188 -2958 1194 -2952
rect 1188 -2964 1194 -2958
rect 1188 -2970 1194 -2964
rect 1188 -2976 1194 -2970
rect 1188 -2982 1194 -2976
rect 1188 -2988 1194 -2982
rect 1188 -2994 1194 -2988
rect 1188 -3000 1194 -2994
rect 1188 -3006 1194 -3000
rect 1188 -3012 1194 -3006
rect 1188 -3018 1194 -3012
rect 1188 -3024 1194 -3018
rect 1188 -3030 1194 -3024
rect 1188 -3108 1194 -3102
rect 1188 -3114 1194 -3108
rect 1188 -3120 1194 -3114
rect 1188 -3126 1194 -3120
rect 1188 -3132 1194 -3126
rect 1188 -3138 1194 -3132
rect 1188 -3144 1194 -3138
rect 1188 -3150 1194 -3144
rect 1188 -3156 1194 -3150
rect 1188 -3162 1194 -3156
rect 1188 -3168 1194 -3162
rect 1188 -3174 1194 -3168
rect 1188 -3180 1194 -3174
rect 1188 -3186 1194 -3180
rect 1188 -3192 1194 -3186
rect 1188 -3198 1194 -3192
rect 1188 -3204 1194 -3198
rect 1188 -3210 1194 -3204
rect 1188 -3216 1194 -3210
rect 1188 -3222 1194 -3216
rect 1188 -3228 1194 -3222
rect 1188 -3234 1194 -3228
rect 1188 -3240 1194 -3234
rect 1188 -3246 1194 -3240
rect 1188 -3324 1194 -3318
rect 1188 -3330 1194 -3324
rect 1188 -3336 1194 -3330
rect 1188 -3342 1194 -3336
rect 1188 -3348 1194 -3342
rect 1188 -3354 1194 -3348
rect 1188 -3360 1194 -3354
rect 1188 -3366 1194 -3360
rect 1188 -3372 1194 -3366
rect 1188 -3378 1194 -3372
rect 1188 -3384 1194 -3378
rect 1188 -3390 1194 -3384
rect 1188 -3396 1194 -3390
rect 1188 -3402 1194 -3396
rect 1188 -3408 1194 -3402
rect 1188 -3414 1194 -3408
rect 1188 -3420 1194 -3414
rect 1188 -3426 1194 -3420
rect 1188 -3432 1194 -3426
rect 1188 -3438 1194 -3432
rect 1188 -3444 1194 -3438
rect 1188 -3450 1194 -3444
rect 1188 -3456 1194 -3450
rect 1188 -3462 1194 -3456
rect 1188 -3468 1194 -3462
rect 1188 -3474 1194 -3468
rect 1188 -3480 1194 -3474
rect 1188 -3486 1194 -3480
rect 1188 -3492 1194 -3486
rect 1188 -3498 1194 -3492
rect 1188 -3504 1194 -3498
rect 1188 -3510 1194 -3504
rect 1188 -3516 1194 -3510
rect 1194 -1104 1200 -1098
rect 1194 -1110 1200 -1104
rect 1194 -1116 1200 -1110
rect 1194 -1122 1200 -1116
rect 1194 -1128 1200 -1122
rect 1194 -1134 1200 -1128
rect 1194 -1140 1200 -1134
rect 1194 -1146 1200 -1140
rect 1194 -1152 1200 -1146
rect 1194 -1158 1200 -1152
rect 1194 -1164 1200 -1158
rect 1194 -1170 1200 -1164
rect 1194 -1176 1200 -1170
rect 1194 -1182 1200 -1176
rect 1194 -1188 1200 -1182
rect 1194 -1194 1200 -1188
rect 1194 -1200 1200 -1194
rect 1194 -1206 1200 -1200
rect 1194 -1212 1200 -1206
rect 1194 -1218 1200 -1212
rect 1194 -1224 1200 -1218
rect 1194 -1230 1200 -1224
rect 1194 -1236 1200 -1230
rect 1194 -1242 1200 -1236
rect 1194 -1248 1200 -1242
rect 1194 -1254 1200 -1248
rect 1194 -1260 1200 -1254
rect 1194 -1266 1200 -1260
rect 1194 -1272 1200 -1266
rect 1194 -1278 1200 -1272
rect 1194 -1284 1200 -1278
rect 1194 -1290 1200 -1284
rect 1194 -1296 1200 -1290
rect 1194 -1302 1200 -1296
rect 1194 -1308 1200 -1302
rect 1194 -1824 1200 -1818
rect 1194 -1830 1200 -1824
rect 1194 -1836 1200 -1830
rect 1194 -1842 1200 -1836
rect 1194 -1848 1200 -1842
rect 1194 -1854 1200 -1848
rect 1194 -1860 1200 -1854
rect 1194 -1866 1200 -1860
rect 1194 -1872 1200 -1866
rect 1194 -1878 1200 -1872
rect 1194 -1884 1200 -1878
rect 1194 -1890 1200 -1884
rect 1194 -1896 1200 -1890
rect 1194 -1902 1200 -1896
rect 1194 -1908 1200 -1902
rect 1194 -1914 1200 -1908
rect 1194 -1920 1200 -1914
rect 1194 -1926 1200 -1920
rect 1194 -1932 1200 -1926
rect 1194 -1938 1200 -1932
rect 1194 -1944 1200 -1938
rect 1194 -1950 1200 -1944
rect 1194 -1956 1200 -1950
rect 1194 -1962 1200 -1956
rect 1194 -1968 1200 -1962
rect 1194 -1974 1200 -1968
rect 1194 -1980 1200 -1974
rect 1194 -1986 1200 -1980
rect 1194 -1992 1200 -1986
rect 1194 -1998 1200 -1992
rect 1194 -2004 1200 -1998
rect 1194 -2010 1200 -2004
rect 1194 -2016 1200 -2010
rect 1194 -2022 1200 -2016
rect 1194 -2028 1200 -2022
rect 1194 -2034 1200 -2028
rect 1194 -2040 1200 -2034
rect 1194 -2046 1200 -2040
rect 1194 -2052 1200 -2046
rect 1194 -2058 1200 -2052
rect 1194 -2064 1200 -2058
rect 1194 -2070 1200 -2064
rect 1194 -2076 1200 -2070
rect 1194 -2082 1200 -2076
rect 1194 -2088 1200 -2082
rect 1194 -2094 1200 -2088
rect 1194 -2100 1200 -2094
rect 1194 -2106 1200 -2100
rect 1194 -2112 1200 -2106
rect 1194 -2118 1200 -2112
rect 1194 -2124 1200 -2118
rect 1194 -2130 1200 -2124
rect 1194 -2136 1200 -2130
rect 1194 -2142 1200 -2136
rect 1194 -2148 1200 -2142
rect 1194 -2154 1200 -2148
rect 1194 -2160 1200 -2154
rect 1194 -2166 1200 -2160
rect 1194 -2172 1200 -2166
rect 1194 -2178 1200 -2172
rect 1194 -2184 1200 -2178
rect 1194 -2190 1200 -2184
rect 1194 -2196 1200 -2190
rect 1194 -2202 1200 -2196
rect 1194 -2208 1200 -2202
rect 1194 -2214 1200 -2208
rect 1194 -2220 1200 -2214
rect 1194 -2226 1200 -2220
rect 1194 -2232 1200 -2226
rect 1194 -2238 1200 -2232
rect 1194 -2244 1200 -2238
rect 1194 -2250 1200 -2244
rect 1194 -2256 1200 -2250
rect 1194 -2262 1200 -2256
rect 1194 -2268 1200 -2262
rect 1194 -2274 1200 -2268
rect 1194 -2280 1200 -2274
rect 1194 -2286 1200 -2280
rect 1194 -2292 1200 -2286
rect 1194 -2298 1200 -2292
rect 1194 -2304 1200 -2298
rect 1194 -2310 1200 -2304
rect 1194 -2316 1200 -2310
rect 1194 -2322 1200 -2316
rect 1194 -2328 1200 -2322
rect 1194 -2334 1200 -2328
rect 1194 -2340 1200 -2334
rect 1194 -2346 1200 -2340
rect 1194 -2352 1200 -2346
rect 1194 -2358 1200 -2352
rect 1194 -2364 1200 -2358
rect 1194 -2370 1200 -2364
rect 1194 -2376 1200 -2370
rect 1194 -2382 1200 -2376
rect 1194 -2388 1200 -2382
rect 1194 -2394 1200 -2388
rect 1194 -2400 1200 -2394
rect 1194 -2406 1200 -2400
rect 1194 -2412 1200 -2406
rect 1194 -2418 1200 -2412
rect 1194 -2424 1200 -2418
rect 1194 -2430 1200 -2424
rect 1194 -2436 1200 -2430
rect 1194 -2442 1200 -2436
rect 1194 -2448 1200 -2442
rect 1194 -2454 1200 -2448
rect 1194 -2460 1200 -2454
rect 1194 -2466 1200 -2460
rect 1194 -2472 1200 -2466
rect 1194 -2478 1200 -2472
rect 1194 -2484 1200 -2478
rect 1194 -2490 1200 -2484
rect 1194 -2496 1200 -2490
rect 1194 -2502 1200 -2496
rect 1194 -2508 1200 -2502
rect 1194 -2514 1200 -2508
rect 1194 -2520 1200 -2514
rect 1194 -2526 1200 -2520
rect 1194 -2532 1200 -2526
rect 1194 -2538 1200 -2532
rect 1194 -2544 1200 -2538
rect 1194 -2550 1200 -2544
rect 1194 -2556 1200 -2550
rect 1194 -2562 1200 -2556
rect 1194 -2568 1200 -2562
rect 1194 -2574 1200 -2568
rect 1194 -2580 1200 -2574
rect 1194 -2586 1200 -2580
rect 1194 -2592 1200 -2586
rect 1194 -2598 1200 -2592
rect 1194 -2604 1200 -2598
rect 1194 -2610 1200 -2604
rect 1194 -2616 1200 -2610
rect 1194 -2706 1200 -2700
rect 1194 -2712 1200 -2706
rect 1194 -2718 1200 -2712
rect 1194 -2724 1200 -2718
rect 1194 -2730 1200 -2724
rect 1194 -2736 1200 -2730
rect 1194 -2742 1200 -2736
rect 1194 -2748 1200 -2742
rect 1194 -2754 1200 -2748
rect 1194 -2760 1200 -2754
rect 1194 -2766 1200 -2760
rect 1194 -2772 1200 -2766
rect 1194 -2778 1200 -2772
rect 1194 -2784 1200 -2778
rect 1194 -2790 1200 -2784
rect 1194 -2796 1200 -2790
rect 1194 -2802 1200 -2796
rect 1194 -2808 1200 -2802
rect 1194 -2814 1200 -2808
rect 1194 -2820 1200 -2814
rect 1194 -2826 1200 -2820
rect 1194 -2832 1200 -2826
rect 1194 -2838 1200 -2832
rect 1194 -2844 1200 -2838
rect 1194 -2850 1200 -2844
rect 1194 -2856 1200 -2850
rect 1194 -2862 1200 -2856
rect 1194 -2868 1200 -2862
rect 1194 -2874 1200 -2868
rect 1194 -2880 1200 -2874
rect 1194 -2886 1200 -2880
rect 1194 -2892 1200 -2886
rect 1194 -2898 1200 -2892
rect 1194 -2904 1200 -2898
rect 1194 -2910 1200 -2904
rect 1194 -2916 1200 -2910
rect 1194 -2922 1200 -2916
rect 1194 -2928 1200 -2922
rect 1194 -2934 1200 -2928
rect 1194 -2940 1200 -2934
rect 1194 -2946 1200 -2940
rect 1194 -2952 1200 -2946
rect 1194 -2958 1200 -2952
rect 1194 -2964 1200 -2958
rect 1194 -2970 1200 -2964
rect 1194 -2976 1200 -2970
rect 1194 -2982 1200 -2976
rect 1194 -2988 1200 -2982
rect 1194 -2994 1200 -2988
rect 1194 -3000 1200 -2994
rect 1194 -3006 1200 -3000
rect 1194 -3012 1200 -3006
rect 1194 -3018 1200 -3012
rect 1194 -3024 1200 -3018
rect 1194 -3102 1200 -3096
rect 1194 -3108 1200 -3102
rect 1194 -3114 1200 -3108
rect 1194 -3120 1200 -3114
rect 1194 -3126 1200 -3120
rect 1194 -3132 1200 -3126
rect 1194 -3138 1200 -3132
rect 1194 -3144 1200 -3138
rect 1194 -3150 1200 -3144
rect 1194 -3156 1200 -3150
rect 1194 -3162 1200 -3156
rect 1194 -3168 1200 -3162
rect 1194 -3174 1200 -3168
rect 1194 -3180 1200 -3174
rect 1194 -3186 1200 -3180
rect 1194 -3192 1200 -3186
rect 1194 -3198 1200 -3192
rect 1194 -3204 1200 -3198
rect 1194 -3210 1200 -3204
rect 1194 -3216 1200 -3210
rect 1194 -3222 1200 -3216
rect 1194 -3228 1200 -3222
rect 1194 -3234 1200 -3228
rect 1194 -3240 1200 -3234
rect 1194 -3246 1200 -3240
rect 1194 -3324 1200 -3318
rect 1194 -3330 1200 -3324
rect 1194 -3336 1200 -3330
rect 1194 -3342 1200 -3336
rect 1194 -3348 1200 -3342
rect 1194 -3354 1200 -3348
rect 1194 -3360 1200 -3354
rect 1194 -3366 1200 -3360
rect 1194 -3372 1200 -3366
rect 1194 -3378 1200 -3372
rect 1194 -3384 1200 -3378
rect 1194 -3390 1200 -3384
rect 1194 -3396 1200 -3390
rect 1194 -3402 1200 -3396
rect 1194 -3408 1200 -3402
rect 1194 -3414 1200 -3408
rect 1194 -3420 1200 -3414
rect 1194 -3426 1200 -3420
rect 1194 -3432 1200 -3426
rect 1194 -3438 1200 -3432
rect 1194 -3444 1200 -3438
rect 1194 -3450 1200 -3444
rect 1194 -3456 1200 -3450
rect 1194 -3462 1200 -3456
rect 1194 -3468 1200 -3462
rect 1194 -3474 1200 -3468
rect 1194 -3480 1200 -3474
rect 1194 -3486 1200 -3480
rect 1194 -3492 1200 -3486
rect 1194 -3498 1200 -3492
rect 1194 -3504 1200 -3498
rect 1194 -3510 1200 -3504
rect 1194 -3516 1200 -3510
rect 1200 -1104 1206 -1098
rect 1200 -1110 1206 -1104
rect 1200 -1116 1206 -1110
rect 1200 -1122 1206 -1116
rect 1200 -1128 1206 -1122
rect 1200 -1134 1206 -1128
rect 1200 -1140 1206 -1134
rect 1200 -1146 1206 -1140
rect 1200 -1152 1206 -1146
rect 1200 -1158 1206 -1152
rect 1200 -1164 1206 -1158
rect 1200 -1170 1206 -1164
rect 1200 -1176 1206 -1170
rect 1200 -1182 1206 -1176
rect 1200 -1188 1206 -1182
rect 1200 -1194 1206 -1188
rect 1200 -1200 1206 -1194
rect 1200 -1206 1206 -1200
rect 1200 -1212 1206 -1206
rect 1200 -1218 1206 -1212
rect 1200 -1224 1206 -1218
rect 1200 -1230 1206 -1224
rect 1200 -1236 1206 -1230
rect 1200 -1242 1206 -1236
rect 1200 -1248 1206 -1242
rect 1200 -1254 1206 -1248
rect 1200 -1260 1206 -1254
rect 1200 -1266 1206 -1260
rect 1200 -1272 1206 -1266
rect 1200 -1278 1206 -1272
rect 1200 -1284 1206 -1278
rect 1200 -1290 1206 -1284
rect 1200 -1296 1206 -1290
rect 1200 -1302 1206 -1296
rect 1200 -1308 1206 -1302
rect 1200 -1812 1206 -1806
rect 1200 -1818 1206 -1812
rect 1200 -1824 1206 -1818
rect 1200 -1830 1206 -1824
rect 1200 -1836 1206 -1830
rect 1200 -1842 1206 -1836
rect 1200 -1848 1206 -1842
rect 1200 -1854 1206 -1848
rect 1200 -1860 1206 -1854
rect 1200 -1866 1206 -1860
rect 1200 -1872 1206 -1866
rect 1200 -1878 1206 -1872
rect 1200 -1884 1206 -1878
rect 1200 -1890 1206 -1884
rect 1200 -1896 1206 -1890
rect 1200 -1902 1206 -1896
rect 1200 -1908 1206 -1902
rect 1200 -1914 1206 -1908
rect 1200 -1920 1206 -1914
rect 1200 -1926 1206 -1920
rect 1200 -1932 1206 -1926
rect 1200 -1938 1206 -1932
rect 1200 -1944 1206 -1938
rect 1200 -1950 1206 -1944
rect 1200 -1956 1206 -1950
rect 1200 -1962 1206 -1956
rect 1200 -1968 1206 -1962
rect 1200 -1974 1206 -1968
rect 1200 -1980 1206 -1974
rect 1200 -1986 1206 -1980
rect 1200 -1992 1206 -1986
rect 1200 -1998 1206 -1992
rect 1200 -2004 1206 -1998
rect 1200 -2010 1206 -2004
rect 1200 -2016 1206 -2010
rect 1200 -2022 1206 -2016
rect 1200 -2028 1206 -2022
rect 1200 -2034 1206 -2028
rect 1200 -2040 1206 -2034
rect 1200 -2046 1206 -2040
rect 1200 -2052 1206 -2046
rect 1200 -2058 1206 -2052
rect 1200 -2064 1206 -2058
rect 1200 -2070 1206 -2064
rect 1200 -2076 1206 -2070
rect 1200 -2082 1206 -2076
rect 1200 -2088 1206 -2082
rect 1200 -2094 1206 -2088
rect 1200 -2100 1206 -2094
rect 1200 -2106 1206 -2100
rect 1200 -2112 1206 -2106
rect 1200 -2118 1206 -2112
rect 1200 -2124 1206 -2118
rect 1200 -2130 1206 -2124
rect 1200 -2136 1206 -2130
rect 1200 -2142 1206 -2136
rect 1200 -2148 1206 -2142
rect 1200 -2154 1206 -2148
rect 1200 -2160 1206 -2154
rect 1200 -2166 1206 -2160
rect 1200 -2172 1206 -2166
rect 1200 -2178 1206 -2172
rect 1200 -2184 1206 -2178
rect 1200 -2190 1206 -2184
rect 1200 -2196 1206 -2190
rect 1200 -2202 1206 -2196
rect 1200 -2208 1206 -2202
rect 1200 -2214 1206 -2208
rect 1200 -2220 1206 -2214
rect 1200 -2226 1206 -2220
rect 1200 -2232 1206 -2226
rect 1200 -2238 1206 -2232
rect 1200 -2244 1206 -2238
rect 1200 -2250 1206 -2244
rect 1200 -2256 1206 -2250
rect 1200 -2262 1206 -2256
rect 1200 -2268 1206 -2262
rect 1200 -2274 1206 -2268
rect 1200 -2280 1206 -2274
rect 1200 -2286 1206 -2280
rect 1200 -2292 1206 -2286
rect 1200 -2298 1206 -2292
rect 1200 -2304 1206 -2298
rect 1200 -2310 1206 -2304
rect 1200 -2316 1206 -2310
rect 1200 -2322 1206 -2316
rect 1200 -2328 1206 -2322
rect 1200 -2334 1206 -2328
rect 1200 -2340 1206 -2334
rect 1200 -2346 1206 -2340
rect 1200 -2352 1206 -2346
rect 1200 -2358 1206 -2352
rect 1200 -2364 1206 -2358
rect 1200 -2370 1206 -2364
rect 1200 -2376 1206 -2370
rect 1200 -2382 1206 -2376
rect 1200 -2388 1206 -2382
rect 1200 -2394 1206 -2388
rect 1200 -2400 1206 -2394
rect 1200 -2406 1206 -2400
rect 1200 -2412 1206 -2406
rect 1200 -2418 1206 -2412
rect 1200 -2424 1206 -2418
rect 1200 -2430 1206 -2424
rect 1200 -2436 1206 -2430
rect 1200 -2442 1206 -2436
rect 1200 -2448 1206 -2442
rect 1200 -2454 1206 -2448
rect 1200 -2460 1206 -2454
rect 1200 -2466 1206 -2460
rect 1200 -2472 1206 -2466
rect 1200 -2478 1206 -2472
rect 1200 -2484 1206 -2478
rect 1200 -2490 1206 -2484
rect 1200 -2496 1206 -2490
rect 1200 -2502 1206 -2496
rect 1200 -2508 1206 -2502
rect 1200 -2514 1206 -2508
rect 1200 -2520 1206 -2514
rect 1200 -2526 1206 -2520
rect 1200 -2532 1206 -2526
rect 1200 -2538 1206 -2532
rect 1200 -2544 1206 -2538
rect 1200 -2550 1206 -2544
rect 1200 -2556 1206 -2550
rect 1200 -2562 1206 -2556
rect 1200 -2568 1206 -2562
rect 1200 -2574 1206 -2568
rect 1200 -2580 1206 -2574
rect 1200 -2586 1206 -2580
rect 1200 -2592 1206 -2586
rect 1200 -2598 1206 -2592
rect 1200 -2604 1206 -2598
rect 1200 -2700 1206 -2694
rect 1200 -2706 1206 -2700
rect 1200 -2712 1206 -2706
rect 1200 -2718 1206 -2712
rect 1200 -2724 1206 -2718
rect 1200 -2730 1206 -2724
rect 1200 -2736 1206 -2730
rect 1200 -2742 1206 -2736
rect 1200 -2748 1206 -2742
rect 1200 -2754 1206 -2748
rect 1200 -2760 1206 -2754
rect 1200 -2766 1206 -2760
rect 1200 -2772 1206 -2766
rect 1200 -2778 1206 -2772
rect 1200 -2784 1206 -2778
rect 1200 -2790 1206 -2784
rect 1200 -2796 1206 -2790
rect 1200 -2802 1206 -2796
rect 1200 -2808 1206 -2802
rect 1200 -2814 1206 -2808
rect 1200 -2820 1206 -2814
rect 1200 -2826 1206 -2820
rect 1200 -2832 1206 -2826
rect 1200 -2838 1206 -2832
rect 1200 -2844 1206 -2838
rect 1200 -2850 1206 -2844
rect 1200 -2856 1206 -2850
rect 1200 -2862 1206 -2856
rect 1200 -2868 1206 -2862
rect 1200 -2874 1206 -2868
rect 1200 -2880 1206 -2874
rect 1200 -2886 1206 -2880
rect 1200 -2892 1206 -2886
rect 1200 -2898 1206 -2892
rect 1200 -2904 1206 -2898
rect 1200 -2910 1206 -2904
rect 1200 -2916 1206 -2910
rect 1200 -2922 1206 -2916
rect 1200 -2928 1206 -2922
rect 1200 -2934 1206 -2928
rect 1200 -2940 1206 -2934
rect 1200 -2946 1206 -2940
rect 1200 -2952 1206 -2946
rect 1200 -2958 1206 -2952
rect 1200 -2964 1206 -2958
rect 1200 -2970 1206 -2964
rect 1200 -2976 1206 -2970
rect 1200 -2982 1206 -2976
rect 1200 -2988 1206 -2982
rect 1200 -2994 1206 -2988
rect 1200 -3000 1206 -2994
rect 1200 -3006 1206 -3000
rect 1200 -3012 1206 -3006
rect 1200 -3018 1206 -3012
rect 1200 -3096 1206 -3090
rect 1200 -3102 1206 -3096
rect 1200 -3108 1206 -3102
rect 1200 -3114 1206 -3108
rect 1200 -3120 1206 -3114
rect 1200 -3126 1206 -3120
rect 1200 -3132 1206 -3126
rect 1200 -3138 1206 -3132
rect 1200 -3144 1206 -3138
rect 1200 -3150 1206 -3144
rect 1200 -3156 1206 -3150
rect 1200 -3162 1206 -3156
rect 1200 -3168 1206 -3162
rect 1200 -3174 1206 -3168
rect 1200 -3180 1206 -3174
rect 1200 -3186 1206 -3180
rect 1200 -3192 1206 -3186
rect 1200 -3198 1206 -3192
rect 1200 -3204 1206 -3198
rect 1200 -3210 1206 -3204
rect 1200 -3216 1206 -3210
rect 1200 -3222 1206 -3216
rect 1200 -3228 1206 -3222
rect 1200 -3234 1206 -3228
rect 1200 -3240 1206 -3234
rect 1200 -3324 1206 -3318
rect 1200 -3330 1206 -3324
rect 1200 -3336 1206 -3330
rect 1200 -3342 1206 -3336
rect 1200 -3348 1206 -3342
rect 1200 -3354 1206 -3348
rect 1200 -3360 1206 -3354
rect 1200 -3366 1206 -3360
rect 1200 -3372 1206 -3366
rect 1200 -3378 1206 -3372
rect 1200 -3384 1206 -3378
rect 1200 -3390 1206 -3384
rect 1200 -3396 1206 -3390
rect 1200 -3402 1206 -3396
rect 1200 -3408 1206 -3402
rect 1200 -3414 1206 -3408
rect 1200 -3420 1206 -3414
rect 1200 -3426 1206 -3420
rect 1200 -3432 1206 -3426
rect 1200 -3438 1206 -3432
rect 1200 -3444 1206 -3438
rect 1200 -3450 1206 -3444
rect 1200 -3456 1206 -3450
rect 1200 -3462 1206 -3456
rect 1200 -3468 1206 -3462
rect 1200 -3474 1206 -3468
rect 1200 -3480 1206 -3474
rect 1200 -3486 1206 -3480
rect 1200 -3492 1206 -3486
rect 1200 -3498 1206 -3492
rect 1200 -3504 1206 -3498
rect 1200 -3510 1206 -3504
rect 1200 -3516 1206 -3510
rect 1206 -1104 1212 -1098
rect 1206 -1110 1212 -1104
rect 1206 -1116 1212 -1110
rect 1206 -1122 1212 -1116
rect 1206 -1128 1212 -1122
rect 1206 -1134 1212 -1128
rect 1206 -1140 1212 -1134
rect 1206 -1146 1212 -1140
rect 1206 -1152 1212 -1146
rect 1206 -1158 1212 -1152
rect 1206 -1164 1212 -1158
rect 1206 -1170 1212 -1164
rect 1206 -1176 1212 -1170
rect 1206 -1182 1212 -1176
rect 1206 -1188 1212 -1182
rect 1206 -1194 1212 -1188
rect 1206 -1200 1212 -1194
rect 1206 -1206 1212 -1200
rect 1206 -1212 1212 -1206
rect 1206 -1218 1212 -1212
rect 1206 -1224 1212 -1218
rect 1206 -1230 1212 -1224
rect 1206 -1236 1212 -1230
rect 1206 -1242 1212 -1236
rect 1206 -1248 1212 -1242
rect 1206 -1254 1212 -1248
rect 1206 -1260 1212 -1254
rect 1206 -1266 1212 -1260
rect 1206 -1272 1212 -1266
rect 1206 -1278 1212 -1272
rect 1206 -1284 1212 -1278
rect 1206 -1290 1212 -1284
rect 1206 -1296 1212 -1290
rect 1206 -1302 1212 -1296
rect 1206 -1308 1212 -1302
rect 1206 -1794 1212 -1788
rect 1206 -1800 1212 -1794
rect 1206 -1806 1212 -1800
rect 1206 -1812 1212 -1806
rect 1206 -1818 1212 -1812
rect 1206 -1824 1212 -1818
rect 1206 -1830 1212 -1824
rect 1206 -1836 1212 -1830
rect 1206 -1842 1212 -1836
rect 1206 -1848 1212 -1842
rect 1206 -1854 1212 -1848
rect 1206 -1860 1212 -1854
rect 1206 -1866 1212 -1860
rect 1206 -1872 1212 -1866
rect 1206 -1878 1212 -1872
rect 1206 -1884 1212 -1878
rect 1206 -1890 1212 -1884
rect 1206 -1896 1212 -1890
rect 1206 -1902 1212 -1896
rect 1206 -1908 1212 -1902
rect 1206 -1914 1212 -1908
rect 1206 -1920 1212 -1914
rect 1206 -1926 1212 -1920
rect 1206 -1932 1212 -1926
rect 1206 -1938 1212 -1932
rect 1206 -1944 1212 -1938
rect 1206 -1950 1212 -1944
rect 1206 -1956 1212 -1950
rect 1206 -1962 1212 -1956
rect 1206 -1968 1212 -1962
rect 1206 -1974 1212 -1968
rect 1206 -1980 1212 -1974
rect 1206 -1986 1212 -1980
rect 1206 -1992 1212 -1986
rect 1206 -1998 1212 -1992
rect 1206 -2004 1212 -1998
rect 1206 -2010 1212 -2004
rect 1206 -2016 1212 -2010
rect 1206 -2022 1212 -2016
rect 1206 -2028 1212 -2022
rect 1206 -2034 1212 -2028
rect 1206 -2040 1212 -2034
rect 1206 -2046 1212 -2040
rect 1206 -2052 1212 -2046
rect 1206 -2058 1212 -2052
rect 1206 -2064 1212 -2058
rect 1206 -2070 1212 -2064
rect 1206 -2076 1212 -2070
rect 1206 -2082 1212 -2076
rect 1206 -2088 1212 -2082
rect 1206 -2094 1212 -2088
rect 1206 -2100 1212 -2094
rect 1206 -2106 1212 -2100
rect 1206 -2112 1212 -2106
rect 1206 -2118 1212 -2112
rect 1206 -2124 1212 -2118
rect 1206 -2130 1212 -2124
rect 1206 -2136 1212 -2130
rect 1206 -2142 1212 -2136
rect 1206 -2148 1212 -2142
rect 1206 -2154 1212 -2148
rect 1206 -2160 1212 -2154
rect 1206 -2166 1212 -2160
rect 1206 -2172 1212 -2166
rect 1206 -2178 1212 -2172
rect 1206 -2184 1212 -2178
rect 1206 -2190 1212 -2184
rect 1206 -2196 1212 -2190
rect 1206 -2202 1212 -2196
rect 1206 -2208 1212 -2202
rect 1206 -2214 1212 -2208
rect 1206 -2220 1212 -2214
rect 1206 -2226 1212 -2220
rect 1206 -2232 1212 -2226
rect 1206 -2238 1212 -2232
rect 1206 -2244 1212 -2238
rect 1206 -2250 1212 -2244
rect 1206 -2256 1212 -2250
rect 1206 -2262 1212 -2256
rect 1206 -2268 1212 -2262
rect 1206 -2274 1212 -2268
rect 1206 -2280 1212 -2274
rect 1206 -2286 1212 -2280
rect 1206 -2292 1212 -2286
rect 1206 -2298 1212 -2292
rect 1206 -2304 1212 -2298
rect 1206 -2310 1212 -2304
rect 1206 -2316 1212 -2310
rect 1206 -2322 1212 -2316
rect 1206 -2328 1212 -2322
rect 1206 -2334 1212 -2328
rect 1206 -2340 1212 -2334
rect 1206 -2346 1212 -2340
rect 1206 -2352 1212 -2346
rect 1206 -2358 1212 -2352
rect 1206 -2364 1212 -2358
rect 1206 -2370 1212 -2364
rect 1206 -2376 1212 -2370
rect 1206 -2382 1212 -2376
rect 1206 -2388 1212 -2382
rect 1206 -2394 1212 -2388
rect 1206 -2400 1212 -2394
rect 1206 -2406 1212 -2400
rect 1206 -2412 1212 -2406
rect 1206 -2418 1212 -2412
rect 1206 -2424 1212 -2418
rect 1206 -2430 1212 -2424
rect 1206 -2436 1212 -2430
rect 1206 -2442 1212 -2436
rect 1206 -2448 1212 -2442
rect 1206 -2454 1212 -2448
rect 1206 -2460 1212 -2454
rect 1206 -2466 1212 -2460
rect 1206 -2472 1212 -2466
rect 1206 -2478 1212 -2472
rect 1206 -2484 1212 -2478
rect 1206 -2490 1212 -2484
rect 1206 -2496 1212 -2490
rect 1206 -2502 1212 -2496
rect 1206 -2508 1212 -2502
rect 1206 -2514 1212 -2508
rect 1206 -2520 1212 -2514
rect 1206 -2526 1212 -2520
rect 1206 -2532 1212 -2526
rect 1206 -2538 1212 -2532
rect 1206 -2544 1212 -2538
rect 1206 -2550 1212 -2544
rect 1206 -2556 1212 -2550
rect 1206 -2562 1212 -2556
rect 1206 -2568 1212 -2562
rect 1206 -2574 1212 -2568
rect 1206 -2580 1212 -2574
rect 1206 -2586 1212 -2580
rect 1206 -2592 1212 -2586
rect 1206 -2598 1212 -2592
rect 1206 -2688 1212 -2682
rect 1206 -2694 1212 -2688
rect 1206 -2700 1212 -2694
rect 1206 -2706 1212 -2700
rect 1206 -2712 1212 -2706
rect 1206 -2718 1212 -2712
rect 1206 -2724 1212 -2718
rect 1206 -2730 1212 -2724
rect 1206 -2736 1212 -2730
rect 1206 -2742 1212 -2736
rect 1206 -2748 1212 -2742
rect 1206 -2754 1212 -2748
rect 1206 -2760 1212 -2754
rect 1206 -2766 1212 -2760
rect 1206 -2772 1212 -2766
rect 1206 -2778 1212 -2772
rect 1206 -2784 1212 -2778
rect 1206 -2790 1212 -2784
rect 1206 -2796 1212 -2790
rect 1206 -2802 1212 -2796
rect 1206 -2808 1212 -2802
rect 1206 -2814 1212 -2808
rect 1206 -2820 1212 -2814
rect 1206 -2826 1212 -2820
rect 1206 -2832 1212 -2826
rect 1206 -2838 1212 -2832
rect 1206 -2844 1212 -2838
rect 1206 -2850 1212 -2844
rect 1206 -2856 1212 -2850
rect 1206 -2862 1212 -2856
rect 1206 -2868 1212 -2862
rect 1206 -2874 1212 -2868
rect 1206 -2880 1212 -2874
rect 1206 -2886 1212 -2880
rect 1206 -2892 1212 -2886
rect 1206 -2898 1212 -2892
rect 1206 -2904 1212 -2898
rect 1206 -2910 1212 -2904
rect 1206 -2916 1212 -2910
rect 1206 -2922 1212 -2916
rect 1206 -2928 1212 -2922
rect 1206 -2934 1212 -2928
rect 1206 -2940 1212 -2934
rect 1206 -2946 1212 -2940
rect 1206 -2952 1212 -2946
rect 1206 -2958 1212 -2952
rect 1206 -2964 1212 -2958
rect 1206 -2970 1212 -2964
rect 1206 -2976 1212 -2970
rect 1206 -2982 1212 -2976
rect 1206 -2988 1212 -2982
rect 1206 -2994 1212 -2988
rect 1206 -3000 1212 -2994
rect 1206 -3006 1212 -3000
rect 1206 -3012 1212 -3006
rect 1206 -3090 1212 -3084
rect 1206 -3096 1212 -3090
rect 1206 -3102 1212 -3096
rect 1206 -3108 1212 -3102
rect 1206 -3114 1212 -3108
rect 1206 -3120 1212 -3114
rect 1206 -3126 1212 -3120
rect 1206 -3132 1212 -3126
rect 1206 -3138 1212 -3132
rect 1206 -3144 1212 -3138
rect 1206 -3150 1212 -3144
rect 1206 -3156 1212 -3150
rect 1206 -3162 1212 -3156
rect 1206 -3168 1212 -3162
rect 1206 -3174 1212 -3168
rect 1206 -3180 1212 -3174
rect 1206 -3186 1212 -3180
rect 1206 -3192 1212 -3186
rect 1206 -3198 1212 -3192
rect 1206 -3204 1212 -3198
rect 1206 -3210 1212 -3204
rect 1206 -3216 1212 -3210
rect 1206 -3222 1212 -3216
rect 1206 -3228 1212 -3222
rect 1206 -3234 1212 -3228
rect 1206 -3240 1212 -3234
rect 1206 -3324 1212 -3318
rect 1206 -3330 1212 -3324
rect 1206 -3336 1212 -3330
rect 1206 -3342 1212 -3336
rect 1206 -3348 1212 -3342
rect 1206 -3354 1212 -3348
rect 1206 -3360 1212 -3354
rect 1206 -3366 1212 -3360
rect 1206 -3372 1212 -3366
rect 1206 -3378 1212 -3372
rect 1206 -3384 1212 -3378
rect 1206 -3390 1212 -3384
rect 1206 -3396 1212 -3390
rect 1206 -3402 1212 -3396
rect 1206 -3408 1212 -3402
rect 1206 -3414 1212 -3408
rect 1206 -3420 1212 -3414
rect 1206 -3426 1212 -3420
rect 1206 -3432 1212 -3426
rect 1206 -3438 1212 -3432
rect 1206 -3444 1212 -3438
rect 1206 -3450 1212 -3444
rect 1206 -3456 1212 -3450
rect 1206 -3462 1212 -3456
rect 1206 -3468 1212 -3462
rect 1206 -3474 1212 -3468
rect 1206 -3480 1212 -3474
rect 1206 -3486 1212 -3480
rect 1206 -3492 1212 -3486
rect 1206 -3498 1212 -3492
rect 1206 -3504 1212 -3498
rect 1206 -3510 1212 -3504
rect 1206 -3516 1212 -3510
rect 1212 -1104 1218 -1098
rect 1212 -1110 1218 -1104
rect 1212 -1116 1218 -1110
rect 1212 -1122 1218 -1116
rect 1212 -1128 1218 -1122
rect 1212 -1134 1218 -1128
rect 1212 -1140 1218 -1134
rect 1212 -1146 1218 -1140
rect 1212 -1152 1218 -1146
rect 1212 -1158 1218 -1152
rect 1212 -1164 1218 -1158
rect 1212 -1170 1218 -1164
rect 1212 -1176 1218 -1170
rect 1212 -1182 1218 -1176
rect 1212 -1188 1218 -1182
rect 1212 -1194 1218 -1188
rect 1212 -1200 1218 -1194
rect 1212 -1206 1218 -1200
rect 1212 -1212 1218 -1206
rect 1212 -1218 1218 -1212
rect 1212 -1224 1218 -1218
rect 1212 -1230 1218 -1224
rect 1212 -1236 1218 -1230
rect 1212 -1242 1218 -1236
rect 1212 -1248 1218 -1242
rect 1212 -1254 1218 -1248
rect 1212 -1260 1218 -1254
rect 1212 -1266 1218 -1260
rect 1212 -1272 1218 -1266
rect 1212 -1278 1218 -1272
rect 1212 -1284 1218 -1278
rect 1212 -1290 1218 -1284
rect 1212 -1296 1218 -1290
rect 1212 -1302 1218 -1296
rect 1212 -1308 1218 -1302
rect 1212 -1782 1218 -1776
rect 1212 -1788 1218 -1782
rect 1212 -1794 1218 -1788
rect 1212 -1800 1218 -1794
rect 1212 -1806 1218 -1800
rect 1212 -1812 1218 -1806
rect 1212 -1818 1218 -1812
rect 1212 -1824 1218 -1818
rect 1212 -1830 1218 -1824
rect 1212 -1836 1218 -1830
rect 1212 -1842 1218 -1836
rect 1212 -1848 1218 -1842
rect 1212 -1854 1218 -1848
rect 1212 -1860 1218 -1854
rect 1212 -1866 1218 -1860
rect 1212 -1872 1218 -1866
rect 1212 -1878 1218 -1872
rect 1212 -1884 1218 -1878
rect 1212 -1890 1218 -1884
rect 1212 -1896 1218 -1890
rect 1212 -1902 1218 -1896
rect 1212 -1908 1218 -1902
rect 1212 -1914 1218 -1908
rect 1212 -1920 1218 -1914
rect 1212 -1926 1218 -1920
rect 1212 -1932 1218 -1926
rect 1212 -1938 1218 -1932
rect 1212 -1944 1218 -1938
rect 1212 -1950 1218 -1944
rect 1212 -1956 1218 -1950
rect 1212 -1962 1218 -1956
rect 1212 -1968 1218 -1962
rect 1212 -1974 1218 -1968
rect 1212 -1980 1218 -1974
rect 1212 -1986 1218 -1980
rect 1212 -1992 1218 -1986
rect 1212 -1998 1218 -1992
rect 1212 -2004 1218 -1998
rect 1212 -2010 1218 -2004
rect 1212 -2016 1218 -2010
rect 1212 -2022 1218 -2016
rect 1212 -2028 1218 -2022
rect 1212 -2034 1218 -2028
rect 1212 -2040 1218 -2034
rect 1212 -2046 1218 -2040
rect 1212 -2052 1218 -2046
rect 1212 -2058 1218 -2052
rect 1212 -2064 1218 -2058
rect 1212 -2070 1218 -2064
rect 1212 -2076 1218 -2070
rect 1212 -2082 1218 -2076
rect 1212 -2088 1218 -2082
rect 1212 -2094 1218 -2088
rect 1212 -2100 1218 -2094
rect 1212 -2106 1218 -2100
rect 1212 -2112 1218 -2106
rect 1212 -2118 1218 -2112
rect 1212 -2124 1218 -2118
rect 1212 -2130 1218 -2124
rect 1212 -2136 1218 -2130
rect 1212 -2142 1218 -2136
rect 1212 -2148 1218 -2142
rect 1212 -2154 1218 -2148
rect 1212 -2160 1218 -2154
rect 1212 -2166 1218 -2160
rect 1212 -2172 1218 -2166
rect 1212 -2178 1218 -2172
rect 1212 -2184 1218 -2178
rect 1212 -2190 1218 -2184
rect 1212 -2196 1218 -2190
rect 1212 -2202 1218 -2196
rect 1212 -2208 1218 -2202
rect 1212 -2214 1218 -2208
rect 1212 -2220 1218 -2214
rect 1212 -2226 1218 -2220
rect 1212 -2232 1218 -2226
rect 1212 -2238 1218 -2232
rect 1212 -2244 1218 -2238
rect 1212 -2250 1218 -2244
rect 1212 -2256 1218 -2250
rect 1212 -2262 1218 -2256
rect 1212 -2268 1218 -2262
rect 1212 -2274 1218 -2268
rect 1212 -2280 1218 -2274
rect 1212 -2286 1218 -2280
rect 1212 -2292 1218 -2286
rect 1212 -2298 1218 -2292
rect 1212 -2304 1218 -2298
rect 1212 -2310 1218 -2304
rect 1212 -2316 1218 -2310
rect 1212 -2322 1218 -2316
rect 1212 -2328 1218 -2322
rect 1212 -2334 1218 -2328
rect 1212 -2340 1218 -2334
rect 1212 -2346 1218 -2340
rect 1212 -2352 1218 -2346
rect 1212 -2358 1218 -2352
rect 1212 -2364 1218 -2358
rect 1212 -2370 1218 -2364
rect 1212 -2376 1218 -2370
rect 1212 -2382 1218 -2376
rect 1212 -2388 1218 -2382
rect 1212 -2394 1218 -2388
rect 1212 -2400 1218 -2394
rect 1212 -2406 1218 -2400
rect 1212 -2412 1218 -2406
rect 1212 -2418 1218 -2412
rect 1212 -2424 1218 -2418
rect 1212 -2430 1218 -2424
rect 1212 -2436 1218 -2430
rect 1212 -2442 1218 -2436
rect 1212 -2448 1218 -2442
rect 1212 -2454 1218 -2448
rect 1212 -2460 1218 -2454
rect 1212 -2466 1218 -2460
rect 1212 -2472 1218 -2466
rect 1212 -2478 1218 -2472
rect 1212 -2484 1218 -2478
rect 1212 -2490 1218 -2484
rect 1212 -2496 1218 -2490
rect 1212 -2502 1218 -2496
rect 1212 -2508 1218 -2502
rect 1212 -2514 1218 -2508
rect 1212 -2520 1218 -2514
rect 1212 -2526 1218 -2520
rect 1212 -2532 1218 -2526
rect 1212 -2538 1218 -2532
rect 1212 -2544 1218 -2538
rect 1212 -2550 1218 -2544
rect 1212 -2556 1218 -2550
rect 1212 -2562 1218 -2556
rect 1212 -2568 1218 -2562
rect 1212 -2574 1218 -2568
rect 1212 -2580 1218 -2574
rect 1212 -2586 1218 -2580
rect 1212 -2682 1218 -2676
rect 1212 -2688 1218 -2682
rect 1212 -2694 1218 -2688
rect 1212 -2700 1218 -2694
rect 1212 -2706 1218 -2700
rect 1212 -2712 1218 -2706
rect 1212 -2718 1218 -2712
rect 1212 -2724 1218 -2718
rect 1212 -2730 1218 -2724
rect 1212 -2736 1218 -2730
rect 1212 -2742 1218 -2736
rect 1212 -2748 1218 -2742
rect 1212 -2754 1218 -2748
rect 1212 -2760 1218 -2754
rect 1212 -2766 1218 -2760
rect 1212 -2772 1218 -2766
rect 1212 -2778 1218 -2772
rect 1212 -2784 1218 -2778
rect 1212 -2790 1218 -2784
rect 1212 -2796 1218 -2790
rect 1212 -2802 1218 -2796
rect 1212 -2808 1218 -2802
rect 1212 -2814 1218 -2808
rect 1212 -2820 1218 -2814
rect 1212 -2826 1218 -2820
rect 1212 -2832 1218 -2826
rect 1212 -2838 1218 -2832
rect 1212 -2844 1218 -2838
rect 1212 -2850 1218 -2844
rect 1212 -2856 1218 -2850
rect 1212 -2862 1218 -2856
rect 1212 -2868 1218 -2862
rect 1212 -2874 1218 -2868
rect 1212 -2880 1218 -2874
rect 1212 -2886 1218 -2880
rect 1212 -2892 1218 -2886
rect 1212 -2898 1218 -2892
rect 1212 -2904 1218 -2898
rect 1212 -2910 1218 -2904
rect 1212 -2916 1218 -2910
rect 1212 -2922 1218 -2916
rect 1212 -2928 1218 -2922
rect 1212 -2934 1218 -2928
rect 1212 -2940 1218 -2934
rect 1212 -2946 1218 -2940
rect 1212 -2952 1218 -2946
rect 1212 -2958 1218 -2952
rect 1212 -2964 1218 -2958
rect 1212 -2970 1218 -2964
rect 1212 -2976 1218 -2970
rect 1212 -2982 1218 -2976
rect 1212 -2988 1218 -2982
rect 1212 -2994 1218 -2988
rect 1212 -3000 1218 -2994
rect 1212 -3006 1218 -3000
rect 1212 -3012 1218 -3006
rect 1212 -3090 1218 -3084
rect 1212 -3096 1218 -3090
rect 1212 -3102 1218 -3096
rect 1212 -3108 1218 -3102
rect 1212 -3114 1218 -3108
rect 1212 -3120 1218 -3114
rect 1212 -3126 1218 -3120
rect 1212 -3132 1218 -3126
rect 1212 -3138 1218 -3132
rect 1212 -3144 1218 -3138
rect 1212 -3150 1218 -3144
rect 1212 -3156 1218 -3150
rect 1212 -3162 1218 -3156
rect 1212 -3168 1218 -3162
rect 1212 -3174 1218 -3168
rect 1212 -3180 1218 -3174
rect 1212 -3186 1218 -3180
rect 1212 -3192 1218 -3186
rect 1212 -3198 1218 -3192
rect 1212 -3204 1218 -3198
rect 1212 -3210 1218 -3204
rect 1212 -3216 1218 -3210
rect 1212 -3222 1218 -3216
rect 1212 -3228 1218 -3222
rect 1212 -3234 1218 -3228
rect 1212 -3240 1218 -3234
rect 1212 -3324 1218 -3318
rect 1212 -3330 1218 -3324
rect 1212 -3336 1218 -3330
rect 1212 -3342 1218 -3336
rect 1212 -3348 1218 -3342
rect 1212 -3354 1218 -3348
rect 1212 -3360 1218 -3354
rect 1212 -3366 1218 -3360
rect 1212 -3372 1218 -3366
rect 1212 -3378 1218 -3372
rect 1212 -3384 1218 -3378
rect 1212 -3390 1218 -3384
rect 1212 -3396 1218 -3390
rect 1212 -3402 1218 -3396
rect 1212 -3408 1218 -3402
rect 1212 -3414 1218 -3408
rect 1212 -3420 1218 -3414
rect 1212 -3426 1218 -3420
rect 1212 -3432 1218 -3426
rect 1212 -3438 1218 -3432
rect 1212 -3444 1218 -3438
rect 1212 -3450 1218 -3444
rect 1212 -3456 1218 -3450
rect 1212 -3462 1218 -3456
rect 1212 -3468 1218 -3462
rect 1212 -3474 1218 -3468
rect 1212 -3480 1218 -3474
rect 1212 -3486 1218 -3480
rect 1212 -3492 1218 -3486
rect 1212 -3498 1218 -3492
rect 1212 -3504 1218 -3498
rect 1212 -3510 1218 -3504
rect 1212 -3516 1218 -3510
rect 1212 -3522 1218 -3516
rect 1218 -1104 1224 -1098
rect 1218 -1110 1224 -1104
rect 1218 -1116 1224 -1110
rect 1218 -1122 1224 -1116
rect 1218 -1128 1224 -1122
rect 1218 -1134 1224 -1128
rect 1218 -1140 1224 -1134
rect 1218 -1146 1224 -1140
rect 1218 -1152 1224 -1146
rect 1218 -1158 1224 -1152
rect 1218 -1164 1224 -1158
rect 1218 -1170 1224 -1164
rect 1218 -1176 1224 -1170
rect 1218 -1182 1224 -1176
rect 1218 -1188 1224 -1182
rect 1218 -1194 1224 -1188
rect 1218 -1200 1224 -1194
rect 1218 -1206 1224 -1200
rect 1218 -1212 1224 -1206
rect 1218 -1218 1224 -1212
rect 1218 -1224 1224 -1218
rect 1218 -1230 1224 -1224
rect 1218 -1236 1224 -1230
rect 1218 -1242 1224 -1236
rect 1218 -1248 1224 -1242
rect 1218 -1254 1224 -1248
rect 1218 -1260 1224 -1254
rect 1218 -1266 1224 -1260
rect 1218 -1272 1224 -1266
rect 1218 -1278 1224 -1272
rect 1218 -1284 1224 -1278
rect 1218 -1290 1224 -1284
rect 1218 -1296 1224 -1290
rect 1218 -1302 1224 -1296
rect 1218 -1308 1224 -1302
rect 1218 -1764 1224 -1758
rect 1218 -1770 1224 -1764
rect 1218 -1776 1224 -1770
rect 1218 -1782 1224 -1776
rect 1218 -1788 1224 -1782
rect 1218 -1794 1224 -1788
rect 1218 -1800 1224 -1794
rect 1218 -1806 1224 -1800
rect 1218 -1812 1224 -1806
rect 1218 -1818 1224 -1812
rect 1218 -1824 1224 -1818
rect 1218 -1830 1224 -1824
rect 1218 -1836 1224 -1830
rect 1218 -1842 1224 -1836
rect 1218 -1848 1224 -1842
rect 1218 -1854 1224 -1848
rect 1218 -1860 1224 -1854
rect 1218 -1866 1224 -1860
rect 1218 -1872 1224 -1866
rect 1218 -1878 1224 -1872
rect 1218 -1884 1224 -1878
rect 1218 -1890 1224 -1884
rect 1218 -1896 1224 -1890
rect 1218 -1902 1224 -1896
rect 1218 -1908 1224 -1902
rect 1218 -1914 1224 -1908
rect 1218 -1920 1224 -1914
rect 1218 -1926 1224 -1920
rect 1218 -1932 1224 -1926
rect 1218 -1938 1224 -1932
rect 1218 -1944 1224 -1938
rect 1218 -1950 1224 -1944
rect 1218 -1956 1224 -1950
rect 1218 -1962 1224 -1956
rect 1218 -1968 1224 -1962
rect 1218 -1974 1224 -1968
rect 1218 -1980 1224 -1974
rect 1218 -1986 1224 -1980
rect 1218 -1992 1224 -1986
rect 1218 -1998 1224 -1992
rect 1218 -2004 1224 -1998
rect 1218 -2010 1224 -2004
rect 1218 -2016 1224 -2010
rect 1218 -2022 1224 -2016
rect 1218 -2028 1224 -2022
rect 1218 -2034 1224 -2028
rect 1218 -2040 1224 -2034
rect 1218 -2046 1224 -2040
rect 1218 -2052 1224 -2046
rect 1218 -2058 1224 -2052
rect 1218 -2064 1224 -2058
rect 1218 -2070 1224 -2064
rect 1218 -2076 1224 -2070
rect 1218 -2082 1224 -2076
rect 1218 -2088 1224 -2082
rect 1218 -2094 1224 -2088
rect 1218 -2100 1224 -2094
rect 1218 -2106 1224 -2100
rect 1218 -2112 1224 -2106
rect 1218 -2118 1224 -2112
rect 1218 -2124 1224 -2118
rect 1218 -2130 1224 -2124
rect 1218 -2136 1224 -2130
rect 1218 -2142 1224 -2136
rect 1218 -2148 1224 -2142
rect 1218 -2154 1224 -2148
rect 1218 -2160 1224 -2154
rect 1218 -2166 1224 -2160
rect 1218 -2172 1224 -2166
rect 1218 -2178 1224 -2172
rect 1218 -2184 1224 -2178
rect 1218 -2190 1224 -2184
rect 1218 -2196 1224 -2190
rect 1218 -2202 1224 -2196
rect 1218 -2208 1224 -2202
rect 1218 -2214 1224 -2208
rect 1218 -2220 1224 -2214
rect 1218 -2226 1224 -2220
rect 1218 -2232 1224 -2226
rect 1218 -2238 1224 -2232
rect 1218 -2244 1224 -2238
rect 1218 -2250 1224 -2244
rect 1218 -2256 1224 -2250
rect 1218 -2262 1224 -2256
rect 1218 -2268 1224 -2262
rect 1218 -2274 1224 -2268
rect 1218 -2280 1224 -2274
rect 1218 -2286 1224 -2280
rect 1218 -2292 1224 -2286
rect 1218 -2298 1224 -2292
rect 1218 -2304 1224 -2298
rect 1218 -2310 1224 -2304
rect 1218 -2316 1224 -2310
rect 1218 -2322 1224 -2316
rect 1218 -2328 1224 -2322
rect 1218 -2334 1224 -2328
rect 1218 -2340 1224 -2334
rect 1218 -2346 1224 -2340
rect 1218 -2352 1224 -2346
rect 1218 -2358 1224 -2352
rect 1218 -2364 1224 -2358
rect 1218 -2370 1224 -2364
rect 1218 -2376 1224 -2370
rect 1218 -2382 1224 -2376
rect 1218 -2388 1224 -2382
rect 1218 -2394 1224 -2388
rect 1218 -2400 1224 -2394
rect 1218 -2406 1224 -2400
rect 1218 -2412 1224 -2406
rect 1218 -2418 1224 -2412
rect 1218 -2424 1224 -2418
rect 1218 -2430 1224 -2424
rect 1218 -2436 1224 -2430
rect 1218 -2442 1224 -2436
rect 1218 -2448 1224 -2442
rect 1218 -2454 1224 -2448
rect 1218 -2460 1224 -2454
rect 1218 -2466 1224 -2460
rect 1218 -2472 1224 -2466
rect 1218 -2478 1224 -2472
rect 1218 -2484 1224 -2478
rect 1218 -2490 1224 -2484
rect 1218 -2496 1224 -2490
rect 1218 -2502 1224 -2496
rect 1218 -2508 1224 -2502
rect 1218 -2514 1224 -2508
rect 1218 -2520 1224 -2514
rect 1218 -2526 1224 -2520
rect 1218 -2532 1224 -2526
rect 1218 -2538 1224 -2532
rect 1218 -2544 1224 -2538
rect 1218 -2550 1224 -2544
rect 1218 -2556 1224 -2550
rect 1218 -2562 1224 -2556
rect 1218 -2568 1224 -2562
rect 1218 -2574 1224 -2568
rect 1218 -2580 1224 -2574
rect 1218 -2670 1224 -2664
rect 1218 -2676 1224 -2670
rect 1218 -2682 1224 -2676
rect 1218 -2688 1224 -2682
rect 1218 -2694 1224 -2688
rect 1218 -2700 1224 -2694
rect 1218 -2706 1224 -2700
rect 1218 -2712 1224 -2706
rect 1218 -2718 1224 -2712
rect 1218 -2724 1224 -2718
rect 1218 -2730 1224 -2724
rect 1218 -2736 1224 -2730
rect 1218 -2742 1224 -2736
rect 1218 -2748 1224 -2742
rect 1218 -2754 1224 -2748
rect 1218 -2760 1224 -2754
rect 1218 -2766 1224 -2760
rect 1218 -2772 1224 -2766
rect 1218 -2778 1224 -2772
rect 1218 -2784 1224 -2778
rect 1218 -2790 1224 -2784
rect 1218 -2796 1224 -2790
rect 1218 -2802 1224 -2796
rect 1218 -2808 1224 -2802
rect 1218 -2814 1224 -2808
rect 1218 -2820 1224 -2814
rect 1218 -2826 1224 -2820
rect 1218 -2832 1224 -2826
rect 1218 -2838 1224 -2832
rect 1218 -2844 1224 -2838
rect 1218 -2850 1224 -2844
rect 1218 -2856 1224 -2850
rect 1218 -2862 1224 -2856
rect 1218 -2868 1224 -2862
rect 1218 -2874 1224 -2868
rect 1218 -2880 1224 -2874
rect 1218 -2886 1224 -2880
rect 1218 -2892 1224 -2886
rect 1218 -2898 1224 -2892
rect 1218 -2904 1224 -2898
rect 1218 -2910 1224 -2904
rect 1218 -2916 1224 -2910
rect 1218 -2922 1224 -2916
rect 1218 -2928 1224 -2922
rect 1218 -2934 1224 -2928
rect 1218 -2940 1224 -2934
rect 1218 -2946 1224 -2940
rect 1218 -2952 1224 -2946
rect 1218 -2958 1224 -2952
rect 1218 -2964 1224 -2958
rect 1218 -2970 1224 -2964
rect 1218 -2976 1224 -2970
rect 1218 -2982 1224 -2976
rect 1218 -2988 1224 -2982
rect 1218 -2994 1224 -2988
rect 1218 -3000 1224 -2994
rect 1218 -3006 1224 -3000
rect 1218 -3084 1224 -3078
rect 1218 -3090 1224 -3084
rect 1218 -3096 1224 -3090
rect 1218 -3102 1224 -3096
rect 1218 -3108 1224 -3102
rect 1218 -3114 1224 -3108
rect 1218 -3120 1224 -3114
rect 1218 -3126 1224 -3120
rect 1218 -3132 1224 -3126
rect 1218 -3138 1224 -3132
rect 1218 -3144 1224 -3138
rect 1218 -3150 1224 -3144
rect 1218 -3156 1224 -3150
rect 1218 -3162 1224 -3156
rect 1218 -3168 1224 -3162
rect 1218 -3174 1224 -3168
rect 1218 -3180 1224 -3174
rect 1218 -3186 1224 -3180
rect 1218 -3192 1224 -3186
rect 1218 -3198 1224 -3192
rect 1218 -3204 1224 -3198
rect 1218 -3210 1224 -3204
rect 1218 -3216 1224 -3210
rect 1218 -3222 1224 -3216
rect 1218 -3228 1224 -3222
rect 1218 -3234 1224 -3228
rect 1218 -3240 1224 -3234
rect 1218 -3324 1224 -3318
rect 1218 -3330 1224 -3324
rect 1218 -3336 1224 -3330
rect 1218 -3342 1224 -3336
rect 1218 -3348 1224 -3342
rect 1218 -3354 1224 -3348
rect 1218 -3360 1224 -3354
rect 1218 -3366 1224 -3360
rect 1218 -3372 1224 -3366
rect 1218 -3378 1224 -3372
rect 1218 -3384 1224 -3378
rect 1218 -3390 1224 -3384
rect 1218 -3396 1224 -3390
rect 1218 -3402 1224 -3396
rect 1218 -3408 1224 -3402
rect 1218 -3414 1224 -3408
rect 1218 -3420 1224 -3414
rect 1218 -3426 1224 -3420
rect 1218 -3432 1224 -3426
rect 1218 -3438 1224 -3432
rect 1218 -3444 1224 -3438
rect 1218 -3450 1224 -3444
rect 1218 -3456 1224 -3450
rect 1218 -3462 1224 -3456
rect 1218 -3468 1224 -3462
rect 1218 -3474 1224 -3468
rect 1218 -3480 1224 -3474
rect 1218 -3486 1224 -3480
rect 1218 -3492 1224 -3486
rect 1218 -3498 1224 -3492
rect 1218 -3504 1224 -3498
rect 1218 -3510 1224 -3504
rect 1218 -3516 1224 -3510
rect 1218 -3522 1224 -3516
rect 1224 -1104 1230 -1098
rect 1224 -1110 1230 -1104
rect 1224 -1116 1230 -1110
rect 1224 -1122 1230 -1116
rect 1224 -1128 1230 -1122
rect 1224 -1134 1230 -1128
rect 1224 -1140 1230 -1134
rect 1224 -1146 1230 -1140
rect 1224 -1152 1230 -1146
rect 1224 -1158 1230 -1152
rect 1224 -1164 1230 -1158
rect 1224 -1170 1230 -1164
rect 1224 -1176 1230 -1170
rect 1224 -1182 1230 -1176
rect 1224 -1188 1230 -1182
rect 1224 -1194 1230 -1188
rect 1224 -1200 1230 -1194
rect 1224 -1206 1230 -1200
rect 1224 -1212 1230 -1206
rect 1224 -1218 1230 -1212
rect 1224 -1224 1230 -1218
rect 1224 -1230 1230 -1224
rect 1224 -1236 1230 -1230
rect 1224 -1242 1230 -1236
rect 1224 -1248 1230 -1242
rect 1224 -1254 1230 -1248
rect 1224 -1260 1230 -1254
rect 1224 -1266 1230 -1260
rect 1224 -1272 1230 -1266
rect 1224 -1278 1230 -1272
rect 1224 -1284 1230 -1278
rect 1224 -1290 1230 -1284
rect 1224 -1296 1230 -1290
rect 1224 -1302 1230 -1296
rect 1224 -1308 1230 -1302
rect 1224 -1752 1230 -1746
rect 1224 -1758 1230 -1752
rect 1224 -1764 1230 -1758
rect 1224 -1770 1230 -1764
rect 1224 -1776 1230 -1770
rect 1224 -1782 1230 -1776
rect 1224 -1788 1230 -1782
rect 1224 -1794 1230 -1788
rect 1224 -1800 1230 -1794
rect 1224 -1806 1230 -1800
rect 1224 -1812 1230 -1806
rect 1224 -1818 1230 -1812
rect 1224 -1824 1230 -1818
rect 1224 -1830 1230 -1824
rect 1224 -1836 1230 -1830
rect 1224 -1842 1230 -1836
rect 1224 -1848 1230 -1842
rect 1224 -1854 1230 -1848
rect 1224 -1860 1230 -1854
rect 1224 -1866 1230 -1860
rect 1224 -1872 1230 -1866
rect 1224 -1878 1230 -1872
rect 1224 -1884 1230 -1878
rect 1224 -1890 1230 -1884
rect 1224 -1896 1230 -1890
rect 1224 -1902 1230 -1896
rect 1224 -1908 1230 -1902
rect 1224 -1914 1230 -1908
rect 1224 -1920 1230 -1914
rect 1224 -1926 1230 -1920
rect 1224 -1932 1230 -1926
rect 1224 -1938 1230 -1932
rect 1224 -1944 1230 -1938
rect 1224 -1950 1230 -1944
rect 1224 -1956 1230 -1950
rect 1224 -1962 1230 -1956
rect 1224 -1968 1230 -1962
rect 1224 -1974 1230 -1968
rect 1224 -1980 1230 -1974
rect 1224 -1986 1230 -1980
rect 1224 -1992 1230 -1986
rect 1224 -1998 1230 -1992
rect 1224 -2004 1230 -1998
rect 1224 -2010 1230 -2004
rect 1224 -2016 1230 -2010
rect 1224 -2022 1230 -2016
rect 1224 -2028 1230 -2022
rect 1224 -2034 1230 -2028
rect 1224 -2040 1230 -2034
rect 1224 -2046 1230 -2040
rect 1224 -2052 1230 -2046
rect 1224 -2058 1230 -2052
rect 1224 -2064 1230 -2058
rect 1224 -2070 1230 -2064
rect 1224 -2076 1230 -2070
rect 1224 -2082 1230 -2076
rect 1224 -2088 1230 -2082
rect 1224 -2094 1230 -2088
rect 1224 -2100 1230 -2094
rect 1224 -2106 1230 -2100
rect 1224 -2112 1230 -2106
rect 1224 -2118 1230 -2112
rect 1224 -2124 1230 -2118
rect 1224 -2130 1230 -2124
rect 1224 -2136 1230 -2130
rect 1224 -2142 1230 -2136
rect 1224 -2148 1230 -2142
rect 1224 -2154 1230 -2148
rect 1224 -2160 1230 -2154
rect 1224 -2166 1230 -2160
rect 1224 -2172 1230 -2166
rect 1224 -2178 1230 -2172
rect 1224 -2184 1230 -2178
rect 1224 -2190 1230 -2184
rect 1224 -2196 1230 -2190
rect 1224 -2202 1230 -2196
rect 1224 -2208 1230 -2202
rect 1224 -2214 1230 -2208
rect 1224 -2220 1230 -2214
rect 1224 -2226 1230 -2220
rect 1224 -2232 1230 -2226
rect 1224 -2238 1230 -2232
rect 1224 -2244 1230 -2238
rect 1224 -2250 1230 -2244
rect 1224 -2256 1230 -2250
rect 1224 -2262 1230 -2256
rect 1224 -2268 1230 -2262
rect 1224 -2274 1230 -2268
rect 1224 -2280 1230 -2274
rect 1224 -2286 1230 -2280
rect 1224 -2292 1230 -2286
rect 1224 -2298 1230 -2292
rect 1224 -2304 1230 -2298
rect 1224 -2310 1230 -2304
rect 1224 -2316 1230 -2310
rect 1224 -2322 1230 -2316
rect 1224 -2328 1230 -2322
rect 1224 -2334 1230 -2328
rect 1224 -2340 1230 -2334
rect 1224 -2346 1230 -2340
rect 1224 -2352 1230 -2346
rect 1224 -2358 1230 -2352
rect 1224 -2364 1230 -2358
rect 1224 -2370 1230 -2364
rect 1224 -2376 1230 -2370
rect 1224 -2382 1230 -2376
rect 1224 -2388 1230 -2382
rect 1224 -2394 1230 -2388
rect 1224 -2400 1230 -2394
rect 1224 -2406 1230 -2400
rect 1224 -2412 1230 -2406
rect 1224 -2418 1230 -2412
rect 1224 -2424 1230 -2418
rect 1224 -2430 1230 -2424
rect 1224 -2436 1230 -2430
rect 1224 -2442 1230 -2436
rect 1224 -2448 1230 -2442
rect 1224 -2454 1230 -2448
rect 1224 -2460 1230 -2454
rect 1224 -2466 1230 -2460
rect 1224 -2472 1230 -2466
rect 1224 -2478 1230 -2472
rect 1224 -2484 1230 -2478
rect 1224 -2490 1230 -2484
rect 1224 -2496 1230 -2490
rect 1224 -2502 1230 -2496
rect 1224 -2508 1230 -2502
rect 1224 -2514 1230 -2508
rect 1224 -2520 1230 -2514
rect 1224 -2526 1230 -2520
rect 1224 -2532 1230 -2526
rect 1224 -2538 1230 -2532
rect 1224 -2544 1230 -2538
rect 1224 -2550 1230 -2544
rect 1224 -2556 1230 -2550
rect 1224 -2562 1230 -2556
rect 1224 -2568 1230 -2562
rect 1224 -2658 1230 -2652
rect 1224 -2664 1230 -2658
rect 1224 -2670 1230 -2664
rect 1224 -2676 1230 -2670
rect 1224 -2682 1230 -2676
rect 1224 -2688 1230 -2682
rect 1224 -2694 1230 -2688
rect 1224 -2700 1230 -2694
rect 1224 -2706 1230 -2700
rect 1224 -2712 1230 -2706
rect 1224 -2718 1230 -2712
rect 1224 -2724 1230 -2718
rect 1224 -2730 1230 -2724
rect 1224 -2736 1230 -2730
rect 1224 -2742 1230 -2736
rect 1224 -2748 1230 -2742
rect 1224 -2754 1230 -2748
rect 1224 -2760 1230 -2754
rect 1224 -2766 1230 -2760
rect 1224 -2772 1230 -2766
rect 1224 -2778 1230 -2772
rect 1224 -2784 1230 -2778
rect 1224 -2790 1230 -2784
rect 1224 -2796 1230 -2790
rect 1224 -2802 1230 -2796
rect 1224 -2808 1230 -2802
rect 1224 -2814 1230 -2808
rect 1224 -2820 1230 -2814
rect 1224 -2826 1230 -2820
rect 1224 -2832 1230 -2826
rect 1224 -2838 1230 -2832
rect 1224 -2844 1230 -2838
rect 1224 -2850 1230 -2844
rect 1224 -2856 1230 -2850
rect 1224 -2862 1230 -2856
rect 1224 -2868 1230 -2862
rect 1224 -2874 1230 -2868
rect 1224 -2880 1230 -2874
rect 1224 -2886 1230 -2880
rect 1224 -2892 1230 -2886
rect 1224 -2898 1230 -2892
rect 1224 -2904 1230 -2898
rect 1224 -2910 1230 -2904
rect 1224 -2916 1230 -2910
rect 1224 -2922 1230 -2916
rect 1224 -2928 1230 -2922
rect 1224 -2934 1230 -2928
rect 1224 -2940 1230 -2934
rect 1224 -2946 1230 -2940
rect 1224 -2952 1230 -2946
rect 1224 -2958 1230 -2952
rect 1224 -2964 1230 -2958
rect 1224 -2970 1230 -2964
rect 1224 -2976 1230 -2970
rect 1224 -2982 1230 -2976
rect 1224 -2988 1230 -2982
rect 1224 -2994 1230 -2988
rect 1224 -3000 1230 -2994
rect 1224 -3078 1230 -3072
rect 1224 -3084 1230 -3078
rect 1224 -3090 1230 -3084
rect 1224 -3096 1230 -3090
rect 1224 -3102 1230 -3096
rect 1224 -3108 1230 -3102
rect 1224 -3114 1230 -3108
rect 1224 -3120 1230 -3114
rect 1224 -3126 1230 -3120
rect 1224 -3132 1230 -3126
rect 1224 -3138 1230 -3132
rect 1224 -3144 1230 -3138
rect 1224 -3150 1230 -3144
rect 1224 -3156 1230 -3150
rect 1224 -3162 1230 -3156
rect 1224 -3168 1230 -3162
rect 1224 -3174 1230 -3168
rect 1224 -3180 1230 -3174
rect 1224 -3186 1230 -3180
rect 1224 -3192 1230 -3186
rect 1224 -3198 1230 -3192
rect 1224 -3204 1230 -3198
rect 1224 -3210 1230 -3204
rect 1224 -3216 1230 -3210
rect 1224 -3222 1230 -3216
rect 1224 -3228 1230 -3222
rect 1224 -3234 1230 -3228
rect 1224 -3240 1230 -3234
rect 1224 -3324 1230 -3318
rect 1224 -3330 1230 -3324
rect 1224 -3336 1230 -3330
rect 1224 -3342 1230 -3336
rect 1224 -3348 1230 -3342
rect 1224 -3354 1230 -3348
rect 1224 -3360 1230 -3354
rect 1224 -3366 1230 -3360
rect 1224 -3372 1230 -3366
rect 1224 -3378 1230 -3372
rect 1224 -3384 1230 -3378
rect 1224 -3390 1230 -3384
rect 1224 -3396 1230 -3390
rect 1224 -3402 1230 -3396
rect 1224 -3408 1230 -3402
rect 1224 -3414 1230 -3408
rect 1224 -3420 1230 -3414
rect 1224 -3426 1230 -3420
rect 1224 -3432 1230 -3426
rect 1224 -3438 1230 -3432
rect 1224 -3444 1230 -3438
rect 1224 -3450 1230 -3444
rect 1224 -3456 1230 -3450
rect 1224 -3462 1230 -3456
rect 1224 -3468 1230 -3462
rect 1224 -3474 1230 -3468
rect 1224 -3480 1230 -3474
rect 1224 -3486 1230 -3480
rect 1224 -3492 1230 -3486
rect 1224 -3498 1230 -3492
rect 1224 -3504 1230 -3498
rect 1224 -3510 1230 -3504
rect 1224 -3516 1230 -3510
rect 1224 -3522 1230 -3516
rect 1230 -1104 1236 -1098
rect 1230 -1110 1236 -1104
rect 1230 -1116 1236 -1110
rect 1230 -1122 1236 -1116
rect 1230 -1128 1236 -1122
rect 1230 -1134 1236 -1128
rect 1230 -1140 1236 -1134
rect 1230 -1146 1236 -1140
rect 1230 -1152 1236 -1146
rect 1230 -1158 1236 -1152
rect 1230 -1164 1236 -1158
rect 1230 -1170 1236 -1164
rect 1230 -1176 1236 -1170
rect 1230 -1182 1236 -1176
rect 1230 -1188 1236 -1182
rect 1230 -1194 1236 -1188
rect 1230 -1200 1236 -1194
rect 1230 -1206 1236 -1200
rect 1230 -1212 1236 -1206
rect 1230 -1218 1236 -1212
rect 1230 -1224 1236 -1218
rect 1230 -1230 1236 -1224
rect 1230 -1236 1236 -1230
rect 1230 -1242 1236 -1236
rect 1230 -1248 1236 -1242
rect 1230 -1254 1236 -1248
rect 1230 -1260 1236 -1254
rect 1230 -1266 1236 -1260
rect 1230 -1272 1236 -1266
rect 1230 -1278 1236 -1272
rect 1230 -1284 1236 -1278
rect 1230 -1290 1236 -1284
rect 1230 -1296 1236 -1290
rect 1230 -1302 1236 -1296
rect 1230 -1308 1236 -1302
rect 1230 -1734 1236 -1728
rect 1230 -1740 1236 -1734
rect 1230 -1746 1236 -1740
rect 1230 -1752 1236 -1746
rect 1230 -1758 1236 -1752
rect 1230 -1764 1236 -1758
rect 1230 -1770 1236 -1764
rect 1230 -1776 1236 -1770
rect 1230 -1782 1236 -1776
rect 1230 -1788 1236 -1782
rect 1230 -1794 1236 -1788
rect 1230 -1800 1236 -1794
rect 1230 -1806 1236 -1800
rect 1230 -1812 1236 -1806
rect 1230 -1818 1236 -1812
rect 1230 -1824 1236 -1818
rect 1230 -1830 1236 -1824
rect 1230 -1836 1236 -1830
rect 1230 -1842 1236 -1836
rect 1230 -1848 1236 -1842
rect 1230 -1854 1236 -1848
rect 1230 -1860 1236 -1854
rect 1230 -1866 1236 -1860
rect 1230 -1872 1236 -1866
rect 1230 -1878 1236 -1872
rect 1230 -1884 1236 -1878
rect 1230 -1890 1236 -1884
rect 1230 -1896 1236 -1890
rect 1230 -1902 1236 -1896
rect 1230 -1908 1236 -1902
rect 1230 -1914 1236 -1908
rect 1230 -1920 1236 -1914
rect 1230 -1926 1236 -1920
rect 1230 -1932 1236 -1926
rect 1230 -1938 1236 -1932
rect 1230 -1944 1236 -1938
rect 1230 -1950 1236 -1944
rect 1230 -1956 1236 -1950
rect 1230 -1962 1236 -1956
rect 1230 -1968 1236 -1962
rect 1230 -1974 1236 -1968
rect 1230 -1980 1236 -1974
rect 1230 -1986 1236 -1980
rect 1230 -1992 1236 -1986
rect 1230 -1998 1236 -1992
rect 1230 -2004 1236 -1998
rect 1230 -2010 1236 -2004
rect 1230 -2016 1236 -2010
rect 1230 -2022 1236 -2016
rect 1230 -2028 1236 -2022
rect 1230 -2034 1236 -2028
rect 1230 -2040 1236 -2034
rect 1230 -2046 1236 -2040
rect 1230 -2052 1236 -2046
rect 1230 -2058 1236 -2052
rect 1230 -2064 1236 -2058
rect 1230 -2070 1236 -2064
rect 1230 -2076 1236 -2070
rect 1230 -2082 1236 -2076
rect 1230 -2088 1236 -2082
rect 1230 -2094 1236 -2088
rect 1230 -2100 1236 -2094
rect 1230 -2106 1236 -2100
rect 1230 -2112 1236 -2106
rect 1230 -2118 1236 -2112
rect 1230 -2124 1236 -2118
rect 1230 -2130 1236 -2124
rect 1230 -2136 1236 -2130
rect 1230 -2142 1236 -2136
rect 1230 -2148 1236 -2142
rect 1230 -2154 1236 -2148
rect 1230 -2160 1236 -2154
rect 1230 -2166 1236 -2160
rect 1230 -2172 1236 -2166
rect 1230 -2178 1236 -2172
rect 1230 -2184 1236 -2178
rect 1230 -2190 1236 -2184
rect 1230 -2196 1236 -2190
rect 1230 -2202 1236 -2196
rect 1230 -2208 1236 -2202
rect 1230 -2214 1236 -2208
rect 1230 -2220 1236 -2214
rect 1230 -2226 1236 -2220
rect 1230 -2232 1236 -2226
rect 1230 -2238 1236 -2232
rect 1230 -2244 1236 -2238
rect 1230 -2250 1236 -2244
rect 1230 -2256 1236 -2250
rect 1230 -2262 1236 -2256
rect 1230 -2268 1236 -2262
rect 1230 -2274 1236 -2268
rect 1230 -2280 1236 -2274
rect 1230 -2286 1236 -2280
rect 1230 -2292 1236 -2286
rect 1230 -2298 1236 -2292
rect 1230 -2304 1236 -2298
rect 1230 -2310 1236 -2304
rect 1230 -2316 1236 -2310
rect 1230 -2322 1236 -2316
rect 1230 -2328 1236 -2322
rect 1230 -2334 1236 -2328
rect 1230 -2340 1236 -2334
rect 1230 -2346 1236 -2340
rect 1230 -2352 1236 -2346
rect 1230 -2358 1236 -2352
rect 1230 -2364 1236 -2358
rect 1230 -2370 1236 -2364
rect 1230 -2376 1236 -2370
rect 1230 -2382 1236 -2376
rect 1230 -2388 1236 -2382
rect 1230 -2394 1236 -2388
rect 1230 -2400 1236 -2394
rect 1230 -2406 1236 -2400
rect 1230 -2412 1236 -2406
rect 1230 -2418 1236 -2412
rect 1230 -2424 1236 -2418
rect 1230 -2430 1236 -2424
rect 1230 -2436 1236 -2430
rect 1230 -2442 1236 -2436
rect 1230 -2448 1236 -2442
rect 1230 -2454 1236 -2448
rect 1230 -2460 1236 -2454
rect 1230 -2466 1236 -2460
rect 1230 -2472 1236 -2466
rect 1230 -2478 1236 -2472
rect 1230 -2484 1236 -2478
rect 1230 -2490 1236 -2484
rect 1230 -2496 1236 -2490
rect 1230 -2502 1236 -2496
rect 1230 -2508 1236 -2502
rect 1230 -2514 1236 -2508
rect 1230 -2520 1236 -2514
rect 1230 -2526 1236 -2520
rect 1230 -2532 1236 -2526
rect 1230 -2538 1236 -2532
rect 1230 -2544 1236 -2538
rect 1230 -2550 1236 -2544
rect 1230 -2556 1236 -2550
rect 1230 -2562 1236 -2556
rect 1230 -2652 1236 -2646
rect 1230 -2658 1236 -2652
rect 1230 -2664 1236 -2658
rect 1230 -2670 1236 -2664
rect 1230 -2676 1236 -2670
rect 1230 -2682 1236 -2676
rect 1230 -2688 1236 -2682
rect 1230 -2694 1236 -2688
rect 1230 -2700 1236 -2694
rect 1230 -2706 1236 -2700
rect 1230 -2712 1236 -2706
rect 1230 -2718 1236 -2712
rect 1230 -2724 1236 -2718
rect 1230 -2730 1236 -2724
rect 1230 -2736 1236 -2730
rect 1230 -2742 1236 -2736
rect 1230 -2748 1236 -2742
rect 1230 -2754 1236 -2748
rect 1230 -2760 1236 -2754
rect 1230 -2766 1236 -2760
rect 1230 -2772 1236 -2766
rect 1230 -2778 1236 -2772
rect 1230 -2784 1236 -2778
rect 1230 -2790 1236 -2784
rect 1230 -2796 1236 -2790
rect 1230 -2802 1236 -2796
rect 1230 -2808 1236 -2802
rect 1230 -2814 1236 -2808
rect 1230 -2820 1236 -2814
rect 1230 -2826 1236 -2820
rect 1230 -2832 1236 -2826
rect 1230 -2838 1236 -2832
rect 1230 -2844 1236 -2838
rect 1230 -2850 1236 -2844
rect 1230 -2856 1236 -2850
rect 1230 -2862 1236 -2856
rect 1230 -2868 1236 -2862
rect 1230 -2874 1236 -2868
rect 1230 -2880 1236 -2874
rect 1230 -2886 1236 -2880
rect 1230 -2892 1236 -2886
rect 1230 -2898 1236 -2892
rect 1230 -2904 1236 -2898
rect 1230 -2910 1236 -2904
rect 1230 -2916 1236 -2910
rect 1230 -2922 1236 -2916
rect 1230 -2928 1236 -2922
rect 1230 -2934 1236 -2928
rect 1230 -2940 1236 -2934
rect 1230 -2946 1236 -2940
rect 1230 -2952 1236 -2946
rect 1230 -2958 1236 -2952
rect 1230 -2964 1236 -2958
rect 1230 -2970 1236 -2964
rect 1230 -2976 1236 -2970
rect 1230 -2982 1236 -2976
rect 1230 -2988 1236 -2982
rect 1230 -2994 1236 -2988
rect 1230 -3078 1236 -3072
rect 1230 -3084 1236 -3078
rect 1230 -3090 1236 -3084
rect 1230 -3096 1236 -3090
rect 1230 -3102 1236 -3096
rect 1230 -3108 1236 -3102
rect 1230 -3114 1236 -3108
rect 1230 -3120 1236 -3114
rect 1230 -3126 1236 -3120
rect 1230 -3132 1236 -3126
rect 1230 -3138 1236 -3132
rect 1230 -3144 1236 -3138
rect 1230 -3150 1236 -3144
rect 1230 -3156 1236 -3150
rect 1230 -3162 1236 -3156
rect 1230 -3168 1236 -3162
rect 1230 -3174 1236 -3168
rect 1230 -3180 1236 -3174
rect 1230 -3186 1236 -3180
rect 1230 -3192 1236 -3186
rect 1230 -3198 1236 -3192
rect 1230 -3204 1236 -3198
rect 1230 -3210 1236 -3204
rect 1230 -3216 1236 -3210
rect 1230 -3222 1236 -3216
rect 1230 -3228 1236 -3222
rect 1230 -3234 1236 -3228
rect 1230 -3240 1236 -3234
rect 1230 -3324 1236 -3318
rect 1230 -3330 1236 -3324
rect 1230 -3336 1236 -3330
rect 1230 -3342 1236 -3336
rect 1230 -3348 1236 -3342
rect 1230 -3354 1236 -3348
rect 1230 -3360 1236 -3354
rect 1230 -3366 1236 -3360
rect 1230 -3372 1236 -3366
rect 1230 -3378 1236 -3372
rect 1230 -3384 1236 -3378
rect 1230 -3390 1236 -3384
rect 1230 -3396 1236 -3390
rect 1230 -3402 1236 -3396
rect 1230 -3408 1236 -3402
rect 1230 -3414 1236 -3408
rect 1230 -3420 1236 -3414
rect 1230 -3426 1236 -3420
rect 1230 -3432 1236 -3426
rect 1230 -3438 1236 -3432
rect 1230 -3444 1236 -3438
rect 1230 -3450 1236 -3444
rect 1230 -3456 1236 -3450
rect 1230 -3462 1236 -3456
rect 1230 -3468 1236 -3462
rect 1230 -3474 1236 -3468
rect 1230 -3480 1236 -3474
rect 1230 -3486 1236 -3480
rect 1230 -3492 1236 -3486
rect 1230 -3498 1236 -3492
rect 1230 -3504 1236 -3498
rect 1230 -3510 1236 -3504
rect 1230 -3516 1236 -3510
rect 1230 -3522 1236 -3516
rect 1236 -1104 1242 -1098
rect 1236 -1110 1242 -1104
rect 1236 -1116 1242 -1110
rect 1236 -1122 1242 -1116
rect 1236 -1128 1242 -1122
rect 1236 -1134 1242 -1128
rect 1236 -1140 1242 -1134
rect 1236 -1146 1242 -1140
rect 1236 -1152 1242 -1146
rect 1236 -1158 1242 -1152
rect 1236 -1164 1242 -1158
rect 1236 -1170 1242 -1164
rect 1236 -1176 1242 -1170
rect 1236 -1182 1242 -1176
rect 1236 -1188 1242 -1182
rect 1236 -1194 1242 -1188
rect 1236 -1200 1242 -1194
rect 1236 -1206 1242 -1200
rect 1236 -1212 1242 -1206
rect 1236 -1218 1242 -1212
rect 1236 -1224 1242 -1218
rect 1236 -1230 1242 -1224
rect 1236 -1236 1242 -1230
rect 1236 -1242 1242 -1236
rect 1236 -1248 1242 -1242
rect 1236 -1254 1242 -1248
rect 1236 -1260 1242 -1254
rect 1236 -1266 1242 -1260
rect 1236 -1272 1242 -1266
rect 1236 -1278 1242 -1272
rect 1236 -1284 1242 -1278
rect 1236 -1290 1242 -1284
rect 1236 -1296 1242 -1290
rect 1236 -1302 1242 -1296
rect 1236 -1308 1242 -1302
rect 1236 -1722 1242 -1716
rect 1236 -1728 1242 -1722
rect 1236 -1734 1242 -1728
rect 1236 -1740 1242 -1734
rect 1236 -1746 1242 -1740
rect 1236 -1752 1242 -1746
rect 1236 -1758 1242 -1752
rect 1236 -1764 1242 -1758
rect 1236 -1770 1242 -1764
rect 1236 -1776 1242 -1770
rect 1236 -1782 1242 -1776
rect 1236 -1788 1242 -1782
rect 1236 -1794 1242 -1788
rect 1236 -1800 1242 -1794
rect 1236 -1806 1242 -1800
rect 1236 -1812 1242 -1806
rect 1236 -1818 1242 -1812
rect 1236 -1824 1242 -1818
rect 1236 -1830 1242 -1824
rect 1236 -1836 1242 -1830
rect 1236 -1842 1242 -1836
rect 1236 -1848 1242 -1842
rect 1236 -1854 1242 -1848
rect 1236 -1860 1242 -1854
rect 1236 -1866 1242 -1860
rect 1236 -1872 1242 -1866
rect 1236 -1878 1242 -1872
rect 1236 -1884 1242 -1878
rect 1236 -1890 1242 -1884
rect 1236 -1896 1242 -1890
rect 1236 -1902 1242 -1896
rect 1236 -1908 1242 -1902
rect 1236 -1914 1242 -1908
rect 1236 -1920 1242 -1914
rect 1236 -1926 1242 -1920
rect 1236 -1932 1242 -1926
rect 1236 -1938 1242 -1932
rect 1236 -1944 1242 -1938
rect 1236 -1950 1242 -1944
rect 1236 -1956 1242 -1950
rect 1236 -1962 1242 -1956
rect 1236 -1968 1242 -1962
rect 1236 -1974 1242 -1968
rect 1236 -1980 1242 -1974
rect 1236 -1986 1242 -1980
rect 1236 -1992 1242 -1986
rect 1236 -1998 1242 -1992
rect 1236 -2004 1242 -1998
rect 1236 -2010 1242 -2004
rect 1236 -2016 1242 -2010
rect 1236 -2022 1242 -2016
rect 1236 -2028 1242 -2022
rect 1236 -2034 1242 -2028
rect 1236 -2040 1242 -2034
rect 1236 -2046 1242 -2040
rect 1236 -2052 1242 -2046
rect 1236 -2058 1242 -2052
rect 1236 -2064 1242 -2058
rect 1236 -2070 1242 -2064
rect 1236 -2076 1242 -2070
rect 1236 -2082 1242 -2076
rect 1236 -2088 1242 -2082
rect 1236 -2094 1242 -2088
rect 1236 -2100 1242 -2094
rect 1236 -2106 1242 -2100
rect 1236 -2112 1242 -2106
rect 1236 -2118 1242 -2112
rect 1236 -2124 1242 -2118
rect 1236 -2130 1242 -2124
rect 1236 -2136 1242 -2130
rect 1236 -2142 1242 -2136
rect 1236 -2148 1242 -2142
rect 1236 -2154 1242 -2148
rect 1236 -2160 1242 -2154
rect 1236 -2166 1242 -2160
rect 1236 -2172 1242 -2166
rect 1236 -2178 1242 -2172
rect 1236 -2184 1242 -2178
rect 1236 -2190 1242 -2184
rect 1236 -2196 1242 -2190
rect 1236 -2202 1242 -2196
rect 1236 -2208 1242 -2202
rect 1236 -2214 1242 -2208
rect 1236 -2220 1242 -2214
rect 1236 -2226 1242 -2220
rect 1236 -2232 1242 -2226
rect 1236 -2238 1242 -2232
rect 1236 -2244 1242 -2238
rect 1236 -2250 1242 -2244
rect 1236 -2256 1242 -2250
rect 1236 -2262 1242 -2256
rect 1236 -2268 1242 -2262
rect 1236 -2274 1242 -2268
rect 1236 -2280 1242 -2274
rect 1236 -2286 1242 -2280
rect 1236 -2292 1242 -2286
rect 1236 -2298 1242 -2292
rect 1236 -2304 1242 -2298
rect 1236 -2310 1242 -2304
rect 1236 -2316 1242 -2310
rect 1236 -2322 1242 -2316
rect 1236 -2328 1242 -2322
rect 1236 -2334 1242 -2328
rect 1236 -2340 1242 -2334
rect 1236 -2346 1242 -2340
rect 1236 -2352 1242 -2346
rect 1236 -2358 1242 -2352
rect 1236 -2364 1242 -2358
rect 1236 -2370 1242 -2364
rect 1236 -2376 1242 -2370
rect 1236 -2382 1242 -2376
rect 1236 -2388 1242 -2382
rect 1236 -2394 1242 -2388
rect 1236 -2400 1242 -2394
rect 1236 -2406 1242 -2400
rect 1236 -2412 1242 -2406
rect 1236 -2418 1242 -2412
rect 1236 -2424 1242 -2418
rect 1236 -2430 1242 -2424
rect 1236 -2436 1242 -2430
rect 1236 -2442 1242 -2436
rect 1236 -2448 1242 -2442
rect 1236 -2454 1242 -2448
rect 1236 -2460 1242 -2454
rect 1236 -2466 1242 -2460
rect 1236 -2472 1242 -2466
rect 1236 -2478 1242 -2472
rect 1236 -2484 1242 -2478
rect 1236 -2490 1242 -2484
rect 1236 -2496 1242 -2490
rect 1236 -2502 1242 -2496
rect 1236 -2508 1242 -2502
rect 1236 -2514 1242 -2508
rect 1236 -2520 1242 -2514
rect 1236 -2526 1242 -2520
rect 1236 -2532 1242 -2526
rect 1236 -2538 1242 -2532
rect 1236 -2544 1242 -2538
rect 1236 -2550 1242 -2544
rect 1236 -2640 1242 -2634
rect 1236 -2646 1242 -2640
rect 1236 -2652 1242 -2646
rect 1236 -2658 1242 -2652
rect 1236 -2664 1242 -2658
rect 1236 -2670 1242 -2664
rect 1236 -2676 1242 -2670
rect 1236 -2682 1242 -2676
rect 1236 -2688 1242 -2682
rect 1236 -2694 1242 -2688
rect 1236 -2700 1242 -2694
rect 1236 -2706 1242 -2700
rect 1236 -2712 1242 -2706
rect 1236 -2718 1242 -2712
rect 1236 -2724 1242 -2718
rect 1236 -2730 1242 -2724
rect 1236 -2736 1242 -2730
rect 1236 -2742 1242 -2736
rect 1236 -2748 1242 -2742
rect 1236 -2754 1242 -2748
rect 1236 -2760 1242 -2754
rect 1236 -2766 1242 -2760
rect 1236 -2772 1242 -2766
rect 1236 -2778 1242 -2772
rect 1236 -2784 1242 -2778
rect 1236 -2790 1242 -2784
rect 1236 -2796 1242 -2790
rect 1236 -2802 1242 -2796
rect 1236 -2808 1242 -2802
rect 1236 -2814 1242 -2808
rect 1236 -2820 1242 -2814
rect 1236 -2826 1242 -2820
rect 1236 -2832 1242 -2826
rect 1236 -2838 1242 -2832
rect 1236 -2844 1242 -2838
rect 1236 -2850 1242 -2844
rect 1236 -2856 1242 -2850
rect 1236 -2862 1242 -2856
rect 1236 -2868 1242 -2862
rect 1236 -2874 1242 -2868
rect 1236 -2880 1242 -2874
rect 1236 -2886 1242 -2880
rect 1236 -2892 1242 -2886
rect 1236 -2898 1242 -2892
rect 1236 -2904 1242 -2898
rect 1236 -2910 1242 -2904
rect 1236 -2916 1242 -2910
rect 1236 -2922 1242 -2916
rect 1236 -2928 1242 -2922
rect 1236 -2934 1242 -2928
rect 1236 -2940 1242 -2934
rect 1236 -2946 1242 -2940
rect 1236 -2952 1242 -2946
rect 1236 -2958 1242 -2952
rect 1236 -2964 1242 -2958
rect 1236 -2970 1242 -2964
rect 1236 -2976 1242 -2970
rect 1236 -2982 1242 -2976
rect 1236 -2988 1242 -2982
rect 1236 -2994 1242 -2988
rect 1236 -3072 1242 -3066
rect 1236 -3078 1242 -3072
rect 1236 -3084 1242 -3078
rect 1236 -3090 1242 -3084
rect 1236 -3096 1242 -3090
rect 1236 -3102 1242 -3096
rect 1236 -3108 1242 -3102
rect 1236 -3114 1242 -3108
rect 1236 -3120 1242 -3114
rect 1236 -3126 1242 -3120
rect 1236 -3132 1242 -3126
rect 1236 -3138 1242 -3132
rect 1236 -3144 1242 -3138
rect 1236 -3150 1242 -3144
rect 1236 -3156 1242 -3150
rect 1236 -3162 1242 -3156
rect 1236 -3168 1242 -3162
rect 1236 -3174 1242 -3168
rect 1236 -3180 1242 -3174
rect 1236 -3186 1242 -3180
rect 1236 -3192 1242 -3186
rect 1236 -3198 1242 -3192
rect 1236 -3204 1242 -3198
rect 1236 -3210 1242 -3204
rect 1236 -3216 1242 -3210
rect 1236 -3222 1242 -3216
rect 1236 -3228 1242 -3222
rect 1236 -3234 1242 -3228
rect 1236 -3240 1242 -3234
rect 1236 -3324 1242 -3318
rect 1236 -3330 1242 -3324
rect 1236 -3336 1242 -3330
rect 1236 -3342 1242 -3336
rect 1236 -3348 1242 -3342
rect 1236 -3354 1242 -3348
rect 1236 -3360 1242 -3354
rect 1236 -3366 1242 -3360
rect 1236 -3372 1242 -3366
rect 1236 -3378 1242 -3372
rect 1236 -3384 1242 -3378
rect 1236 -3390 1242 -3384
rect 1236 -3396 1242 -3390
rect 1236 -3402 1242 -3396
rect 1236 -3408 1242 -3402
rect 1236 -3414 1242 -3408
rect 1236 -3420 1242 -3414
rect 1236 -3426 1242 -3420
rect 1236 -3432 1242 -3426
rect 1236 -3438 1242 -3432
rect 1236 -3444 1242 -3438
rect 1236 -3450 1242 -3444
rect 1236 -3456 1242 -3450
rect 1236 -3462 1242 -3456
rect 1236 -3468 1242 -3462
rect 1236 -3474 1242 -3468
rect 1236 -3480 1242 -3474
rect 1236 -3486 1242 -3480
rect 1236 -3492 1242 -3486
rect 1236 -3498 1242 -3492
rect 1236 -3504 1242 -3498
rect 1236 -3510 1242 -3504
rect 1236 -3516 1242 -3510
rect 1236 -3522 1242 -3516
rect 1242 -1104 1248 -1098
rect 1242 -1110 1248 -1104
rect 1242 -1116 1248 -1110
rect 1242 -1122 1248 -1116
rect 1242 -1128 1248 -1122
rect 1242 -1134 1248 -1128
rect 1242 -1140 1248 -1134
rect 1242 -1146 1248 -1140
rect 1242 -1152 1248 -1146
rect 1242 -1158 1248 -1152
rect 1242 -1164 1248 -1158
rect 1242 -1170 1248 -1164
rect 1242 -1176 1248 -1170
rect 1242 -1182 1248 -1176
rect 1242 -1188 1248 -1182
rect 1242 -1194 1248 -1188
rect 1242 -1200 1248 -1194
rect 1242 -1206 1248 -1200
rect 1242 -1212 1248 -1206
rect 1242 -1218 1248 -1212
rect 1242 -1224 1248 -1218
rect 1242 -1230 1248 -1224
rect 1242 -1236 1248 -1230
rect 1242 -1242 1248 -1236
rect 1242 -1248 1248 -1242
rect 1242 -1254 1248 -1248
rect 1242 -1260 1248 -1254
rect 1242 -1266 1248 -1260
rect 1242 -1272 1248 -1266
rect 1242 -1278 1248 -1272
rect 1242 -1284 1248 -1278
rect 1242 -1290 1248 -1284
rect 1242 -1296 1248 -1290
rect 1242 -1302 1248 -1296
rect 1242 -1308 1248 -1302
rect 1242 -1704 1248 -1698
rect 1242 -1710 1248 -1704
rect 1242 -1716 1248 -1710
rect 1242 -1722 1248 -1716
rect 1242 -1728 1248 -1722
rect 1242 -1734 1248 -1728
rect 1242 -1740 1248 -1734
rect 1242 -1746 1248 -1740
rect 1242 -1752 1248 -1746
rect 1242 -1758 1248 -1752
rect 1242 -1764 1248 -1758
rect 1242 -1770 1248 -1764
rect 1242 -1776 1248 -1770
rect 1242 -1782 1248 -1776
rect 1242 -1788 1248 -1782
rect 1242 -1794 1248 -1788
rect 1242 -1800 1248 -1794
rect 1242 -1806 1248 -1800
rect 1242 -1812 1248 -1806
rect 1242 -1818 1248 -1812
rect 1242 -1824 1248 -1818
rect 1242 -1830 1248 -1824
rect 1242 -1836 1248 -1830
rect 1242 -1842 1248 -1836
rect 1242 -1848 1248 -1842
rect 1242 -1854 1248 -1848
rect 1242 -1860 1248 -1854
rect 1242 -1866 1248 -1860
rect 1242 -1872 1248 -1866
rect 1242 -1878 1248 -1872
rect 1242 -1884 1248 -1878
rect 1242 -1890 1248 -1884
rect 1242 -1896 1248 -1890
rect 1242 -1902 1248 -1896
rect 1242 -1908 1248 -1902
rect 1242 -1914 1248 -1908
rect 1242 -1920 1248 -1914
rect 1242 -1926 1248 -1920
rect 1242 -1932 1248 -1926
rect 1242 -1938 1248 -1932
rect 1242 -1944 1248 -1938
rect 1242 -1950 1248 -1944
rect 1242 -1956 1248 -1950
rect 1242 -1962 1248 -1956
rect 1242 -1968 1248 -1962
rect 1242 -1974 1248 -1968
rect 1242 -1980 1248 -1974
rect 1242 -1986 1248 -1980
rect 1242 -1992 1248 -1986
rect 1242 -1998 1248 -1992
rect 1242 -2004 1248 -1998
rect 1242 -2010 1248 -2004
rect 1242 -2016 1248 -2010
rect 1242 -2022 1248 -2016
rect 1242 -2028 1248 -2022
rect 1242 -2034 1248 -2028
rect 1242 -2040 1248 -2034
rect 1242 -2046 1248 -2040
rect 1242 -2052 1248 -2046
rect 1242 -2058 1248 -2052
rect 1242 -2064 1248 -2058
rect 1242 -2070 1248 -2064
rect 1242 -2076 1248 -2070
rect 1242 -2082 1248 -2076
rect 1242 -2088 1248 -2082
rect 1242 -2094 1248 -2088
rect 1242 -2100 1248 -2094
rect 1242 -2106 1248 -2100
rect 1242 -2112 1248 -2106
rect 1242 -2118 1248 -2112
rect 1242 -2124 1248 -2118
rect 1242 -2130 1248 -2124
rect 1242 -2136 1248 -2130
rect 1242 -2142 1248 -2136
rect 1242 -2148 1248 -2142
rect 1242 -2154 1248 -2148
rect 1242 -2160 1248 -2154
rect 1242 -2166 1248 -2160
rect 1242 -2172 1248 -2166
rect 1242 -2178 1248 -2172
rect 1242 -2184 1248 -2178
rect 1242 -2190 1248 -2184
rect 1242 -2196 1248 -2190
rect 1242 -2202 1248 -2196
rect 1242 -2208 1248 -2202
rect 1242 -2214 1248 -2208
rect 1242 -2220 1248 -2214
rect 1242 -2226 1248 -2220
rect 1242 -2232 1248 -2226
rect 1242 -2238 1248 -2232
rect 1242 -2244 1248 -2238
rect 1242 -2250 1248 -2244
rect 1242 -2256 1248 -2250
rect 1242 -2262 1248 -2256
rect 1242 -2268 1248 -2262
rect 1242 -2274 1248 -2268
rect 1242 -2280 1248 -2274
rect 1242 -2286 1248 -2280
rect 1242 -2292 1248 -2286
rect 1242 -2298 1248 -2292
rect 1242 -2304 1248 -2298
rect 1242 -2310 1248 -2304
rect 1242 -2316 1248 -2310
rect 1242 -2322 1248 -2316
rect 1242 -2328 1248 -2322
rect 1242 -2334 1248 -2328
rect 1242 -2340 1248 -2334
rect 1242 -2346 1248 -2340
rect 1242 -2352 1248 -2346
rect 1242 -2358 1248 -2352
rect 1242 -2364 1248 -2358
rect 1242 -2370 1248 -2364
rect 1242 -2376 1248 -2370
rect 1242 -2382 1248 -2376
rect 1242 -2388 1248 -2382
rect 1242 -2394 1248 -2388
rect 1242 -2400 1248 -2394
rect 1242 -2406 1248 -2400
rect 1242 -2412 1248 -2406
rect 1242 -2418 1248 -2412
rect 1242 -2424 1248 -2418
rect 1242 -2430 1248 -2424
rect 1242 -2436 1248 -2430
rect 1242 -2442 1248 -2436
rect 1242 -2448 1248 -2442
rect 1242 -2454 1248 -2448
rect 1242 -2460 1248 -2454
rect 1242 -2466 1248 -2460
rect 1242 -2472 1248 -2466
rect 1242 -2478 1248 -2472
rect 1242 -2484 1248 -2478
rect 1242 -2490 1248 -2484
rect 1242 -2496 1248 -2490
rect 1242 -2502 1248 -2496
rect 1242 -2508 1248 -2502
rect 1242 -2514 1248 -2508
rect 1242 -2520 1248 -2514
rect 1242 -2526 1248 -2520
rect 1242 -2532 1248 -2526
rect 1242 -2538 1248 -2532
rect 1242 -2544 1248 -2538
rect 1242 -2634 1248 -2628
rect 1242 -2640 1248 -2634
rect 1242 -2646 1248 -2640
rect 1242 -2652 1248 -2646
rect 1242 -2658 1248 -2652
rect 1242 -2664 1248 -2658
rect 1242 -2670 1248 -2664
rect 1242 -2676 1248 -2670
rect 1242 -2682 1248 -2676
rect 1242 -2688 1248 -2682
rect 1242 -2694 1248 -2688
rect 1242 -2700 1248 -2694
rect 1242 -2706 1248 -2700
rect 1242 -2712 1248 -2706
rect 1242 -2718 1248 -2712
rect 1242 -2724 1248 -2718
rect 1242 -2730 1248 -2724
rect 1242 -2736 1248 -2730
rect 1242 -2742 1248 -2736
rect 1242 -2748 1248 -2742
rect 1242 -2754 1248 -2748
rect 1242 -2760 1248 -2754
rect 1242 -2766 1248 -2760
rect 1242 -2772 1248 -2766
rect 1242 -2778 1248 -2772
rect 1242 -2784 1248 -2778
rect 1242 -2790 1248 -2784
rect 1242 -2796 1248 -2790
rect 1242 -2802 1248 -2796
rect 1242 -2808 1248 -2802
rect 1242 -2814 1248 -2808
rect 1242 -2820 1248 -2814
rect 1242 -2826 1248 -2820
rect 1242 -2832 1248 -2826
rect 1242 -2838 1248 -2832
rect 1242 -2844 1248 -2838
rect 1242 -2850 1248 -2844
rect 1242 -2856 1248 -2850
rect 1242 -2862 1248 -2856
rect 1242 -2868 1248 -2862
rect 1242 -2874 1248 -2868
rect 1242 -2880 1248 -2874
rect 1242 -2886 1248 -2880
rect 1242 -2892 1248 -2886
rect 1242 -2898 1248 -2892
rect 1242 -2904 1248 -2898
rect 1242 -2910 1248 -2904
rect 1242 -2916 1248 -2910
rect 1242 -2922 1248 -2916
rect 1242 -2928 1248 -2922
rect 1242 -2934 1248 -2928
rect 1242 -2940 1248 -2934
rect 1242 -2946 1248 -2940
rect 1242 -2952 1248 -2946
rect 1242 -2958 1248 -2952
rect 1242 -2964 1248 -2958
rect 1242 -2970 1248 -2964
rect 1242 -2976 1248 -2970
rect 1242 -2982 1248 -2976
rect 1242 -2988 1248 -2982
rect 1242 -3066 1248 -3060
rect 1242 -3072 1248 -3066
rect 1242 -3078 1248 -3072
rect 1242 -3084 1248 -3078
rect 1242 -3090 1248 -3084
rect 1242 -3096 1248 -3090
rect 1242 -3102 1248 -3096
rect 1242 -3108 1248 -3102
rect 1242 -3114 1248 -3108
rect 1242 -3120 1248 -3114
rect 1242 -3126 1248 -3120
rect 1242 -3132 1248 -3126
rect 1242 -3138 1248 -3132
rect 1242 -3144 1248 -3138
rect 1242 -3150 1248 -3144
rect 1242 -3156 1248 -3150
rect 1242 -3162 1248 -3156
rect 1242 -3168 1248 -3162
rect 1242 -3174 1248 -3168
rect 1242 -3180 1248 -3174
rect 1242 -3186 1248 -3180
rect 1242 -3192 1248 -3186
rect 1242 -3198 1248 -3192
rect 1242 -3204 1248 -3198
rect 1242 -3210 1248 -3204
rect 1242 -3216 1248 -3210
rect 1242 -3222 1248 -3216
rect 1242 -3228 1248 -3222
rect 1242 -3234 1248 -3228
rect 1242 -3318 1248 -3312
rect 1242 -3324 1248 -3318
rect 1242 -3330 1248 -3324
rect 1242 -3336 1248 -3330
rect 1242 -3342 1248 -3336
rect 1242 -3348 1248 -3342
rect 1242 -3354 1248 -3348
rect 1242 -3360 1248 -3354
rect 1242 -3366 1248 -3360
rect 1242 -3372 1248 -3366
rect 1242 -3378 1248 -3372
rect 1242 -3384 1248 -3378
rect 1242 -3390 1248 -3384
rect 1242 -3396 1248 -3390
rect 1242 -3402 1248 -3396
rect 1242 -3408 1248 -3402
rect 1242 -3414 1248 -3408
rect 1242 -3420 1248 -3414
rect 1242 -3426 1248 -3420
rect 1242 -3432 1248 -3426
rect 1242 -3438 1248 -3432
rect 1242 -3444 1248 -3438
rect 1242 -3450 1248 -3444
rect 1242 -3456 1248 -3450
rect 1242 -3462 1248 -3456
rect 1242 -3468 1248 -3462
rect 1242 -3474 1248 -3468
rect 1242 -3480 1248 -3474
rect 1242 -3486 1248 -3480
rect 1242 -3492 1248 -3486
rect 1242 -3498 1248 -3492
rect 1242 -3504 1248 -3498
rect 1242 -3510 1248 -3504
rect 1242 -3516 1248 -3510
rect 1242 -3522 1248 -3516
rect 1248 -1104 1254 -1098
rect 1248 -1110 1254 -1104
rect 1248 -1116 1254 -1110
rect 1248 -1122 1254 -1116
rect 1248 -1128 1254 -1122
rect 1248 -1134 1254 -1128
rect 1248 -1140 1254 -1134
rect 1248 -1146 1254 -1140
rect 1248 -1152 1254 -1146
rect 1248 -1158 1254 -1152
rect 1248 -1164 1254 -1158
rect 1248 -1170 1254 -1164
rect 1248 -1176 1254 -1170
rect 1248 -1182 1254 -1176
rect 1248 -1188 1254 -1182
rect 1248 -1194 1254 -1188
rect 1248 -1200 1254 -1194
rect 1248 -1206 1254 -1200
rect 1248 -1212 1254 -1206
rect 1248 -1218 1254 -1212
rect 1248 -1224 1254 -1218
rect 1248 -1230 1254 -1224
rect 1248 -1236 1254 -1230
rect 1248 -1242 1254 -1236
rect 1248 -1248 1254 -1242
rect 1248 -1254 1254 -1248
rect 1248 -1260 1254 -1254
rect 1248 -1266 1254 -1260
rect 1248 -1272 1254 -1266
rect 1248 -1278 1254 -1272
rect 1248 -1284 1254 -1278
rect 1248 -1290 1254 -1284
rect 1248 -1296 1254 -1290
rect 1248 -1302 1254 -1296
rect 1248 -1308 1254 -1302
rect 1248 -1692 1254 -1686
rect 1248 -1698 1254 -1692
rect 1248 -1704 1254 -1698
rect 1248 -1710 1254 -1704
rect 1248 -1716 1254 -1710
rect 1248 -1722 1254 -1716
rect 1248 -1728 1254 -1722
rect 1248 -1734 1254 -1728
rect 1248 -1740 1254 -1734
rect 1248 -1746 1254 -1740
rect 1248 -1752 1254 -1746
rect 1248 -1758 1254 -1752
rect 1248 -1764 1254 -1758
rect 1248 -1770 1254 -1764
rect 1248 -1776 1254 -1770
rect 1248 -1782 1254 -1776
rect 1248 -1788 1254 -1782
rect 1248 -1794 1254 -1788
rect 1248 -1800 1254 -1794
rect 1248 -1806 1254 -1800
rect 1248 -1812 1254 -1806
rect 1248 -1818 1254 -1812
rect 1248 -1824 1254 -1818
rect 1248 -1830 1254 -1824
rect 1248 -1836 1254 -1830
rect 1248 -1842 1254 -1836
rect 1248 -1848 1254 -1842
rect 1248 -1854 1254 -1848
rect 1248 -1860 1254 -1854
rect 1248 -1866 1254 -1860
rect 1248 -1872 1254 -1866
rect 1248 -1878 1254 -1872
rect 1248 -1884 1254 -1878
rect 1248 -1890 1254 -1884
rect 1248 -1896 1254 -1890
rect 1248 -1902 1254 -1896
rect 1248 -1908 1254 -1902
rect 1248 -1914 1254 -1908
rect 1248 -1920 1254 -1914
rect 1248 -1926 1254 -1920
rect 1248 -1932 1254 -1926
rect 1248 -1938 1254 -1932
rect 1248 -1944 1254 -1938
rect 1248 -1950 1254 -1944
rect 1248 -1956 1254 -1950
rect 1248 -1962 1254 -1956
rect 1248 -1968 1254 -1962
rect 1248 -1974 1254 -1968
rect 1248 -1980 1254 -1974
rect 1248 -1986 1254 -1980
rect 1248 -1992 1254 -1986
rect 1248 -1998 1254 -1992
rect 1248 -2004 1254 -1998
rect 1248 -2010 1254 -2004
rect 1248 -2016 1254 -2010
rect 1248 -2022 1254 -2016
rect 1248 -2028 1254 -2022
rect 1248 -2034 1254 -2028
rect 1248 -2040 1254 -2034
rect 1248 -2046 1254 -2040
rect 1248 -2052 1254 -2046
rect 1248 -2058 1254 -2052
rect 1248 -2064 1254 -2058
rect 1248 -2070 1254 -2064
rect 1248 -2076 1254 -2070
rect 1248 -2082 1254 -2076
rect 1248 -2088 1254 -2082
rect 1248 -2094 1254 -2088
rect 1248 -2100 1254 -2094
rect 1248 -2106 1254 -2100
rect 1248 -2112 1254 -2106
rect 1248 -2118 1254 -2112
rect 1248 -2124 1254 -2118
rect 1248 -2130 1254 -2124
rect 1248 -2136 1254 -2130
rect 1248 -2142 1254 -2136
rect 1248 -2148 1254 -2142
rect 1248 -2154 1254 -2148
rect 1248 -2160 1254 -2154
rect 1248 -2166 1254 -2160
rect 1248 -2172 1254 -2166
rect 1248 -2178 1254 -2172
rect 1248 -2184 1254 -2178
rect 1248 -2190 1254 -2184
rect 1248 -2196 1254 -2190
rect 1248 -2202 1254 -2196
rect 1248 -2208 1254 -2202
rect 1248 -2214 1254 -2208
rect 1248 -2220 1254 -2214
rect 1248 -2226 1254 -2220
rect 1248 -2232 1254 -2226
rect 1248 -2238 1254 -2232
rect 1248 -2244 1254 -2238
rect 1248 -2250 1254 -2244
rect 1248 -2256 1254 -2250
rect 1248 -2262 1254 -2256
rect 1248 -2268 1254 -2262
rect 1248 -2274 1254 -2268
rect 1248 -2280 1254 -2274
rect 1248 -2286 1254 -2280
rect 1248 -2292 1254 -2286
rect 1248 -2298 1254 -2292
rect 1248 -2304 1254 -2298
rect 1248 -2310 1254 -2304
rect 1248 -2316 1254 -2310
rect 1248 -2322 1254 -2316
rect 1248 -2328 1254 -2322
rect 1248 -2334 1254 -2328
rect 1248 -2340 1254 -2334
rect 1248 -2346 1254 -2340
rect 1248 -2352 1254 -2346
rect 1248 -2358 1254 -2352
rect 1248 -2364 1254 -2358
rect 1248 -2370 1254 -2364
rect 1248 -2376 1254 -2370
rect 1248 -2382 1254 -2376
rect 1248 -2388 1254 -2382
rect 1248 -2394 1254 -2388
rect 1248 -2400 1254 -2394
rect 1248 -2406 1254 -2400
rect 1248 -2412 1254 -2406
rect 1248 -2418 1254 -2412
rect 1248 -2424 1254 -2418
rect 1248 -2430 1254 -2424
rect 1248 -2436 1254 -2430
rect 1248 -2442 1254 -2436
rect 1248 -2448 1254 -2442
rect 1248 -2454 1254 -2448
rect 1248 -2460 1254 -2454
rect 1248 -2466 1254 -2460
rect 1248 -2472 1254 -2466
rect 1248 -2478 1254 -2472
rect 1248 -2484 1254 -2478
rect 1248 -2490 1254 -2484
rect 1248 -2496 1254 -2490
rect 1248 -2502 1254 -2496
rect 1248 -2508 1254 -2502
rect 1248 -2514 1254 -2508
rect 1248 -2520 1254 -2514
rect 1248 -2526 1254 -2520
rect 1248 -2532 1254 -2526
rect 1248 -2622 1254 -2616
rect 1248 -2628 1254 -2622
rect 1248 -2634 1254 -2628
rect 1248 -2640 1254 -2634
rect 1248 -2646 1254 -2640
rect 1248 -2652 1254 -2646
rect 1248 -2658 1254 -2652
rect 1248 -2664 1254 -2658
rect 1248 -2670 1254 -2664
rect 1248 -2676 1254 -2670
rect 1248 -2682 1254 -2676
rect 1248 -2688 1254 -2682
rect 1248 -2694 1254 -2688
rect 1248 -2700 1254 -2694
rect 1248 -2706 1254 -2700
rect 1248 -2712 1254 -2706
rect 1248 -2718 1254 -2712
rect 1248 -2724 1254 -2718
rect 1248 -2730 1254 -2724
rect 1248 -2736 1254 -2730
rect 1248 -2742 1254 -2736
rect 1248 -2748 1254 -2742
rect 1248 -2754 1254 -2748
rect 1248 -2760 1254 -2754
rect 1248 -2766 1254 -2760
rect 1248 -2772 1254 -2766
rect 1248 -2778 1254 -2772
rect 1248 -2784 1254 -2778
rect 1248 -2790 1254 -2784
rect 1248 -2796 1254 -2790
rect 1248 -2802 1254 -2796
rect 1248 -2808 1254 -2802
rect 1248 -2814 1254 -2808
rect 1248 -2820 1254 -2814
rect 1248 -2826 1254 -2820
rect 1248 -2832 1254 -2826
rect 1248 -2838 1254 -2832
rect 1248 -2844 1254 -2838
rect 1248 -2850 1254 -2844
rect 1248 -2856 1254 -2850
rect 1248 -2862 1254 -2856
rect 1248 -2868 1254 -2862
rect 1248 -2874 1254 -2868
rect 1248 -2880 1254 -2874
rect 1248 -2886 1254 -2880
rect 1248 -2892 1254 -2886
rect 1248 -2898 1254 -2892
rect 1248 -2904 1254 -2898
rect 1248 -2910 1254 -2904
rect 1248 -2916 1254 -2910
rect 1248 -2922 1254 -2916
rect 1248 -2928 1254 -2922
rect 1248 -2934 1254 -2928
rect 1248 -2940 1254 -2934
rect 1248 -2946 1254 -2940
rect 1248 -2952 1254 -2946
rect 1248 -2958 1254 -2952
rect 1248 -2964 1254 -2958
rect 1248 -2970 1254 -2964
rect 1248 -2976 1254 -2970
rect 1248 -2982 1254 -2976
rect 1248 -3066 1254 -3060
rect 1248 -3072 1254 -3066
rect 1248 -3078 1254 -3072
rect 1248 -3084 1254 -3078
rect 1248 -3090 1254 -3084
rect 1248 -3096 1254 -3090
rect 1248 -3102 1254 -3096
rect 1248 -3108 1254 -3102
rect 1248 -3114 1254 -3108
rect 1248 -3120 1254 -3114
rect 1248 -3126 1254 -3120
rect 1248 -3132 1254 -3126
rect 1248 -3138 1254 -3132
rect 1248 -3144 1254 -3138
rect 1248 -3150 1254 -3144
rect 1248 -3156 1254 -3150
rect 1248 -3162 1254 -3156
rect 1248 -3168 1254 -3162
rect 1248 -3174 1254 -3168
rect 1248 -3180 1254 -3174
rect 1248 -3186 1254 -3180
rect 1248 -3192 1254 -3186
rect 1248 -3198 1254 -3192
rect 1248 -3204 1254 -3198
rect 1248 -3210 1254 -3204
rect 1248 -3216 1254 -3210
rect 1248 -3222 1254 -3216
rect 1248 -3228 1254 -3222
rect 1248 -3234 1254 -3228
rect 1248 -3318 1254 -3312
rect 1248 -3324 1254 -3318
rect 1248 -3330 1254 -3324
rect 1248 -3336 1254 -3330
rect 1248 -3342 1254 -3336
rect 1248 -3348 1254 -3342
rect 1248 -3354 1254 -3348
rect 1248 -3360 1254 -3354
rect 1248 -3366 1254 -3360
rect 1248 -3372 1254 -3366
rect 1248 -3378 1254 -3372
rect 1248 -3384 1254 -3378
rect 1248 -3390 1254 -3384
rect 1248 -3396 1254 -3390
rect 1248 -3402 1254 -3396
rect 1248 -3408 1254 -3402
rect 1248 -3414 1254 -3408
rect 1248 -3420 1254 -3414
rect 1248 -3426 1254 -3420
rect 1248 -3432 1254 -3426
rect 1248 -3438 1254 -3432
rect 1248 -3444 1254 -3438
rect 1248 -3450 1254 -3444
rect 1248 -3456 1254 -3450
rect 1248 -3462 1254 -3456
rect 1248 -3468 1254 -3462
rect 1248 -3474 1254 -3468
rect 1248 -3480 1254 -3474
rect 1248 -3486 1254 -3480
rect 1248 -3492 1254 -3486
rect 1248 -3498 1254 -3492
rect 1248 -3504 1254 -3498
rect 1248 -3510 1254 -3504
rect 1248 -3516 1254 -3510
rect 1248 -3522 1254 -3516
rect 1254 -1104 1260 -1098
rect 1254 -1110 1260 -1104
rect 1254 -1116 1260 -1110
rect 1254 -1122 1260 -1116
rect 1254 -1128 1260 -1122
rect 1254 -1134 1260 -1128
rect 1254 -1140 1260 -1134
rect 1254 -1146 1260 -1140
rect 1254 -1152 1260 -1146
rect 1254 -1158 1260 -1152
rect 1254 -1164 1260 -1158
rect 1254 -1170 1260 -1164
rect 1254 -1176 1260 -1170
rect 1254 -1182 1260 -1176
rect 1254 -1188 1260 -1182
rect 1254 -1194 1260 -1188
rect 1254 -1200 1260 -1194
rect 1254 -1206 1260 -1200
rect 1254 -1212 1260 -1206
rect 1254 -1218 1260 -1212
rect 1254 -1224 1260 -1218
rect 1254 -1230 1260 -1224
rect 1254 -1236 1260 -1230
rect 1254 -1242 1260 -1236
rect 1254 -1248 1260 -1242
rect 1254 -1254 1260 -1248
rect 1254 -1260 1260 -1254
rect 1254 -1266 1260 -1260
rect 1254 -1272 1260 -1266
rect 1254 -1278 1260 -1272
rect 1254 -1284 1260 -1278
rect 1254 -1290 1260 -1284
rect 1254 -1296 1260 -1290
rect 1254 -1302 1260 -1296
rect 1254 -1308 1260 -1302
rect 1254 -1680 1260 -1674
rect 1254 -1686 1260 -1680
rect 1254 -1692 1260 -1686
rect 1254 -1698 1260 -1692
rect 1254 -1704 1260 -1698
rect 1254 -1710 1260 -1704
rect 1254 -1716 1260 -1710
rect 1254 -1722 1260 -1716
rect 1254 -1728 1260 -1722
rect 1254 -1734 1260 -1728
rect 1254 -1740 1260 -1734
rect 1254 -1746 1260 -1740
rect 1254 -1752 1260 -1746
rect 1254 -1758 1260 -1752
rect 1254 -1764 1260 -1758
rect 1254 -1770 1260 -1764
rect 1254 -1776 1260 -1770
rect 1254 -1782 1260 -1776
rect 1254 -1788 1260 -1782
rect 1254 -1794 1260 -1788
rect 1254 -1800 1260 -1794
rect 1254 -1806 1260 -1800
rect 1254 -1812 1260 -1806
rect 1254 -1818 1260 -1812
rect 1254 -1824 1260 -1818
rect 1254 -1830 1260 -1824
rect 1254 -1836 1260 -1830
rect 1254 -1842 1260 -1836
rect 1254 -1848 1260 -1842
rect 1254 -1854 1260 -1848
rect 1254 -1860 1260 -1854
rect 1254 -1866 1260 -1860
rect 1254 -1872 1260 -1866
rect 1254 -1878 1260 -1872
rect 1254 -1884 1260 -1878
rect 1254 -1890 1260 -1884
rect 1254 -1896 1260 -1890
rect 1254 -1902 1260 -1896
rect 1254 -1908 1260 -1902
rect 1254 -1914 1260 -1908
rect 1254 -1920 1260 -1914
rect 1254 -1926 1260 -1920
rect 1254 -1932 1260 -1926
rect 1254 -1938 1260 -1932
rect 1254 -1944 1260 -1938
rect 1254 -1950 1260 -1944
rect 1254 -1956 1260 -1950
rect 1254 -1962 1260 -1956
rect 1254 -1968 1260 -1962
rect 1254 -1974 1260 -1968
rect 1254 -1980 1260 -1974
rect 1254 -1986 1260 -1980
rect 1254 -1992 1260 -1986
rect 1254 -1998 1260 -1992
rect 1254 -2004 1260 -1998
rect 1254 -2010 1260 -2004
rect 1254 -2016 1260 -2010
rect 1254 -2022 1260 -2016
rect 1254 -2028 1260 -2022
rect 1254 -2034 1260 -2028
rect 1254 -2040 1260 -2034
rect 1254 -2046 1260 -2040
rect 1254 -2052 1260 -2046
rect 1254 -2058 1260 -2052
rect 1254 -2064 1260 -2058
rect 1254 -2070 1260 -2064
rect 1254 -2076 1260 -2070
rect 1254 -2082 1260 -2076
rect 1254 -2088 1260 -2082
rect 1254 -2094 1260 -2088
rect 1254 -2100 1260 -2094
rect 1254 -2106 1260 -2100
rect 1254 -2112 1260 -2106
rect 1254 -2118 1260 -2112
rect 1254 -2124 1260 -2118
rect 1254 -2130 1260 -2124
rect 1254 -2136 1260 -2130
rect 1254 -2142 1260 -2136
rect 1254 -2148 1260 -2142
rect 1254 -2154 1260 -2148
rect 1254 -2160 1260 -2154
rect 1254 -2166 1260 -2160
rect 1254 -2172 1260 -2166
rect 1254 -2178 1260 -2172
rect 1254 -2184 1260 -2178
rect 1254 -2190 1260 -2184
rect 1254 -2196 1260 -2190
rect 1254 -2202 1260 -2196
rect 1254 -2208 1260 -2202
rect 1254 -2214 1260 -2208
rect 1254 -2220 1260 -2214
rect 1254 -2226 1260 -2220
rect 1254 -2232 1260 -2226
rect 1254 -2238 1260 -2232
rect 1254 -2244 1260 -2238
rect 1254 -2250 1260 -2244
rect 1254 -2256 1260 -2250
rect 1254 -2262 1260 -2256
rect 1254 -2268 1260 -2262
rect 1254 -2274 1260 -2268
rect 1254 -2280 1260 -2274
rect 1254 -2286 1260 -2280
rect 1254 -2292 1260 -2286
rect 1254 -2298 1260 -2292
rect 1254 -2304 1260 -2298
rect 1254 -2310 1260 -2304
rect 1254 -2316 1260 -2310
rect 1254 -2322 1260 -2316
rect 1254 -2328 1260 -2322
rect 1254 -2334 1260 -2328
rect 1254 -2340 1260 -2334
rect 1254 -2346 1260 -2340
rect 1254 -2352 1260 -2346
rect 1254 -2358 1260 -2352
rect 1254 -2364 1260 -2358
rect 1254 -2370 1260 -2364
rect 1254 -2376 1260 -2370
rect 1254 -2382 1260 -2376
rect 1254 -2388 1260 -2382
rect 1254 -2394 1260 -2388
rect 1254 -2400 1260 -2394
rect 1254 -2406 1260 -2400
rect 1254 -2412 1260 -2406
rect 1254 -2418 1260 -2412
rect 1254 -2424 1260 -2418
rect 1254 -2430 1260 -2424
rect 1254 -2436 1260 -2430
rect 1254 -2442 1260 -2436
rect 1254 -2448 1260 -2442
rect 1254 -2454 1260 -2448
rect 1254 -2460 1260 -2454
rect 1254 -2466 1260 -2460
rect 1254 -2472 1260 -2466
rect 1254 -2478 1260 -2472
rect 1254 -2484 1260 -2478
rect 1254 -2490 1260 -2484
rect 1254 -2496 1260 -2490
rect 1254 -2502 1260 -2496
rect 1254 -2508 1260 -2502
rect 1254 -2514 1260 -2508
rect 1254 -2520 1260 -2514
rect 1254 -2526 1260 -2520
rect 1254 -2616 1260 -2610
rect 1254 -2622 1260 -2616
rect 1254 -2628 1260 -2622
rect 1254 -2634 1260 -2628
rect 1254 -2640 1260 -2634
rect 1254 -2646 1260 -2640
rect 1254 -2652 1260 -2646
rect 1254 -2658 1260 -2652
rect 1254 -2664 1260 -2658
rect 1254 -2670 1260 -2664
rect 1254 -2676 1260 -2670
rect 1254 -2682 1260 -2676
rect 1254 -2688 1260 -2682
rect 1254 -2694 1260 -2688
rect 1254 -2700 1260 -2694
rect 1254 -2706 1260 -2700
rect 1254 -2712 1260 -2706
rect 1254 -2718 1260 -2712
rect 1254 -2724 1260 -2718
rect 1254 -2730 1260 -2724
rect 1254 -2736 1260 -2730
rect 1254 -2742 1260 -2736
rect 1254 -2748 1260 -2742
rect 1254 -2754 1260 -2748
rect 1254 -2760 1260 -2754
rect 1254 -2766 1260 -2760
rect 1254 -2772 1260 -2766
rect 1254 -2778 1260 -2772
rect 1254 -2784 1260 -2778
rect 1254 -2790 1260 -2784
rect 1254 -2796 1260 -2790
rect 1254 -2802 1260 -2796
rect 1254 -2808 1260 -2802
rect 1254 -2814 1260 -2808
rect 1254 -2820 1260 -2814
rect 1254 -2826 1260 -2820
rect 1254 -2832 1260 -2826
rect 1254 -2838 1260 -2832
rect 1254 -2844 1260 -2838
rect 1254 -2850 1260 -2844
rect 1254 -2856 1260 -2850
rect 1254 -2862 1260 -2856
rect 1254 -2868 1260 -2862
rect 1254 -2874 1260 -2868
rect 1254 -2880 1260 -2874
rect 1254 -2886 1260 -2880
rect 1254 -2892 1260 -2886
rect 1254 -2898 1260 -2892
rect 1254 -2904 1260 -2898
rect 1254 -2910 1260 -2904
rect 1254 -2916 1260 -2910
rect 1254 -2922 1260 -2916
rect 1254 -2928 1260 -2922
rect 1254 -2934 1260 -2928
rect 1254 -2940 1260 -2934
rect 1254 -2946 1260 -2940
rect 1254 -2952 1260 -2946
rect 1254 -2958 1260 -2952
rect 1254 -2964 1260 -2958
rect 1254 -2970 1260 -2964
rect 1254 -2976 1260 -2970
rect 1254 -3060 1260 -3054
rect 1254 -3066 1260 -3060
rect 1254 -3072 1260 -3066
rect 1254 -3078 1260 -3072
rect 1254 -3084 1260 -3078
rect 1254 -3090 1260 -3084
rect 1254 -3096 1260 -3090
rect 1254 -3102 1260 -3096
rect 1254 -3108 1260 -3102
rect 1254 -3114 1260 -3108
rect 1254 -3120 1260 -3114
rect 1254 -3126 1260 -3120
rect 1254 -3132 1260 -3126
rect 1254 -3138 1260 -3132
rect 1254 -3144 1260 -3138
rect 1254 -3150 1260 -3144
rect 1254 -3156 1260 -3150
rect 1254 -3162 1260 -3156
rect 1254 -3168 1260 -3162
rect 1254 -3174 1260 -3168
rect 1254 -3180 1260 -3174
rect 1254 -3186 1260 -3180
rect 1254 -3192 1260 -3186
rect 1254 -3198 1260 -3192
rect 1254 -3204 1260 -3198
rect 1254 -3210 1260 -3204
rect 1254 -3216 1260 -3210
rect 1254 -3222 1260 -3216
rect 1254 -3228 1260 -3222
rect 1254 -3234 1260 -3228
rect 1254 -3318 1260 -3312
rect 1254 -3324 1260 -3318
rect 1254 -3330 1260 -3324
rect 1254 -3336 1260 -3330
rect 1254 -3342 1260 -3336
rect 1254 -3348 1260 -3342
rect 1254 -3354 1260 -3348
rect 1254 -3360 1260 -3354
rect 1254 -3366 1260 -3360
rect 1254 -3372 1260 -3366
rect 1254 -3378 1260 -3372
rect 1254 -3384 1260 -3378
rect 1254 -3390 1260 -3384
rect 1254 -3396 1260 -3390
rect 1254 -3402 1260 -3396
rect 1254 -3408 1260 -3402
rect 1254 -3414 1260 -3408
rect 1254 -3420 1260 -3414
rect 1254 -3426 1260 -3420
rect 1254 -3432 1260 -3426
rect 1254 -3438 1260 -3432
rect 1254 -3444 1260 -3438
rect 1254 -3450 1260 -3444
rect 1254 -3456 1260 -3450
rect 1254 -3462 1260 -3456
rect 1254 -3468 1260 -3462
rect 1254 -3474 1260 -3468
rect 1254 -3480 1260 -3474
rect 1254 -3486 1260 -3480
rect 1254 -3492 1260 -3486
rect 1254 -3498 1260 -3492
rect 1254 -3504 1260 -3498
rect 1254 -3510 1260 -3504
rect 1254 -3516 1260 -3510
rect 1254 -3522 1260 -3516
rect 1260 -1104 1266 -1098
rect 1260 -1110 1266 -1104
rect 1260 -1116 1266 -1110
rect 1260 -1122 1266 -1116
rect 1260 -1128 1266 -1122
rect 1260 -1134 1266 -1128
rect 1260 -1140 1266 -1134
rect 1260 -1146 1266 -1140
rect 1260 -1152 1266 -1146
rect 1260 -1158 1266 -1152
rect 1260 -1164 1266 -1158
rect 1260 -1170 1266 -1164
rect 1260 -1176 1266 -1170
rect 1260 -1182 1266 -1176
rect 1260 -1188 1266 -1182
rect 1260 -1194 1266 -1188
rect 1260 -1200 1266 -1194
rect 1260 -1206 1266 -1200
rect 1260 -1212 1266 -1206
rect 1260 -1218 1266 -1212
rect 1260 -1224 1266 -1218
rect 1260 -1230 1266 -1224
rect 1260 -1236 1266 -1230
rect 1260 -1242 1266 -1236
rect 1260 -1248 1266 -1242
rect 1260 -1254 1266 -1248
rect 1260 -1260 1266 -1254
rect 1260 -1266 1266 -1260
rect 1260 -1272 1266 -1266
rect 1260 -1278 1266 -1272
rect 1260 -1284 1266 -1278
rect 1260 -1290 1266 -1284
rect 1260 -1296 1266 -1290
rect 1260 -1302 1266 -1296
rect 1260 -1308 1266 -1302
rect 1260 -1662 1266 -1656
rect 1260 -1668 1266 -1662
rect 1260 -1674 1266 -1668
rect 1260 -1680 1266 -1674
rect 1260 -1686 1266 -1680
rect 1260 -1692 1266 -1686
rect 1260 -1698 1266 -1692
rect 1260 -1704 1266 -1698
rect 1260 -1710 1266 -1704
rect 1260 -1716 1266 -1710
rect 1260 -1722 1266 -1716
rect 1260 -1728 1266 -1722
rect 1260 -1734 1266 -1728
rect 1260 -1740 1266 -1734
rect 1260 -1746 1266 -1740
rect 1260 -1752 1266 -1746
rect 1260 -1758 1266 -1752
rect 1260 -1764 1266 -1758
rect 1260 -1770 1266 -1764
rect 1260 -1776 1266 -1770
rect 1260 -1782 1266 -1776
rect 1260 -1788 1266 -1782
rect 1260 -1794 1266 -1788
rect 1260 -1800 1266 -1794
rect 1260 -1806 1266 -1800
rect 1260 -1812 1266 -1806
rect 1260 -1818 1266 -1812
rect 1260 -1824 1266 -1818
rect 1260 -1830 1266 -1824
rect 1260 -1836 1266 -1830
rect 1260 -1842 1266 -1836
rect 1260 -1848 1266 -1842
rect 1260 -1854 1266 -1848
rect 1260 -1860 1266 -1854
rect 1260 -1866 1266 -1860
rect 1260 -1872 1266 -1866
rect 1260 -1878 1266 -1872
rect 1260 -1884 1266 -1878
rect 1260 -1890 1266 -1884
rect 1260 -1896 1266 -1890
rect 1260 -1902 1266 -1896
rect 1260 -1908 1266 -1902
rect 1260 -1914 1266 -1908
rect 1260 -1920 1266 -1914
rect 1260 -1926 1266 -1920
rect 1260 -1932 1266 -1926
rect 1260 -1938 1266 -1932
rect 1260 -1944 1266 -1938
rect 1260 -1950 1266 -1944
rect 1260 -1956 1266 -1950
rect 1260 -1962 1266 -1956
rect 1260 -1968 1266 -1962
rect 1260 -1974 1266 -1968
rect 1260 -1980 1266 -1974
rect 1260 -1986 1266 -1980
rect 1260 -1992 1266 -1986
rect 1260 -1998 1266 -1992
rect 1260 -2004 1266 -1998
rect 1260 -2010 1266 -2004
rect 1260 -2016 1266 -2010
rect 1260 -2022 1266 -2016
rect 1260 -2028 1266 -2022
rect 1260 -2034 1266 -2028
rect 1260 -2040 1266 -2034
rect 1260 -2046 1266 -2040
rect 1260 -2052 1266 -2046
rect 1260 -2058 1266 -2052
rect 1260 -2064 1266 -2058
rect 1260 -2070 1266 -2064
rect 1260 -2076 1266 -2070
rect 1260 -2082 1266 -2076
rect 1260 -2088 1266 -2082
rect 1260 -2094 1266 -2088
rect 1260 -2100 1266 -2094
rect 1260 -2106 1266 -2100
rect 1260 -2112 1266 -2106
rect 1260 -2118 1266 -2112
rect 1260 -2124 1266 -2118
rect 1260 -2130 1266 -2124
rect 1260 -2136 1266 -2130
rect 1260 -2142 1266 -2136
rect 1260 -2148 1266 -2142
rect 1260 -2154 1266 -2148
rect 1260 -2160 1266 -2154
rect 1260 -2166 1266 -2160
rect 1260 -2172 1266 -2166
rect 1260 -2178 1266 -2172
rect 1260 -2184 1266 -2178
rect 1260 -2190 1266 -2184
rect 1260 -2196 1266 -2190
rect 1260 -2202 1266 -2196
rect 1260 -2208 1266 -2202
rect 1260 -2214 1266 -2208
rect 1260 -2220 1266 -2214
rect 1260 -2226 1266 -2220
rect 1260 -2232 1266 -2226
rect 1260 -2238 1266 -2232
rect 1260 -2244 1266 -2238
rect 1260 -2250 1266 -2244
rect 1260 -2256 1266 -2250
rect 1260 -2262 1266 -2256
rect 1260 -2268 1266 -2262
rect 1260 -2274 1266 -2268
rect 1260 -2280 1266 -2274
rect 1260 -2286 1266 -2280
rect 1260 -2292 1266 -2286
rect 1260 -2298 1266 -2292
rect 1260 -2304 1266 -2298
rect 1260 -2310 1266 -2304
rect 1260 -2316 1266 -2310
rect 1260 -2322 1266 -2316
rect 1260 -2328 1266 -2322
rect 1260 -2334 1266 -2328
rect 1260 -2340 1266 -2334
rect 1260 -2346 1266 -2340
rect 1260 -2352 1266 -2346
rect 1260 -2358 1266 -2352
rect 1260 -2364 1266 -2358
rect 1260 -2370 1266 -2364
rect 1260 -2376 1266 -2370
rect 1260 -2382 1266 -2376
rect 1260 -2388 1266 -2382
rect 1260 -2394 1266 -2388
rect 1260 -2400 1266 -2394
rect 1260 -2406 1266 -2400
rect 1260 -2412 1266 -2406
rect 1260 -2418 1266 -2412
rect 1260 -2424 1266 -2418
rect 1260 -2430 1266 -2424
rect 1260 -2436 1266 -2430
rect 1260 -2442 1266 -2436
rect 1260 -2448 1266 -2442
rect 1260 -2454 1266 -2448
rect 1260 -2460 1266 -2454
rect 1260 -2466 1266 -2460
rect 1260 -2472 1266 -2466
rect 1260 -2478 1266 -2472
rect 1260 -2484 1266 -2478
rect 1260 -2490 1266 -2484
rect 1260 -2496 1266 -2490
rect 1260 -2502 1266 -2496
rect 1260 -2508 1266 -2502
rect 1260 -2514 1266 -2508
rect 1260 -2604 1266 -2598
rect 1260 -2610 1266 -2604
rect 1260 -2616 1266 -2610
rect 1260 -2622 1266 -2616
rect 1260 -2628 1266 -2622
rect 1260 -2634 1266 -2628
rect 1260 -2640 1266 -2634
rect 1260 -2646 1266 -2640
rect 1260 -2652 1266 -2646
rect 1260 -2658 1266 -2652
rect 1260 -2664 1266 -2658
rect 1260 -2670 1266 -2664
rect 1260 -2676 1266 -2670
rect 1260 -2682 1266 -2676
rect 1260 -2688 1266 -2682
rect 1260 -2694 1266 -2688
rect 1260 -2700 1266 -2694
rect 1260 -2706 1266 -2700
rect 1260 -2712 1266 -2706
rect 1260 -2718 1266 -2712
rect 1260 -2724 1266 -2718
rect 1260 -2730 1266 -2724
rect 1260 -2736 1266 -2730
rect 1260 -2742 1266 -2736
rect 1260 -2748 1266 -2742
rect 1260 -2754 1266 -2748
rect 1260 -2760 1266 -2754
rect 1260 -2766 1266 -2760
rect 1260 -2772 1266 -2766
rect 1260 -2778 1266 -2772
rect 1260 -2784 1266 -2778
rect 1260 -2790 1266 -2784
rect 1260 -2796 1266 -2790
rect 1260 -2802 1266 -2796
rect 1260 -2808 1266 -2802
rect 1260 -2814 1266 -2808
rect 1260 -2820 1266 -2814
rect 1260 -2826 1266 -2820
rect 1260 -2832 1266 -2826
rect 1260 -2838 1266 -2832
rect 1260 -2844 1266 -2838
rect 1260 -2850 1266 -2844
rect 1260 -2856 1266 -2850
rect 1260 -2862 1266 -2856
rect 1260 -2868 1266 -2862
rect 1260 -2874 1266 -2868
rect 1260 -2880 1266 -2874
rect 1260 -2886 1266 -2880
rect 1260 -2892 1266 -2886
rect 1260 -2898 1266 -2892
rect 1260 -2904 1266 -2898
rect 1260 -2910 1266 -2904
rect 1260 -2916 1266 -2910
rect 1260 -2922 1266 -2916
rect 1260 -2928 1266 -2922
rect 1260 -2934 1266 -2928
rect 1260 -2940 1266 -2934
rect 1260 -2946 1266 -2940
rect 1260 -2952 1266 -2946
rect 1260 -2958 1266 -2952
rect 1260 -2964 1266 -2958
rect 1260 -2970 1266 -2964
rect 1260 -2976 1266 -2970
rect 1260 -3054 1266 -3048
rect 1260 -3060 1266 -3054
rect 1260 -3066 1266 -3060
rect 1260 -3072 1266 -3066
rect 1260 -3078 1266 -3072
rect 1260 -3084 1266 -3078
rect 1260 -3090 1266 -3084
rect 1260 -3096 1266 -3090
rect 1260 -3102 1266 -3096
rect 1260 -3108 1266 -3102
rect 1260 -3114 1266 -3108
rect 1260 -3120 1266 -3114
rect 1260 -3126 1266 -3120
rect 1260 -3132 1266 -3126
rect 1260 -3138 1266 -3132
rect 1260 -3144 1266 -3138
rect 1260 -3150 1266 -3144
rect 1260 -3156 1266 -3150
rect 1260 -3162 1266 -3156
rect 1260 -3168 1266 -3162
rect 1260 -3174 1266 -3168
rect 1260 -3180 1266 -3174
rect 1260 -3186 1266 -3180
rect 1260 -3192 1266 -3186
rect 1260 -3198 1266 -3192
rect 1260 -3204 1266 -3198
rect 1260 -3210 1266 -3204
rect 1260 -3216 1266 -3210
rect 1260 -3222 1266 -3216
rect 1260 -3228 1266 -3222
rect 1260 -3234 1266 -3228
rect 1260 -3318 1266 -3312
rect 1260 -3324 1266 -3318
rect 1260 -3330 1266 -3324
rect 1260 -3336 1266 -3330
rect 1260 -3342 1266 -3336
rect 1260 -3348 1266 -3342
rect 1260 -3354 1266 -3348
rect 1260 -3360 1266 -3354
rect 1260 -3366 1266 -3360
rect 1260 -3372 1266 -3366
rect 1260 -3378 1266 -3372
rect 1260 -3384 1266 -3378
rect 1260 -3390 1266 -3384
rect 1260 -3396 1266 -3390
rect 1260 -3402 1266 -3396
rect 1260 -3408 1266 -3402
rect 1260 -3414 1266 -3408
rect 1260 -3420 1266 -3414
rect 1260 -3426 1266 -3420
rect 1260 -3432 1266 -3426
rect 1260 -3438 1266 -3432
rect 1260 -3444 1266 -3438
rect 1260 -3450 1266 -3444
rect 1260 -3456 1266 -3450
rect 1260 -3462 1266 -3456
rect 1260 -3468 1266 -3462
rect 1260 -3474 1266 -3468
rect 1260 -3480 1266 -3474
rect 1260 -3486 1266 -3480
rect 1260 -3492 1266 -3486
rect 1260 -3498 1266 -3492
rect 1260 -3504 1266 -3498
rect 1260 -3510 1266 -3504
rect 1260 -3516 1266 -3510
rect 1260 -3522 1266 -3516
rect 1266 -1104 1272 -1098
rect 1266 -1110 1272 -1104
rect 1266 -1116 1272 -1110
rect 1266 -1122 1272 -1116
rect 1266 -1128 1272 -1122
rect 1266 -1134 1272 -1128
rect 1266 -1140 1272 -1134
rect 1266 -1146 1272 -1140
rect 1266 -1152 1272 -1146
rect 1266 -1158 1272 -1152
rect 1266 -1164 1272 -1158
rect 1266 -1170 1272 -1164
rect 1266 -1176 1272 -1170
rect 1266 -1182 1272 -1176
rect 1266 -1188 1272 -1182
rect 1266 -1194 1272 -1188
rect 1266 -1200 1272 -1194
rect 1266 -1206 1272 -1200
rect 1266 -1212 1272 -1206
rect 1266 -1218 1272 -1212
rect 1266 -1224 1272 -1218
rect 1266 -1230 1272 -1224
rect 1266 -1236 1272 -1230
rect 1266 -1242 1272 -1236
rect 1266 -1248 1272 -1242
rect 1266 -1254 1272 -1248
rect 1266 -1260 1272 -1254
rect 1266 -1266 1272 -1260
rect 1266 -1272 1272 -1266
rect 1266 -1278 1272 -1272
rect 1266 -1284 1272 -1278
rect 1266 -1290 1272 -1284
rect 1266 -1296 1272 -1290
rect 1266 -1302 1272 -1296
rect 1266 -1308 1272 -1302
rect 1266 -1650 1272 -1644
rect 1266 -1656 1272 -1650
rect 1266 -1662 1272 -1656
rect 1266 -1668 1272 -1662
rect 1266 -1674 1272 -1668
rect 1266 -1680 1272 -1674
rect 1266 -1686 1272 -1680
rect 1266 -1692 1272 -1686
rect 1266 -1698 1272 -1692
rect 1266 -1704 1272 -1698
rect 1266 -1710 1272 -1704
rect 1266 -1716 1272 -1710
rect 1266 -1722 1272 -1716
rect 1266 -1728 1272 -1722
rect 1266 -1734 1272 -1728
rect 1266 -1740 1272 -1734
rect 1266 -1746 1272 -1740
rect 1266 -1752 1272 -1746
rect 1266 -1758 1272 -1752
rect 1266 -1764 1272 -1758
rect 1266 -1770 1272 -1764
rect 1266 -1776 1272 -1770
rect 1266 -1782 1272 -1776
rect 1266 -1788 1272 -1782
rect 1266 -1794 1272 -1788
rect 1266 -1800 1272 -1794
rect 1266 -1806 1272 -1800
rect 1266 -1812 1272 -1806
rect 1266 -1818 1272 -1812
rect 1266 -1824 1272 -1818
rect 1266 -1830 1272 -1824
rect 1266 -1836 1272 -1830
rect 1266 -1842 1272 -1836
rect 1266 -1848 1272 -1842
rect 1266 -1854 1272 -1848
rect 1266 -1860 1272 -1854
rect 1266 -1866 1272 -1860
rect 1266 -1872 1272 -1866
rect 1266 -1878 1272 -1872
rect 1266 -1884 1272 -1878
rect 1266 -1890 1272 -1884
rect 1266 -1896 1272 -1890
rect 1266 -1902 1272 -1896
rect 1266 -1908 1272 -1902
rect 1266 -1914 1272 -1908
rect 1266 -1920 1272 -1914
rect 1266 -1926 1272 -1920
rect 1266 -1932 1272 -1926
rect 1266 -1938 1272 -1932
rect 1266 -1944 1272 -1938
rect 1266 -1950 1272 -1944
rect 1266 -1956 1272 -1950
rect 1266 -1962 1272 -1956
rect 1266 -1968 1272 -1962
rect 1266 -1974 1272 -1968
rect 1266 -1980 1272 -1974
rect 1266 -1986 1272 -1980
rect 1266 -1992 1272 -1986
rect 1266 -1998 1272 -1992
rect 1266 -2004 1272 -1998
rect 1266 -2010 1272 -2004
rect 1266 -2016 1272 -2010
rect 1266 -2022 1272 -2016
rect 1266 -2028 1272 -2022
rect 1266 -2034 1272 -2028
rect 1266 -2040 1272 -2034
rect 1266 -2046 1272 -2040
rect 1266 -2052 1272 -2046
rect 1266 -2058 1272 -2052
rect 1266 -2064 1272 -2058
rect 1266 -2070 1272 -2064
rect 1266 -2076 1272 -2070
rect 1266 -2082 1272 -2076
rect 1266 -2088 1272 -2082
rect 1266 -2094 1272 -2088
rect 1266 -2100 1272 -2094
rect 1266 -2106 1272 -2100
rect 1266 -2112 1272 -2106
rect 1266 -2118 1272 -2112
rect 1266 -2124 1272 -2118
rect 1266 -2130 1272 -2124
rect 1266 -2136 1272 -2130
rect 1266 -2142 1272 -2136
rect 1266 -2148 1272 -2142
rect 1266 -2154 1272 -2148
rect 1266 -2160 1272 -2154
rect 1266 -2166 1272 -2160
rect 1266 -2172 1272 -2166
rect 1266 -2178 1272 -2172
rect 1266 -2184 1272 -2178
rect 1266 -2190 1272 -2184
rect 1266 -2196 1272 -2190
rect 1266 -2202 1272 -2196
rect 1266 -2208 1272 -2202
rect 1266 -2214 1272 -2208
rect 1266 -2220 1272 -2214
rect 1266 -2226 1272 -2220
rect 1266 -2232 1272 -2226
rect 1266 -2238 1272 -2232
rect 1266 -2244 1272 -2238
rect 1266 -2250 1272 -2244
rect 1266 -2256 1272 -2250
rect 1266 -2262 1272 -2256
rect 1266 -2268 1272 -2262
rect 1266 -2274 1272 -2268
rect 1266 -2280 1272 -2274
rect 1266 -2286 1272 -2280
rect 1266 -2292 1272 -2286
rect 1266 -2298 1272 -2292
rect 1266 -2304 1272 -2298
rect 1266 -2310 1272 -2304
rect 1266 -2316 1272 -2310
rect 1266 -2322 1272 -2316
rect 1266 -2328 1272 -2322
rect 1266 -2334 1272 -2328
rect 1266 -2340 1272 -2334
rect 1266 -2346 1272 -2340
rect 1266 -2352 1272 -2346
rect 1266 -2358 1272 -2352
rect 1266 -2364 1272 -2358
rect 1266 -2370 1272 -2364
rect 1266 -2376 1272 -2370
rect 1266 -2382 1272 -2376
rect 1266 -2388 1272 -2382
rect 1266 -2394 1272 -2388
rect 1266 -2400 1272 -2394
rect 1266 -2406 1272 -2400
rect 1266 -2412 1272 -2406
rect 1266 -2418 1272 -2412
rect 1266 -2424 1272 -2418
rect 1266 -2430 1272 -2424
rect 1266 -2436 1272 -2430
rect 1266 -2442 1272 -2436
rect 1266 -2448 1272 -2442
rect 1266 -2454 1272 -2448
rect 1266 -2460 1272 -2454
rect 1266 -2466 1272 -2460
rect 1266 -2472 1272 -2466
rect 1266 -2478 1272 -2472
rect 1266 -2484 1272 -2478
rect 1266 -2490 1272 -2484
rect 1266 -2496 1272 -2490
rect 1266 -2502 1272 -2496
rect 1266 -2508 1272 -2502
rect 1266 -2598 1272 -2592
rect 1266 -2604 1272 -2598
rect 1266 -2610 1272 -2604
rect 1266 -2616 1272 -2610
rect 1266 -2622 1272 -2616
rect 1266 -2628 1272 -2622
rect 1266 -2634 1272 -2628
rect 1266 -2640 1272 -2634
rect 1266 -2646 1272 -2640
rect 1266 -2652 1272 -2646
rect 1266 -2658 1272 -2652
rect 1266 -2664 1272 -2658
rect 1266 -2670 1272 -2664
rect 1266 -2676 1272 -2670
rect 1266 -2682 1272 -2676
rect 1266 -2688 1272 -2682
rect 1266 -2694 1272 -2688
rect 1266 -2700 1272 -2694
rect 1266 -2706 1272 -2700
rect 1266 -2712 1272 -2706
rect 1266 -2718 1272 -2712
rect 1266 -2724 1272 -2718
rect 1266 -2730 1272 -2724
rect 1266 -2736 1272 -2730
rect 1266 -2742 1272 -2736
rect 1266 -2748 1272 -2742
rect 1266 -2754 1272 -2748
rect 1266 -2760 1272 -2754
rect 1266 -2766 1272 -2760
rect 1266 -2772 1272 -2766
rect 1266 -2778 1272 -2772
rect 1266 -2784 1272 -2778
rect 1266 -2790 1272 -2784
rect 1266 -2796 1272 -2790
rect 1266 -2802 1272 -2796
rect 1266 -2808 1272 -2802
rect 1266 -2814 1272 -2808
rect 1266 -2820 1272 -2814
rect 1266 -2826 1272 -2820
rect 1266 -2832 1272 -2826
rect 1266 -2838 1272 -2832
rect 1266 -2844 1272 -2838
rect 1266 -2850 1272 -2844
rect 1266 -2856 1272 -2850
rect 1266 -2862 1272 -2856
rect 1266 -2868 1272 -2862
rect 1266 -2874 1272 -2868
rect 1266 -2880 1272 -2874
rect 1266 -2886 1272 -2880
rect 1266 -2892 1272 -2886
rect 1266 -2898 1272 -2892
rect 1266 -2904 1272 -2898
rect 1266 -2910 1272 -2904
rect 1266 -2916 1272 -2910
rect 1266 -2922 1272 -2916
rect 1266 -2928 1272 -2922
rect 1266 -2934 1272 -2928
rect 1266 -2940 1272 -2934
rect 1266 -2946 1272 -2940
rect 1266 -2952 1272 -2946
rect 1266 -2958 1272 -2952
rect 1266 -2964 1272 -2958
rect 1266 -2970 1272 -2964
rect 1266 -3048 1272 -3042
rect 1266 -3054 1272 -3048
rect 1266 -3060 1272 -3054
rect 1266 -3066 1272 -3060
rect 1266 -3072 1272 -3066
rect 1266 -3078 1272 -3072
rect 1266 -3084 1272 -3078
rect 1266 -3090 1272 -3084
rect 1266 -3096 1272 -3090
rect 1266 -3102 1272 -3096
rect 1266 -3108 1272 -3102
rect 1266 -3114 1272 -3108
rect 1266 -3120 1272 -3114
rect 1266 -3126 1272 -3120
rect 1266 -3132 1272 -3126
rect 1266 -3138 1272 -3132
rect 1266 -3144 1272 -3138
rect 1266 -3150 1272 -3144
rect 1266 -3156 1272 -3150
rect 1266 -3162 1272 -3156
rect 1266 -3168 1272 -3162
rect 1266 -3174 1272 -3168
rect 1266 -3180 1272 -3174
rect 1266 -3186 1272 -3180
rect 1266 -3192 1272 -3186
rect 1266 -3198 1272 -3192
rect 1266 -3204 1272 -3198
rect 1266 -3210 1272 -3204
rect 1266 -3216 1272 -3210
rect 1266 -3222 1272 -3216
rect 1266 -3228 1272 -3222
rect 1266 -3234 1272 -3228
rect 1266 -3318 1272 -3312
rect 1266 -3324 1272 -3318
rect 1266 -3330 1272 -3324
rect 1266 -3336 1272 -3330
rect 1266 -3342 1272 -3336
rect 1266 -3348 1272 -3342
rect 1266 -3354 1272 -3348
rect 1266 -3360 1272 -3354
rect 1266 -3366 1272 -3360
rect 1266 -3372 1272 -3366
rect 1266 -3378 1272 -3372
rect 1266 -3384 1272 -3378
rect 1266 -3390 1272 -3384
rect 1266 -3396 1272 -3390
rect 1266 -3402 1272 -3396
rect 1266 -3408 1272 -3402
rect 1266 -3414 1272 -3408
rect 1266 -3420 1272 -3414
rect 1266 -3426 1272 -3420
rect 1266 -3432 1272 -3426
rect 1266 -3438 1272 -3432
rect 1266 -3444 1272 -3438
rect 1266 -3450 1272 -3444
rect 1266 -3456 1272 -3450
rect 1266 -3462 1272 -3456
rect 1266 -3468 1272 -3462
rect 1266 -3474 1272 -3468
rect 1266 -3480 1272 -3474
rect 1266 -3486 1272 -3480
rect 1266 -3492 1272 -3486
rect 1266 -3498 1272 -3492
rect 1266 -3504 1272 -3498
rect 1266 -3510 1272 -3504
rect 1266 -3516 1272 -3510
rect 1266 -3522 1272 -3516
rect 1272 -1104 1278 -1098
rect 1272 -1110 1278 -1104
rect 1272 -1116 1278 -1110
rect 1272 -1122 1278 -1116
rect 1272 -1128 1278 -1122
rect 1272 -1134 1278 -1128
rect 1272 -1140 1278 -1134
rect 1272 -1146 1278 -1140
rect 1272 -1152 1278 -1146
rect 1272 -1158 1278 -1152
rect 1272 -1164 1278 -1158
rect 1272 -1170 1278 -1164
rect 1272 -1176 1278 -1170
rect 1272 -1182 1278 -1176
rect 1272 -1188 1278 -1182
rect 1272 -1194 1278 -1188
rect 1272 -1200 1278 -1194
rect 1272 -1206 1278 -1200
rect 1272 -1212 1278 -1206
rect 1272 -1218 1278 -1212
rect 1272 -1224 1278 -1218
rect 1272 -1230 1278 -1224
rect 1272 -1236 1278 -1230
rect 1272 -1242 1278 -1236
rect 1272 -1248 1278 -1242
rect 1272 -1254 1278 -1248
rect 1272 -1260 1278 -1254
rect 1272 -1266 1278 -1260
rect 1272 -1272 1278 -1266
rect 1272 -1278 1278 -1272
rect 1272 -1284 1278 -1278
rect 1272 -1290 1278 -1284
rect 1272 -1296 1278 -1290
rect 1272 -1302 1278 -1296
rect 1272 -1308 1278 -1302
rect 1272 -1632 1278 -1626
rect 1272 -1638 1278 -1632
rect 1272 -1644 1278 -1638
rect 1272 -1650 1278 -1644
rect 1272 -1656 1278 -1650
rect 1272 -1662 1278 -1656
rect 1272 -1668 1278 -1662
rect 1272 -1674 1278 -1668
rect 1272 -1680 1278 -1674
rect 1272 -1686 1278 -1680
rect 1272 -1692 1278 -1686
rect 1272 -1698 1278 -1692
rect 1272 -1704 1278 -1698
rect 1272 -1710 1278 -1704
rect 1272 -1716 1278 -1710
rect 1272 -1722 1278 -1716
rect 1272 -1728 1278 -1722
rect 1272 -1734 1278 -1728
rect 1272 -1740 1278 -1734
rect 1272 -1746 1278 -1740
rect 1272 -1752 1278 -1746
rect 1272 -1758 1278 -1752
rect 1272 -1764 1278 -1758
rect 1272 -1770 1278 -1764
rect 1272 -1776 1278 -1770
rect 1272 -1782 1278 -1776
rect 1272 -1788 1278 -1782
rect 1272 -1794 1278 -1788
rect 1272 -1800 1278 -1794
rect 1272 -1806 1278 -1800
rect 1272 -1812 1278 -1806
rect 1272 -1818 1278 -1812
rect 1272 -1824 1278 -1818
rect 1272 -1830 1278 -1824
rect 1272 -1836 1278 -1830
rect 1272 -1842 1278 -1836
rect 1272 -1848 1278 -1842
rect 1272 -1854 1278 -1848
rect 1272 -1860 1278 -1854
rect 1272 -1866 1278 -1860
rect 1272 -1872 1278 -1866
rect 1272 -1878 1278 -1872
rect 1272 -1884 1278 -1878
rect 1272 -1890 1278 -1884
rect 1272 -1896 1278 -1890
rect 1272 -1902 1278 -1896
rect 1272 -1908 1278 -1902
rect 1272 -1914 1278 -1908
rect 1272 -1920 1278 -1914
rect 1272 -1926 1278 -1920
rect 1272 -1932 1278 -1926
rect 1272 -1938 1278 -1932
rect 1272 -1944 1278 -1938
rect 1272 -1950 1278 -1944
rect 1272 -1956 1278 -1950
rect 1272 -1962 1278 -1956
rect 1272 -1968 1278 -1962
rect 1272 -1974 1278 -1968
rect 1272 -1980 1278 -1974
rect 1272 -1986 1278 -1980
rect 1272 -1992 1278 -1986
rect 1272 -1998 1278 -1992
rect 1272 -2004 1278 -1998
rect 1272 -2010 1278 -2004
rect 1272 -2016 1278 -2010
rect 1272 -2022 1278 -2016
rect 1272 -2028 1278 -2022
rect 1272 -2034 1278 -2028
rect 1272 -2040 1278 -2034
rect 1272 -2046 1278 -2040
rect 1272 -2052 1278 -2046
rect 1272 -2058 1278 -2052
rect 1272 -2064 1278 -2058
rect 1272 -2070 1278 -2064
rect 1272 -2076 1278 -2070
rect 1272 -2082 1278 -2076
rect 1272 -2088 1278 -2082
rect 1272 -2094 1278 -2088
rect 1272 -2100 1278 -2094
rect 1272 -2106 1278 -2100
rect 1272 -2112 1278 -2106
rect 1272 -2118 1278 -2112
rect 1272 -2124 1278 -2118
rect 1272 -2130 1278 -2124
rect 1272 -2136 1278 -2130
rect 1272 -2142 1278 -2136
rect 1272 -2148 1278 -2142
rect 1272 -2154 1278 -2148
rect 1272 -2160 1278 -2154
rect 1272 -2166 1278 -2160
rect 1272 -2172 1278 -2166
rect 1272 -2178 1278 -2172
rect 1272 -2184 1278 -2178
rect 1272 -2190 1278 -2184
rect 1272 -2196 1278 -2190
rect 1272 -2202 1278 -2196
rect 1272 -2208 1278 -2202
rect 1272 -2214 1278 -2208
rect 1272 -2220 1278 -2214
rect 1272 -2226 1278 -2220
rect 1272 -2232 1278 -2226
rect 1272 -2238 1278 -2232
rect 1272 -2244 1278 -2238
rect 1272 -2250 1278 -2244
rect 1272 -2256 1278 -2250
rect 1272 -2262 1278 -2256
rect 1272 -2268 1278 -2262
rect 1272 -2274 1278 -2268
rect 1272 -2280 1278 -2274
rect 1272 -2286 1278 -2280
rect 1272 -2292 1278 -2286
rect 1272 -2298 1278 -2292
rect 1272 -2304 1278 -2298
rect 1272 -2310 1278 -2304
rect 1272 -2316 1278 -2310
rect 1272 -2322 1278 -2316
rect 1272 -2328 1278 -2322
rect 1272 -2334 1278 -2328
rect 1272 -2340 1278 -2334
rect 1272 -2346 1278 -2340
rect 1272 -2352 1278 -2346
rect 1272 -2358 1278 -2352
rect 1272 -2364 1278 -2358
rect 1272 -2370 1278 -2364
rect 1272 -2376 1278 -2370
rect 1272 -2382 1278 -2376
rect 1272 -2388 1278 -2382
rect 1272 -2394 1278 -2388
rect 1272 -2400 1278 -2394
rect 1272 -2406 1278 -2400
rect 1272 -2412 1278 -2406
rect 1272 -2418 1278 -2412
rect 1272 -2424 1278 -2418
rect 1272 -2430 1278 -2424
rect 1272 -2436 1278 -2430
rect 1272 -2442 1278 -2436
rect 1272 -2448 1278 -2442
rect 1272 -2454 1278 -2448
rect 1272 -2460 1278 -2454
rect 1272 -2466 1278 -2460
rect 1272 -2472 1278 -2466
rect 1272 -2478 1278 -2472
rect 1272 -2484 1278 -2478
rect 1272 -2490 1278 -2484
rect 1272 -2496 1278 -2490
rect 1272 -2502 1278 -2496
rect 1272 -2586 1278 -2580
rect 1272 -2592 1278 -2586
rect 1272 -2598 1278 -2592
rect 1272 -2604 1278 -2598
rect 1272 -2610 1278 -2604
rect 1272 -2616 1278 -2610
rect 1272 -2622 1278 -2616
rect 1272 -2628 1278 -2622
rect 1272 -2634 1278 -2628
rect 1272 -2640 1278 -2634
rect 1272 -2646 1278 -2640
rect 1272 -2652 1278 -2646
rect 1272 -2658 1278 -2652
rect 1272 -2664 1278 -2658
rect 1272 -2670 1278 -2664
rect 1272 -2676 1278 -2670
rect 1272 -2682 1278 -2676
rect 1272 -2688 1278 -2682
rect 1272 -2694 1278 -2688
rect 1272 -2700 1278 -2694
rect 1272 -2706 1278 -2700
rect 1272 -2712 1278 -2706
rect 1272 -2718 1278 -2712
rect 1272 -2724 1278 -2718
rect 1272 -2730 1278 -2724
rect 1272 -2736 1278 -2730
rect 1272 -2742 1278 -2736
rect 1272 -2748 1278 -2742
rect 1272 -2754 1278 -2748
rect 1272 -2760 1278 -2754
rect 1272 -2766 1278 -2760
rect 1272 -2772 1278 -2766
rect 1272 -2778 1278 -2772
rect 1272 -2784 1278 -2778
rect 1272 -2790 1278 -2784
rect 1272 -2796 1278 -2790
rect 1272 -2802 1278 -2796
rect 1272 -2808 1278 -2802
rect 1272 -2814 1278 -2808
rect 1272 -2820 1278 -2814
rect 1272 -2826 1278 -2820
rect 1272 -2832 1278 -2826
rect 1272 -2838 1278 -2832
rect 1272 -2844 1278 -2838
rect 1272 -2850 1278 -2844
rect 1272 -2856 1278 -2850
rect 1272 -2862 1278 -2856
rect 1272 -2868 1278 -2862
rect 1272 -2874 1278 -2868
rect 1272 -2880 1278 -2874
rect 1272 -2886 1278 -2880
rect 1272 -2892 1278 -2886
rect 1272 -2898 1278 -2892
rect 1272 -2904 1278 -2898
rect 1272 -2910 1278 -2904
rect 1272 -2916 1278 -2910
rect 1272 -2922 1278 -2916
rect 1272 -2928 1278 -2922
rect 1272 -2934 1278 -2928
rect 1272 -2940 1278 -2934
rect 1272 -2946 1278 -2940
rect 1272 -2952 1278 -2946
rect 1272 -2958 1278 -2952
rect 1272 -2964 1278 -2958
rect 1272 -3048 1278 -3042
rect 1272 -3054 1278 -3048
rect 1272 -3060 1278 -3054
rect 1272 -3066 1278 -3060
rect 1272 -3072 1278 -3066
rect 1272 -3078 1278 -3072
rect 1272 -3084 1278 -3078
rect 1272 -3090 1278 -3084
rect 1272 -3096 1278 -3090
rect 1272 -3102 1278 -3096
rect 1272 -3108 1278 -3102
rect 1272 -3114 1278 -3108
rect 1272 -3120 1278 -3114
rect 1272 -3126 1278 -3120
rect 1272 -3132 1278 -3126
rect 1272 -3138 1278 -3132
rect 1272 -3144 1278 -3138
rect 1272 -3150 1278 -3144
rect 1272 -3156 1278 -3150
rect 1272 -3162 1278 -3156
rect 1272 -3168 1278 -3162
rect 1272 -3174 1278 -3168
rect 1272 -3180 1278 -3174
rect 1272 -3186 1278 -3180
rect 1272 -3192 1278 -3186
rect 1272 -3198 1278 -3192
rect 1272 -3204 1278 -3198
rect 1272 -3210 1278 -3204
rect 1272 -3216 1278 -3210
rect 1272 -3222 1278 -3216
rect 1272 -3228 1278 -3222
rect 1272 -3234 1278 -3228
rect 1272 -3318 1278 -3312
rect 1272 -3324 1278 -3318
rect 1272 -3330 1278 -3324
rect 1272 -3336 1278 -3330
rect 1272 -3342 1278 -3336
rect 1272 -3348 1278 -3342
rect 1272 -3354 1278 -3348
rect 1272 -3360 1278 -3354
rect 1272 -3366 1278 -3360
rect 1272 -3372 1278 -3366
rect 1272 -3378 1278 -3372
rect 1272 -3384 1278 -3378
rect 1272 -3390 1278 -3384
rect 1272 -3396 1278 -3390
rect 1272 -3402 1278 -3396
rect 1272 -3408 1278 -3402
rect 1272 -3414 1278 -3408
rect 1272 -3420 1278 -3414
rect 1272 -3426 1278 -3420
rect 1272 -3432 1278 -3426
rect 1272 -3438 1278 -3432
rect 1272 -3444 1278 -3438
rect 1272 -3450 1278 -3444
rect 1272 -3456 1278 -3450
rect 1272 -3462 1278 -3456
rect 1272 -3468 1278 -3462
rect 1272 -3474 1278 -3468
rect 1272 -3480 1278 -3474
rect 1272 -3486 1278 -3480
rect 1272 -3492 1278 -3486
rect 1272 -3498 1278 -3492
rect 1272 -3504 1278 -3498
rect 1272 -3510 1278 -3504
rect 1272 -3516 1278 -3510
rect 1272 -3522 1278 -3516
rect 1278 -1104 1284 -1098
rect 1278 -1110 1284 -1104
rect 1278 -1116 1284 -1110
rect 1278 -1122 1284 -1116
rect 1278 -1128 1284 -1122
rect 1278 -1134 1284 -1128
rect 1278 -1140 1284 -1134
rect 1278 -1146 1284 -1140
rect 1278 -1152 1284 -1146
rect 1278 -1158 1284 -1152
rect 1278 -1164 1284 -1158
rect 1278 -1170 1284 -1164
rect 1278 -1176 1284 -1170
rect 1278 -1182 1284 -1176
rect 1278 -1188 1284 -1182
rect 1278 -1194 1284 -1188
rect 1278 -1200 1284 -1194
rect 1278 -1206 1284 -1200
rect 1278 -1212 1284 -1206
rect 1278 -1218 1284 -1212
rect 1278 -1224 1284 -1218
rect 1278 -1230 1284 -1224
rect 1278 -1236 1284 -1230
rect 1278 -1242 1284 -1236
rect 1278 -1248 1284 -1242
rect 1278 -1254 1284 -1248
rect 1278 -1260 1284 -1254
rect 1278 -1266 1284 -1260
rect 1278 -1272 1284 -1266
rect 1278 -1278 1284 -1272
rect 1278 -1284 1284 -1278
rect 1278 -1290 1284 -1284
rect 1278 -1296 1284 -1290
rect 1278 -1302 1284 -1296
rect 1278 -1308 1284 -1302
rect 1278 -1620 1284 -1614
rect 1278 -1626 1284 -1620
rect 1278 -1632 1284 -1626
rect 1278 -1638 1284 -1632
rect 1278 -1644 1284 -1638
rect 1278 -1650 1284 -1644
rect 1278 -1656 1284 -1650
rect 1278 -1662 1284 -1656
rect 1278 -1668 1284 -1662
rect 1278 -1674 1284 -1668
rect 1278 -1680 1284 -1674
rect 1278 -1686 1284 -1680
rect 1278 -1692 1284 -1686
rect 1278 -1698 1284 -1692
rect 1278 -1704 1284 -1698
rect 1278 -1710 1284 -1704
rect 1278 -1716 1284 -1710
rect 1278 -1722 1284 -1716
rect 1278 -1728 1284 -1722
rect 1278 -1734 1284 -1728
rect 1278 -1740 1284 -1734
rect 1278 -1746 1284 -1740
rect 1278 -1752 1284 -1746
rect 1278 -1758 1284 -1752
rect 1278 -1764 1284 -1758
rect 1278 -1770 1284 -1764
rect 1278 -1776 1284 -1770
rect 1278 -1782 1284 -1776
rect 1278 -1788 1284 -1782
rect 1278 -1794 1284 -1788
rect 1278 -1800 1284 -1794
rect 1278 -1806 1284 -1800
rect 1278 -1812 1284 -1806
rect 1278 -1818 1284 -1812
rect 1278 -1824 1284 -1818
rect 1278 -1830 1284 -1824
rect 1278 -1836 1284 -1830
rect 1278 -1842 1284 -1836
rect 1278 -1848 1284 -1842
rect 1278 -1854 1284 -1848
rect 1278 -1860 1284 -1854
rect 1278 -1866 1284 -1860
rect 1278 -1872 1284 -1866
rect 1278 -1878 1284 -1872
rect 1278 -1884 1284 -1878
rect 1278 -1890 1284 -1884
rect 1278 -1896 1284 -1890
rect 1278 -1902 1284 -1896
rect 1278 -1908 1284 -1902
rect 1278 -1914 1284 -1908
rect 1278 -1920 1284 -1914
rect 1278 -1926 1284 -1920
rect 1278 -1932 1284 -1926
rect 1278 -1938 1284 -1932
rect 1278 -1944 1284 -1938
rect 1278 -1950 1284 -1944
rect 1278 -1956 1284 -1950
rect 1278 -1962 1284 -1956
rect 1278 -1968 1284 -1962
rect 1278 -1974 1284 -1968
rect 1278 -1980 1284 -1974
rect 1278 -1986 1284 -1980
rect 1278 -1992 1284 -1986
rect 1278 -1998 1284 -1992
rect 1278 -2004 1284 -1998
rect 1278 -2010 1284 -2004
rect 1278 -2016 1284 -2010
rect 1278 -2022 1284 -2016
rect 1278 -2028 1284 -2022
rect 1278 -2034 1284 -2028
rect 1278 -2040 1284 -2034
rect 1278 -2046 1284 -2040
rect 1278 -2052 1284 -2046
rect 1278 -2058 1284 -2052
rect 1278 -2064 1284 -2058
rect 1278 -2070 1284 -2064
rect 1278 -2076 1284 -2070
rect 1278 -2082 1284 -2076
rect 1278 -2088 1284 -2082
rect 1278 -2094 1284 -2088
rect 1278 -2100 1284 -2094
rect 1278 -2106 1284 -2100
rect 1278 -2112 1284 -2106
rect 1278 -2118 1284 -2112
rect 1278 -2124 1284 -2118
rect 1278 -2130 1284 -2124
rect 1278 -2136 1284 -2130
rect 1278 -2142 1284 -2136
rect 1278 -2148 1284 -2142
rect 1278 -2154 1284 -2148
rect 1278 -2160 1284 -2154
rect 1278 -2166 1284 -2160
rect 1278 -2172 1284 -2166
rect 1278 -2178 1284 -2172
rect 1278 -2184 1284 -2178
rect 1278 -2190 1284 -2184
rect 1278 -2196 1284 -2190
rect 1278 -2202 1284 -2196
rect 1278 -2208 1284 -2202
rect 1278 -2214 1284 -2208
rect 1278 -2220 1284 -2214
rect 1278 -2226 1284 -2220
rect 1278 -2232 1284 -2226
rect 1278 -2238 1284 -2232
rect 1278 -2244 1284 -2238
rect 1278 -2250 1284 -2244
rect 1278 -2256 1284 -2250
rect 1278 -2262 1284 -2256
rect 1278 -2268 1284 -2262
rect 1278 -2274 1284 -2268
rect 1278 -2280 1284 -2274
rect 1278 -2286 1284 -2280
rect 1278 -2292 1284 -2286
rect 1278 -2298 1284 -2292
rect 1278 -2304 1284 -2298
rect 1278 -2310 1284 -2304
rect 1278 -2316 1284 -2310
rect 1278 -2322 1284 -2316
rect 1278 -2328 1284 -2322
rect 1278 -2334 1284 -2328
rect 1278 -2340 1284 -2334
rect 1278 -2346 1284 -2340
rect 1278 -2352 1284 -2346
rect 1278 -2358 1284 -2352
rect 1278 -2364 1284 -2358
rect 1278 -2370 1284 -2364
rect 1278 -2376 1284 -2370
rect 1278 -2382 1284 -2376
rect 1278 -2388 1284 -2382
rect 1278 -2394 1284 -2388
rect 1278 -2400 1284 -2394
rect 1278 -2406 1284 -2400
rect 1278 -2412 1284 -2406
rect 1278 -2418 1284 -2412
rect 1278 -2424 1284 -2418
rect 1278 -2430 1284 -2424
rect 1278 -2436 1284 -2430
rect 1278 -2442 1284 -2436
rect 1278 -2448 1284 -2442
rect 1278 -2454 1284 -2448
rect 1278 -2460 1284 -2454
rect 1278 -2466 1284 -2460
rect 1278 -2472 1284 -2466
rect 1278 -2478 1284 -2472
rect 1278 -2484 1284 -2478
rect 1278 -2490 1284 -2484
rect 1278 -2580 1284 -2574
rect 1278 -2586 1284 -2580
rect 1278 -2592 1284 -2586
rect 1278 -2598 1284 -2592
rect 1278 -2604 1284 -2598
rect 1278 -2610 1284 -2604
rect 1278 -2616 1284 -2610
rect 1278 -2622 1284 -2616
rect 1278 -2628 1284 -2622
rect 1278 -2634 1284 -2628
rect 1278 -2640 1284 -2634
rect 1278 -2646 1284 -2640
rect 1278 -2652 1284 -2646
rect 1278 -2658 1284 -2652
rect 1278 -2664 1284 -2658
rect 1278 -2670 1284 -2664
rect 1278 -2676 1284 -2670
rect 1278 -2682 1284 -2676
rect 1278 -2688 1284 -2682
rect 1278 -2694 1284 -2688
rect 1278 -2700 1284 -2694
rect 1278 -2706 1284 -2700
rect 1278 -2712 1284 -2706
rect 1278 -2718 1284 -2712
rect 1278 -2724 1284 -2718
rect 1278 -2730 1284 -2724
rect 1278 -2736 1284 -2730
rect 1278 -2742 1284 -2736
rect 1278 -2748 1284 -2742
rect 1278 -2754 1284 -2748
rect 1278 -2760 1284 -2754
rect 1278 -2766 1284 -2760
rect 1278 -2772 1284 -2766
rect 1278 -2778 1284 -2772
rect 1278 -2784 1284 -2778
rect 1278 -2790 1284 -2784
rect 1278 -2796 1284 -2790
rect 1278 -2802 1284 -2796
rect 1278 -2808 1284 -2802
rect 1278 -2814 1284 -2808
rect 1278 -2820 1284 -2814
rect 1278 -2826 1284 -2820
rect 1278 -2832 1284 -2826
rect 1278 -2838 1284 -2832
rect 1278 -2844 1284 -2838
rect 1278 -2850 1284 -2844
rect 1278 -2856 1284 -2850
rect 1278 -2862 1284 -2856
rect 1278 -2868 1284 -2862
rect 1278 -2874 1284 -2868
rect 1278 -2880 1284 -2874
rect 1278 -2886 1284 -2880
rect 1278 -2892 1284 -2886
rect 1278 -2898 1284 -2892
rect 1278 -2904 1284 -2898
rect 1278 -2910 1284 -2904
rect 1278 -2916 1284 -2910
rect 1278 -2922 1284 -2916
rect 1278 -2928 1284 -2922
rect 1278 -2934 1284 -2928
rect 1278 -2940 1284 -2934
rect 1278 -2946 1284 -2940
rect 1278 -2952 1284 -2946
rect 1278 -2958 1284 -2952
rect 1278 -3042 1284 -3036
rect 1278 -3048 1284 -3042
rect 1278 -3054 1284 -3048
rect 1278 -3060 1284 -3054
rect 1278 -3066 1284 -3060
rect 1278 -3072 1284 -3066
rect 1278 -3078 1284 -3072
rect 1278 -3084 1284 -3078
rect 1278 -3090 1284 -3084
rect 1278 -3096 1284 -3090
rect 1278 -3102 1284 -3096
rect 1278 -3108 1284 -3102
rect 1278 -3114 1284 -3108
rect 1278 -3120 1284 -3114
rect 1278 -3126 1284 -3120
rect 1278 -3132 1284 -3126
rect 1278 -3138 1284 -3132
rect 1278 -3144 1284 -3138
rect 1278 -3150 1284 -3144
rect 1278 -3156 1284 -3150
rect 1278 -3162 1284 -3156
rect 1278 -3168 1284 -3162
rect 1278 -3174 1284 -3168
rect 1278 -3180 1284 -3174
rect 1278 -3186 1284 -3180
rect 1278 -3192 1284 -3186
rect 1278 -3198 1284 -3192
rect 1278 -3204 1284 -3198
rect 1278 -3210 1284 -3204
rect 1278 -3216 1284 -3210
rect 1278 -3222 1284 -3216
rect 1278 -3228 1284 -3222
rect 1278 -3234 1284 -3228
rect 1278 -3318 1284 -3312
rect 1278 -3324 1284 -3318
rect 1278 -3330 1284 -3324
rect 1278 -3336 1284 -3330
rect 1278 -3342 1284 -3336
rect 1278 -3348 1284 -3342
rect 1278 -3354 1284 -3348
rect 1278 -3360 1284 -3354
rect 1278 -3366 1284 -3360
rect 1278 -3372 1284 -3366
rect 1278 -3378 1284 -3372
rect 1278 -3384 1284 -3378
rect 1278 -3390 1284 -3384
rect 1278 -3396 1284 -3390
rect 1278 -3402 1284 -3396
rect 1278 -3408 1284 -3402
rect 1278 -3414 1284 -3408
rect 1278 -3420 1284 -3414
rect 1278 -3426 1284 -3420
rect 1278 -3432 1284 -3426
rect 1278 -3438 1284 -3432
rect 1278 -3444 1284 -3438
rect 1278 -3450 1284 -3444
rect 1278 -3456 1284 -3450
rect 1278 -3462 1284 -3456
rect 1278 -3468 1284 -3462
rect 1278 -3474 1284 -3468
rect 1278 -3480 1284 -3474
rect 1278 -3486 1284 -3480
rect 1278 -3492 1284 -3486
rect 1278 -3498 1284 -3492
rect 1278 -3504 1284 -3498
rect 1278 -3510 1284 -3504
rect 1278 -3516 1284 -3510
rect 1278 -3522 1284 -3516
rect 1284 -1104 1290 -1098
rect 1284 -1110 1290 -1104
rect 1284 -1116 1290 -1110
rect 1284 -1122 1290 -1116
rect 1284 -1128 1290 -1122
rect 1284 -1134 1290 -1128
rect 1284 -1140 1290 -1134
rect 1284 -1146 1290 -1140
rect 1284 -1152 1290 -1146
rect 1284 -1158 1290 -1152
rect 1284 -1164 1290 -1158
rect 1284 -1170 1290 -1164
rect 1284 -1176 1290 -1170
rect 1284 -1182 1290 -1176
rect 1284 -1188 1290 -1182
rect 1284 -1194 1290 -1188
rect 1284 -1200 1290 -1194
rect 1284 -1206 1290 -1200
rect 1284 -1212 1290 -1206
rect 1284 -1218 1290 -1212
rect 1284 -1224 1290 -1218
rect 1284 -1230 1290 -1224
rect 1284 -1236 1290 -1230
rect 1284 -1242 1290 -1236
rect 1284 -1248 1290 -1242
rect 1284 -1254 1290 -1248
rect 1284 -1260 1290 -1254
rect 1284 -1266 1290 -1260
rect 1284 -1272 1290 -1266
rect 1284 -1278 1290 -1272
rect 1284 -1284 1290 -1278
rect 1284 -1290 1290 -1284
rect 1284 -1296 1290 -1290
rect 1284 -1302 1290 -1296
rect 1284 -1308 1290 -1302
rect 1284 -1608 1290 -1602
rect 1284 -1614 1290 -1608
rect 1284 -1620 1290 -1614
rect 1284 -1626 1290 -1620
rect 1284 -1632 1290 -1626
rect 1284 -1638 1290 -1632
rect 1284 -1644 1290 -1638
rect 1284 -1650 1290 -1644
rect 1284 -1656 1290 -1650
rect 1284 -1662 1290 -1656
rect 1284 -1668 1290 -1662
rect 1284 -1674 1290 -1668
rect 1284 -1680 1290 -1674
rect 1284 -1686 1290 -1680
rect 1284 -1692 1290 -1686
rect 1284 -1698 1290 -1692
rect 1284 -1704 1290 -1698
rect 1284 -1710 1290 -1704
rect 1284 -1716 1290 -1710
rect 1284 -1722 1290 -1716
rect 1284 -1728 1290 -1722
rect 1284 -1734 1290 -1728
rect 1284 -1740 1290 -1734
rect 1284 -1746 1290 -1740
rect 1284 -1752 1290 -1746
rect 1284 -1758 1290 -1752
rect 1284 -1764 1290 -1758
rect 1284 -1770 1290 -1764
rect 1284 -1776 1290 -1770
rect 1284 -1782 1290 -1776
rect 1284 -1788 1290 -1782
rect 1284 -1794 1290 -1788
rect 1284 -1800 1290 -1794
rect 1284 -1806 1290 -1800
rect 1284 -1812 1290 -1806
rect 1284 -1818 1290 -1812
rect 1284 -1824 1290 -1818
rect 1284 -1830 1290 -1824
rect 1284 -1836 1290 -1830
rect 1284 -1842 1290 -1836
rect 1284 -1848 1290 -1842
rect 1284 -1854 1290 -1848
rect 1284 -1860 1290 -1854
rect 1284 -1866 1290 -1860
rect 1284 -1872 1290 -1866
rect 1284 -1878 1290 -1872
rect 1284 -1884 1290 -1878
rect 1284 -1890 1290 -1884
rect 1284 -1896 1290 -1890
rect 1284 -1902 1290 -1896
rect 1284 -1908 1290 -1902
rect 1284 -1914 1290 -1908
rect 1284 -1920 1290 -1914
rect 1284 -1926 1290 -1920
rect 1284 -1932 1290 -1926
rect 1284 -1938 1290 -1932
rect 1284 -1944 1290 -1938
rect 1284 -1950 1290 -1944
rect 1284 -1956 1290 -1950
rect 1284 -1962 1290 -1956
rect 1284 -1968 1290 -1962
rect 1284 -1974 1290 -1968
rect 1284 -1980 1290 -1974
rect 1284 -1986 1290 -1980
rect 1284 -1992 1290 -1986
rect 1284 -1998 1290 -1992
rect 1284 -2004 1290 -1998
rect 1284 -2010 1290 -2004
rect 1284 -2016 1290 -2010
rect 1284 -2022 1290 -2016
rect 1284 -2028 1290 -2022
rect 1284 -2034 1290 -2028
rect 1284 -2040 1290 -2034
rect 1284 -2046 1290 -2040
rect 1284 -2052 1290 -2046
rect 1284 -2058 1290 -2052
rect 1284 -2064 1290 -2058
rect 1284 -2070 1290 -2064
rect 1284 -2076 1290 -2070
rect 1284 -2082 1290 -2076
rect 1284 -2088 1290 -2082
rect 1284 -2094 1290 -2088
rect 1284 -2100 1290 -2094
rect 1284 -2106 1290 -2100
rect 1284 -2112 1290 -2106
rect 1284 -2118 1290 -2112
rect 1284 -2124 1290 -2118
rect 1284 -2130 1290 -2124
rect 1284 -2136 1290 -2130
rect 1284 -2142 1290 -2136
rect 1284 -2148 1290 -2142
rect 1284 -2154 1290 -2148
rect 1284 -2160 1290 -2154
rect 1284 -2166 1290 -2160
rect 1284 -2172 1290 -2166
rect 1284 -2178 1290 -2172
rect 1284 -2184 1290 -2178
rect 1284 -2190 1290 -2184
rect 1284 -2196 1290 -2190
rect 1284 -2202 1290 -2196
rect 1284 -2208 1290 -2202
rect 1284 -2214 1290 -2208
rect 1284 -2220 1290 -2214
rect 1284 -2226 1290 -2220
rect 1284 -2232 1290 -2226
rect 1284 -2238 1290 -2232
rect 1284 -2244 1290 -2238
rect 1284 -2250 1290 -2244
rect 1284 -2256 1290 -2250
rect 1284 -2262 1290 -2256
rect 1284 -2268 1290 -2262
rect 1284 -2274 1290 -2268
rect 1284 -2280 1290 -2274
rect 1284 -2286 1290 -2280
rect 1284 -2292 1290 -2286
rect 1284 -2298 1290 -2292
rect 1284 -2304 1290 -2298
rect 1284 -2310 1290 -2304
rect 1284 -2316 1290 -2310
rect 1284 -2322 1290 -2316
rect 1284 -2328 1290 -2322
rect 1284 -2334 1290 -2328
rect 1284 -2340 1290 -2334
rect 1284 -2346 1290 -2340
rect 1284 -2352 1290 -2346
rect 1284 -2358 1290 -2352
rect 1284 -2364 1290 -2358
rect 1284 -2370 1290 -2364
rect 1284 -2376 1290 -2370
rect 1284 -2382 1290 -2376
rect 1284 -2388 1290 -2382
rect 1284 -2394 1290 -2388
rect 1284 -2400 1290 -2394
rect 1284 -2406 1290 -2400
rect 1284 -2412 1290 -2406
rect 1284 -2418 1290 -2412
rect 1284 -2424 1290 -2418
rect 1284 -2430 1290 -2424
rect 1284 -2436 1290 -2430
rect 1284 -2442 1290 -2436
rect 1284 -2448 1290 -2442
rect 1284 -2454 1290 -2448
rect 1284 -2460 1290 -2454
rect 1284 -2466 1290 -2460
rect 1284 -2472 1290 -2466
rect 1284 -2478 1290 -2472
rect 1284 -2484 1290 -2478
rect 1284 -2568 1290 -2562
rect 1284 -2574 1290 -2568
rect 1284 -2580 1290 -2574
rect 1284 -2586 1290 -2580
rect 1284 -2592 1290 -2586
rect 1284 -2598 1290 -2592
rect 1284 -2604 1290 -2598
rect 1284 -2610 1290 -2604
rect 1284 -2616 1290 -2610
rect 1284 -2622 1290 -2616
rect 1284 -2628 1290 -2622
rect 1284 -2634 1290 -2628
rect 1284 -2640 1290 -2634
rect 1284 -2646 1290 -2640
rect 1284 -2652 1290 -2646
rect 1284 -2658 1290 -2652
rect 1284 -2664 1290 -2658
rect 1284 -2670 1290 -2664
rect 1284 -2676 1290 -2670
rect 1284 -2682 1290 -2676
rect 1284 -2688 1290 -2682
rect 1284 -2694 1290 -2688
rect 1284 -2700 1290 -2694
rect 1284 -2706 1290 -2700
rect 1284 -2712 1290 -2706
rect 1284 -2718 1290 -2712
rect 1284 -2724 1290 -2718
rect 1284 -2730 1290 -2724
rect 1284 -2736 1290 -2730
rect 1284 -2742 1290 -2736
rect 1284 -2748 1290 -2742
rect 1284 -2754 1290 -2748
rect 1284 -2760 1290 -2754
rect 1284 -2766 1290 -2760
rect 1284 -2772 1290 -2766
rect 1284 -2778 1290 -2772
rect 1284 -2784 1290 -2778
rect 1284 -2790 1290 -2784
rect 1284 -2796 1290 -2790
rect 1284 -2802 1290 -2796
rect 1284 -2808 1290 -2802
rect 1284 -2814 1290 -2808
rect 1284 -2820 1290 -2814
rect 1284 -2826 1290 -2820
rect 1284 -2832 1290 -2826
rect 1284 -2838 1290 -2832
rect 1284 -2844 1290 -2838
rect 1284 -2850 1290 -2844
rect 1284 -2856 1290 -2850
rect 1284 -2862 1290 -2856
rect 1284 -2868 1290 -2862
rect 1284 -2874 1290 -2868
rect 1284 -2880 1290 -2874
rect 1284 -2886 1290 -2880
rect 1284 -2892 1290 -2886
rect 1284 -2898 1290 -2892
rect 1284 -2904 1290 -2898
rect 1284 -2910 1290 -2904
rect 1284 -2916 1290 -2910
rect 1284 -2922 1290 -2916
rect 1284 -2928 1290 -2922
rect 1284 -2934 1290 -2928
rect 1284 -2940 1290 -2934
rect 1284 -2946 1290 -2940
rect 1284 -2952 1290 -2946
rect 1284 -2958 1290 -2952
rect 1284 -3036 1290 -3030
rect 1284 -3042 1290 -3036
rect 1284 -3048 1290 -3042
rect 1284 -3054 1290 -3048
rect 1284 -3060 1290 -3054
rect 1284 -3066 1290 -3060
rect 1284 -3072 1290 -3066
rect 1284 -3078 1290 -3072
rect 1284 -3084 1290 -3078
rect 1284 -3090 1290 -3084
rect 1284 -3096 1290 -3090
rect 1284 -3102 1290 -3096
rect 1284 -3108 1290 -3102
rect 1284 -3114 1290 -3108
rect 1284 -3120 1290 -3114
rect 1284 -3126 1290 -3120
rect 1284 -3132 1290 -3126
rect 1284 -3138 1290 -3132
rect 1284 -3144 1290 -3138
rect 1284 -3150 1290 -3144
rect 1284 -3156 1290 -3150
rect 1284 -3162 1290 -3156
rect 1284 -3168 1290 -3162
rect 1284 -3174 1290 -3168
rect 1284 -3180 1290 -3174
rect 1284 -3186 1290 -3180
rect 1284 -3192 1290 -3186
rect 1284 -3198 1290 -3192
rect 1284 -3204 1290 -3198
rect 1284 -3210 1290 -3204
rect 1284 -3216 1290 -3210
rect 1284 -3222 1290 -3216
rect 1284 -3228 1290 -3222
rect 1284 -3234 1290 -3228
rect 1284 -3318 1290 -3312
rect 1284 -3324 1290 -3318
rect 1284 -3330 1290 -3324
rect 1284 -3336 1290 -3330
rect 1284 -3342 1290 -3336
rect 1284 -3348 1290 -3342
rect 1284 -3354 1290 -3348
rect 1284 -3360 1290 -3354
rect 1284 -3366 1290 -3360
rect 1284 -3372 1290 -3366
rect 1284 -3378 1290 -3372
rect 1284 -3384 1290 -3378
rect 1284 -3390 1290 -3384
rect 1284 -3396 1290 -3390
rect 1284 -3402 1290 -3396
rect 1284 -3408 1290 -3402
rect 1284 -3414 1290 -3408
rect 1284 -3420 1290 -3414
rect 1284 -3426 1290 -3420
rect 1284 -3432 1290 -3426
rect 1284 -3438 1290 -3432
rect 1284 -3444 1290 -3438
rect 1284 -3450 1290 -3444
rect 1284 -3456 1290 -3450
rect 1284 -3462 1290 -3456
rect 1284 -3468 1290 -3462
rect 1284 -3474 1290 -3468
rect 1284 -3480 1290 -3474
rect 1284 -3486 1290 -3480
rect 1284 -3492 1290 -3486
rect 1284 -3498 1290 -3492
rect 1284 -3504 1290 -3498
rect 1284 -3510 1290 -3504
rect 1284 -3516 1290 -3510
rect 1290 -1110 1296 -1104
rect 1290 -1116 1296 -1110
rect 1290 -1122 1296 -1116
rect 1290 -1128 1296 -1122
rect 1290 -1134 1296 -1128
rect 1290 -1140 1296 -1134
rect 1290 -1146 1296 -1140
rect 1290 -1152 1296 -1146
rect 1290 -1158 1296 -1152
rect 1290 -1164 1296 -1158
rect 1290 -1170 1296 -1164
rect 1290 -1176 1296 -1170
rect 1290 -1182 1296 -1176
rect 1290 -1188 1296 -1182
rect 1290 -1194 1296 -1188
rect 1290 -1200 1296 -1194
rect 1290 -1206 1296 -1200
rect 1290 -1212 1296 -1206
rect 1290 -1218 1296 -1212
rect 1290 -1224 1296 -1218
rect 1290 -1230 1296 -1224
rect 1290 -1236 1296 -1230
rect 1290 -1242 1296 -1236
rect 1290 -1248 1296 -1242
rect 1290 -1254 1296 -1248
rect 1290 -1260 1296 -1254
rect 1290 -1266 1296 -1260
rect 1290 -1272 1296 -1266
rect 1290 -1278 1296 -1272
rect 1290 -1284 1296 -1278
rect 1290 -1290 1296 -1284
rect 1290 -1296 1296 -1290
rect 1290 -1302 1296 -1296
rect 1290 -1308 1296 -1302
rect 1290 -1596 1296 -1590
rect 1290 -1602 1296 -1596
rect 1290 -1608 1296 -1602
rect 1290 -1614 1296 -1608
rect 1290 -1620 1296 -1614
rect 1290 -1626 1296 -1620
rect 1290 -1632 1296 -1626
rect 1290 -1638 1296 -1632
rect 1290 -1644 1296 -1638
rect 1290 -1650 1296 -1644
rect 1290 -1656 1296 -1650
rect 1290 -1662 1296 -1656
rect 1290 -1668 1296 -1662
rect 1290 -1674 1296 -1668
rect 1290 -1680 1296 -1674
rect 1290 -1686 1296 -1680
rect 1290 -1692 1296 -1686
rect 1290 -1698 1296 -1692
rect 1290 -1704 1296 -1698
rect 1290 -1710 1296 -1704
rect 1290 -1716 1296 -1710
rect 1290 -1722 1296 -1716
rect 1290 -1728 1296 -1722
rect 1290 -1734 1296 -1728
rect 1290 -1740 1296 -1734
rect 1290 -1746 1296 -1740
rect 1290 -1752 1296 -1746
rect 1290 -1758 1296 -1752
rect 1290 -1764 1296 -1758
rect 1290 -1770 1296 -1764
rect 1290 -1776 1296 -1770
rect 1290 -1782 1296 -1776
rect 1290 -1788 1296 -1782
rect 1290 -1794 1296 -1788
rect 1290 -1800 1296 -1794
rect 1290 -1806 1296 -1800
rect 1290 -1812 1296 -1806
rect 1290 -1818 1296 -1812
rect 1290 -1824 1296 -1818
rect 1290 -1830 1296 -1824
rect 1290 -1836 1296 -1830
rect 1290 -1842 1296 -1836
rect 1290 -1848 1296 -1842
rect 1290 -1854 1296 -1848
rect 1290 -1860 1296 -1854
rect 1290 -1866 1296 -1860
rect 1290 -1872 1296 -1866
rect 1290 -1878 1296 -1872
rect 1290 -1884 1296 -1878
rect 1290 -1890 1296 -1884
rect 1290 -1896 1296 -1890
rect 1290 -1902 1296 -1896
rect 1290 -1908 1296 -1902
rect 1290 -1914 1296 -1908
rect 1290 -1920 1296 -1914
rect 1290 -1926 1296 -1920
rect 1290 -1932 1296 -1926
rect 1290 -1938 1296 -1932
rect 1290 -1944 1296 -1938
rect 1290 -1950 1296 -1944
rect 1290 -1956 1296 -1950
rect 1290 -1962 1296 -1956
rect 1290 -1968 1296 -1962
rect 1290 -1974 1296 -1968
rect 1290 -1980 1296 -1974
rect 1290 -1986 1296 -1980
rect 1290 -1992 1296 -1986
rect 1290 -1998 1296 -1992
rect 1290 -2004 1296 -1998
rect 1290 -2010 1296 -2004
rect 1290 -2016 1296 -2010
rect 1290 -2022 1296 -2016
rect 1290 -2028 1296 -2022
rect 1290 -2034 1296 -2028
rect 1290 -2040 1296 -2034
rect 1290 -2046 1296 -2040
rect 1290 -2052 1296 -2046
rect 1290 -2058 1296 -2052
rect 1290 -2064 1296 -2058
rect 1290 -2070 1296 -2064
rect 1290 -2076 1296 -2070
rect 1290 -2082 1296 -2076
rect 1290 -2088 1296 -2082
rect 1290 -2094 1296 -2088
rect 1290 -2100 1296 -2094
rect 1290 -2106 1296 -2100
rect 1290 -2112 1296 -2106
rect 1290 -2118 1296 -2112
rect 1290 -2124 1296 -2118
rect 1290 -2130 1296 -2124
rect 1290 -2136 1296 -2130
rect 1290 -2142 1296 -2136
rect 1290 -2148 1296 -2142
rect 1290 -2154 1296 -2148
rect 1290 -2160 1296 -2154
rect 1290 -2166 1296 -2160
rect 1290 -2172 1296 -2166
rect 1290 -2178 1296 -2172
rect 1290 -2184 1296 -2178
rect 1290 -2190 1296 -2184
rect 1290 -2196 1296 -2190
rect 1290 -2202 1296 -2196
rect 1290 -2208 1296 -2202
rect 1290 -2214 1296 -2208
rect 1290 -2220 1296 -2214
rect 1290 -2226 1296 -2220
rect 1290 -2232 1296 -2226
rect 1290 -2238 1296 -2232
rect 1290 -2244 1296 -2238
rect 1290 -2250 1296 -2244
rect 1290 -2256 1296 -2250
rect 1290 -2262 1296 -2256
rect 1290 -2268 1296 -2262
rect 1290 -2274 1296 -2268
rect 1290 -2280 1296 -2274
rect 1290 -2286 1296 -2280
rect 1290 -2292 1296 -2286
rect 1290 -2298 1296 -2292
rect 1290 -2304 1296 -2298
rect 1290 -2310 1296 -2304
rect 1290 -2316 1296 -2310
rect 1290 -2322 1296 -2316
rect 1290 -2328 1296 -2322
rect 1290 -2334 1296 -2328
rect 1290 -2340 1296 -2334
rect 1290 -2346 1296 -2340
rect 1290 -2352 1296 -2346
rect 1290 -2358 1296 -2352
rect 1290 -2364 1296 -2358
rect 1290 -2370 1296 -2364
rect 1290 -2376 1296 -2370
rect 1290 -2382 1296 -2376
rect 1290 -2388 1296 -2382
rect 1290 -2394 1296 -2388
rect 1290 -2400 1296 -2394
rect 1290 -2406 1296 -2400
rect 1290 -2412 1296 -2406
rect 1290 -2418 1296 -2412
rect 1290 -2424 1296 -2418
rect 1290 -2430 1296 -2424
rect 1290 -2436 1296 -2430
rect 1290 -2442 1296 -2436
rect 1290 -2448 1296 -2442
rect 1290 -2454 1296 -2448
rect 1290 -2460 1296 -2454
rect 1290 -2466 1296 -2460
rect 1290 -2472 1296 -2466
rect 1290 -2562 1296 -2556
rect 1290 -2568 1296 -2562
rect 1290 -2574 1296 -2568
rect 1290 -2580 1296 -2574
rect 1290 -2586 1296 -2580
rect 1290 -2592 1296 -2586
rect 1290 -2598 1296 -2592
rect 1290 -2604 1296 -2598
rect 1290 -2610 1296 -2604
rect 1290 -2616 1296 -2610
rect 1290 -2622 1296 -2616
rect 1290 -2628 1296 -2622
rect 1290 -2634 1296 -2628
rect 1290 -2640 1296 -2634
rect 1290 -2646 1296 -2640
rect 1290 -2652 1296 -2646
rect 1290 -2658 1296 -2652
rect 1290 -2664 1296 -2658
rect 1290 -2670 1296 -2664
rect 1290 -2676 1296 -2670
rect 1290 -2682 1296 -2676
rect 1290 -2688 1296 -2682
rect 1290 -2694 1296 -2688
rect 1290 -2700 1296 -2694
rect 1290 -2706 1296 -2700
rect 1290 -2712 1296 -2706
rect 1290 -2718 1296 -2712
rect 1290 -2724 1296 -2718
rect 1290 -2730 1296 -2724
rect 1290 -2736 1296 -2730
rect 1290 -2742 1296 -2736
rect 1290 -2748 1296 -2742
rect 1290 -2754 1296 -2748
rect 1290 -2760 1296 -2754
rect 1290 -2766 1296 -2760
rect 1290 -2772 1296 -2766
rect 1290 -2778 1296 -2772
rect 1290 -2784 1296 -2778
rect 1290 -2790 1296 -2784
rect 1290 -2796 1296 -2790
rect 1290 -2802 1296 -2796
rect 1290 -2808 1296 -2802
rect 1290 -2814 1296 -2808
rect 1290 -2820 1296 -2814
rect 1290 -2826 1296 -2820
rect 1290 -2832 1296 -2826
rect 1290 -2838 1296 -2832
rect 1290 -2844 1296 -2838
rect 1290 -2850 1296 -2844
rect 1290 -2856 1296 -2850
rect 1290 -2862 1296 -2856
rect 1290 -2868 1296 -2862
rect 1290 -2874 1296 -2868
rect 1290 -2880 1296 -2874
rect 1290 -2886 1296 -2880
rect 1290 -2892 1296 -2886
rect 1290 -2898 1296 -2892
rect 1290 -2904 1296 -2898
rect 1290 -2910 1296 -2904
rect 1290 -2916 1296 -2910
rect 1290 -2922 1296 -2916
rect 1290 -2928 1296 -2922
rect 1290 -2934 1296 -2928
rect 1290 -2940 1296 -2934
rect 1290 -2946 1296 -2940
rect 1290 -2952 1296 -2946
rect 1290 -3036 1296 -3030
rect 1290 -3042 1296 -3036
rect 1290 -3048 1296 -3042
rect 1290 -3054 1296 -3048
rect 1290 -3060 1296 -3054
rect 1290 -3066 1296 -3060
rect 1290 -3072 1296 -3066
rect 1290 -3078 1296 -3072
rect 1290 -3084 1296 -3078
rect 1290 -3090 1296 -3084
rect 1290 -3096 1296 -3090
rect 1290 -3102 1296 -3096
rect 1290 -3108 1296 -3102
rect 1290 -3114 1296 -3108
rect 1290 -3120 1296 -3114
rect 1290 -3126 1296 -3120
rect 1290 -3132 1296 -3126
rect 1290 -3138 1296 -3132
rect 1290 -3144 1296 -3138
rect 1290 -3150 1296 -3144
rect 1290 -3156 1296 -3150
rect 1290 -3162 1296 -3156
rect 1290 -3168 1296 -3162
rect 1290 -3174 1296 -3168
rect 1290 -3180 1296 -3174
rect 1290 -3186 1296 -3180
rect 1290 -3192 1296 -3186
rect 1290 -3198 1296 -3192
rect 1290 -3204 1296 -3198
rect 1290 -3210 1296 -3204
rect 1290 -3216 1296 -3210
rect 1290 -3222 1296 -3216
rect 1290 -3228 1296 -3222
rect 1290 -3234 1296 -3228
rect 1290 -3318 1296 -3312
rect 1290 -3324 1296 -3318
rect 1290 -3330 1296 -3324
rect 1290 -3336 1296 -3330
rect 1290 -3342 1296 -3336
rect 1290 -3348 1296 -3342
rect 1290 -3354 1296 -3348
rect 1290 -3360 1296 -3354
rect 1290 -3366 1296 -3360
rect 1290 -3372 1296 -3366
rect 1290 -3378 1296 -3372
rect 1290 -3384 1296 -3378
rect 1290 -3390 1296 -3384
rect 1290 -3396 1296 -3390
rect 1290 -3402 1296 -3396
rect 1290 -3408 1296 -3402
rect 1290 -3414 1296 -3408
rect 1290 -3420 1296 -3414
rect 1290 -3426 1296 -3420
rect 1290 -3432 1296 -3426
rect 1290 -3438 1296 -3432
rect 1290 -3444 1296 -3438
rect 1290 -3450 1296 -3444
rect 1290 -3456 1296 -3450
rect 1290 -3462 1296 -3456
rect 1290 -3468 1296 -3462
rect 1290 -3474 1296 -3468
rect 1290 -3480 1296 -3474
rect 1290 -3486 1296 -3480
rect 1290 -3492 1296 -3486
rect 1290 -3498 1296 -3492
rect 1290 -3504 1296 -3498
rect 1290 -3510 1296 -3504
rect 1290 -3516 1296 -3510
rect 1296 -1110 1302 -1104
rect 1296 -1116 1302 -1110
rect 1296 -1122 1302 -1116
rect 1296 -1128 1302 -1122
rect 1296 -1134 1302 -1128
rect 1296 -1140 1302 -1134
rect 1296 -1146 1302 -1140
rect 1296 -1152 1302 -1146
rect 1296 -1158 1302 -1152
rect 1296 -1164 1302 -1158
rect 1296 -1170 1302 -1164
rect 1296 -1176 1302 -1170
rect 1296 -1182 1302 -1176
rect 1296 -1188 1302 -1182
rect 1296 -1194 1302 -1188
rect 1296 -1200 1302 -1194
rect 1296 -1206 1302 -1200
rect 1296 -1212 1302 -1206
rect 1296 -1218 1302 -1212
rect 1296 -1224 1302 -1218
rect 1296 -1230 1302 -1224
rect 1296 -1236 1302 -1230
rect 1296 -1242 1302 -1236
rect 1296 -1248 1302 -1242
rect 1296 -1254 1302 -1248
rect 1296 -1260 1302 -1254
rect 1296 -1266 1302 -1260
rect 1296 -1272 1302 -1266
rect 1296 -1278 1302 -1272
rect 1296 -1284 1302 -1278
rect 1296 -1290 1302 -1284
rect 1296 -1296 1302 -1290
rect 1296 -1302 1302 -1296
rect 1296 -1308 1302 -1302
rect 1296 -1578 1302 -1572
rect 1296 -1584 1302 -1578
rect 1296 -1590 1302 -1584
rect 1296 -1596 1302 -1590
rect 1296 -1602 1302 -1596
rect 1296 -1608 1302 -1602
rect 1296 -1614 1302 -1608
rect 1296 -1620 1302 -1614
rect 1296 -1626 1302 -1620
rect 1296 -1632 1302 -1626
rect 1296 -1638 1302 -1632
rect 1296 -1644 1302 -1638
rect 1296 -1650 1302 -1644
rect 1296 -1656 1302 -1650
rect 1296 -1662 1302 -1656
rect 1296 -1668 1302 -1662
rect 1296 -1674 1302 -1668
rect 1296 -1680 1302 -1674
rect 1296 -1686 1302 -1680
rect 1296 -1692 1302 -1686
rect 1296 -1698 1302 -1692
rect 1296 -1704 1302 -1698
rect 1296 -1710 1302 -1704
rect 1296 -1716 1302 -1710
rect 1296 -1722 1302 -1716
rect 1296 -1728 1302 -1722
rect 1296 -1734 1302 -1728
rect 1296 -1740 1302 -1734
rect 1296 -1746 1302 -1740
rect 1296 -1752 1302 -1746
rect 1296 -1758 1302 -1752
rect 1296 -1764 1302 -1758
rect 1296 -1770 1302 -1764
rect 1296 -1776 1302 -1770
rect 1296 -1782 1302 -1776
rect 1296 -1788 1302 -1782
rect 1296 -1794 1302 -1788
rect 1296 -1800 1302 -1794
rect 1296 -1806 1302 -1800
rect 1296 -1812 1302 -1806
rect 1296 -1818 1302 -1812
rect 1296 -1824 1302 -1818
rect 1296 -1830 1302 -1824
rect 1296 -1836 1302 -1830
rect 1296 -1842 1302 -1836
rect 1296 -1848 1302 -1842
rect 1296 -1854 1302 -1848
rect 1296 -1860 1302 -1854
rect 1296 -1866 1302 -1860
rect 1296 -1872 1302 -1866
rect 1296 -1878 1302 -1872
rect 1296 -1884 1302 -1878
rect 1296 -1890 1302 -1884
rect 1296 -1896 1302 -1890
rect 1296 -1902 1302 -1896
rect 1296 -1908 1302 -1902
rect 1296 -1914 1302 -1908
rect 1296 -1920 1302 -1914
rect 1296 -1926 1302 -1920
rect 1296 -1932 1302 -1926
rect 1296 -1938 1302 -1932
rect 1296 -1944 1302 -1938
rect 1296 -1950 1302 -1944
rect 1296 -1956 1302 -1950
rect 1296 -1962 1302 -1956
rect 1296 -1968 1302 -1962
rect 1296 -1974 1302 -1968
rect 1296 -1980 1302 -1974
rect 1296 -1986 1302 -1980
rect 1296 -1992 1302 -1986
rect 1296 -1998 1302 -1992
rect 1296 -2004 1302 -1998
rect 1296 -2010 1302 -2004
rect 1296 -2016 1302 -2010
rect 1296 -2022 1302 -2016
rect 1296 -2028 1302 -2022
rect 1296 -2034 1302 -2028
rect 1296 -2040 1302 -2034
rect 1296 -2046 1302 -2040
rect 1296 -2052 1302 -2046
rect 1296 -2058 1302 -2052
rect 1296 -2064 1302 -2058
rect 1296 -2070 1302 -2064
rect 1296 -2076 1302 -2070
rect 1296 -2082 1302 -2076
rect 1296 -2088 1302 -2082
rect 1296 -2094 1302 -2088
rect 1296 -2100 1302 -2094
rect 1296 -2106 1302 -2100
rect 1296 -2112 1302 -2106
rect 1296 -2118 1302 -2112
rect 1296 -2124 1302 -2118
rect 1296 -2130 1302 -2124
rect 1296 -2136 1302 -2130
rect 1296 -2142 1302 -2136
rect 1296 -2148 1302 -2142
rect 1296 -2154 1302 -2148
rect 1296 -2160 1302 -2154
rect 1296 -2166 1302 -2160
rect 1296 -2172 1302 -2166
rect 1296 -2178 1302 -2172
rect 1296 -2184 1302 -2178
rect 1296 -2190 1302 -2184
rect 1296 -2196 1302 -2190
rect 1296 -2202 1302 -2196
rect 1296 -2208 1302 -2202
rect 1296 -2214 1302 -2208
rect 1296 -2220 1302 -2214
rect 1296 -2226 1302 -2220
rect 1296 -2232 1302 -2226
rect 1296 -2238 1302 -2232
rect 1296 -2244 1302 -2238
rect 1296 -2250 1302 -2244
rect 1296 -2256 1302 -2250
rect 1296 -2262 1302 -2256
rect 1296 -2268 1302 -2262
rect 1296 -2274 1302 -2268
rect 1296 -2280 1302 -2274
rect 1296 -2286 1302 -2280
rect 1296 -2292 1302 -2286
rect 1296 -2298 1302 -2292
rect 1296 -2304 1302 -2298
rect 1296 -2310 1302 -2304
rect 1296 -2316 1302 -2310
rect 1296 -2322 1302 -2316
rect 1296 -2328 1302 -2322
rect 1296 -2334 1302 -2328
rect 1296 -2340 1302 -2334
rect 1296 -2346 1302 -2340
rect 1296 -2352 1302 -2346
rect 1296 -2358 1302 -2352
rect 1296 -2364 1302 -2358
rect 1296 -2370 1302 -2364
rect 1296 -2376 1302 -2370
rect 1296 -2382 1302 -2376
rect 1296 -2388 1302 -2382
rect 1296 -2394 1302 -2388
rect 1296 -2400 1302 -2394
rect 1296 -2406 1302 -2400
rect 1296 -2412 1302 -2406
rect 1296 -2418 1302 -2412
rect 1296 -2424 1302 -2418
rect 1296 -2430 1302 -2424
rect 1296 -2436 1302 -2430
rect 1296 -2442 1302 -2436
rect 1296 -2448 1302 -2442
rect 1296 -2454 1302 -2448
rect 1296 -2460 1302 -2454
rect 1296 -2466 1302 -2460
rect 1296 -2550 1302 -2544
rect 1296 -2556 1302 -2550
rect 1296 -2562 1302 -2556
rect 1296 -2568 1302 -2562
rect 1296 -2574 1302 -2568
rect 1296 -2580 1302 -2574
rect 1296 -2586 1302 -2580
rect 1296 -2592 1302 -2586
rect 1296 -2598 1302 -2592
rect 1296 -2604 1302 -2598
rect 1296 -2610 1302 -2604
rect 1296 -2616 1302 -2610
rect 1296 -2622 1302 -2616
rect 1296 -2628 1302 -2622
rect 1296 -2634 1302 -2628
rect 1296 -2640 1302 -2634
rect 1296 -2646 1302 -2640
rect 1296 -2652 1302 -2646
rect 1296 -2658 1302 -2652
rect 1296 -2664 1302 -2658
rect 1296 -2670 1302 -2664
rect 1296 -2676 1302 -2670
rect 1296 -2682 1302 -2676
rect 1296 -2688 1302 -2682
rect 1296 -2694 1302 -2688
rect 1296 -2700 1302 -2694
rect 1296 -2706 1302 -2700
rect 1296 -2712 1302 -2706
rect 1296 -2718 1302 -2712
rect 1296 -2724 1302 -2718
rect 1296 -2730 1302 -2724
rect 1296 -2736 1302 -2730
rect 1296 -2742 1302 -2736
rect 1296 -2748 1302 -2742
rect 1296 -2754 1302 -2748
rect 1296 -2760 1302 -2754
rect 1296 -2766 1302 -2760
rect 1296 -2772 1302 -2766
rect 1296 -2778 1302 -2772
rect 1296 -2784 1302 -2778
rect 1296 -2790 1302 -2784
rect 1296 -2796 1302 -2790
rect 1296 -2802 1302 -2796
rect 1296 -2808 1302 -2802
rect 1296 -2814 1302 -2808
rect 1296 -2820 1302 -2814
rect 1296 -2826 1302 -2820
rect 1296 -2832 1302 -2826
rect 1296 -2838 1302 -2832
rect 1296 -2844 1302 -2838
rect 1296 -2850 1302 -2844
rect 1296 -2856 1302 -2850
rect 1296 -2862 1302 -2856
rect 1296 -2868 1302 -2862
rect 1296 -2874 1302 -2868
rect 1296 -2880 1302 -2874
rect 1296 -2886 1302 -2880
rect 1296 -2892 1302 -2886
rect 1296 -2898 1302 -2892
rect 1296 -2904 1302 -2898
rect 1296 -2910 1302 -2904
rect 1296 -2916 1302 -2910
rect 1296 -2922 1302 -2916
rect 1296 -2928 1302 -2922
rect 1296 -2934 1302 -2928
rect 1296 -2940 1302 -2934
rect 1296 -2946 1302 -2940
rect 1296 -3030 1302 -3024
rect 1296 -3036 1302 -3030
rect 1296 -3042 1302 -3036
rect 1296 -3048 1302 -3042
rect 1296 -3054 1302 -3048
rect 1296 -3060 1302 -3054
rect 1296 -3066 1302 -3060
rect 1296 -3072 1302 -3066
rect 1296 -3078 1302 -3072
rect 1296 -3084 1302 -3078
rect 1296 -3090 1302 -3084
rect 1296 -3096 1302 -3090
rect 1296 -3102 1302 -3096
rect 1296 -3108 1302 -3102
rect 1296 -3114 1302 -3108
rect 1296 -3120 1302 -3114
rect 1296 -3126 1302 -3120
rect 1296 -3132 1302 -3126
rect 1296 -3138 1302 -3132
rect 1296 -3144 1302 -3138
rect 1296 -3150 1302 -3144
rect 1296 -3156 1302 -3150
rect 1296 -3162 1302 -3156
rect 1296 -3168 1302 -3162
rect 1296 -3174 1302 -3168
rect 1296 -3180 1302 -3174
rect 1296 -3186 1302 -3180
rect 1296 -3192 1302 -3186
rect 1296 -3198 1302 -3192
rect 1296 -3204 1302 -3198
rect 1296 -3210 1302 -3204
rect 1296 -3216 1302 -3210
rect 1296 -3222 1302 -3216
rect 1296 -3228 1302 -3222
rect 1296 -3234 1302 -3228
rect 1296 -3318 1302 -3312
rect 1296 -3324 1302 -3318
rect 1296 -3330 1302 -3324
rect 1296 -3336 1302 -3330
rect 1296 -3342 1302 -3336
rect 1296 -3348 1302 -3342
rect 1296 -3354 1302 -3348
rect 1296 -3360 1302 -3354
rect 1296 -3366 1302 -3360
rect 1296 -3372 1302 -3366
rect 1296 -3378 1302 -3372
rect 1296 -3384 1302 -3378
rect 1296 -3390 1302 -3384
rect 1296 -3396 1302 -3390
rect 1296 -3402 1302 -3396
rect 1296 -3408 1302 -3402
rect 1296 -3414 1302 -3408
rect 1296 -3420 1302 -3414
rect 1296 -3426 1302 -3420
rect 1296 -3432 1302 -3426
rect 1296 -3438 1302 -3432
rect 1296 -3444 1302 -3438
rect 1296 -3450 1302 -3444
rect 1296 -3456 1302 -3450
rect 1296 -3462 1302 -3456
rect 1296 -3468 1302 -3462
rect 1296 -3474 1302 -3468
rect 1296 -3480 1302 -3474
rect 1296 -3486 1302 -3480
rect 1296 -3492 1302 -3486
rect 1296 -3498 1302 -3492
rect 1296 -3504 1302 -3498
rect 1296 -3510 1302 -3504
rect 1296 -3516 1302 -3510
rect 1302 -1110 1308 -1104
rect 1302 -1116 1308 -1110
rect 1302 -1122 1308 -1116
rect 1302 -1128 1308 -1122
rect 1302 -1134 1308 -1128
rect 1302 -1140 1308 -1134
rect 1302 -1146 1308 -1140
rect 1302 -1152 1308 -1146
rect 1302 -1158 1308 -1152
rect 1302 -1164 1308 -1158
rect 1302 -1170 1308 -1164
rect 1302 -1176 1308 -1170
rect 1302 -1182 1308 -1176
rect 1302 -1188 1308 -1182
rect 1302 -1194 1308 -1188
rect 1302 -1200 1308 -1194
rect 1302 -1206 1308 -1200
rect 1302 -1212 1308 -1206
rect 1302 -1218 1308 -1212
rect 1302 -1224 1308 -1218
rect 1302 -1230 1308 -1224
rect 1302 -1236 1308 -1230
rect 1302 -1242 1308 -1236
rect 1302 -1248 1308 -1242
rect 1302 -1254 1308 -1248
rect 1302 -1260 1308 -1254
rect 1302 -1266 1308 -1260
rect 1302 -1272 1308 -1266
rect 1302 -1278 1308 -1272
rect 1302 -1284 1308 -1278
rect 1302 -1290 1308 -1284
rect 1302 -1296 1308 -1290
rect 1302 -1302 1308 -1296
rect 1302 -1308 1308 -1302
rect 1302 -1566 1308 -1560
rect 1302 -1572 1308 -1566
rect 1302 -1578 1308 -1572
rect 1302 -1584 1308 -1578
rect 1302 -1590 1308 -1584
rect 1302 -1596 1308 -1590
rect 1302 -1602 1308 -1596
rect 1302 -1608 1308 -1602
rect 1302 -1614 1308 -1608
rect 1302 -1620 1308 -1614
rect 1302 -1626 1308 -1620
rect 1302 -1632 1308 -1626
rect 1302 -1638 1308 -1632
rect 1302 -1644 1308 -1638
rect 1302 -1650 1308 -1644
rect 1302 -1656 1308 -1650
rect 1302 -1662 1308 -1656
rect 1302 -1668 1308 -1662
rect 1302 -1674 1308 -1668
rect 1302 -1680 1308 -1674
rect 1302 -1686 1308 -1680
rect 1302 -1692 1308 -1686
rect 1302 -1698 1308 -1692
rect 1302 -1704 1308 -1698
rect 1302 -1710 1308 -1704
rect 1302 -1716 1308 -1710
rect 1302 -1722 1308 -1716
rect 1302 -1728 1308 -1722
rect 1302 -1734 1308 -1728
rect 1302 -1740 1308 -1734
rect 1302 -1746 1308 -1740
rect 1302 -1752 1308 -1746
rect 1302 -1758 1308 -1752
rect 1302 -1764 1308 -1758
rect 1302 -1770 1308 -1764
rect 1302 -1776 1308 -1770
rect 1302 -1782 1308 -1776
rect 1302 -1788 1308 -1782
rect 1302 -1794 1308 -1788
rect 1302 -1800 1308 -1794
rect 1302 -1806 1308 -1800
rect 1302 -1812 1308 -1806
rect 1302 -1818 1308 -1812
rect 1302 -1824 1308 -1818
rect 1302 -1830 1308 -1824
rect 1302 -1836 1308 -1830
rect 1302 -1842 1308 -1836
rect 1302 -1848 1308 -1842
rect 1302 -1854 1308 -1848
rect 1302 -1860 1308 -1854
rect 1302 -1866 1308 -1860
rect 1302 -1872 1308 -1866
rect 1302 -1878 1308 -1872
rect 1302 -1884 1308 -1878
rect 1302 -1890 1308 -1884
rect 1302 -1896 1308 -1890
rect 1302 -1902 1308 -1896
rect 1302 -1908 1308 -1902
rect 1302 -1914 1308 -1908
rect 1302 -1920 1308 -1914
rect 1302 -1926 1308 -1920
rect 1302 -1932 1308 -1926
rect 1302 -1938 1308 -1932
rect 1302 -1944 1308 -1938
rect 1302 -1950 1308 -1944
rect 1302 -1956 1308 -1950
rect 1302 -1962 1308 -1956
rect 1302 -1968 1308 -1962
rect 1302 -1974 1308 -1968
rect 1302 -1980 1308 -1974
rect 1302 -1986 1308 -1980
rect 1302 -1992 1308 -1986
rect 1302 -1998 1308 -1992
rect 1302 -2004 1308 -1998
rect 1302 -2010 1308 -2004
rect 1302 -2016 1308 -2010
rect 1302 -2022 1308 -2016
rect 1302 -2028 1308 -2022
rect 1302 -2034 1308 -2028
rect 1302 -2040 1308 -2034
rect 1302 -2046 1308 -2040
rect 1302 -2052 1308 -2046
rect 1302 -2058 1308 -2052
rect 1302 -2064 1308 -2058
rect 1302 -2070 1308 -2064
rect 1302 -2076 1308 -2070
rect 1302 -2082 1308 -2076
rect 1302 -2088 1308 -2082
rect 1302 -2094 1308 -2088
rect 1302 -2100 1308 -2094
rect 1302 -2106 1308 -2100
rect 1302 -2112 1308 -2106
rect 1302 -2118 1308 -2112
rect 1302 -2124 1308 -2118
rect 1302 -2130 1308 -2124
rect 1302 -2136 1308 -2130
rect 1302 -2142 1308 -2136
rect 1302 -2148 1308 -2142
rect 1302 -2154 1308 -2148
rect 1302 -2160 1308 -2154
rect 1302 -2166 1308 -2160
rect 1302 -2172 1308 -2166
rect 1302 -2178 1308 -2172
rect 1302 -2184 1308 -2178
rect 1302 -2190 1308 -2184
rect 1302 -2196 1308 -2190
rect 1302 -2202 1308 -2196
rect 1302 -2208 1308 -2202
rect 1302 -2214 1308 -2208
rect 1302 -2220 1308 -2214
rect 1302 -2226 1308 -2220
rect 1302 -2232 1308 -2226
rect 1302 -2238 1308 -2232
rect 1302 -2244 1308 -2238
rect 1302 -2250 1308 -2244
rect 1302 -2256 1308 -2250
rect 1302 -2262 1308 -2256
rect 1302 -2268 1308 -2262
rect 1302 -2274 1308 -2268
rect 1302 -2280 1308 -2274
rect 1302 -2286 1308 -2280
rect 1302 -2292 1308 -2286
rect 1302 -2298 1308 -2292
rect 1302 -2304 1308 -2298
rect 1302 -2310 1308 -2304
rect 1302 -2316 1308 -2310
rect 1302 -2322 1308 -2316
rect 1302 -2328 1308 -2322
rect 1302 -2334 1308 -2328
rect 1302 -2340 1308 -2334
rect 1302 -2346 1308 -2340
rect 1302 -2352 1308 -2346
rect 1302 -2358 1308 -2352
rect 1302 -2364 1308 -2358
rect 1302 -2370 1308 -2364
rect 1302 -2376 1308 -2370
rect 1302 -2382 1308 -2376
rect 1302 -2388 1308 -2382
rect 1302 -2394 1308 -2388
rect 1302 -2400 1308 -2394
rect 1302 -2406 1308 -2400
rect 1302 -2412 1308 -2406
rect 1302 -2418 1308 -2412
rect 1302 -2424 1308 -2418
rect 1302 -2430 1308 -2424
rect 1302 -2436 1308 -2430
rect 1302 -2442 1308 -2436
rect 1302 -2448 1308 -2442
rect 1302 -2454 1308 -2448
rect 1302 -2544 1308 -2538
rect 1302 -2550 1308 -2544
rect 1302 -2556 1308 -2550
rect 1302 -2562 1308 -2556
rect 1302 -2568 1308 -2562
rect 1302 -2574 1308 -2568
rect 1302 -2580 1308 -2574
rect 1302 -2586 1308 -2580
rect 1302 -2592 1308 -2586
rect 1302 -2598 1308 -2592
rect 1302 -2604 1308 -2598
rect 1302 -2610 1308 -2604
rect 1302 -2616 1308 -2610
rect 1302 -2622 1308 -2616
rect 1302 -2628 1308 -2622
rect 1302 -2634 1308 -2628
rect 1302 -2640 1308 -2634
rect 1302 -2646 1308 -2640
rect 1302 -2652 1308 -2646
rect 1302 -2658 1308 -2652
rect 1302 -2664 1308 -2658
rect 1302 -2670 1308 -2664
rect 1302 -2676 1308 -2670
rect 1302 -2682 1308 -2676
rect 1302 -2688 1308 -2682
rect 1302 -2694 1308 -2688
rect 1302 -2700 1308 -2694
rect 1302 -2706 1308 -2700
rect 1302 -2712 1308 -2706
rect 1302 -2718 1308 -2712
rect 1302 -2724 1308 -2718
rect 1302 -2730 1308 -2724
rect 1302 -2736 1308 -2730
rect 1302 -2742 1308 -2736
rect 1302 -2748 1308 -2742
rect 1302 -2754 1308 -2748
rect 1302 -2760 1308 -2754
rect 1302 -2766 1308 -2760
rect 1302 -2772 1308 -2766
rect 1302 -2778 1308 -2772
rect 1302 -2784 1308 -2778
rect 1302 -2790 1308 -2784
rect 1302 -2796 1308 -2790
rect 1302 -2802 1308 -2796
rect 1302 -2808 1308 -2802
rect 1302 -2814 1308 -2808
rect 1302 -2820 1308 -2814
rect 1302 -2826 1308 -2820
rect 1302 -2832 1308 -2826
rect 1302 -2838 1308 -2832
rect 1302 -2844 1308 -2838
rect 1302 -2850 1308 -2844
rect 1302 -2856 1308 -2850
rect 1302 -2862 1308 -2856
rect 1302 -2868 1308 -2862
rect 1302 -2874 1308 -2868
rect 1302 -2880 1308 -2874
rect 1302 -2886 1308 -2880
rect 1302 -2892 1308 -2886
rect 1302 -2898 1308 -2892
rect 1302 -2904 1308 -2898
rect 1302 -2910 1308 -2904
rect 1302 -2916 1308 -2910
rect 1302 -2922 1308 -2916
rect 1302 -2928 1308 -2922
rect 1302 -2934 1308 -2928
rect 1302 -2940 1308 -2934
rect 1302 -2946 1308 -2940
rect 1302 -3024 1308 -3018
rect 1302 -3030 1308 -3024
rect 1302 -3036 1308 -3030
rect 1302 -3042 1308 -3036
rect 1302 -3048 1308 -3042
rect 1302 -3054 1308 -3048
rect 1302 -3060 1308 -3054
rect 1302 -3066 1308 -3060
rect 1302 -3072 1308 -3066
rect 1302 -3078 1308 -3072
rect 1302 -3084 1308 -3078
rect 1302 -3090 1308 -3084
rect 1302 -3096 1308 -3090
rect 1302 -3102 1308 -3096
rect 1302 -3108 1308 -3102
rect 1302 -3114 1308 -3108
rect 1302 -3120 1308 -3114
rect 1302 -3126 1308 -3120
rect 1302 -3132 1308 -3126
rect 1302 -3138 1308 -3132
rect 1302 -3144 1308 -3138
rect 1302 -3150 1308 -3144
rect 1302 -3156 1308 -3150
rect 1302 -3162 1308 -3156
rect 1302 -3168 1308 -3162
rect 1302 -3174 1308 -3168
rect 1302 -3180 1308 -3174
rect 1302 -3186 1308 -3180
rect 1302 -3192 1308 -3186
rect 1302 -3198 1308 -3192
rect 1302 -3204 1308 -3198
rect 1302 -3210 1308 -3204
rect 1302 -3216 1308 -3210
rect 1302 -3222 1308 -3216
rect 1302 -3228 1308 -3222
rect 1302 -3234 1308 -3228
rect 1302 -3318 1308 -3312
rect 1302 -3324 1308 -3318
rect 1302 -3330 1308 -3324
rect 1302 -3336 1308 -3330
rect 1302 -3342 1308 -3336
rect 1302 -3348 1308 -3342
rect 1302 -3354 1308 -3348
rect 1302 -3360 1308 -3354
rect 1302 -3366 1308 -3360
rect 1302 -3372 1308 -3366
rect 1302 -3378 1308 -3372
rect 1302 -3384 1308 -3378
rect 1302 -3390 1308 -3384
rect 1302 -3396 1308 -3390
rect 1302 -3402 1308 -3396
rect 1302 -3408 1308 -3402
rect 1302 -3414 1308 -3408
rect 1302 -3420 1308 -3414
rect 1302 -3426 1308 -3420
rect 1302 -3432 1308 -3426
rect 1302 -3438 1308 -3432
rect 1302 -3444 1308 -3438
rect 1302 -3450 1308 -3444
rect 1302 -3456 1308 -3450
rect 1302 -3462 1308 -3456
rect 1302 -3468 1308 -3462
rect 1302 -3474 1308 -3468
rect 1302 -3480 1308 -3474
rect 1302 -3486 1308 -3480
rect 1302 -3492 1308 -3486
rect 1302 -3498 1308 -3492
rect 1302 -3504 1308 -3498
rect 1302 -3510 1308 -3504
rect 1302 -3516 1308 -3510
rect 1308 -1110 1314 -1104
rect 1308 -1116 1314 -1110
rect 1308 -1122 1314 -1116
rect 1308 -1128 1314 -1122
rect 1308 -1134 1314 -1128
rect 1308 -1140 1314 -1134
rect 1308 -1146 1314 -1140
rect 1308 -1152 1314 -1146
rect 1308 -1158 1314 -1152
rect 1308 -1164 1314 -1158
rect 1308 -1170 1314 -1164
rect 1308 -1176 1314 -1170
rect 1308 -1182 1314 -1176
rect 1308 -1188 1314 -1182
rect 1308 -1194 1314 -1188
rect 1308 -1200 1314 -1194
rect 1308 -1206 1314 -1200
rect 1308 -1212 1314 -1206
rect 1308 -1218 1314 -1212
rect 1308 -1224 1314 -1218
rect 1308 -1230 1314 -1224
rect 1308 -1236 1314 -1230
rect 1308 -1242 1314 -1236
rect 1308 -1248 1314 -1242
rect 1308 -1254 1314 -1248
rect 1308 -1260 1314 -1254
rect 1308 -1266 1314 -1260
rect 1308 -1272 1314 -1266
rect 1308 -1278 1314 -1272
rect 1308 -1284 1314 -1278
rect 1308 -1290 1314 -1284
rect 1308 -1296 1314 -1290
rect 1308 -1302 1314 -1296
rect 1308 -1308 1314 -1302
rect 1308 -1554 1314 -1548
rect 1308 -1560 1314 -1554
rect 1308 -1566 1314 -1560
rect 1308 -1572 1314 -1566
rect 1308 -1578 1314 -1572
rect 1308 -1584 1314 -1578
rect 1308 -1590 1314 -1584
rect 1308 -1596 1314 -1590
rect 1308 -1602 1314 -1596
rect 1308 -1608 1314 -1602
rect 1308 -1614 1314 -1608
rect 1308 -1620 1314 -1614
rect 1308 -1626 1314 -1620
rect 1308 -1632 1314 -1626
rect 1308 -1638 1314 -1632
rect 1308 -1644 1314 -1638
rect 1308 -1650 1314 -1644
rect 1308 -1656 1314 -1650
rect 1308 -1662 1314 -1656
rect 1308 -1668 1314 -1662
rect 1308 -1674 1314 -1668
rect 1308 -1680 1314 -1674
rect 1308 -1686 1314 -1680
rect 1308 -1692 1314 -1686
rect 1308 -1698 1314 -1692
rect 1308 -1704 1314 -1698
rect 1308 -1710 1314 -1704
rect 1308 -1716 1314 -1710
rect 1308 -1722 1314 -1716
rect 1308 -1728 1314 -1722
rect 1308 -1734 1314 -1728
rect 1308 -1740 1314 -1734
rect 1308 -1746 1314 -1740
rect 1308 -1752 1314 -1746
rect 1308 -1758 1314 -1752
rect 1308 -1764 1314 -1758
rect 1308 -1770 1314 -1764
rect 1308 -1776 1314 -1770
rect 1308 -1782 1314 -1776
rect 1308 -1788 1314 -1782
rect 1308 -1794 1314 -1788
rect 1308 -1800 1314 -1794
rect 1308 -1806 1314 -1800
rect 1308 -1812 1314 -1806
rect 1308 -1818 1314 -1812
rect 1308 -1824 1314 -1818
rect 1308 -1830 1314 -1824
rect 1308 -1836 1314 -1830
rect 1308 -1842 1314 -1836
rect 1308 -1848 1314 -1842
rect 1308 -1854 1314 -1848
rect 1308 -1860 1314 -1854
rect 1308 -1866 1314 -1860
rect 1308 -1872 1314 -1866
rect 1308 -1878 1314 -1872
rect 1308 -1884 1314 -1878
rect 1308 -1890 1314 -1884
rect 1308 -1896 1314 -1890
rect 1308 -1902 1314 -1896
rect 1308 -1908 1314 -1902
rect 1308 -1914 1314 -1908
rect 1308 -1920 1314 -1914
rect 1308 -1926 1314 -1920
rect 1308 -1932 1314 -1926
rect 1308 -1938 1314 -1932
rect 1308 -1944 1314 -1938
rect 1308 -1950 1314 -1944
rect 1308 -1956 1314 -1950
rect 1308 -1962 1314 -1956
rect 1308 -1968 1314 -1962
rect 1308 -1974 1314 -1968
rect 1308 -1980 1314 -1974
rect 1308 -1986 1314 -1980
rect 1308 -1992 1314 -1986
rect 1308 -1998 1314 -1992
rect 1308 -2004 1314 -1998
rect 1308 -2010 1314 -2004
rect 1308 -2016 1314 -2010
rect 1308 -2022 1314 -2016
rect 1308 -2028 1314 -2022
rect 1308 -2034 1314 -2028
rect 1308 -2040 1314 -2034
rect 1308 -2046 1314 -2040
rect 1308 -2052 1314 -2046
rect 1308 -2058 1314 -2052
rect 1308 -2064 1314 -2058
rect 1308 -2070 1314 -2064
rect 1308 -2076 1314 -2070
rect 1308 -2082 1314 -2076
rect 1308 -2088 1314 -2082
rect 1308 -2094 1314 -2088
rect 1308 -2100 1314 -2094
rect 1308 -2106 1314 -2100
rect 1308 -2112 1314 -2106
rect 1308 -2118 1314 -2112
rect 1308 -2124 1314 -2118
rect 1308 -2130 1314 -2124
rect 1308 -2136 1314 -2130
rect 1308 -2142 1314 -2136
rect 1308 -2148 1314 -2142
rect 1308 -2154 1314 -2148
rect 1308 -2160 1314 -2154
rect 1308 -2166 1314 -2160
rect 1308 -2172 1314 -2166
rect 1308 -2178 1314 -2172
rect 1308 -2184 1314 -2178
rect 1308 -2190 1314 -2184
rect 1308 -2196 1314 -2190
rect 1308 -2202 1314 -2196
rect 1308 -2208 1314 -2202
rect 1308 -2214 1314 -2208
rect 1308 -2220 1314 -2214
rect 1308 -2226 1314 -2220
rect 1308 -2232 1314 -2226
rect 1308 -2238 1314 -2232
rect 1308 -2244 1314 -2238
rect 1308 -2250 1314 -2244
rect 1308 -2256 1314 -2250
rect 1308 -2262 1314 -2256
rect 1308 -2268 1314 -2262
rect 1308 -2274 1314 -2268
rect 1308 -2280 1314 -2274
rect 1308 -2286 1314 -2280
rect 1308 -2292 1314 -2286
rect 1308 -2298 1314 -2292
rect 1308 -2304 1314 -2298
rect 1308 -2310 1314 -2304
rect 1308 -2316 1314 -2310
rect 1308 -2322 1314 -2316
rect 1308 -2328 1314 -2322
rect 1308 -2334 1314 -2328
rect 1308 -2340 1314 -2334
rect 1308 -2346 1314 -2340
rect 1308 -2352 1314 -2346
rect 1308 -2358 1314 -2352
rect 1308 -2364 1314 -2358
rect 1308 -2370 1314 -2364
rect 1308 -2376 1314 -2370
rect 1308 -2382 1314 -2376
rect 1308 -2388 1314 -2382
rect 1308 -2394 1314 -2388
rect 1308 -2400 1314 -2394
rect 1308 -2406 1314 -2400
rect 1308 -2412 1314 -2406
rect 1308 -2418 1314 -2412
rect 1308 -2424 1314 -2418
rect 1308 -2430 1314 -2424
rect 1308 -2436 1314 -2430
rect 1308 -2442 1314 -2436
rect 1308 -2448 1314 -2442
rect 1308 -2532 1314 -2526
rect 1308 -2538 1314 -2532
rect 1308 -2544 1314 -2538
rect 1308 -2550 1314 -2544
rect 1308 -2556 1314 -2550
rect 1308 -2562 1314 -2556
rect 1308 -2568 1314 -2562
rect 1308 -2574 1314 -2568
rect 1308 -2580 1314 -2574
rect 1308 -2586 1314 -2580
rect 1308 -2592 1314 -2586
rect 1308 -2598 1314 -2592
rect 1308 -2604 1314 -2598
rect 1308 -2610 1314 -2604
rect 1308 -2616 1314 -2610
rect 1308 -2622 1314 -2616
rect 1308 -2628 1314 -2622
rect 1308 -2634 1314 -2628
rect 1308 -2640 1314 -2634
rect 1308 -2646 1314 -2640
rect 1308 -2652 1314 -2646
rect 1308 -2658 1314 -2652
rect 1308 -2664 1314 -2658
rect 1308 -2670 1314 -2664
rect 1308 -2676 1314 -2670
rect 1308 -2682 1314 -2676
rect 1308 -2688 1314 -2682
rect 1308 -2694 1314 -2688
rect 1308 -2700 1314 -2694
rect 1308 -2706 1314 -2700
rect 1308 -2712 1314 -2706
rect 1308 -2718 1314 -2712
rect 1308 -2724 1314 -2718
rect 1308 -2730 1314 -2724
rect 1308 -2736 1314 -2730
rect 1308 -2742 1314 -2736
rect 1308 -2748 1314 -2742
rect 1308 -2754 1314 -2748
rect 1308 -2760 1314 -2754
rect 1308 -2766 1314 -2760
rect 1308 -2772 1314 -2766
rect 1308 -2778 1314 -2772
rect 1308 -2784 1314 -2778
rect 1308 -2790 1314 -2784
rect 1308 -2796 1314 -2790
rect 1308 -2802 1314 -2796
rect 1308 -2808 1314 -2802
rect 1308 -2814 1314 -2808
rect 1308 -2820 1314 -2814
rect 1308 -2826 1314 -2820
rect 1308 -2832 1314 -2826
rect 1308 -2838 1314 -2832
rect 1308 -2844 1314 -2838
rect 1308 -2850 1314 -2844
rect 1308 -2856 1314 -2850
rect 1308 -2862 1314 -2856
rect 1308 -2868 1314 -2862
rect 1308 -2874 1314 -2868
rect 1308 -2880 1314 -2874
rect 1308 -2886 1314 -2880
rect 1308 -2892 1314 -2886
rect 1308 -2898 1314 -2892
rect 1308 -2904 1314 -2898
rect 1308 -2910 1314 -2904
rect 1308 -2916 1314 -2910
rect 1308 -2922 1314 -2916
rect 1308 -2928 1314 -2922
rect 1308 -2934 1314 -2928
rect 1308 -2940 1314 -2934
rect 1308 -3024 1314 -3018
rect 1308 -3030 1314 -3024
rect 1308 -3036 1314 -3030
rect 1308 -3042 1314 -3036
rect 1308 -3048 1314 -3042
rect 1308 -3054 1314 -3048
rect 1308 -3060 1314 -3054
rect 1308 -3066 1314 -3060
rect 1308 -3072 1314 -3066
rect 1308 -3078 1314 -3072
rect 1308 -3084 1314 -3078
rect 1308 -3090 1314 -3084
rect 1308 -3096 1314 -3090
rect 1308 -3102 1314 -3096
rect 1308 -3108 1314 -3102
rect 1308 -3114 1314 -3108
rect 1308 -3120 1314 -3114
rect 1308 -3126 1314 -3120
rect 1308 -3132 1314 -3126
rect 1308 -3138 1314 -3132
rect 1308 -3144 1314 -3138
rect 1308 -3150 1314 -3144
rect 1308 -3156 1314 -3150
rect 1308 -3162 1314 -3156
rect 1308 -3168 1314 -3162
rect 1308 -3174 1314 -3168
rect 1308 -3180 1314 -3174
rect 1308 -3186 1314 -3180
rect 1308 -3192 1314 -3186
rect 1308 -3198 1314 -3192
rect 1308 -3204 1314 -3198
rect 1308 -3210 1314 -3204
rect 1308 -3216 1314 -3210
rect 1308 -3222 1314 -3216
rect 1308 -3228 1314 -3222
rect 1308 -3234 1314 -3228
rect 1308 -3318 1314 -3312
rect 1308 -3324 1314 -3318
rect 1308 -3330 1314 -3324
rect 1308 -3336 1314 -3330
rect 1308 -3342 1314 -3336
rect 1308 -3348 1314 -3342
rect 1308 -3354 1314 -3348
rect 1308 -3360 1314 -3354
rect 1308 -3366 1314 -3360
rect 1308 -3372 1314 -3366
rect 1308 -3378 1314 -3372
rect 1308 -3384 1314 -3378
rect 1308 -3390 1314 -3384
rect 1308 -3396 1314 -3390
rect 1308 -3402 1314 -3396
rect 1308 -3408 1314 -3402
rect 1308 -3414 1314 -3408
rect 1308 -3420 1314 -3414
rect 1308 -3426 1314 -3420
rect 1308 -3432 1314 -3426
rect 1308 -3438 1314 -3432
rect 1308 -3444 1314 -3438
rect 1308 -3450 1314 -3444
rect 1308 -3456 1314 -3450
rect 1308 -3462 1314 -3456
rect 1308 -3468 1314 -3462
rect 1308 -3474 1314 -3468
rect 1308 -3480 1314 -3474
rect 1308 -3486 1314 -3480
rect 1308 -3492 1314 -3486
rect 1308 -3498 1314 -3492
rect 1308 -3504 1314 -3498
rect 1308 -3510 1314 -3504
rect 1308 -3516 1314 -3510
rect 1314 -1110 1320 -1104
rect 1314 -1116 1320 -1110
rect 1314 -1122 1320 -1116
rect 1314 -1128 1320 -1122
rect 1314 -1134 1320 -1128
rect 1314 -1140 1320 -1134
rect 1314 -1146 1320 -1140
rect 1314 -1152 1320 -1146
rect 1314 -1158 1320 -1152
rect 1314 -1164 1320 -1158
rect 1314 -1170 1320 -1164
rect 1314 -1176 1320 -1170
rect 1314 -1182 1320 -1176
rect 1314 -1188 1320 -1182
rect 1314 -1194 1320 -1188
rect 1314 -1200 1320 -1194
rect 1314 -1206 1320 -1200
rect 1314 -1212 1320 -1206
rect 1314 -1218 1320 -1212
rect 1314 -1224 1320 -1218
rect 1314 -1230 1320 -1224
rect 1314 -1236 1320 -1230
rect 1314 -1242 1320 -1236
rect 1314 -1248 1320 -1242
rect 1314 -1254 1320 -1248
rect 1314 -1260 1320 -1254
rect 1314 -1266 1320 -1260
rect 1314 -1272 1320 -1266
rect 1314 -1278 1320 -1272
rect 1314 -1284 1320 -1278
rect 1314 -1290 1320 -1284
rect 1314 -1296 1320 -1290
rect 1314 -1302 1320 -1296
rect 1314 -1308 1320 -1302
rect 1314 -1542 1320 -1536
rect 1314 -1548 1320 -1542
rect 1314 -1554 1320 -1548
rect 1314 -1560 1320 -1554
rect 1314 -1566 1320 -1560
rect 1314 -1572 1320 -1566
rect 1314 -1578 1320 -1572
rect 1314 -1584 1320 -1578
rect 1314 -1590 1320 -1584
rect 1314 -1596 1320 -1590
rect 1314 -1602 1320 -1596
rect 1314 -1608 1320 -1602
rect 1314 -1614 1320 -1608
rect 1314 -1620 1320 -1614
rect 1314 -1626 1320 -1620
rect 1314 -1632 1320 -1626
rect 1314 -1638 1320 -1632
rect 1314 -1644 1320 -1638
rect 1314 -1650 1320 -1644
rect 1314 -1656 1320 -1650
rect 1314 -1662 1320 -1656
rect 1314 -1668 1320 -1662
rect 1314 -1674 1320 -1668
rect 1314 -1680 1320 -1674
rect 1314 -1686 1320 -1680
rect 1314 -1692 1320 -1686
rect 1314 -1698 1320 -1692
rect 1314 -1704 1320 -1698
rect 1314 -1710 1320 -1704
rect 1314 -1716 1320 -1710
rect 1314 -1722 1320 -1716
rect 1314 -1728 1320 -1722
rect 1314 -1734 1320 -1728
rect 1314 -1740 1320 -1734
rect 1314 -1746 1320 -1740
rect 1314 -1752 1320 -1746
rect 1314 -1758 1320 -1752
rect 1314 -1764 1320 -1758
rect 1314 -1770 1320 -1764
rect 1314 -1776 1320 -1770
rect 1314 -1782 1320 -1776
rect 1314 -1788 1320 -1782
rect 1314 -1794 1320 -1788
rect 1314 -1800 1320 -1794
rect 1314 -1806 1320 -1800
rect 1314 -1812 1320 -1806
rect 1314 -1818 1320 -1812
rect 1314 -1824 1320 -1818
rect 1314 -1830 1320 -1824
rect 1314 -1836 1320 -1830
rect 1314 -1842 1320 -1836
rect 1314 -1848 1320 -1842
rect 1314 -1854 1320 -1848
rect 1314 -1860 1320 -1854
rect 1314 -1866 1320 -1860
rect 1314 -1872 1320 -1866
rect 1314 -1878 1320 -1872
rect 1314 -1884 1320 -1878
rect 1314 -1890 1320 -1884
rect 1314 -1896 1320 -1890
rect 1314 -1902 1320 -1896
rect 1314 -1908 1320 -1902
rect 1314 -1914 1320 -1908
rect 1314 -1920 1320 -1914
rect 1314 -1926 1320 -1920
rect 1314 -1932 1320 -1926
rect 1314 -1938 1320 -1932
rect 1314 -1944 1320 -1938
rect 1314 -1950 1320 -1944
rect 1314 -1956 1320 -1950
rect 1314 -1962 1320 -1956
rect 1314 -1968 1320 -1962
rect 1314 -1974 1320 -1968
rect 1314 -1980 1320 -1974
rect 1314 -1986 1320 -1980
rect 1314 -1992 1320 -1986
rect 1314 -1998 1320 -1992
rect 1314 -2004 1320 -1998
rect 1314 -2010 1320 -2004
rect 1314 -2016 1320 -2010
rect 1314 -2022 1320 -2016
rect 1314 -2028 1320 -2022
rect 1314 -2034 1320 -2028
rect 1314 -2040 1320 -2034
rect 1314 -2046 1320 -2040
rect 1314 -2052 1320 -2046
rect 1314 -2058 1320 -2052
rect 1314 -2064 1320 -2058
rect 1314 -2070 1320 -2064
rect 1314 -2076 1320 -2070
rect 1314 -2082 1320 -2076
rect 1314 -2088 1320 -2082
rect 1314 -2094 1320 -2088
rect 1314 -2100 1320 -2094
rect 1314 -2106 1320 -2100
rect 1314 -2112 1320 -2106
rect 1314 -2118 1320 -2112
rect 1314 -2124 1320 -2118
rect 1314 -2130 1320 -2124
rect 1314 -2136 1320 -2130
rect 1314 -2142 1320 -2136
rect 1314 -2148 1320 -2142
rect 1314 -2154 1320 -2148
rect 1314 -2160 1320 -2154
rect 1314 -2166 1320 -2160
rect 1314 -2172 1320 -2166
rect 1314 -2178 1320 -2172
rect 1314 -2184 1320 -2178
rect 1314 -2190 1320 -2184
rect 1314 -2196 1320 -2190
rect 1314 -2202 1320 -2196
rect 1314 -2208 1320 -2202
rect 1314 -2214 1320 -2208
rect 1314 -2220 1320 -2214
rect 1314 -2226 1320 -2220
rect 1314 -2232 1320 -2226
rect 1314 -2238 1320 -2232
rect 1314 -2244 1320 -2238
rect 1314 -2250 1320 -2244
rect 1314 -2256 1320 -2250
rect 1314 -2262 1320 -2256
rect 1314 -2268 1320 -2262
rect 1314 -2274 1320 -2268
rect 1314 -2280 1320 -2274
rect 1314 -2286 1320 -2280
rect 1314 -2292 1320 -2286
rect 1314 -2298 1320 -2292
rect 1314 -2304 1320 -2298
rect 1314 -2310 1320 -2304
rect 1314 -2316 1320 -2310
rect 1314 -2322 1320 -2316
rect 1314 -2328 1320 -2322
rect 1314 -2334 1320 -2328
rect 1314 -2340 1320 -2334
rect 1314 -2346 1320 -2340
rect 1314 -2352 1320 -2346
rect 1314 -2358 1320 -2352
rect 1314 -2364 1320 -2358
rect 1314 -2370 1320 -2364
rect 1314 -2376 1320 -2370
rect 1314 -2382 1320 -2376
rect 1314 -2388 1320 -2382
rect 1314 -2394 1320 -2388
rect 1314 -2400 1320 -2394
rect 1314 -2406 1320 -2400
rect 1314 -2412 1320 -2406
rect 1314 -2418 1320 -2412
rect 1314 -2424 1320 -2418
rect 1314 -2430 1320 -2424
rect 1314 -2436 1320 -2430
rect 1314 -2442 1320 -2436
rect 1314 -2526 1320 -2520
rect 1314 -2532 1320 -2526
rect 1314 -2538 1320 -2532
rect 1314 -2544 1320 -2538
rect 1314 -2550 1320 -2544
rect 1314 -2556 1320 -2550
rect 1314 -2562 1320 -2556
rect 1314 -2568 1320 -2562
rect 1314 -2574 1320 -2568
rect 1314 -2580 1320 -2574
rect 1314 -2586 1320 -2580
rect 1314 -2592 1320 -2586
rect 1314 -2598 1320 -2592
rect 1314 -2604 1320 -2598
rect 1314 -2610 1320 -2604
rect 1314 -2616 1320 -2610
rect 1314 -2622 1320 -2616
rect 1314 -2628 1320 -2622
rect 1314 -2634 1320 -2628
rect 1314 -2640 1320 -2634
rect 1314 -2646 1320 -2640
rect 1314 -2652 1320 -2646
rect 1314 -2658 1320 -2652
rect 1314 -2664 1320 -2658
rect 1314 -2670 1320 -2664
rect 1314 -2676 1320 -2670
rect 1314 -2682 1320 -2676
rect 1314 -2688 1320 -2682
rect 1314 -2694 1320 -2688
rect 1314 -2700 1320 -2694
rect 1314 -2706 1320 -2700
rect 1314 -2712 1320 -2706
rect 1314 -2718 1320 -2712
rect 1314 -2724 1320 -2718
rect 1314 -2730 1320 -2724
rect 1314 -2736 1320 -2730
rect 1314 -2742 1320 -2736
rect 1314 -2748 1320 -2742
rect 1314 -2754 1320 -2748
rect 1314 -2760 1320 -2754
rect 1314 -2766 1320 -2760
rect 1314 -2772 1320 -2766
rect 1314 -2778 1320 -2772
rect 1314 -2784 1320 -2778
rect 1314 -2790 1320 -2784
rect 1314 -2796 1320 -2790
rect 1314 -2802 1320 -2796
rect 1314 -2808 1320 -2802
rect 1314 -2814 1320 -2808
rect 1314 -2820 1320 -2814
rect 1314 -2826 1320 -2820
rect 1314 -2832 1320 -2826
rect 1314 -2838 1320 -2832
rect 1314 -2844 1320 -2838
rect 1314 -2850 1320 -2844
rect 1314 -2856 1320 -2850
rect 1314 -2862 1320 -2856
rect 1314 -2868 1320 -2862
rect 1314 -2874 1320 -2868
rect 1314 -2880 1320 -2874
rect 1314 -2886 1320 -2880
rect 1314 -2892 1320 -2886
rect 1314 -2898 1320 -2892
rect 1314 -2904 1320 -2898
rect 1314 -2910 1320 -2904
rect 1314 -2916 1320 -2910
rect 1314 -2922 1320 -2916
rect 1314 -2928 1320 -2922
rect 1314 -2934 1320 -2928
rect 1314 -3018 1320 -3012
rect 1314 -3024 1320 -3018
rect 1314 -3030 1320 -3024
rect 1314 -3036 1320 -3030
rect 1314 -3042 1320 -3036
rect 1314 -3048 1320 -3042
rect 1314 -3054 1320 -3048
rect 1314 -3060 1320 -3054
rect 1314 -3066 1320 -3060
rect 1314 -3072 1320 -3066
rect 1314 -3078 1320 -3072
rect 1314 -3084 1320 -3078
rect 1314 -3090 1320 -3084
rect 1314 -3096 1320 -3090
rect 1314 -3102 1320 -3096
rect 1314 -3108 1320 -3102
rect 1314 -3114 1320 -3108
rect 1314 -3120 1320 -3114
rect 1314 -3126 1320 -3120
rect 1314 -3132 1320 -3126
rect 1314 -3138 1320 -3132
rect 1314 -3144 1320 -3138
rect 1314 -3150 1320 -3144
rect 1314 -3156 1320 -3150
rect 1314 -3162 1320 -3156
rect 1314 -3168 1320 -3162
rect 1314 -3174 1320 -3168
rect 1314 -3180 1320 -3174
rect 1314 -3186 1320 -3180
rect 1314 -3192 1320 -3186
rect 1314 -3198 1320 -3192
rect 1314 -3204 1320 -3198
rect 1314 -3210 1320 -3204
rect 1314 -3216 1320 -3210
rect 1314 -3222 1320 -3216
rect 1314 -3228 1320 -3222
rect 1314 -3234 1320 -3228
rect 1314 -3318 1320 -3312
rect 1314 -3324 1320 -3318
rect 1314 -3330 1320 -3324
rect 1314 -3336 1320 -3330
rect 1314 -3342 1320 -3336
rect 1314 -3348 1320 -3342
rect 1314 -3354 1320 -3348
rect 1314 -3360 1320 -3354
rect 1314 -3366 1320 -3360
rect 1314 -3372 1320 -3366
rect 1314 -3378 1320 -3372
rect 1314 -3384 1320 -3378
rect 1314 -3390 1320 -3384
rect 1314 -3396 1320 -3390
rect 1314 -3402 1320 -3396
rect 1314 -3408 1320 -3402
rect 1314 -3414 1320 -3408
rect 1314 -3420 1320 -3414
rect 1314 -3426 1320 -3420
rect 1314 -3432 1320 -3426
rect 1314 -3438 1320 -3432
rect 1314 -3444 1320 -3438
rect 1314 -3450 1320 -3444
rect 1314 -3456 1320 -3450
rect 1314 -3462 1320 -3456
rect 1314 -3468 1320 -3462
rect 1314 -3474 1320 -3468
rect 1314 -3480 1320 -3474
rect 1314 -3486 1320 -3480
rect 1314 -3492 1320 -3486
rect 1314 -3498 1320 -3492
rect 1314 -3504 1320 -3498
rect 1314 -3510 1320 -3504
rect 1314 -3516 1320 -3510
rect 1320 -1110 1326 -1104
rect 1320 -1116 1326 -1110
rect 1320 -1122 1326 -1116
rect 1320 -1128 1326 -1122
rect 1320 -1134 1326 -1128
rect 1320 -1140 1326 -1134
rect 1320 -1146 1326 -1140
rect 1320 -1152 1326 -1146
rect 1320 -1158 1326 -1152
rect 1320 -1164 1326 -1158
rect 1320 -1170 1326 -1164
rect 1320 -1176 1326 -1170
rect 1320 -1182 1326 -1176
rect 1320 -1188 1326 -1182
rect 1320 -1194 1326 -1188
rect 1320 -1200 1326 -1194
rect 1320 -1206 1326 -1200
rect 1320 -1212 1326 -1206
rect 1320 -1218 1326 -1212
rect 1320 -1224 1326 -1218
rect 1320 -1230 1326 -1224
rect 1320 -1236 1326 -1230
rect 1320 -1242 1326 -1236
rect 1320 -1248 1326 -1242
rect 1320 -1254 1326 -1248
rect 1320 -1260 1326 -1254
rect 1320 -1266 1326 -1260
rect 1320 -1272 1326 -1266
rect 1320 -1278 1326 -1272
rect 1320 -1284 1326 -1278
rect 1320 -1290 1326 -1284
rect 1320 -1296 1326 -1290
rect 1320 -1302 1326 -1296
rect 1320 -1308 1326 -1302
rect 1320 -1524 1326 -1518
rect 1320 -1530 1326 -1524
rect 1320 -1536 1326 -1530
rect 1320 -1542 1326 -1536
rect 1320 -1548 1326 -1542
rect 1320 -1554 1326 -1548
rect 1320 -1560 1326 -1554
rect 1320 -1566 1326 -1560
rect 1320 -1572 1326 -1566
rect 1320 -1578 1326 -1572
rect 1320 -1584 1326 -1578
rect 1320 -1590 1326 -1584
rect 1320 -1596 1326 -1590
rect 1320 -1602 1326 -1596
rect 1320 -1608 1326 -1602
rect 1320 -1614 1326 -1608
rect 1320 -1620 1326 -1614
rect 1320 -1626 1326 -1620
rect 1320 -1632 1326 -1626
rect 1320 -1638 1326 -1632
rect 1320 -1644 1326 -1638
rect 1320 -1650 1326 -1644
rect 1320 -1656 1326 -1650
rect 1320 -1662 1326 -1656
rect 1320 -1668 1326 -1662
rect 1320 -1674 1326 -1668
rect 1320 -1680 1326 -1674
rect 1320 -1686 1326 -1680
rect 1320 -1692 1326 -1686
rect 1320 -1698 1326 -1692
rect 1320 -1704 1326 -1698
rect 1320 -1710 1326 -1704
rect 1320 -1716 1326 -1710
rect 1320 -1722 1326 -1716
rect 1320 -1728 1326 -1722
rect 1320 -1734 1326 -1728
rect 1320 -1740 1326 -1734
rect 1320 -1746 1326 -1740
rect 1320 -1752 1326 -1746
rect 1320 -1758 1326 -1752
rect 1320 -1764 1326 -1758
rect 1320 -1770 1326 -1764
rect 1320 -1776 1326 -1770
rect 1320 -1782 1326 -1776
rect 1320 -1788 1326 -1782
rect 1320 -1794 1326 -1788
rect 1320 -1800 1326 -1794
rect 1320 -1806 1326 -1800
rect 1320 -1812 1326 -1806
rect 1320 -1818 1326 -1812
rect 1320 -1824 1326 -1818
rect 1320 -1830 1326 -1824
rect 1320 -1836 1326 -1830
rect 1320 -1842 1326 -1836
rect 1320 -1848 1326 -1842
rect 1320 -1854 1326 -1848
rect 1320 -1860 1326 -1854
rect 1320 -1866 1326 -1860
rect 1320 -1872 1326 -1866
rect 1320 -1878 1326 -1872
rect 1320 -1884 1326 -1878
rect 1320 -1890 1326 -1884
rect 1320 -1896 1326 -1890
rect 1320 -1902 1326 -1896
rect 1320 -1908 1326 -1902
rect 1320 -1914 1326 -1908
rect 1320 -1920 1326 -1914
rect 1320 -1926 1326 -1920
rect 1320 -1932 1326 -1926
rect 1320 -1938 1326 -1932
rect 1320 -1944 1326 -1938
rect 1320 -1950 1326 -1944
rect 1320 -1956 1326 -1950
rect 1320 -1962 1326 -1956
rect 1320 -1968 1326 -1962
rect 1320 -1974 1326 -1968
rect 1320 -1980 1326 -1974
rect 1320 -1986 1326 -1980
rect 1320 -1992 1326 -1986
rect 1320 -1998 1326 -1992
rect 1320 -2004 1326 -1998
rect 1320 -2010 1326 -2004
rect 1320 -2016 1326 -2010
rect 1320 -2022 1326 -2016
rect 1320 -2028 1326 -2022
rect 1320 -2034 1326 -2028
rect 1320 -2040 1326 -2034
rect 1320 -2046 1326 -2040
rect 1320 -2052 1326 -2046
rect 1320 -2058 1326 -2052
rect 1320 -2064 1326 -2058
rect 1320 -2070 1326 -2064
rect 1320 -2076 1326 -2070
rect 1320 -2082 1326 -2076
rect 1320 -2088 1326 -2082
rect 1320 -2094 1326 -2088
rect 1320 -2100 1326 -2094
rect 1320 -2106 1326 -2100
rect 1320 -2112 1326 -2106
rect 1320 -2118 1326 -2112
rect 1320 -2124 1326 -2118
rect 1320 -2130 1326 -2124
rect 1320 -2136 1326 -2130
rect 1320 -2142 1326 -2136
rect 1320 -2148 1326 -2142
rect 1320 -2154 1326 -2148
rect 1320 -2160 1326 -2154
rect 1320 -2166 1326 -2160
rect 1320 -2172 1326 -2166
rect 1320 -2178 1326 -2172
rect 1320 -2184 1326 -2178
rect 1320 -2190 1326 -2184
rect 1320 -2196 1326 -2190
rect 1320 -2202 1326 -2196
rect 1320 -2208 1326 -2202
rect 1320 -2214 1326 -2208
rect 1320 -2220 1326 -2214
rect 1320 -2226 1326 -2220
rect 1320 -2232 1326 -2226
rect 1320 -2238 1326 -2232
rect 1320 -2244 1326 -2238
rect 1320 -2250 1326 -2244
rect 1320 -2256 1326 -2250
rect 1320 -2262 1326 -2256
rect 1320 -2268 1326 -2262
rect 1320 -2274 1326 -2268
rect 1320 -2280 1326 -2274
rect 1320 -2286 1326 -2280
rect 1320 -2292 1326 -2286
rect 1320 -2298 1326 -2292
rect 1320 -2304 1326 -2298
rect 1320 -2310 1326 -2304
rect 1320 -2316 1326 -2310
rect 1320 -2322 1326 -2316
rect 1320 -2328 1326 -2322
rect 1320 -2334 1326 -2328
rect 1320 -2340 1326 -2334
rect 1320 -2346 1326 -2340
rect 1320 -2352 1326 -2346
rect 1320 -2358 1326 -2352
rect 1320 -2364 1326 -2358
rect 1320 -2370 1326 -2364
rect 1320 -2376 1326 -2370
rect 1320 -2382 1326 -2376
rect 1320 -2388 1326 -2382
rect 1320 -2394 1326 -2388
rect 1320 -2400 1326 -2394
rect 1320 -2406 1326 -2400
rect 1320 -2412 1326 -2406
rect 1320 -2418 1326 -2412
rect 1320 -2424 1326 -2418
rect 1320 -2430 1326 -2424
rect 1320 -2514 1326 -2508
rect 1320 -2520 1326 -2514
rect 1320 -2526 1326 -2520
rect 1320 -2532 1326 -2526
rect 1320 -2538 1326 -2532
rect 1320 -2544 1326 -2538
rect 1320 -2550 1326 -2544
rect 1320 -2556 1326 -2550
rect 1320 -2562 1326 -2556
rect 1320 -2568 1326 -2562
rect 1320 -2574 1326 -2568
rect 1320 -2580 1326 -2574
rect 1320 -2586 1326 -2580
rect 1320 -2592 1326 -2586
rect 1320 -2598 1326 -2592
rect 1320 -2604 1326 -2598
rect 1320 -2610 1326 -2604
rect 1320 -2616 1326 -2610
rect 1320 -2622 1326 -2616
rect 1320 -2628 1326 -2622
rect 1320 -2634 1326 -2628
rect 1320 -2640 1326 -2634
rect 1320 -2646 1326 -2640
rect 1320 -2652 1326 -2646
rect 1320 -2658 1326 -2652
rect 1320 -2664 1326 -2658
rect 1320 -2670 1326 -2664
rect 1320 -2676 1326 -2670
rect 1320 -2682 1326 -2676
rect 1320 -2688 1326 -2682
rect 1320 -2694 1326 -2688
rect 1320 -2700 1326 -2694
rect 1320 -2706 1326 -2700
rect 1320 -2712 1326 -2706
rect 1320 -2718 1326 -2712
rect 1320 -2724 1326 -2718
rect 1320 -2730 1326 -2724
rect 1320 -2736 1326 -2730
rect 1320 -2742 1326 -2736
rect 1320 -2748 1326 -2742
rect 1320 -2754 1326 -2748
rect 1320 -2760 1326 -2754
rect 1320 -2766 1326 -2760
rect 1320 -2772 1326 -2766
rect 1320 -2778 1326 -2772
rect 1320 -2784 1326 -2778
rect 1320 -2790 1326 -2784
rect 1320 -2796 1326 -2790
rect 1320 -2802 1326 -2796
rect 1320 -2808 1326 -2802
rect 1320 -2814 1326 -2808
rect 1320 -2820 1326 -2814
rect 1320 -2826 1326 -2820
rect 1320 -2832 1326 -2826
rect 1320 -2838 1326 -2832
rect 1320 -2844 1326 -2838
rect 1320 -2850 1326 -2844
rect 1320 -2856 1326 -2850
rect 1320 -2862 1326 -2856
rect 1320 -2868 1326 -2862
rect 1320 -2874 1326 -2868
rect 1320 -2880 1326 -2874
rect 1320 -2886 1326 -2880
rect 1320 -2892 1326 -2886
rect 1320 -2898 1326 -2892
rect 1320 -2904 1326 -2898
rect 1320 -2910 1326 -2904
rect 1320 -2916 1326 -2910
rect 1320 -2922 1326 -2916
rect 1320 -2928 1326 -2922
rect 1320 -3012 1326 -3006
rect 1320 -3018 1326 -3012
rect 1320 -3024 1326 -3018
rect 1320 -3030 1326 -3024
rect 1320 -3036 1326 -3030
rect 1320 -3042 1326 -3036
rect 1320 -3048 1326 -3042
rect 1320 -3054 1326 -3048
rect 1320 -3060 1326 -3054
rect 1320 -3066 1326 -3060
rect 1320 -3072 1326 -3066
rect 1320 -3078 1326 -3072
rect 1320 -3084 1326 -3078
rect 1320 -3090 1326 -3084
rect 1320 -3096 1326 -3090
rect 1320 -3102 1326 -3096
rect 1320 -3108 1326 -3102
rect 1320 -3114 1326 -3108
rect 1320 -3120 1326 -3114
rect 1320 -3126 1326 -3120
rect 1320 -3132 1326 -3126
rect 1320 -3138 1326 -3132
rect 1320 -3144 1326 -3138
rect 1320 -3150 1326 -3144
rect 1320 -3156 1326 -3150
rect 1320 -3162 1326 -3156
rect 1320 -3168 1326 -3162
rect 1320 -3174 1326 -3168
rect 1320 -3180 1326 -3174
rect 1320 -3186 1326 -3180
rect 1320 -3192 1326 -3186
rect 1320 -3198 1326 -3192
rect 1320 -3204 1326 -3198
rect 1320 -3210 1326 -3204
rect 1320 -3216 1326 -3210
rect 1320 -3222 1326 -3216
rect 1320 -3228 1326 -3222
rect 1320 -3234 1326 -3228
rect 1320 -3318 1326 -3312
rect 1320 -3324 1326 -3318
rect 1320 -3330 1326 -3324
rect 1320 -3336 1326 -3330
rect 1320 -3342 1326 -3336
rect 1320 -3348 1326 -3342
rect 1320 -3354 1326 -3348
rect 1320 -3360 1326 -3354
rect 1320 -3366 1326 -3360
rect 1320 -3372 1326 -3366
rect 1320 -3378 1326 -3372
rect 1320 -3384 1326 -3378
rect 1320 -3390 1326 -3384
rect 1320 -3396 1326 -3390
rect 1320 -3402 1326 -3396
rect 1320 -3408 1326 -3402
rect 1320 -3414 1326 -3408
rect 1320 -3420 1326 -3414
rect 1320 -3426 1326 -3420
rect 1320 -3432 1326 -3426
rect 1320 -3438 1326 -3432
rect 1320 -3444 1326 -3438
rect 1320 -3450 1326 -3444
rect 1320 -3456 1326 -3450
rect 1320 -3462 1326 -3456
rect 1320 -3468 1326 -3462
rect 1320 -3474 1326 -3468
rect 1320 -3480 1326 -3474
rect 1320 -3486 1326 -3480
rect 1320 -3492 1326 -3486
rect 1320 -3498 1326 -3492
rect 1320 -3504 1326 -3498
rect 1320 -3510 1326 -3504
rect 1320 -3516 1326 -3510
rect 1326 -1110 1332 -1104
rect 1326 -1116 1332 -1110
rect 1326 -1122 1332 -1116
rect 1326 -1128 1332 -1122
rect 1326 -1134 1332 -1128
rect 1326 -1140 1332 -1134
rect 1326 -1146 1332 -1140
rect 1326 -1152 1332 -1146
rect 1326 -1158 1332 -1152
rect 1326 -1164 1332 -1158
rect 1326 -1170 1332 -1164
rect 1326 -1176 1332 -1170
rect 1326 -1182 1332 -1176
rect 1326 -1188 1332 -1182
rect 1326 -1194 1332 -1188
rect 1326 -1200 1332 -1194
rect 1326 -1206 1332 -1200
rect 1326 -1212 1332 -1206
rect 1326 -1218 1332 -1212
rect 1326 -1224 1332 -1218
rect 1326 -1230 1332 -1224
rect 1326 -1236 1332 -1230
rect 1326 -1242 1332 -1236
rect 1326 -1248 1332 -1242
rect 1326 -1254 1332 -1248
rect 1326 -1260 1332 -1254
rect 1326 -1266 1332 -1260
rect 1326 -1272 1332 -1266
rect 1326 -1278 1332 -1272
rect 1326 -1284 1332 -1278
rect 1326 -1290 1332 -1284
rect 1326 -1296 1332 -1290
rect 1326 -1302 1332 -1296
rect 1326 -1308 1332 -1302
rect 1326 -1314 1332 -1308
rect 1326 -1512 1332 -1506
rect 1326 -1518 1332 -1512
rect 1326 -1524 1332 -1518
rect 1326 -1530 1332 -1524
rect 1326 -1536 1332 -1530
rect 1326 -1542 1332 -1536
rect 1326 -1548 1332 -1542
rect 1326 -1554 1332 -1548
rect 1326 -1560 1332 -1554
rect 1326 -1566 1332 -1560
rect 1326 -1572 1332 -1566
rect 1326 -1578 1332 -1572
rect 1326 -1584 1332 -1578
rect 1326 -1590 1332 -1584
rect 1326 -1596 1332 -1590
rect 1326 -1602 1332 -1596
rect 1326 -1608 1332 -1602
rect 1326 -1614 1332 -1608
rect 1326 -1620 1332 -1614
rect 1326 -1626 1332 -1620
rect 1326 -1632 1332 -1626
rect 1326 -1638 1332 -1632
rect 1326 -1644 1332 -1638
rect 1326 -1650 1332 -1644
rect 1326 -1656 1332 -1650
rect 1326 -1662 1332 -1656
rect 1326 -1668 1332 -1662
rect 1326 -1674 1332 -1668
rect 1326 -1680 1332 -1674
rect 1326 -1686 1332 -1680
rect 1326 -1692 1332 -1686
rect 1326 -1698 1332 -1692
rect 1326 -1704 1332 -1698
rect 1326 -1710 1332 -1704
rect 1326 -1716 1332 -1710
rect 1326 -1722 1332 -1716
rect 1326 -1728 1332 -1722
rect 1326 -1734 1332 -1728
rect 1326 -1740 1332 -1734
rect 1326 -1746 1332 -1740
rect 1326 -1752 1332 -1746
rect 1326 -1758 1332 -1752
rect 1326 -1764 1332 -1758
rect 1326 -1770 1332 -1764
rect 1326 -1776 1332 -1770
rect 1326 -1782 1332 -1776
rect 1326 -1788 1332 -1782
rect 1326 -1794 1332 -1788
rect 1326 -1800 1332 -1794
rect 1326 -1806 1332 -1800
rect 1326 -1812 1332 -1806
rect 1326 -1818 1332 -1812
rect 1326 -1824 1332 -1818
rect 1326 -1830 1332 -1824
rect 1326 -1836 1332 -1830
rect 1326 -1842 1332 -1836
rect 1326 -1848 1332 -1842
rect 1326 -1854 1332 -1848
rect 1326 -1860 1332 -1854
rect 1326 -1866 1332 -1860
rect 1326 -1872 1332 -1866
rect 1326 -1878 1332 -1872
rect 1326 -1884 1332 -1878
rect 1326 -1890 1332 -1884
rect 1326 -1896 1332 -1890
rect 1326 -1902 1332 -1896
rect 1326 -1908 1332 -1902
rect 1326 -1914 1332 -1908
rect 1326 -1920 1332 -1914
rect 1326 -1926 1332 -1920
rect 1326 -1932 1332 -1926
rect 1326 -1938 1332 -1932
rect 1326 -1944 1332 -1938
rect 1326 -1950 1332 -1944
rect 1326 -1956 1332 -1950
rect 1326 -1962 1332 -1956
rect 1326 -1968 1332 -1962
rect 1326 -1974 1332 -1968
rect 1326 -1980 1332 -1974
rect 1326 -1986 1332 -1980
rect 1326 -1992 1332 -1986
rect 1326 -1998 1332 -1992
rect 1326 -2004 1332 -1998
rect 1326 -2010 1332 -2004
rect 1326 -2016 1332 -2010
rect 1326 -2022 1332 -2016
rect 1326 -2028 1332 -2022
rect 1326 -2034 1332 -2028
rect 1326 -2040 1332 -2034
rect 1326 -2046 1332 -2040
rect 1326 -2052 1332 -2046
rect 1326 -2058 1332 -2052
rect 1326 -2064 1332 -2058
rect 1326 -2070 1332 -2064
rect 1326 -2076 1332 -2070
rect 1326 -2082 1332 -2076
rect 1326 -2088 1332 -2082
rect 1326 -2094 1332 -2088
rect 1326 -2100 1332 -2094
rect 1326 -2106 1332 -2100
rect 1326 -2112 1332 -2106
rect 1326 -2118 1332 -2112
rect 1326 -2124 1332 -2118
rect 1326 -2130 1332 -2124
rect 1326 -2136 1332 -2130
rect 1326 -2142 1332 -2136
rect 1326 -2148 1332 -2142
rect 1326 -2154 1332 -2148
rect 1326 -2160 1332 -2154
rect 1326 -2166 1332 -2160
rect 1326 -2172 1332 -2166
rect 1326 -2178 1332 -2172
rect 1326 -2184 1332 -2178
rect 1326 -2190 1332 -2184
rect 1326 -2196 1332 -2190
rect 1326 -2202 1332 -2196
rect 1326 -2208 1332 -2202
rect 1326 -2214 1332 -2208
rect 1326 -2220 1332 -2214
rect 1326 -2226 1332 -2220
rect 1326 -2232 1332 -2226
rect 1326 -2238 1332 -2232
rect 1326 -2244 1332 -2238
rect 1326 -2250 1332 -2244
rect 1326 -2256 1332 -2250
rect 1326 -2262 1332 -2256
rect 1326 -2268 1332 -2262
rect 1326 -2274 1332 -2268
rect 1326 -2280 1332 -2274
rect 1326 -2286 1332 -2280
rect 1326 -2292 1332 -2286
rect 1326 -2298 1332 -2292
rect 1326 -2304 1332 -2298
rect 1326 -2310 1332 -2304
rect 1326 -2316 1332 -2310
rect 1326 -2322 1332 -2316
rect 1326 -2328 1332 -2322
rect 1326 -2334 1332 -2328
rect 1326 -2340 1332 -2334
rect 1326 -2346 1332 -2340
rect 1326 -2352 1332 -2346
rect 1326 -2358 1332 -2352
rect 1326 -2364 1332 -2358
rect 1326 -2370 1332 -2364
rect 1326 -2376 1332 -2370
rect 1326 -2382 1332 -2376
rect 1326 -2388 1332 -2382
rect 1326 -2394 1332 -2388
rect 1326 -2400 1332 -2394
rect 1326 -2406 1332 -2400
rect 1326 -2412 1332 -2406
rect 1326 -2418 1332 -2412
rect 1326 -2424 1332 -2418
rect 1326 -2508 1332 -2502
rect 1326 -2514 1332 -2508
rect 1326 -2520 1332 -2514
rect 1326 -2526 1332 -2520
rect 1326 -2532 1332 -2526
rect 1326 -2538 1332 -2532
rect 1326 -2544 1332 -2538
rect 1326 -2550 1332 -2544
rect 1326 -2556 1332 -2550
rect 1326 -2562 1332 -2556
rect 1326 -2568 1332 -2562
rect 1326 -2574 1332 -2568
rect 1326 -2580 1332 -2574
rect 1326 -2586 1332 -2580
rect 1326 -2592 1332 -2586
rect 1326 -2598 1332 -2592
rect 1326 -2604 1332 -2598
rect 1326 -2610 1332 -2604
rect 1326 -2616 1332 -2610
rect 1326 -2622 1332 -2616
rect 1326 -2628 1332 -2622
rect 1326 -2634 1332 -2628
rect 1326 -2640 1332 -2634
rect 1326 -2646 1332 -2640
rect 1326 -2652 1332 -2646
rect 1326 -2658 1332 -2652
rect 1326 -2664 1332 -2658
rect 1326 -2670 1332 -2664
rect 1326 -2676 1332 -2670
rect 1326 -2682 1332 -2676
rect 1326 -2688 1332 -2682
rect 1326 -2694 1332 -2688
rect 1326 -2700 1332 -2694
rect 1326 -2706 1332 -2700
rect 1326 -2712 1332 -2706
rect 1326 -2718 1332 -2712
rect 1326 -2724 1332 -2718
rect 1326 -2730 1332 -2724
rect 1326 -2736 1332 -2730
rect 1326 -2742 1332 -2736
rect 1326 -2748 1332 -2742
rect 1326 -2754 1332 -2748
rect 1326 -2760 1332 -2754
rect 1326 -2766 1332 -2760
rect 1326 -2772 1332 -2766
rect 1326 -2778 1332 -2772
rect 1326 -2784 1332 -2778
rect 1326 -2790 1332 -2784
rect 1326 -2796 1332 -2790
rect 1326 -2802 1332 -2796
rect 1326 -2808 1332 -2802
rect 1326 -2814 1332 -2808
rect 1326 -2820 1332 -2814
rect 1326 -2826 1332 -2820
rect 1326 -2832 1332 -2826
rect 1326 -2838 1332 -2832
rect 1326 -2844 1332 -2838
rect 1326 -2850 1332 -2844
rect 1326 -2856 1332 -2850
rect 1326 -2862 1332 -2856
rect 1326 -2868 1332 -2862
rect 1326 -2874 1332 -2868
rect 1326 -2880 1332 -2874
rect 1326 -2886 1332 -2880
rect 1326 -2892 1332 -2886
rect 1326 -2898 1332 -2892
rect 1326 -2904 1332 -2898
rect 1326 -2910 1332 -2904
rect 1326 -2916 1332 -2910
rect 1326 -2922 1332 -2916
rect 1326 -2928 1332 -2922
rect 1326 -3012 1332 -3006
rect 1326 -3018 1332 -3012
rect 1326 -3024 1332 -3018
rect 1326 -3030 1332 -3024
rect 1326 -3036 1332 -3030
rect 1326 -3042 1332 -3036
rect 1326 -3048 1332 -3042
rect 1326 -3054 1332 -3048
rect 1326 -3060 1332 -3054
rect 1326 -3066 1332 -3060
rect 1326 -3072 1332 -3066
rect 1326 -3078 1332 -3072
rect 1326 -3084 1332 -3078
rect 1326 -3090 1332 -3084
rect 1326 -3096 1332 -3090
rect 1326 -3102 1332 -3096
rect 1326 -3108 1332 -3102
rect 1326 -3114 1332 -3108
rect 1326 -3120 1332 -3114
rect 1326 -3126 1332 -3120
rect 1326 -3132 1332 -3126
rect 1326 -3138 1332 -3132
rect 1326 -3144 1332 -3138
rect 1326 -3150 1332 -3144
rect 1326 -3156 1332 -3150
rect 1326 -3162 1332 -3156
rect 1326 -3168 1332 -3162
rect 1326 -3174 1332 -3168
rect 1326 -3180 1332 -3174
rect 1326 -3186 1332 -3180
rect 1326 -3192 1332 -3186
rect 1326 -3198 1332 -3192
rect 1326 -3204 1332 -3198
rect 1326 -3210 1332 -3204
rect 1326 -3216 1332 -3210
rect 1326 -3222 1332 -3216
rect 1326 -3228 1332 -3222
rect 1326 -3234 1332 -3228
rect 1326 -3312 1332 -3306
rect 1326 -3318 1332 -3312
rect 1326 -3324 1332 -3318
rect 1326 -3330 1332 -3324
rect 1326 -3336 1332 -3330
rect 1326 -3342 1332 -3336
rect 1326 -3348 1332 -3342
rect 1326 -3354 1332 -3348
rect 1326 -3360 1332 -3354
rect 1326 -3366 1332 -3360
rect 1326 -3372 1332 -3366
rect 1326 -3378 1332 -3372
rect 1326 -3384 1332 -3378
rect 1326 -3390 1332 -3384
rect 1326 -3396 1332 -3390
rect 1326 -3402 1332 -3396
rect 1326 -3408 1332 -3402
rect 1326 -3414 1332 -3408
rect 1326 -3420 1332 -3414
rect 1326 -3426 1332 -3420
rect 1326 -3432 1332 -3426
rect 1326 -3438 1332 -3432
rect 1326 -3444 1332 -3438
rect 1326 -3450 1332 -3444
rect 1326 -3456 1332 -3450
rect 1326 -3462 1332 -3456
rect 1326 -3468 1332 -3462
rect 1326 -3474 1332 -3468
rect 1326 -3480 1332 -3474
rect 1326 -3486 1332 -3480
rect 1326 -3492 1332 -3486
rect 1326 -3498 1332 -3492
rect 1326 -3504 1332 -3498
rect 1326 -3510 1332 -3504
rect 1326 -3516 1332 -3510
rect 1332 -1110 1338 -1104
rect 1332 -1116 1338 -1110
rect 1332 -1122 1338 -1116
rect 1332 -1128 1338 -1122
rect 1332 -1134 1338 -1128
rect 1332 -1140 1338 -1134
rect 1332 -1146 1338 -1140
rect 1332 -1152 1338 -1146
rect 1332 -1158 1338 -1152
rect 1332 -1164 1338 -1158
rect 1332 -1170 1338 -1164
rect 1332 -1176 1338 -1170
rect 1332 -1182 1338 -1176
rect 1332 -1188 1338 -1182
rect 1332 -1194 1338 -1188
rect 1332 -1200 1338 -1194
rect 1332 -1206 1338 -1200
rect 1332 -1212 1338 -1206
rect 1332 -1218 1338 -1212
rect 1332 -1224 1338 -1218
rect 1332 -1230 1338 -1224
rect 1332 -1236 1338 -1230
rect 1332 -1242 1338 -1236
rect 1332 -1248 1338 -1242
rect 1332 -1254 1338 -1248
rect 1332 -1260 1338 -1254
rect 1332 -1266 1338 -1260
rect 1332 -1272 1338 -1266
rect 1332 -1278 1338 -1272
rect 1332 -1284 1338 -1278
rect 1332 -1290 1338 -1284
rect 1332 -1296 1338 -1290
rect 1332 -1302 1338 -1296
rect 1332 -1308 1338 -1302
rect 1332 -1314 1338 -1308
rect 1332 -1500 1338 -1494
rect 1332 -1506 1338 -1500
rect 1332 -1512 1338 -1506
rect 1332 -1518 1338 -1512
rect 1332 -1524 1338 -1518
rect 1332 -1530 1338 -1524
rect 1332 -1536 1338 -1530
rect 1332 -1542 1338 -1536
rect 1332 -1548 1338 -1542
rect 1332 -1554 1338 -1548
rect 1332 -1560 1338 -1554
rect 1332 -1566 1338 -1560
rect 1332 -1572 1338 -1566
rect 1332 -1578 1338 -1572
rect 1332 -1584 1338 -1578
rect 1332 -1590 1338 -1584
rect 1332 -1596 1338 -1590
rect 1332 -1602 1338 -1596
rect 1332 -1608 1338 -1602
rect 1332 -1614 1338 -1608
rect 1332 -1620 1338 -1614
rect 1332 -1626 1338 -1620
rect 1332 -1632 1338 -1626
rect 1332 -1638 1338 -1632
rect 1332 -1644 1338 -1638
rect 1332 -1650 1338 -1644
rect 1332 -1656 1338 -1650
rect 1332 -1662 1338 -1656
rect 1332 -1668 1338 -1662
rect 1332 -1674 1338 -1668
rect 1332 -1680 1338 -1674
rect 1332 -1686 1338 -1680
rect 1332 -1692 1338 -1686
rect 1332 -1698 1338 -1692
rect 1332 -1704 1338 -1698
rect 1332 -1710 1338 -1704
rect 1332 -1716 1338 -1710
rect 1332 -1722 1338 -1716
rect 1332 -1728 1338 -1722
rect 1332 -1734 1338 -1728
rect 1332 -1740 1338 -1734
rect 1332 -1746 1338 -1740
rect 1332 -1752 1338 -1746
rect 1332 -1758 1338 -1752
rect 1332 -1764 1338 -1758
rect 1332 -1770 1338 -1764
rect 1332 -1776 1338 -1770
rect 1332 -1782 1338 -1776
rect 1332 -1788 1338 -1782
rect 1332 -1794 1338 -1788
rect 1332 -1800 1338 -1794
rect 1332 -1806 1338 -1800
rect 1332 -1812 1338 -1806
rect 1332 -1818 1338 -1812
rect 1332 -1824 1338 -1818
rect 1332 -1830 1338 -1824
rect 1332 -1836 1338 -1830
rect 1332 -1842 1338 -1836
rect 1332 -1848 1338 -1842
rect 1332 -1854 1338 -1848
rect 1332 -1860 1338 -1854
rect 1332 -1866 1338 -1860
rect 1332 -1872 1338 -1866
rect 1332 -1878 1338 -1872
rect 1332 -1884 1338 -1878
rect 1332 -1890 1338 -1884
rect 1332 -1896 1338 -1890
rect 1332 -1902 1338 -1896
rect 1332 -1908 1338 -1902
rect 1332 -1914 1338 -1908
rect 1332 -1920 1338 -1914
rect 1332 -1926 1338 -1920
rect 1332 -1932 1338 -1926
rect 1332 -1938 1338 -1932
rect 1332 -1944 1338 -1938
rect 1332 -1950 1338 -1944
rect 1332 -1956 1338 -1950
rect 1332 -1962 1338 -1956
rect 1332 -1968 1338 -1962
rect 1332 -1974 1338 -1968
rect 1332 -1980 1338 -1974
rect 1332 -1986 1338 -1980
rect 1332 -1992 1338 -1986
rect 1332 -1998 1338 -1992
rect 1332 -2004 1338 -1998
rect 1332 -2010 1338 -2004
rect 1332 -2016 1338 -2010
rect 1332 -2022 1338 -2016
rect 1332 -2028 1338 -2022
rect 1332 -2034 1338 -2028
rect 1332 -2040 1338 -2034
rect 1332 -2046 1338 -2040
rect 1332 -2052 1338 -2046
rect 1332 -2058 1338 -2052
rect 1332 -2064 1338 -2058
rect 1332 -2070 1338 -2064
rect 1332 -2076 1338 -2070
rect 1332 -2082 1338 -2076
rect 1332 -2088 1338 -2082
rect 1332 -2094 1338 -2088
rect 1332 -2100 1338 -2094
rect 1332 -2106 1338 -2100
rect 1332 -2112 1338 -2106
rect 1332 -2118 1338 -2112
rect 1332 -2124 1338 -2118
rect 1332 -2130 1338 -2124
rect 1332 -2136 1338 -2130
rect 1332 -2142 1338 -2136
rect 1332 -2148 1338 -2142
rect 1332 -2154 1338 -2148
rect 1332 -2160 1338 -2154
rect 1332 -2166 1338 -2160
rect 1332 -2172 1338 -2166
rect 1332 -2178 1338 -2172
rect 1332 -2184 1338 -2178
rect 1332 -2190 1338 -2184
rect 1332 -2196 1338 -2190
rect 1332 -2202 1338 -2196
rect 1332 -2208 1338 -2202
rect 1332 -2214 1338 -2208
rect 1332 -2220 1338 -2214
rect 1332 -2226 1338 -2220
rect 1332 -2232 1338 -2226
rect 1332 -2238 1338 -2232
rect 1332 -2244 1338 -2238
rect 1332 -2250 1338 -2244
rect 1332 -2256 1338 -2250
rect 1332 -2262 1338 -2256
rect 1332 -2268 1338 -2262
rect 1332 -2274 1338 -2268
rect 1332 -2280 1338 -2274
rect 1332 -2286 1338 -2280
rect 1332 -2292 1338 -2286
rect 1332 -2298 1338 -2292
rect 1332 -2304 1338 -2298
rect 1332 -2310 1338 -2304
rect 1332 -2316 1338 -2310
rect 1332 -2322 1338 -2316
rect 1332 -2328 1338 -2322
rect 1332 -2334 1338 -2328
rect 1332 -2340 1338 -2334
rect 1332 -2346 1338 -2340
rect 1332 -2352 1338 -2346
rect 1332 -2358 1338 -2352
rect 1332 -2364 1338 -2358
rect 1332 -2370 1338 -2364
rect 1332 -2376 1338 -2370
rect 1332 -2382 1338 -2376
rect 1332 -2388 1338 -2382
rect 1332 -2394 1338 -2388
rect 1332 -2400 1338 -2394
rect 1332 -2406 1338 -2400
rect 1332 -2412 1338 -2406
rect 1332 -2418 1338 -2412
rect 1332 -2496 1338 -2490
rect 1332 -2502 1338 -2496
rect 1332 -2508 1338 -2502
rect 1332 -2514 1338 -2508
rect 1332 -2520 1338 -2514
rect 1332 -2526 1338 -2520
rect 1332 -2532 1338 -2526
rect 1332 -2538 1338 -2532
rect 1332 -2544 1338 -2538
rect 1332 -2550 1338 -2544
rect 1332 -2556 1338 -2550
rect 1332 -2562 1338 -2556
rect 1332 -2568 1338 -2562
rect 1332 -2574 1338 -2568
rect 1332 -2580 1338 -2574
rect 1332 -2586 1338 -2580
rect 1332 -2592 1338 -2586
rect 1332 -2598 1338 -2592
rect 1332 -2604 1338 -2598
rect 1332 -2610 1338 -2604
rect 1332 -2616 1338 -2610
rect 1332 -2622 1338 -2616
rect 1332 -2628 1338 -2622
rect 1332 -2634 1338 -2628
rect 1332 -2640 1338 -2634
rect 1332 -2646 1338 -2640
rect 1332 -2652 1338 -2646
rect 1332 -2658 1338 -2652
rect 1332 -2664 1338 -2658
rect 1332 -2670 1338 -2664
rect 1332 -2676 1338 -2670
rect 1332 -2682 1338 -2676
rect 1332 -2688 1338 -2682
rect 1332 -2694 1338 -2688
rect 1332 -2700 1338 -2694
rect 1332 -2706 1338 -2700
rect 1332 -2712 1338 -2706
rect 1332 -2718 1338 -2712
rect 1332 -2724 1338 -2718
rect 1332 -2730 1338 -2724
rect 1332 -2736 1338 -2730
rect 1332 -2742 1338 -2736
rect 1332 -2748 1338 -2742
rect 1332 -2754 1338 -2748
rect 1332 -2760 1338 -2754
rect 1332 -2766 1338 -2760
rect 1332 -2772 1338 -2766
rect 1332 -2778 1338 -2772
rect 1332 -2784 1338 -2778
rect 1332 -2790 1338 -2784
rect 1332 -2796 1338 -2790
rect 1332 -2802 1338 -2796
rect 1332 -2808 1338 -2802
rect 1332 -2814 1338 -2808
rect 1332 -2820 1338 -2814
rect 1332 -2826 1338 -2820
rect 1332 -2832 1338 -2826
rect 1332 -2838 1338 -2832
rect 1332 -2844 1338 -2838
rect 1332 -2850 1338 -2844
rect 1332 -2856 1338 -2850
rect 1332 -2862 1338 -2856
rect 1332 -2868 1338 -2862
rect 1332 -2874 1338 -2868
rect 1332 -2880 1338 -2874
rect 1332 -2886 1338 -2880
rect 1332 -2892 1338 -2886
rect 1332 -2898 1338 -2892
rect 1332 -2904 1338 -2898
rect 1332 -2910 1338 -2904
rect 1332 -2916 1338 -2910
rect 1332 -2922 1338 -2916
rect 1332 -3006 1338 -3000
rect 1332 -3012 1338 -3006
rect 1332 -3018 1338 -3012
rect 1332 -3024 1338 -3018
rect 1332 -3030 1338 -3024
rect 1332 -3036 1338 -3030
rect 1332 -3042 1338 -3036
rect 1332 -3048 1338 -3042
rect 1332 -3054 1338 -3048
rect 1332 -3060 1338 -3054
rect 1332 -3066 1338 -3060
rect 1332 -3072 1338 -3066
rect 1332 -3078 1338 -3072
rect 1332 -3084 1338 -3078
rect 1332 -3090 1338 -3084
rect 1332 -3096 1338 -3090
rect 1332 -3102 1338 -3096
rect 1332 -3108 1338 -3102
rect 1332 -3114 1338 -3108
rect 1332 -3120 1338 -3114
rect 1332 -3126 1338 -3120
rect 1332 -3132 1338 -3126
rect 1332 -3138 1338 -3132
rect 1332 -3144 1338 -3138
rect 1332 -3150 1338 -3144
rect 1332 -3156 1338 -3150
rect 1332 -3162 1338 -3156
rect 1332 -3168 1338 -3162
rect 1332 -3174 1338 -3168
rect 1332 -3180 1338 -3174
rect 1332 -3186 1338 -3180
rect 1332 -3192 1338 -3186
rect 1332 -3198 1338 -3192
rect 1332 -3204 1338 -3198
rect 1332 -3210 1338 -3204
rect 1332 -3216 1338 -3210
rect 1332 -3222 1338 -3216
rect 1332 -3228 1338 -3222
rect 1332 -3234 1338 -3228
rect 1332 -3312 1338 -3306
rect 1332 -3318 1338 -3312
rect 1332 -3324 1338 -3318
rect 1332 -3330 1338 -3324
rect 1332 -3336 1338 -3330
rect 1332 -3342 1338 -3336
rect 1332 -3348 1338 -3342
rect 1332 -3354 1338 -3348
rect 1332 -3360 1338 -3354
rect 1332 -3366 1338 -3360
rect 1332 -3372 1338 -3366
rect 1332 -3378 1338 -3372
rect 1332 -3384 1338 -3378
rect 1332 -3390 1338 -3384
rect 1332 -3396 1338 -3390
rect 1332 -3402 1338 -3396
rect 1332 -3408 1338 -3402
rect 1332 -3414 1338 -3408
rect 1332 -3420 1338 -3414
rect 1332 -3426 1338 -3420
rect 1332 -3432 1338 -3426
rect 1332 -3438 1338 -3432
rect 1332 -3444 1338 -3438
rect 1332 -3450 1338 -3444
rect 1332 -3456 1338 -3450
rect 1332 -3462 1338 -3456
rect 1332 -3468 1338 -3462
rect 1332 -3474 1338 -3468
rect 1332 -3480 1338 -3474
rect 1332 -3486 1338 -3480
rect 1332 -3492 1338 -3486
rect 1332 -3498 1338 -3492
rect 1332 -3504 1338 -3498
rect 1332 -3510 1338 -3504
rect 1332 -3516 1338 -3510
rect 1338 -1110 1344 -1104
rect 1338 -1116 1344 -1110
rect 1338 -1122 1344 -1116
rect 1338 -1128 1344 -1122
rect 1338 -1134 1344 -1128
rect 1338 -1140 1344 -1134
rect 1338 -1146 1344 -1140
rect 1338 -1152 1344 -1146
rect 1338 -1158 1344 -1152
rect 1338 -1164 1344 -1158
rect 1338 -1170 1344 -1164
rect 1338 -1176 1344 -1170
rect 1338 -1182 1344 -1176
rect 1338 -1188 1344 -1182
rect 1338 -1194 1344 -1188
rect 1338 -1200 1344 -1194
rect 1338 -1206 1344 -1200
rect 1338 -1212 1344 -1206
rect 1338 -1218 1344 -1212
rect 1338 -1224 1344 -1218
rect 1338 -1230 1344 -1224
rect 1338 -1236 1344 -1230
rect 1338 -1242 1344 -1236
rect 1338 -1248 1344 -1242
rect 1338 -1254 1344 -1248
rect 1338 -1260 1344 -1254
rect 1338 -1266 1344 -1260
rect 1338 -1272 1344 -1266
rect 1338 -1278 1344 -1272
rect 1338 -1284 1344 -1278
rect 1338 -1290 1344 -1284
rect 1338 -1296 1344 -1290
rect 1338 -1302 1344 -1296
rect 1338 -1308 1344 -1302
rect 1338 -1314 1344 -1308
rect 1338 -1488 1344 -1482
rect 1338 -1494 1344 -1488
rect 1338 -1500 1344 -1494
rect 1338 -1506 1344 -1500
rect 1338 -1512 1344 -1506
rect 1338 -1518 1344 -1512
rect 1338 -1524 1344 -1518
rect 1338 -1530 1344 -1524
rect 1338 -1536 1344 -1530
rect 1338 -1542 1344 -1536
rect 1338 -1548 1344 -1542
rect 1338 -1554 1344 -1548
rect 1338 -1560 1344 -1554
rect 1338 -1566 1344 -1560
rect 1338 -1572 1344 -1566
rect 1338 -1578 1344 -1572
rect 1338 -1584 1344 -1578
rect 1338 -1590 1344 -1584
rect 1338 -1596 1344 -1590
rect 1338 -1602 1344 -1596
rect 1338 -1608 1344 -1602
rect 1338 -1614 1344 -1608
rect 1338 -1620 1344 -1614
rect 1338 -1626 1344 -1620
rect 1338 -1632 1344 -1626
rect 1338 -1638 1344 -1632
rect 1338 -1644 1344 -1638
rect 1338 -1650 1344 -1644
rect 1338 -1656 1344 -1650
rect 1338 -1662 1344 -1656
rect 1338 -1668 1344 -1662
rect 1338 -1674 1344 -1668
rect 1338 -1680 1344 -1674
rect 1338 -1686 1344 -1680
rect 1338 -1692 1344 -1686
rect 1338 -1698 1344 -1692
rect 1338 -1704 1344 -1698
rect 1338 -1710 1344 -1704
rect 1338 -1716 1344 -1710
rect 1338 -1722 1344 -1716
rect 1338 -1728 1344 -1722
rect 1338 -1734 1344 -1728
rect 1338 -1740 1344 -1734
rect 1338 -1746 1344 -1740
rect 1338 -1752 1344 -1746
rect 1338 -1758 1344 -1752
rect 1338 -1764 1344 -1758
rect 1338 -1770 1344 -1764
rect 1338 -1776 1344 -1770
rect 1338 -1782 1344 -1776
rect 1338 -1788 1344 -1782
rect 1338 -1794 1344 -1788
rect 1338 -1800 1344 -1794
rect 1338 -1806 1344 -1800
rect 1338 -1812 1344 -1806
rect 1338 -1818 1344 -1812
rect 1338 -1824 1344 -1818
rect 1338 -1830 1344 -1824
rect 1338 -1836 1344 -1830
rect 1338 -1842 1344 -1836
rect 1338 -1848 1344 -1842
rect 1338 -1854 1344 -1848
rect 1338 -1860 1344 -1854
rect 1338 -1866 1344 -1860
rect 1338 -1872 1344 -1866
rect 1338 -1878 1344 -1872
rect 1338 -1884 1344 -1878
rect 1338 -1890 1344 -1884
rect 1338 -1896 1344 -1890
rect 1338 -1902 1344 -1896
rect 1338 -1908 1344 -1902
rect 1338 -1914 1344 -1908
rect 1338 -1920 1344 -1914
rect 1338 -1926 1344 -1920
rect 1338 -1932 1344 -1926
rect 1338 -1938 1344 -1932
rect 1338 -1944 1344 -1938
rect 1338 -1950 1344 -1944
rect 1338 -1956 1344 -1950
rect 1338 -1962 1344 -1956
rect 1338 -1968 1344 -1962
rect 1338 -1974 1344 -1968
rect 1338 -1980 1344 -1974
rect 1338 -1986 1344 -1980
rect 1338 -1992 1344 -1986
rect 1338 -1998 1344 -1992
rect 1338 -2004 1344 -1998
rect 1338 -2010 1344 -2004
rect 1338 -2016 1344 -2010
rect 1338 -2022 1344 -2016
rect 1338 -2028 1344 -2022
rect 1338 -2034 1344 -2028
rect 1338 -2040 1344 -2034
rect 1338 -2046 1344 -2040
rect 1338 -2052 1344 -2046
rect 1338 -2058 1344 -2052
rect 1338 -2064 1344 -2058
rect 1338 -2070 1344 -2064
rect 1338 -2076 1344 -2070
rect 1338 -2082 1344 -2076
rect 1338 -2088 1344 -2082
rect 1338 -2094 1344 -2088
rect 1338 -2100 1344 -2094
rect 1338 -2106 1344 -2100
rect 1338 -2112 1344 -2106
rect 1338 -2118 1344 -2112
rect 1338 -2124 1344 -2118
rect 1338 -2130 1344 -2124
rect 1338 -2136 1344 -2130
rect 1338 -2142 1344 -2136
rect 1338 -2148 1344 -2142
rect 1338 -2154 1344 -2148
rect 1338 -2160 1344 -2154
rect 1338 -2166 1344 -2160
rect 1338 -2172 1344 -2166
rect 1338 -2178 1344 -2172
rect 1338 -2184 1344 -2178
rect 1338 -2190 1344 -2184
rect 1338 -2196 1344 -2190
rect 1338 -2202 1344 -2196
rect 1338 -2208 1344 -2202
rect 1338 -2214 1344 -2208
rect 1338 -2220 1344 -2214
rect 1338 -2226 1344 -2220
rect 1338 -2232 1344 -2226
rect 1338 -2238 1344 -2232
rect 1338 -2244 1344 -2238
rect 1338 -2250 1344 -2244
rect 1338 -2256 1344 -2250
rect 1338 -2262 1344 -2256
rect 1338 -2268 1344 -2262
rect 1338 -2274 1344 -2268
rect 1338 -2280 1344 -2274
rect 1338 -2286 1344 -2280
rect 1338 -2292 1344 -2286
rect 1338 -2298 1344 -2292
rect 1338 -2304 1344 -2298
rect 1338 -2310 1344 -2304
rect 1338 -2316 1344 -2310
rect 1338 -2322 1344 -2316
rect 1338 -2328 1344 -2322
rect 1338 -2334 1344 -2328
rect 1338 -2340 1344 -2334
rect 1338 -2346 1344 -2340
rect 1338 -2352 1344 -2346
rect 1338 -2358 1344 -2352
rect 1338 -2364 1344 -2358
rect 1338 -2370 1344 -2364
rect 1338 -2376 1344 -2370
rect 1338 -2382 1344 -2376
rect 1338 -2388 1344 -2382
rect 1338 -2394 1344 -2388
rect 1338 -2400 1344 -2394
rect 1338 -2406 1344 -2400
rect 1338 -2490 1344 -2484
rect 1338 -2496 1344 -2490
rect 1338 -2502 1344 -2496
rect 1338 -2508 1344 -2502
rect 1338 -2514 1344 -2508
rect 1338 -2520 1344 -2514
rect 1338 -2526 1344 -2520
rect 1338 -2532 1344 -2526
rect 1338 -2538 1344 -2532
rect 1338 -2544 1344 -2538
rect 1338 -2550 1344 -2544
rect 1338 -2556 1344 -2550
rect 1338 -2562 1344 -2556
rect 1338 -2568 1344 -2562
rect 1338 -2574 1344 -2568
rect 1338 -2580 1344 -2574
rect 1338 -2586 1344 -2580
rect 1338 -2592 1344 -2586
rect 1338 -2598 1344 -2592
rect 1338 -2604 1344 -2598
rect 1338 -2610 1344 -2604
rect 1338 -2616 1344 -2610
rect 1338 -2622 1344 -2616
rect 1338 -2628 1344 -2622
rect 1338 -2634 1344 -2628
rect 1338 -2640 1344 -2634
rect 1338 -2646 1344 -2640
rect 1338 -2652 1344 -2646
rect 1338 -2658 1344 -2652
rect 1338 -2664 1344 -2658
rect 1338 -2670 1344 -2664
rect 1338 -2676 1344 -2670
rect 1338 -2682 1344 -2676
rect 1338 -2688 1344 -2682
rect 1338 -2694 1344 -2688
rect 1338 -2700 1344 -2694
rect 1338 -2706 1344 -2700
rect 1338 -2712 1344 -2706
rect 1338 -2718 1344 -2712
rect 1338 -2724 1344 -2718
rect 1338 -2730 1344 -2724
rect 1338 -2736 1344 -2730
rect 1338 -2742 1344 -2736
rect 1338 -2748 1344 -2742
rect 1338 -2754 1344 -2748
rect 1338 -2760 1344 -2754
rect 1338 -2766 1344 -2760
rect 1338 -2772 1344 -2766
rect 1338 -2778 1344 -2772
rect 1338 -2784 1344 -2778
rect 1338 -2790 1344 -2784
rect 1338 -2796 1344 -2790
rect 1338 -2802 1344 -2796
rect 1338 -2808 1344 -2802
rect 1338 -2814 1344 -2808
rect 1338 -2820 1344 -2814
rect 1338 -2826 1344 -2820
rect 1338 -2832 1344 -2826
rect 1338 -2838 1344 -2832
rect 1338 -2844 1344 -2838
rect 1338 -2850 1344 -2844
rect 1338 -2856 1344 -2850
rect 1338 -2862 1344 -2856
rect 1338 -2868 1344 -2862
rect 1338 -2874 1344 -2868
rect 1338 -2880 1344 -2874
rect 1338 -2886 1344 -2880
rect 1338 -2892 1344 -2886
rect 1338 -2898 1344 -2892
rect 1338 -2904 1344 -2898
rect 1338 -2910 1344 -2904
rect 1338 -2916 1344 -2910
rect 1338 -3000 1344 -2994
rect 1338 -3006 1344 -3000
rect 1338 -3012 1344 -3006
rect 1338 -3018 1344 -3012
rect 1338 -3024 1344 -3018
rect 1338 -3030 1344 -3024
rect 1338 -3036 1344 -3030
rect 1338 -3042 1344 -3036
rect 1338 -3048 1344 -3042
rect 1338 -3054 1344 -3048
rect 1338 -3060 1344 -3054
rect 1338 -3066 1344 -3060
rect 1338 -3072 1344 -3066
rect 1338 -3078 1344 -3072
rect 1338 -3084 1344 -3078
rect 1338 -3090 1344 -3084
rect 1338 -3096 1344 -3090
rect 1338 -3102 1344 -3096
rect 1338 -3108 1344 -3102
rect 1338 -3114 1344 -3108
rect 1338 -3120 1344 -3114
rect 1338 -3126 1344 -3120
rect 1338 -3132 1344 -3126
rect 1338 -3138 1344 -3132
rect 1338 -3144 1344 -3138
rect 1338 -3150 1344 -3144
rect 1338 -3156 1344 -3150
rect 1338 -3162 1344 -3156
rect 1338 -3168 1344 -3162
rect 1338 -3174 1344 -3168
rect 1338 -3180 1344 -3174
rect 1338 -3186 1344 -3180
rect 1338 -3192 1344 -3186
rect 1338 -3198 1344 -3192
rect 1338 -3204 1344 -3198
rect 1338 -3210 1344 -3204
rect 1338 -3216 1344 -3210
rect 1338 -3222 1344 -3216
rect 1338 -3228 1344 -3222
rect 1338 -3234 1344 -3228
rect 1338 -3312 1344 -3306
rect 1338 -3318 1344 -3312
rect 1338 -3324 1344 -3318
rect 1338 -3330 1344 -3324
rect 1338 -3336 1344 -3330
rect 1338 -3342 1344 -3336
rect 1338 -3348 1344 -3342
rect 1338 -3354 1344 -3348
rect 1338 -3360 1344 -3354
rect 1338 -3366 1344 -3360
rect 1338 -3372 1344 -3366
rect 1338 -3378 1344 -3372
rect 1338 -3384 1344 -3378
rect 1338 -3390 1344 -3384
rect 1338 -3396 1344 -3390
rect 1338 -3402 1344 -3396
rect 1338 -3408 1344 -3402
rect 1338 -3414 1344 -3408
rect 1338 -3420 1344 -3414
rect 1338 -3426 1344 -3420
rect 1338 -3432 1344 -3426
rect 1338 -3438 1344 -3432
rect 1338 -3444 1344 -3438
rect 1338 -3450 1344 -3444
rect 1338 -3456 1344 -3450
rect 1338 -3462 1344 -3456
rect 1338 -3468 1344 -3462
rect 1338 -3474 1344 -3468
rect 1338 -3480 1344 -3474
rect 1338 -3486 1344 -3480
rect 1338 -3492 1344 -3486
rect 1338 -3498 1344 -3492
rect 1338 -3504 1344 -3498
rect 1338 -3510 1344 -3504
rect 1338 -3516 1344 -3510
rect 1344 -1110 1350 -1104
rect 1344 -1116 1350 -1110
rect 1344 -1122 1350 -1116
rect 1344 -1128 1350 -1122
rect 1344 -1134 1350 -1128
rect 1344 -1140 1350 -1134
rect 1344 -1146 1350 -1140
rect 1344 -1152 1350 -1146
rect 1344 -1158 1350 -1152
rect 1344 -1164 1350 -1158
rect 1344 -1170 1350 -1164
rect 1344 -1176 1350 -1170
rect 1344 -1182 1350 -1176
rect 1344 -1188 1350 -1182
rect 1344 -1194 1350 -1188
rect 1344 -1200 1350 -1194
rect 1344 -1206 1350 -1200
rect 1344 -1212 1350 -1206
rect 1344 -1218 1350 -1212
rect 1344 -1224 1350 -1218
rect 1344 -1230 1350 -1224
rect 1344 -1236 1350 -1230
rect 1344 -1242 1350 -1236
rect 1344 -1248 1350 -1242
rect 1344 -1254 1350 -1248
rect 1344 -1260 1350 -1254
rect 1344 -1266 1350 -1260
rect 1344 -1272 1350 -1266
rect 1344 -1278 1350 -1272
rect 1344 -1284 1350 -1278
rect 1344 -1290 1350 -1284
rect 1344 -1296 1350 -1290
rect 1344 -1302 1350 -1296
rect 1344 -1308 1350 -1302
rect 1344 -1314 1350 -1308
rect 1344 -1476 1350 -1470
rect 1344 -1482 1350 -1476
rect 1344 -1488 1350 -1482
rect 1344 -1494 1350 -1488
rect 1344 -1500 1350 -1494
rect 1344 -1506 1350 -1500
rect 1344 -1512 1350 -1506
rect 1344 -1518 1350 -1512
rect 1344 -1524 1350 -1518
rect 1344 -1530 1350 -1524
rect 1344 -1536 1350 -1530
rect 1344 -1542 1350 -1536
rect 1344 -1548 1350 -1542
rect 1344 -1554 1350 -1548
rect 1344 -1560 1350 -1554
rect 1344 -1566 1350 -1560
rect 1344 -1572 1350 -1566
rect 1344 -1578 1350 -1572
rect 1344 -1584 1350 -1578
rect 1344 -1590 1350 -1584
rect 1344 -1596 1350 -1590
rect 1344 -1602 1350 -1596
rect 1344 -1608 1350 -1602
rect 1344 -1614 1350 -1608
rect 1344 -1620 1350 -1614
rect 1344 -1626 1350 -1620
rect 1344 -1632 1350 -1626
rect 1344 -1638 1350 -1632
rect 1344 -1644 1350 -1638
rect 1344 -1650 1350 -1644
rect 1344 -1656 1350 -1650
rect 1344 -1662 1350 -1656
rect 1344 -1668 1350 -1662
rect 1344 -1674 1350 -1668
rect 1344 -1680 1350 -1674
rect 1344 -1686 1350 -1680
rect 1344 -1692 1350 -1686
rect 1344 -1698 1350 -1692
rect 1344 -1704 1350 -1698
rect 1344 -1710 1350 -1704
rect 1344 -1716 1350 -1710
rect 1344 -1722 1350 -1716
rect 1344 -1728 1350 -1722
rect 1344 -1734 1350 -1728
rect 1344 -1740 1350 -1734
rect 1344 -1746 1350 -1740
rect 1344 -1752 1350 -1746
rect 1344 -1758 1350 -1752
rect 1344 -1764 1350 -1758
rect 1344 -1770 1350 -1764
rect 1344 -1776 1350 -1770
rect 1344 -1782 1350 -1776
rect 1344 -1788 1350 -1782
rect 1344 -1794 1350 -1788
rect 1344 -1800 1350 -1794
rect 1344 -1806 1350 -1800
rect 1344 -1812 1350 -1806
rect 1344 -1818 1350 -1812
rect 1344 -1824 1350 -1818
rect 1344 -1830 1350 -1824
rect 1344 -1836 1350 -1830
rect 1344 -1842 1350 -1836
rect 1344 -1848 1350 -1842
rect 1344 -1854 1350 -1848
rect 1344 -1860 1350 -1854
rect 1344 -1866 1350 -1860
rect 1344 -1872 1350 -1866
rect 1344 -1878 1350 -1872
rect 1344 -1884 1350 -1878
rect 1344 -1890 1350 -1884
rect 1344 -1896 1350 -1890
rect 1344 -1902 1350 -1896
rect 1344 -1908 1350 -1902
rect 1344 -1914 1350 -1908
rect 1344 -1920 1350 -1914
rect 1344 -1926 1350 -1920
rect 1344 -1932 1350 -1926
rect 1344 -1938 1350 -1932
rect 1344 -1944 1350 -1938
rect 1344 -1950 1350 -1944
rect 1344 -1956 1350 -1950
rect 1344 -1962 1350 -1956
rect 1344 -1968 1350 -1962
rect 1344 -1974 1350 -1968
rect 1344 -1980 1350 -1974
rect 1344 -1986 1350 -1980
rect 1344 -1992 1350 -1986
rect 1344 -1998 1350 -1992
rect 1344 -2004 1350 -1998
rect 1344 -2010 1350 -2004
rect 1344 -2016 1350 -2010
rect 1344 -2022 1350 -2016
rect 1344 -2028 1350 -2022
rect 1344 -2034 1350 -2028
rect 1344 -2040 1350 -2034
rect 1344 -2046 1350 -2040
rect 1344 -2052 1350 -2046
rect 1344 -2058 1350 -2052
rect 1344 -2064 1350 -2058
rect 1344 -2070 1350 -2064
rect 1344 -2076 1350 -2070
rect 1344 -2082 1350 -2076
rect 1344 -2088 1350 -2082
rect 1344 -2094 1350 -2088
rect 1344 -2100 1350 -2094
rect 1344 -2106 1350 -2100
rect 1344 -2112 1350 -2106
rect 1344 -2118 1350 -2112
rect 1344 -2124 1350 -2118
rect 1344 -2130 1350 -2124
rect 1344 -2136 1350 -2130
rect 1344 -2142 1350 -2136
rect 1344 -2148 1350 -2142
rect 1344 -2154 1350 -2148
rect 1344 -2160 1350 -2154
rect 1344 -2166 1350 -2160
rect 1344 -2172 1350 -2166
rect 1344 -2178 1350 -2172
rect 1344 -2184 1350 -2178
rect 1344 -2190 1350 -2184
rect 1344 -2196 1350 -2190
rect 1344 -2202 1350 -2196
rect 1344 -2208 1350 -2202
rect 1344 -2214 1350 -2208
rect 1344 -2220 1350 -2214
rect 1344 -2226 1350 -2220
rect 1344 -2232 1350 -2226
rect 1344 -2238 1350 -2232
rect 1344 -2244 1350 -2238
rect 1344 -2250 1350 -2244
rect 1344 -2256 1350 -2250
rect 1344 -2262 1350 -2256
rect 1344 -2268 1350 -2262
rect 1344 -2274 1350 -2268
rect 1344 -2280 1350 -2274
rect 1344 -2286 1350 -2280
rect 1344 -2292 1350 -2286
rect 1344 -2298 1350 -2292
rect 1344 -2304 1350 -2298
rect 1344 -2310 1350 -2304
rect 1344 -2316 1350 -2310
rect 1344 -2322 1350 -2316
rect 1344 -2328 1350 -2322
rect 1344 -2334 1350 -2328
rect 1344 -2340 1350 -2334
rect 1344 -2346 1350 -2340
rect 1344 -2352 1350 -2346
rect 1344 -2358 1350 -2352
rect 1344 -2364 1350 -2358
rect 1344 -2370 1350 -2364
rect 1344 -2376 1350 -2370
rect 1344 -2382 1350 -2376
rect 1344 -2388 1350 -2382
rect 1344 -2394 1350 -2388
rect 1344 -2400 1350 -2394
rect 1344 -2478 1350 -2472
rect 1344 -2484 1350 -2478
rect 1344 -2490 1350 -2484
rect 1344 -2496 1350 -2490
rect 1344 -2502 1350 -2496
rect 1344 -2508 1350 -2502
rect 1344 -2514 1350 -2508
rect 1344 -2520 1350 -2514
rect 1344 -2526 1350 -2520
rect 1344 -2532 1350 -2526
rect 1344 -2538 1350 -2532
rect 1344 -2544 1350 -2538
rect 1344 -2550 1350 -2544
rect 1344 -2556 1350 -2550
rect 1344 -2562 1350 -2556
rect 1344 -2568 1350 -2562
rect 1344 -2574 1350 -2568
rect 1344 -2580 1350 -2574
rect 1344 -2586 1350 -2580
rect 1344 -2592 1350 -2586
rect 1344 -2598 1350 -2592
rect 1344 -2604 1350 -2598
rect 1344 -2610 1350 -2604
rect 1344 -2616 1350 -2610
rect 1344 -2622 1350 -2616
rect 1344 -2628 1350 -2622
rect 1344 -2634 1350 -2628
rect 1344 -2640 1350 -2634
rect 1344 -2646 1350 -2640
rect 1344 -2652 1350 -2646
rect 1344 -2658 1350 -2652
rect 1344 -2664 1350 -2658
rect 1344 -2670 1350 -2664
rect 1344 -2676 1350 -2670
rect 1344 -2682 1350 -2676
rect 1344 -2688 1350 -2682
rect 1344 -2694 1350 -2688
rect 1344 -2700 1350 -2694
rect 1344 -2706 1350 -2700
rect 1344 -2712 1350 -2706
rect 1344 -2718 1350 -2712
rect 1344 -2724 1350 -2718
rect 1344 -2730 1350 -2724
rect 1344 -2736 1350 -2730
rect 1344 -2742 1350 -2736
rect 1344 -2748 1350 -2742
rect 1344 -2754 1350 -2748
rect 1344 -2760 1350 -2754
rect 1344 -2766 1350 -2760
rect 1344 -2772 1350 -2766
rect 1344 -2778 1350 -2772
rect 1344 -2784 1350 -2778
rect 1344 -2790 1350 -2784
rect 1344 -2796 1350 -2790
rect 1344 -2802 1350 -2796
rect 1344 -2808 1350 -2802
rect 1344 -2814 1350 -2808
rect 1344 -2820 1350 -2814
rect 1344 -2826 1350 -2820
rect 1344 -2832 1350 -2826
rect 1344 -2838 1350 -2832
rect 1344 -2844 1350 -2838
rect 1344 -2850 1350 -2844
rect 1344 -2856 1350 -2850
rect 1344 -2862 1350 -2856
rect 1344 -2868 1350 -2862
rect 1344 -2874 1350 -2868
rect 1344 -2880 1350 -2874
rect 1344 -2886 1350 -2880
rect 1344 -2892 1350 -2886
rect 1344 -2898 1350 -2892
rect 1344 -2904 1350 -2898
rect 1344 -2910 1350 -2904
rect 1344 -2916 1350 -2910
rect 1344 -3000 1350 -2994
rect 1344 -3006 1350 -3000
rect 1344 -3012 1350 -3006
rect 1344 -3018 1350 -3012
rect 1344 -3024 1350 -3018
rect 1344 -3030 1350 -3024
rect 1344 -3036 1350 -3030
rect 1344 -3042 1350 -3036
rect 1344 -3048 1350 -3042
rect 1344 -3054 1350 -3048
rect 1344 -3060 1350 -3054
rect 1344 -3066 1350 -3060
rect 1344 -3072 1350 -3066
rect 1344 -3078 1350 -3072
rect 1344 -3084 1350 -3078
rect 1344 -3090 1350 -3084
rect 1344 -3096 1350 -3090
rect 1344 -3102 1350 -3096
rect 1344 -3108 1350 -3102
rect 1344 -3114 1350 -3108
rect 1344 -3120 1350 -3114
rect 1344 -3126 1350 -3120
rect 1344 -3132 1350 -3126
rect 1344 -3138 1350 -3132
rect 1344 -3144 1350 -3138
rect 1344 -3150 1350 -3144
rect 1344 -3156 1350 -3150
rect 1344 -3162 1350 -3156
rect 1344 -3168 1350 -3162
rect 1344 -3174 1350 -3168
rect 1344 -3180 1350 -3174
rect 1344 -3186 1350 -3180
rect 1344 -3192 1350 -3186
rect 1344 -3198 1350 -3192
rect 1344 -3204 1350 -3198
rect 1344 -3210 1350 -3204
rect 1344 -3216 1350 -3210
rect 1344 -3222 1350 -3216
rect 1344 -3228 1350 -3222
rect 1344 -3234 1350 -3228
rect 1344 -3312 1350 -3306
rect 1344 -3318 1350 -3312
rect 1344 -3324 1350 -3318
rect 1344 -3330 1350 -3324
rect 1344 -3336 1350 -3330
rect 1344 -3342 1350 -3336
rect 1344 -3348 1350 -3342
rect 1344 -3354 1350 -3348
rect 1344 -3360 1350 -3354
rect 1344 -3366 1350 -3360
rect 1344 -3372 1350 -3366
rect 1344 -3378 1350 -3372
rect 1344 -3384 1350 -3378
rect 1344 -3390 1350 -3384
rect 1344 -3396 1350 -3390
rect 1344 -3402 1350 -3396
rect 1344 -3408 1350 -3402
rect 1344 -3414 1350 -3408
rect 1344 -3420 1350 -3414
rect 1344 -3426 1350 -3420
rect 1344 -3432 1350 -3426
rect 1344 -3438 1350 -3432
rect 1344 -3444 1350 -3438
rect 1344 -3450 1350 -3444
rect 1344 -3456 1350 -3450
rect 1344 -3462 1350 -3456
rect 1344 -3468 1350 -3462
rect 1344 -3474 1350 -3468
rect 1344 -3480 1350 -3474
rect 1344 -3486 1350 -3480
rect 1344 -3492 1350 -3486
rect 1344 -3498 1350 -3492
rect 1344 -3504 1350 -3498
rect 1344 -3510 1350 -3504
rect 1344 -3516 1350 -3510
rect 1350 -1110 1356 -1104
rect 1350 -1116 1356 -1110
rect 1350 -1122 1356 -1116
rect 1350 -1128 1356 -1122
rect 1350 -1134 1356 -1128
rect 1350 -1140 1356 -1134
rect 1350 -1146 1356 -1140
rect 1350 -1152 1356 -1146
rect 1350 -1158 1356 -1152
rect 1350 -1164 1356 -1158
rect 1350 -1170 1356 -1164
rect 1350 -1176 1356 -1170
rect 1350 -1182 1356 -1176
rect 1350 -1188 1356 -1182
rect 1350 -1194 1356 -1188
rect 1350 -1200 1356 -1194
rect 1350 -1206 1356 -1200
rect 1350 -1212 1356 -1206
rect 1350 -1218 1356 -1212
rect 1350 -1224 1356 -1218
rect 1350 -1230 1356 -1224
rect 1350 -1236 1356 -1230
rect 1350 -1242 1356 -1236
rect 1350 -1248 1356 -1242
rect 1350 -1254 1356 -1248
rect 1350 -1260 1356 -1254
rect 1350 -1266 1356 -1260
rect 1350 -1272 1356 -1266
rect 1350 -1278 1356 -1272
rect 1350 -1284 1356 -1278
rect 1350 -1290 1356 -1284
rect 1350 -1296 1356 -1290
rect 1350 -1302 1356 -1296
rect 1350 -1308 1356 -1302
rect 1350 -1314 1356 -1308
rect 1350 -1464 1356 -1458
rect 1350 -1470 1356 -1464
rect 1350 -1476 1356 -1470
rect 1350 -1482 1356 -1476
rect 1350 -1488 1356 -1482
rect 1350 -1494 1356 -1488
rect 1350 -1500 1356 -1494
rect 1350 -1506 1356 -1500
rect 1350 -1512 1356 -1506
rect 1350 -1518 1356 -1512
rect 1350 -1524 1356 -1518
rect 1350 -1530 1356 -1524
rect 1350 -1536 1356 -1530
rect 1350 -1542 1356 -1536
rect 1350 -1548 1356 -1542
rect 1350 -1554 1356 -1548
rect 1350 -1560 1356 -1554
rect 1350 -1566 1356 -1560
rect 1350 -1572 1356 -1566
rect 1350 -1578 1356 -1572
rect 1350 -1584 1356 -1578
rect 1350 -1590 1356 -1584
rect 1350 -1596 1356 -1590
rect 1350 -1602 1356 -1596
rect 1350 -1608 1356 -1602
rect 1350 -1614 1356 -1608
rect 1350 -1620 1356 -1614
rect 1350 -1626 1356 -1620
rect 1350 -1632 1356 -1626
rect 1350 -1638 1356 -1632
rect 1350 -1644 1356 -1638
rect 1350 -1650 1356 -1644
rect 1350 -1656 1356 -1650
rect 1350 -1662 1356 -1656
rect 1350 -1668 1356 -1662
rect 1350 -1674 1356 -1668
rect 1350 -1680 1356 -1674
rect 1350 -1686 1356 -1680
rect 1350 -1692 1356 -1686
rect 1350 -1698 1356 -1692
rect 1350 -1704 1356 -1698
rect 1350 -1710 1356 -1704
rect 1350 -1716 1356 -1710
rect 1350 -1722 1356 -1716
rect 1350 -1728 1356 -1722
rect 1350 -1734 1356 -1728
rect 1350 -1740 1356 -1734
rect 1350 -1746 1356 -1740
rect 1350 -1752 1356 -1746
rect 1350 -1758 1356 -1752
rect 1350 -1764 1356 -1758
rect 1350 -1770 1356 -1764
rect 1350 -1776 1356 -1770
rect 1350 -1782 1356 -1776
rect 1350 -1788 1356 -1782
rect 1350 -1794 1356 -1788
rect 1350 -1800 1356 -1794
rect 1350 -1806 1356 -1800
rect 1350 -1812 1356 -1806
rect 1350 -1818 1356 -1812
rect 1350 -1824 1356 -1818
rect 1350 -1830 1356 -1824
rect 1350 -1836 1356 -1830
rect 1350 -1842 1356 -1836
rect 1350 -1848 1356 -1842
rect 1350 -1854 1356 -1848
rect 1350 -1860 1356 -1854
rect 1350 -1866 1356 -1860
rect 1350 -1872 1356 -1866
rect 1350 -1878 1356 -1872
rect 1350 -1884 1356 -1878
rect 1350 -1890 1356 -1884
rect 1350 -1896 1356 -1890
rect 1350 -1902 1356 -1896
rect 1350 -1908 1356 -1902
rect 1350 -1914 1356 -1908
rect 1350 -1920 1356 -1914
rect 1350 -1926 1356 -1920
rect 1350 -1932 1356 -1926
rect 1350 -1938 1356 -1932
rect 1350 -1944 1356 -1938
rect 1350 -1950 1356 -1944
rect 1350 -1956 1356 -1950
rect 1350 -1962 1356 -1956
rect 1350 -1968 1356 -1962
rect 1350 -1974 1356 -1968
rect 1350 -1980 1356 -1974
rect 1350 -1986 1356 -1980
rect 1350 -1992 1356 -1986
rect 1350 -1998 1356 -1992
rect 1350 -2004 1356 -1998
rect 1350 -2010 1356 -2004
rect 1350 -2016 1356 -2010
rect 1350 -2022 1356 -2016
rect 1350 -2028 1356 -2022
rect 1350 -2034 1356 -2028
rect 1350 -2040 1356 -2034
rect 1350 -2046 1356 -2040
rect 1350 -2052 1356 -2046
rect 1350 -2058 1356 -2052
rect 1350 -2064 1356 -2058
rect 1350 -2070 1356 -2064
rect 1350 -2076 1356 -2070
rect 1350 -2082 1356 -2076
rect 1350 -2088 1356 -2082
rect 1350 -2094 1356 -2088
rect 1350 -2100 1356 -2094
rect 1350 -2106 1356 -2100
rect 1350 -2112 1356 -2106
rect 1350 -2118 1356 -2112
rect 1350 -2124 1356 -2118
rect 1350 -2130 1356 -2124
rect 1350 -2136 1356 -2130
rect 1350 -2142 1356 -2136
rect 1350 -2148 1356 -2142
rect 1350 -2154 1356 -2148
rect 1350 -2160 1356 -2154
rect 1350 -2166 1356 -2160
rect 1350 -2172 1356 -2166
rect 1350 -2178 1356 -2172
rect 1350 -2184 1356 -2178
rect 1350 -2190 1356 -2184
rect 1350 -2196 1356 -2190
rect 1350 -2202 1356 -2196
rect 1350 -2208 1356 -2202
rect 1350 -2214 1356 -2208
rect 1350 -2220 1356 -2214
rect 1350 -2226 1356 -2220
rect 1350 -2232 1356 -2226
rect 1350 -2238 1356 -2232
rect 1350 -2244 1356 -2238
rect 1350 -2250 1356 -2244
rect 1350 -2256 1356 -2250
rect 1350 -2262 1356 -2256
rect 1350 -2268 1356 -2262
rect 1350 -2274 1356 -2268
rect 1350 -2280 1356 -2274
rect 1350 -2286 1356 -2280
rect 1350 -2292 1356 -2286
rect 1350 -2298 1356 -2292
rect 1350 -2304 1356 -2298
rect 1350 -2310 1356 -2304
rect 1350 -2316 1356 -2310
rect 1350 -2322 1356 -2316
rect 1350 -2328 1356 -2322
rect 1350 -2334 1356 -2328
rect 1350 -2340 1356 -2334
rect 1350 -2346 1356 -2340
rect 1350 -2352 1356 -2346
rect 1350 -2358 1356 -2352
rect 1350 -2364 1356 -2358
rect 1350 -2370 1356 -2364
rect 1350 -2376 1356 -2370
rect 1350 -2382 1356 -2376
rect 1350 -2388 1356 -2382
rect 1350 -2472 1356 -2466
rect 1350 -2478 1356 -2472
rect 1350 -2484 1356 -2478
rect 1350 -2490 1356 -2484
rect 1350 -2496 1356 -2490
rect 1350 -2502 1356 -2496
rect 1350 -2508 1356 -2502
rect 1350 -2514 1356 -2508
rect 1350 -2520 1356 -2514
rect 1350 -2526 1356 -2520
rect 1350 -2532 1356 -2526
rect 1350 -2538 1356 -2532
rect 1350 -2544 1356 -2538
rect 1350 -2550 1356 -2544
rect 1350 -2556 1356 -2550
rect 1350 -2562 1356 -2556
rect 1350 -2568 1356 -2562
rect 1350 -2574 1356 -2568
rect 1350 -2580 1356 -2574
rect 1350 -2586 1356 -2580
rect 1350 -2592 1356 -2586
rect 1350 -2598 1356 -2592
rect 1350 -2604 1356 -2598
rect 1350 -2610 1356 -2604
rect 1350 -2616 1356 -2610
rect 1350 -2622 1356 -2616
rect 1350 -2628 1356 -2622
rect 1350 -2634 1356 -2628
rect 1350 -2640 1356 -2634
rect 1350 -2646 1356 -2640
rect 1350 -2652 1356 -2646
rect 1350 -2658 1356 -2652
rect 1350 -2664 1356 -2658
rect 1350 -2670 1356 -2664
rect 1350 -2676 1356 -2670
rect 1350 -2682 1356 -2676
rect 1350 -2688 1356 -2682
rect 1350 -2694 1356 -2688
rect 1350 -2700 1356 -2694
rect 1350 -2706 1356 -2700
rect 1350 -2712 1356 -2706
rect 1350 -2718 1356 -2712
rect 1350 -2724 1356 -2718
rect 1350 -2730 1356 -2724
rect 1350 -2736 1356 -2730
rect 1350 -2742 1356 -2736
rect 1350 -2748 1356 -2742
rect 1350 -2754 1356 -2748
rect 1350 -2760 1356 -2754
rect 1350 -2766 1356 -2760
rect 1350 -2772 1356 -2766
rect 1350 -2778 1356 -2772
rect 1350 -2784 1356 -2778
rect 1350 -2790 1356 -2784
rect 1350 -2796 1356 -2790
rect 1350 -2802 1356 -2796
rect 1350 -2808 1356 -2802
rect 1350 -2814 1356 -2808
rect 1350 -2820 1356 -2814
rect 1350 -2826 1356 -2820
rect 1350 -2832 1356 -2826
rect 1350 -2838 1356 -2832
rect 1350 -2844 1356 -2838
rect 1350 -2850 1356 -2844
rect 1350 -2856 1356 -2850
rect 1350 -2862 1356 -2856
rect 1350 -2868 1356 -2862
rect 1350 -2874 1356 -2868
rect 1350 -2880 1356 -2874
rect 1350 -2886 1356 -2880
rect 1350 -2892 1356 -2886
rect 1350 -2898 1356 -2892
rect 1350 -2904 1356 -2898
rect 1350 -2910 1356 -2904
rect 1350 -2994 1356 -2988
rect 1350 -3000 1356 -2994
rect 1350 -3006 1356 -3000
rect 1350 -3012 1356 -3006
rect 1350 -3018 1356 -3012
rect 1350 -3024 1356 -3018
rect 1350 -3030 1356 -3024
rect 1350 -3036 1356 -3030
rect 1350 -3042 1356 -3036
rect 1350 -3048 1356 -3042
rect 1350 -3054 1356 -3048
rect 1350 -3060 1356 -3054
rect 1350 -3066 1356 -3060
rect 1350 -3072 1356 -3066
rect 1350 -3078 1356 -3072
rect 1350 -3084 1356 -3078
rect 1350 -3090 1356 -3084
rect 1350 -3096 1356 -3090
rect 1350 -3102 1356 -3096
rect 1350 -3108 1356 -3102
rect 1350 -3114 1356 -3108
rect 1350 -3120 1356 -3114
rect 1350 -3126 1356 -3120
rect 1350 -3132 1356 -3126
rect 1350 -3138 1356 -3132
rect 1350 -3144 1356 -3138
rect 1350 -3150 1356 -3144
rect 1350 -3156 1356 -3150
rect 1350 -3162 1356 -3156
rect 1350 -3168 1356 -3162
rect 1350 -3174 1356 -3168
rect 1350 -3180 1356 -3174
rect 1350 -3186 1356 -3180
rect 1350 -3192 1356 -3186
rect 1350 -3198 1356 -3192
rect 1350 -3204 1356 -3198
rect 1350 -3210 1356 -3204
rect 1350 -3216 1356 -3210
rect 1350 -3222 1356 -3216
rect 1350 -3228 1356 -3222
rect 1350 -3234 1356 -3228
rect 1350 -3312 1356 -3306
rect 1350 -3318 1356 -3312
rect 1350 -3324 1356 -3318
rect 1350 -3330 1356 -3324
rect 1350 -3336 1356 -3330
rect 1350 -3342 1356 -3336
rect 1350 -3348 1356 -3342
rect 1350 -3354 1356 -3348
rect 1350 -3360 1356 -3354
rect 1350 -3366 1356 -3360
rect 1350 -3372 1356 -3366
rect 1350 -3378 1356 -3372
rect 1350 -3384 1356 -3378
rect 1350 -3390 1356 -3384
rect 1350 -3396 1356 -3390
rect 1350 -3402 1356 -3396
rect 1350 -3408 1356 -3402
rect 1350 -3414 1356 -3408
rect 1350 -3420 1356 -3414
rect 1350 -3426 1356 -3420
rect 1350 -3432 1356 -3426
rect 1350 -3438 1356 -3432
rect 1350 -3444 1356 -3438
rect 1350 -3450 1356 -3444
rect 1350 -3456 1356 -3450
rect 1350 -3462 1356 -3456
rect 1350 -3468 1356 -3462
rect 1350 -3474 1356 -3468
rect 1350 -3480 1356 -3474
rect 1350 -3486 1356 -3480
rect 1350 -3492 1356 -3486
rect 1350 -3498 1356 -3492
rect 1350 -3504 1356 -3498
rect 1350 -3510 1356 -3504
rect 1350 -3516 1356 -3510
rect 1356 -1110 1362 -1104
rect 1356 -1116 1362 -1110
rect 1356 -1122 1362 -1116
rect 1356 -1128 1362 -1122
rect 1356 -1134 1362 -1128
rect 1356 -1140 1362 -1134
rect 1356 -1146 1362 -1140
rect 1356 -1152 1362 -1146
rect 1356 -1158 1362 -1152
rect 1356 -1164 1362 -1158
rect 1356 -1170 1362 -1164
rect 1356 -1176 1362 -1170
rect 1356 -1182 1362 -1176
rect 1356 -1188 1362 -1182
rect 1356 -1194 1362 -1188
rect 1356 -1200 1362 -1194
rect 1356 -1206 1362 -1200
rect 1356 -1212 1362 -1206
rect 1356 -1218 1362 -1212
rect 1356 -1224 1362 -1218
rect 1356 -1230 1362 -1224
rect 1356 -1236 1362 -1230
rect 1356 -1242 1362 -1236
rect 1356 -1248 1362 -1242
rect 1356 -1254 1362 -1248
rect 1356 -1260 1362 -1254
rect 1356 -1266 1362 -1260
rect 1356 -1272 1362 -1266
rect 1356 -1278 1362 -1272
rect 1356 -1284 1362 -1278
rect 1356 -1290 1362 -1284
rect 1356 -1296 1362 -1290
rect 1356 -1302 1362 -1296
rect 1356 -1308 1362 -1302
rect 1356 -1314 1362 -1308
rect 1356 -1452 1362 -1446
rect 1356 -1458 1362 -1452
rect 1356 -1464 1362 -1458
rect 1356 -1470 1362 -1464
rect 1356 -1476 1362 -1470
rect 1356 -1482 1362 -1476
rect 1356 -1488 1362 -1482
rect 1356 -1494 1362 -1488
rect 1356 -1500 1362 -1494
rect 1356 -1506 1362 -1500
rect 1356 -1512 1362 -1506
rect 1356 -1518 1362 -1512
rect 1356 -1524 1362 -1518
rect 1356 -1530 1362 -1524
rect 1356 -1536 1362 -1530
rect 1356 -1542 1362 -1536
rect 1356 -1548 1362 -1542
rect 1356 -1554 1362 -1548
rect 1356 -1560 1362 -1554
rect 1356 -1566 1362 -1560
rect 1356 -1572 1362 -1566
rect 1356 -1578 1362 -1572
rect 1356 -1584 1362 -1578
rect 1356 -1590 1362 -1584
rect 1356 -1596 1362 -1590
rect 1356 -1602 1362 -1596
rect 1356 -1608 1362 -1602
rect 1356 -1614 1362 -1608
rect 1356 -1620 1362 -1614
rect 1356 -1626 1362 -1620
rect 1356 -1632 1362 -1626
rect 1356 -1638 1362 -1632
rect 1356 -1644 1362 -1638
rect 1356 -1650 1362 -1644
rect 1356 -1656 1362 -1650
rect 1356 -1662 1362 -1656
rect 1356 -1668 1362 -1662
rect 1356 -1674 1362 -1668
rect 1356 -1680 1362 -1674
rect 1356 -1686 1362 -1680
rect 1356 -1692 1362 -1686
rect 1356 -1698 1362 -1692
rect 1356 -1704 1362 -1698
rect 1356 -1710 1362 -1704
rect 1356 -1716 1362 -1710
rect 1356 -1722 1362 -1716
rect 1356 -1728 1362 -1722
rect 1356 -1734 1362 -1728
rect 1356 -1740 1362 -1734
rect 1356 -1746 1362 -1740
rect 1356 -1752 1362 -1746
rect 1356 -1758 1362 -1752
rect 1356 -1764 1362 -1758
rect 1356 -1770 1362 -1764
rect 1356 -1776 1362 -1770
rect 1356 -1782 1362 -1776
rect 1356 -1788 1362 -1782
rect 1356 -1794 1362 -1788
rect 1356 -1800 1362 -1794
rect 1356 -1806 1362 -1800
rect 1356 -1812 1362 -1806
rect 1356 -1818 1362 -1812
rect 1356 -1824 1362 -1818
rect 1356 -1830 1362 -1824
rect 1356 -1836 1362 -1830
rect 1356 -1842 1362 -1836
rect 1356 -1848 1362 -1842
rect 1356 -1854 1362 -1848
rect 1356 -1860 1362 -1854
rect 1356 -1866 1362 -1860
rect 1356 -1872 1362 -1866
rect 1356 -1878 1362 -1872
rect 1356 -1884 1362 -1878
rect 1356 -1890 1362 -1884
rect 1356 -1896 1362 -1890
rect 1356 -1902 1362 -1896
rect 1356 -1908 1362 -1902
rect 1356 -1914 1362 -1908
rect 1356 -1920 1362 -1914
rect 1356 -1926 1362 -1920
rect 1356 -1932 1362 -1926
rect 1356 -1938 1362 -1932
rect 1356 -1944 1362 -1938
rect 1356 -1950 1362 -1944
rect 1356 -1956 1362 -1950
rect 1356 -1962 1362 -1956
rect 1356 -1968 1362 -1962
rect 1356 -1974 1362 -1968
rect 1356 -1980 1362 -1974
rect 1356 -1986 1362 -1980
rect 1356 -1992 1362 -1986
rect 1356 -1998 1362 -1992
rect 1356 -2004 1362 -1998
rect 1356 -2010 1362 -2004
rect 1356 -2016 1362 -2010
rect 1356 -2022 1362 -2016
rect 1356 -2028 1362 -2022
rect 1356 -2034 1362 -2028
rect 1356 -2040 1362 -2034
rect 1356 -2046 1362 -2040
rect 1356 -2052 1362 -2046
rect 1356 -2058 1362 -2052
rect 1356 -2064 1362 -2058
rect 1356 -2070 1362 -2064
rect 1356 -2076 1362 -2070
rect 1356 -2082 1362 -2076
rect 1356 -2088 1362 -2082
rect 1356 -2094 1362 -2088
rect 1356 -2100 1362 -2094
rect 1356 -2106 1362 -2100
rect 1356 -2112 1362 -2106
rect 1356 -2118 1362 -2112
rect 1356 -2124 1362 -2118
rect 1356 -2130 1362 -2124
rect 1356 -2136 1362 -2130
rect 1356 -2142 1362 -2136
rect 1356 -2148 1362 -2142
rect 1356 -2154 1362 -2148
rect 1356 -2160 1362 -2154
rect 1356 -2166 1362 -2160
rect 1356 -2172 1362 -2166
rect 1356 -2178 1362 -2172
rect 1356 -2184 1362 -2178
rect 1356 -2190 1362 -2184
rect 1356 -2196 1362 -2190
rect 1356 -2202 1362 -2196
rect 1356 -2208 1362 -2202
rect 1356 -2214 1362 -2208
rect 1356 -2220 1362 -2214
rect 1356 -2226 1362 -2220
rect 1356 -2232 1362 -2226
rect 1356 -2238 1362 -2232
rect 1356 -2244 1362 -2238
rect 1356 -2250 1362 -2244
rect 1356 -2256 1362 -2250
rect 1356 -2262 1362 -2256
rect 1356 -2268 1362 -2262
rect 1356 -2274 1362 -2268
rect 1356 -2280 1362 -2274
rect 1356 -2286 1362 -2280
rect 1356 -2292 1362 -2286
rect 1356 -2298 1362 -2292
rect 1356 -2304 1362 -2298
rect 1356 -2310 1362 -2304
rect 1356 -2316 1362 -2310
rect 1356 -2322 1362 -2316
rect 1356 -2328 1362 -2322
rect 1356 -2334 1362 -2328
rect 1356 -2340 1362 -2334
rect 1356 -2346 1362 -2340
rect 1356 -2352 1362 -2346
rect 1356 -2358 1362 -2352
rect 1356 -2364 1362 -2358
rect 1356 -2370 1362 -2364
rect 1356 -2376 1362 -2370
rect 1356 -2382 1362 -2376
rect 1356 -2460 1362 -2454
rect 1356 -2466 1362 -2460
rect 1356 -2472 1362 -2466
rect 1356 -2478 1362 -2472
rect 1356 -2484 1362 -2478
rect 1356 -2490 1362 -2484
rect 1356 -2496 1362 -2490
rect 1356 -2502 1362 -2496
rect 1356 -2508 1362 -2502
rect 1356 -2514 1362 -2508
rect 1356 -2520 1362 -2514
rect 1356 -2526 1362 -2520
rect 1356 -2532 1362 -2526
rect 1356 -2538 1362 -2532
rect 1356 -2544 1362 -2538
rect 1356 -2550 1362 -2544
rect 1356 -2556 1362 -2550
rect 1356 -2562 1362 -2556
rect 1356 -2568 1362 -2562
rect 1356 -2574 1362 -2568
rect 1356 -2580 1362 -2574
rect 1356 -2586 1362 -2580
rect 1356 -2592 1362 -2586
rect 1356 -2598 1362 -2592
rect 1356 -2604 1362 -2598
rect 1356 -2610 1362 -2604
rect 1356 -2616 1362 -2610
rect 1356 -2622 1362 -2616
rect 1356 -2628 1362 -2622
rect 1356 -2634 1362 -2628
rect 1356 -2640 1362 -2634
rect 1356 -2646 1362 -2640
rect 1356 -2652 1362 -2646
rect 1356 -2658 1362 -2652
rect 1356 -2664 1362 -2658
rect 1356 -2670 1362 -2664
rect 1356 -2676 1362 -2670
rect 1356 -2682 1362 -2676
rect 1356 -2688 1362 -2682
rect 1356 -2694 1362 -2688
rect 1356 -2700 1362 -2694
rect 1356 -2706 1362 -2700
rect 1356 -2712 1362 -2706
rect 1356 -2718 1362 -2712
rect 1356 -2724 1362 -2718
rect 1356 -2730 1362 -2724
rect 1356 -2736 1362 -2730
rect 1356 -2742 1362 -2736
rect 1356 -2748 1362 -2742
rect 1356 -2754 1362 -2748
rect 1356 -2760 1362 -2754
rect 1356 -2766 1362 -2760
rect 1356 -2772 1362 -2766
rect 1356 -2778 1362 -2772
rect 1356 -2784 1362 -2778
rect 1356 -2790 1362 -2784
rect 1356 -2796 1362 -2790
rect 1356 -2802 1362 -2796
rect 1356 -2808 1362 -2802
rect 1356 -2814 1362 -2808
rect 1356 -2820 1362 -2814
rect 1356 -2826 1362 -2820
rect 1356 -2832 1362 -2826
rect 1356 -2838 1362 -2832
rect 1356 -2844 1362 -2838
rect 1356 -2850 1362 -2844
rect 1356 -2856 1362 -2850
rect 1356 -2862 1362 -2856
rect 1356 -2868 1362 -2862
rect 1356 -2874 1362 -2868
rect 1356 -2880 1362 -2874
rect 1356 -2886 1362 -2880
rect 1356 -2892 1362 -2886
rect 1356 -2898 1362 -2892
rect 1356 -2904 1362 -2898
rect 1356 -2988 1362 -2982
rect 1356 -2994 1362 -2988
rect 1356 -3000 1362 -2994
rect 1356 -3006 1362 -3000
rect 1356 -3012 1362 -3006
rect 1356 -3018 1362 -3012
rect 1356 -3024 1362 -3018
rect 1356 -3030 1362 -3024
rect 1356 -3036 1362 -3030
rect 1356 -3042 1362 -3036
rect 1356 -3048 1362 -3042
rect 1356 -3054 1362 -3048
rect 1356 -3060 1362 -3054
rect 1356 -3066 1362 -3060
rect 1356 -3072 1362 -3066
rect 1356 -3078 1362 -3072
rect 1356 -3084 1362 -3078
rect 1356 -3090 1362 -3084
rect 1356 -3096 1362 -3090
rect 1356 -3102 1362 -3096
rect 1356 -3108 1362 -3102
rect 1356 -3114 1362 -3108
rect 1356 -3120 1362 -3114
rect 1356 -3126 1362 -3120
rect 1356 -3132 1362 -3126
rect 1356 -3138 1362 -3132
rect 1356 -3144 1362 -3138
rect 1356 -3150 1362 -3144
rect 1356 -3156 1362 -3150
rect 1356 -3162 1362 -3156
rect 1356 -3168 1362 -3162
rect 1356 -3174 1362 -3168
rect 1356 -3180 1362 -3174
rect 1356 -3186 1362 -3180
rect 1356 -3192 1362 -3186
rect 1356 -3198 1362 -3192
rect 1356 -3204 1362 -3198
rect 1356 -3210 1362 -3204
rect 1356 -3216 1362 -3210
rect 1356 -3222 1362 -3216
rect 1356 -3228 1362 -3222
rect 1356 -3234 1362 -3228
rect 1356 -3312 1362 -3306
rect 1356 -3318 1362 -3312
rect 1356 -3324 1362 -3318
rect 1356 -3330 1362 -3324
rect 1356 -3336 1362 -3330
rect 1356 -3342 1362 -3336
rect 1356 -3348 1362 -3342
rect 1356 -3354 1362 -3348
rect 1356 -3360 1362 -3354
rect 1356 -3366 1362 -3360
rect 1356 -3372 1362 -3366
rect 1356 -3378 1362 -3372
rect 1356 -3384 1362 -3378
rect 1356 -3390 1362 -3384
rect 1356 -3396 1362 -3390
rect 1356 -3402 1362 -3396
rect 1356 -3408 1362 -3402
rect 1356 -3414 1362 -3408
rect 1356 -3420 1362 -3414
rect 1356 -3426 1362 -3420
rect 1356 -3432 1362 -3426
rect 1356 -3438 1362 -3432
rect 1356 -3444 1362 -3438
rect 1356 -3450 1362 -3444
rect 1356 -3456 1362 -3450
rect 1356 -3462 1362 -3456
rect 1356 -3468 1362 -3462
rect 1356 -3474 1362 -3468
rect 1356 -3480 1362 -3474
rect 1356 -3486 1362 -3480
rect 1356 -3492 1362 -3486
rect 1356 -3498 1362 -3492
rect 1356 -3504 1362 -3498
rect 1356 -3510 1362 -3504
rect 1356 -3516 1362 -3510
rect 1362 -1110 1368 -1104
rect 1362 -1116 1368 -1110
rect 1362 -1122 1368 -1116
rect 1362 -1128 1368 -1122
rect 1362 -1134 1368 -1128
rect 1362 -1140 1368 -1134
rect 1362 -1146 1368 -1140
rect 1362 -1152 1368 -1146
rect 1362 -1158 1368 -1152
rect 1362 -1164 1368 -1158
rect 1362 -1170 1368 -1164
rect 1362 -1176 1368 -1170
rect 1362 -1182 1368 -1176
rect 1362 -1188 1368 -1182
rect 1362 -1194 1368 -1188
rect 1362 -1200 1368 -1194
rect 1362 -1206 1368 -1200
rect 1362 -1212 1368 -1206
rect 1362 -1218 1368 -1212
rect 1362 -1224 1368 -1218
rect 1362 -1230 1368 -1224
rect 1362 -1236 1368 -1230
rect 1362 -1242 1368 -1236
rect 1362 -1248 1368 -1242
rect 1362 -1254 1368 -1248
rect 1362 -1260 1368 -1254
rect 1362 -1266 1368 -1260
rect 1362 -1272 1368 -1266
rect 1362 -1278 1368 -1272
rect 1362 -1284 1368 -1278
rect 1362 -1290 1368 -1284
rect 1362 -1296 1368 -1290
rect 1362 -1302 1368 -1296
rect 1362 -1308 1368 -1302
rect 1362 -1314 1368 -1308
rect 1362 -1440 1368 -1434
rect 1362 -1446 1368 -1440
rect 1362 -1452 1368 -1446
rect 1362 -1458 1368 -1452
rect 1362 -1464 1368 -1458
rect 1362 -1470 1368 -1464
rect 1362 -1476 1368 -1470
rect 1362 -1482 1368 -1476
rect 1362 -1488 1368 -1482
rect 1362 -1494 1368 -1488
rect 1362 -1500 1368 -1494
rect 1362 -1506 1368 -1500
rect 1362 -1512 1368 -1506
rect 1362 -1518 1368 -1512
rect 1362 -1524 1368 -1518
rect 1362 -1530 1368 -1524
rect 1362 -1536 1368 -1530
rect 1362 -1542 1368 -1536
rect 1362 -1548 1368 -1542
rect 1362 -1554 1368 -1548
rect 1362 -1560 1368 -1554
rect 1362 -1566 1368 -1560
rect 1362 -1572 1368 -1566
rect 1362 -1578 1368 -1572
rect 1362 -1584 1368 -1578
rect 1362 -1590 1368 -1584
rect 1362 -1596 1368 -1590
rect 1362 -1602 1368 -1596
rect 1362 -1608 1368 -1602
rect 1362 -1614 1368 -1608
rect 1362 -1620 1368 -1614
rect 1362 -1626 1368 -1620
rect 1362 -1632 1368 -1626
rect 1362 -1638 1368 -1632
rect 1362 -1644 1368 -1638
rect 1362 -1650 1368 -1644
rect 1362 -1656 1368 -1650
rect 1362 -1662 1368 -1656
rect 1362 -1668 1368 -1662
rect 1362 -1674 1368 -1668
rect 1362 -1680 1368 -1674
rect 1362 -1686 1368 -1680
rect 1362 -1692 1368 -1686
rect 1362 -1698 1368 -1692
rect 1362 -1704 1368 -1698
rect 1362 -1710 1368 -1704
rect 1362 -1716 1368 -1710
rect 1362 -1722 1368 -1716
rect 1362 -1728 1368 -1722
rect 1362 -1734 1368 -1728
rect 1362 -1740 1368 -1734
rect 1362 -1746 1368 -1740
rect 1362 -1752 1368 -1746
rect 1362 -1758 1368 -1752
rect 1362 -1764 1368 -1758
rect 1362 -1770 1368 -1764
rect 1362 -1776 1368 -1770
rect 1362 -1782 1368 -1776
rect 1362 -1788 1368 -1782
rect 1362 -1794 1368 -1788
rect 1362 -1800 1368 -1794
rect 1362 -1806 1368 -1800
rect 1362 -1812 1368 -1806
rect 1362 -1818 1368 -1812
rect 1362 -1824 1368 -1818
rect 1362 -1830 1368 -1824
rect 1362 -1836 1368 -1830
rect 1362 -1842 1368 -1836
rect 1362 -1848 1368 -1842
rect 1362 -1854 1368 -1848
rect 1362 -1860 1368 -1854
rect 1362 -1866 1368 -1860
rect 1362 -1872 1368 -1866
rect 1362 -1878 1368 -1872
rect 1362 -1884 1368 -1878
rect 1362 -1890 1368 -1884
rect 1362 -1896 1368 -1890
rect 1362 -1902 1368 -1896
rect 1362 -1908 1368 -1902
rect 1362 -1914 1368 -1908
rect 1362 -1920 1368 -1914
rect 1362 -1926 1368 -1920
rect 1362 -1932 1368 -1926
rect 1362 -1938 1368 -1932
rect 1362 -1944 1368 -1938
rect 1362 -1950 1368 -1944
rect 1362 -1956 1368 -1950
rect 1362 -1962 1368 -1956
rect 1362 -1968 1368 -1962
rect 1362 -1974 1368 -1968
rect 1362 -1980 1368 -1974
rect 1362 -1986 1368 -1980
rect 1362 -1992 1368 -1986
rect 1362 -1998 1368 -1992
rect 1362 -2004 1368 -1998
rect 1362 -2010 1368 -2004
rect 1362 -2016 1368 -2010
rect 1362 -2022 1368 -2016
rect 1362 -2028 1368 -2022
rect 1362 -2034 1368 -2028
rect 1362 -2040 1368 -2034
rect 1362 -2046 1368 -2040
rect 1362 -2052 1368 -2046
rect 1362 -2058 1368 -2052
rect 1362 -2064 1368 -2058
rect 1362 -2070 1368 -2064
rect 1362 -2076 1368 -2070
rect 1362 -2082 1368 -2076
rect 1362 -2088 1368 -2082
rect 1362 -2094 1368 -2088
rect 1362 -2100 1368 -2094
rect 1362 -2106 1368 -2100
rect 1362 -2112 1368 -2106
rect 1362 -2118 1368 -2112
rect 1362 -2124 1368 -2118
rect 1362 -2130 1368 -2124
rect 1362 -2136 1368 -2130
rect 1362 -2142 1368 -2136
rect 1362 -2148 1368 -2142
rect 1362 -2154 1368 -2148
rect 1362 -2160 1368 -2154
rect 1362 -2166 1368 -2160
rect 1362 -2172 1368 -2166
rect 1362 -2178 1368 -2172
rect 1362 -2184 1368 -2178
rect 1362 -2190 1368 -2184
rect 1362 -2196 1368 -2190
rect 1362 -2202 1368 -2196
rect 1362 -2208 1368 -2202
rect 1362 -2214 1368 -2208
rect 1362 -2220 1368 -2214
rect 1362 -2226 1368 -2220
rect 1362 -2232 1368 -2226
rect 1362 -2238 1368 -2232
rect 1362 -2244 1368 -2238
rect 1362 -2250 1368 -2244
rect 1362 -2256 1368 -2250
rect 1362 -2262 1368 -2256
rect 1362 -2268 1368 -2262
rect 1362 -2274 1368 -2268
rect 1362 -2280 1368 -2274
rect 1362 -2286 1368 -2280
rect 1362 -2292 1368 -2286
rect 1362 -2298 1368 -2292
rect 1362 -2304 1368 -2298
rect 1362 -2310 1368 -2304
rect 1362 -2316 1368 -2310
rect 1362 -2322 1368 -2316
rect 1362 -2328 1368 -2322
rect 1362 -2334 1368 -2328
rect 1362 -2340 1368 -2334
rect 1362 -2346 1368 -2340
rect 1362 -2352 1368 -2346
rect 1362 -2358 1368 -2352
rect 1362 -2364 1368 -2358
rect 1362 -2370 1368 -2364
rect 1362 -2376 1368 -2370
rect 1362 -2454 1368 -2448
rect 1362 -2460 1368 -2454
rect 1362 -2466 1368 -2460
rect 1362 -2472 1368 -2466
rect 1362 -2478 1368 -2472
rect 1362 -2484 1368 -2478
rect 1362 -2490 1368 -2484
rect 1362 -2496 1368 -2490
rect 1362 -2502 1368 -2496
rect 1362 -2508 1368 -2502
rect 1362 -2514 1368 -2508
rect 1362 -2520 1368 -2514
rect 1362 -2526 1368 -2520
rect 1362 -2532 1368 -2526
rect 1362 -2538 1368 -2532
rect 1362 -2544 1368 -2538
rect 1362 -2550 1368 -2544
rect 1362 -2556 1368 -2550
rect 1362 -2562 1368 -2556
rect 1362 -2568 1368 -2562
rect 1362 -2574 1368 -2568
rect 1362 -2580 1368 -2574
rect 1362 -2586 1368 -2580
rect 1362 -2592 1368 -2586
rect 1362 -2598 1368 -2592
rect 1362 -2604 1368 -2598
rect 1362 -2610 1368 -2604
rect 1362 -2616 1368 -2610
rect 1362 -2622 1368 -2616
rect 1362 -2628 1368 -2622
rect 1362 -2634 1368 -2628
rect 1362 -2640 1368 -2634
rect 1362 -2646 1368 -2640
rect 1362 -2652 1368 -2646
rect 1362 -2658 1368 -2652
rect 1362 -2664 1368 -2658
rect 1362 -2670 1368 -2664
rect 1362 -2676 1368 -2670
rect 1362 -2682 1368 -2676
rect 1362 -2688 1368 -2682
rect 1362 -2694 1368 -2688
rect 1362 -2700 1368 -2694
rect 1362 -2706 1368 -2700
rect 1362 -2712 1368 -2706
rect 1362 -2718 1368 -2712
rect 1362 -2724 1368 -2718
rect 1362 -2730 1368 -2724
rect 1362 -2736 1368 -2730
rect 1362 -2742 1368 -2736
rect 1362 -2748 1368 -2742
rect 1362 -2754 1368 -2748
rect 1362 -2760 1368 -2754
rect 1362 -2766 1368 -2760
rect 1362 -2772 1368 -2766
rect 1362 -2778 1368 -2772
rect 1362 -2784 1368 -2778
rect 1362 -2790 1368 -2784
rect 1362 -2796 1368 -2790
rect 1362 -2802 1368 -2796
rect 1362 -2808 1368 -2802
rect 1362 -2814 1368 -2808
rect 1362 -2820 1368 -2814
rect 1362 -2826 1368 -2820
rect 1362 -2832 1368 -2826
rect 1362 -2838 1368 -2832
rect 1362 -2844 1368 -2838
rect 1362 -2850 1368 -2844
rect 1362 -2856 1368 -2850
rect 1362 -2862 1368 -2856
rect 1362 -2868 1368 -2862
rect 1362 -2874 1368 -2868
rect 1362 -2880 1368 -2874
rect 1362 -2886 1368 -2880
rect 1362 -2892 1368 -2886
rect 1362 -2898 1368 -2892
rect 1362 -2904 1368 -2898
rect 1362 -2988 1368 -2982
rect 1362 -2994 1368 -2988
rect 1362 -3000 1368 -2994
rect 1362 -3006 1368 -3000
rect 1362 -3012 1368 -3006
rect 1362 -3018 1368 -3012
rect 1362 -3024 1368 -3018
rect 1362 -3030 1368 -3024
rect 1362 -3036 1368 -3030
rect 1362 -3042 1368 -3036
rect 1362 -3048 1368 -3042
rect 1362 -3054 1368 -3048
rect 1362 -3060 1368 -3054
rect 1362 -3066 1368 -3060
rect 1362 -3072 1368 -3066
rect 1362 -3078 1368 -3072
rect 1362 -3084 1368 -3078
rect 1362 -3090 1368 -3084
rect 1362 -3096 1368 -3090
rect 1362 -3102 1368 -3096
rect 1362 -3108 1368 -3102
rect 1362 -3114 1368 -3108
rect 1362 -3120 1368 -3114
rect 1362 -3126 1368 -3120
rect 1362 -3132 1368 -3126
rect 1362 -3138 1368 -3132
rect 1362 -3144 1368 -3138
rect 1362 -3150 1368 -3144
rect 1362 -3156 1368 -3150
rect 1362 -3162 1368 -3156
rect 1362 -3168 1368 -3162
rect 1362 -3174 1368 -3168
rect 1362 -3180 1368 -3174
rect 1362 -3186 1368 -3180
rect 1362 -3192 1368 -3186
rect 1362 -3198 1368 -3192
rect 1362 -3204 1368 -3198
rect 1362 -3210 1368 -3204
rect 1362 -3216 1368 -3210
rect 1362 -3222 1368 -3216
rect 1362 -3228 1368 -3222
rect 1362 -3234 1368 -3228
rect 1362 -3312 1368 -3306
rect 1362 -3318 1368 -3312
rect 1362 -3324 1368 -3318
rect 1362 -3330 1368 -3324
rect 1362 -3336 1368 -3330
rect 1362 -3342 1368 -3336
rect 1362 -3348 1368 -3342
rect 1362 -3354 1368 -3348
rect 1362 -3360 1368 -3354
rect 1362 -3366 1368 -3360
rect 1362 -3372 1368 -3366
rect 1362 -3378 1368 -3372
rect 1362 -3384 1368 -3378
rect 1362 -3390 1368 -3384
rect 1362 -3396 1368 -3390
rect 1362 -3402 1368 -3396
rect 1362 -3408 1368 -3402
rect 1362 -3414 1368 -3408
rect 1362 -3420 1368 -3414
rect 1362 -3426 1368 -3420
rect 1362 -3432 1368 -3426
rect 1362 -3438 1368 -3432
rect 1362 -3444 1368 -3438
rect 1362 -3450 1368 -3444
rect 1362 -3456 1368 -3450
rect 1362 -3462 1368 -3456
rect 1362 -3468 1368 -3462
rect 1362 -3474 1368 -3468
rect 1362 -3480 1368 -3474
rect 1362 -3486 1368 -3480
rect 1362 -3492 1368 -3486
rect 1362 -3498 1368 -3492
rect 1362 -3504 1368 -3498
rect 1362 -3510 1368 -3504
rect 1362 -3516 1368 -3510
rect 1368 -1116 1374 -1110
rect 1368 -1122 1374 -1116
rect 1368 -1128 1374 -1122
rect 1368 -1134 1374 -1128
rect 1368 -1140 1374 -1134
rect 1368 -1146 1374 -1140
rect 1368 -1152 1374 -1146
rect 1368 -1158 1374 -1152
rect 1368 -1164 1374 -1158
rect 1368 -1170 1374 -1164
rect 1368 -1176 1374 -1170
rect 1368 -1182 1374 -1176
rect 1368 -1188 1374 -1182
rect 1368 -1194 1374 -1188
rect 1368 -1200 1374 -1194
rect 1368 -1206 1374 -1200
rect 1368 -1212 1374 -1206
rect 1368 -1218 1374 -1212
rect 1368 -1224 1374 -1218
rect 1368 -1230 1374 -1224
rect 1368 -1236 1374 -1230
rect 1368 -1242 1374 -1236
rect 1368 -1248 1374 -1242
rect 1368 -1254 1374 -1248
rect 1368 -1260 1374 -1254
rect 1368 -1266 1374 -1260
rect 1368 -1272 1374 -1266
rect 1368 -1278 1374 -1272
rect 1368 -1284 1374 -1278
rect 1368 -1290 1374 -1284
rect 1368 -1296 1374 -1290
rect 1368 -1302 1374 -1296
rect 1368 -1308 1374 -1302
rect 1368 -1428 1374 -1422
rect 1368 -1434 1374 -1428
rect 1368 -1440 1374 -1434
rect 1368 -1446 1374 -1440
rect 1368 -1452 1374 -1446
rect 1368 -1458 1374 -1452
rect 1368 -1464 1374 -1458
rect 1368 -1470 1374 -1464
rect 1368 -1476 1374 -1470
rect 1368 -1482 1374 -1476
rect 1368 -1488 1374 -1482
rect 1368 -1494 1374 -1488
rect 1368 -1500 1374 -1494
rect 1368 -1506 1374 -1500
rect 1368 -1512 1374 -1506
rect 1368 -1518 1374 -1512
rect 1368 -1524 1374 -1518
rect 1368 -1530 1374 -1524
rect 1368 -1536 1374 -1530
rect 1368 -1542 1374 -1536
rect 1368 -1548 1374 -1542
rect 1368 -1554 1374 -1548
rect 1368 -1560 1374 -1554
rect 1368 -1566 1374 -1560
rect 1368 -1572 1374 -1566
rect 1368 -1578 1374 -1572
rect 1368 -1584 1374 -1578
rect 1368 -1590 1374 -1584
rect 1368 -1596 1374 -1590
rect 1368 -1602 1374 -1596
rect 1368 -1608 1374 -1602
rect 1368 -1614 1374 -1608
rect 1368 -1620 1374 -1614
rect 1368 -1626 1374 -1620
rect 1368 -1632 1374 -1626
rect 1368 -1638 1374 -1632
rect 1368 -1644 1374 -1638
rect 1368 -1650 1374 -1644
rect 1368 -1656 1374 -1650
rect 1368 -1662 1374 -1656
rect 1368 -1668 1374 -1662
rect 1368 -1674 1374 -1668
rect 1368 -1680 1374 -1674
rect 1368 -1686 1374 -1680
rect 1368 -1692 1374 -1686
rect 1368 -1698 1374 -1692
rect 1368 -1704 1374 -1698
rect 1368 -1710 1374 -1704
rect 1368 -1716 1374 -1710
rect 1368 -1722 1374 -1716
rect 1368 -1728 1374 -1722
rect 1368 -1734 1374 -1728
rect 1368 -1740 1374 -1734
rect 1368 -1746 1374 -1740
rect 1368 -1752 1374 -1746
rect 1368 -1758 1374 -1752
rect 1368 -1764 1374 -1758
rect 1368 -1770 1374 -1764
rect 1368 -1776 1374 -1770
rect 1368 -1782 1374 -1776
rect 1368 -1788 1374 -1782
rect 1368 -1794 1374 -1788
rect 1368 -1800 1374 -1794
rect 1368 -1806 1374 -1800
rect 1368 -1812 1374 -1806
rect 1368 -1818 1374 -1812
rect 1368 -1824 1374 -1818
rect 1368 -1830 1374 -1824
rect 1368 -1836 1374 -1830
rect 1368 -1842 1374 -1836
rect 1368 -1848 1374 -1842
rect 1368 -1854 1374 -1848
rect 1368 -1860 1374 -1854
rect 1368 -1866 1374 -1860
rect 1368 -1872 1374 -1866
rect 1368 -1878 1374 -1872
rect 1368 -1884 1374 -1878
rect 1368 -1890 1374 -1884
rect 1368 -1896 1374 -1890
rect 1368 -1902 1374 -1896
rect 1368 -1908 1374 -1902
rect 1368 -1914 1374 -1908
rect 1368 -1920 1374 -1914
rect 1368 -1926 1374 -1920
rect 1368 -1932 1374 -1926
rect 1368 -1938 1374 -1932
rect 1368 -1944 1374 -1938
rect 1368 -1950 1374 -1944
rect 1368 -1956 1374 -1950
rect 1368 -1962 1374 -1956
rect 1368 -1968 1374 -1962
rect 1368 -1974 1374 -1968
rect 1368 -1980 1374 -1974
rect 1368 -1986 1374 -1980
rect 1368 -1992 1374 -1986
rect 1368 -1998 1374 -1992
rect 1368 -2004 1374 -1998
rect 1368 -2010 1374 -2004
rect 1368 -2016 1374 -2010
rect 1368 -2022 1374 -2016
rect 1368 -2028 1374 -2022
rect 1368 -2034 1374 -2028
rect 1368 -2040 1374 -2034
rect 1368 -2046 1374 -2040
rect 1368 -2052 1374 -2046
rect 1368 -2058 1374 -2052
rect 1368 -2064 1374 -2058
rect 1368 -2070 1374 -2064
rect 1368 -2076 1374 -2070
rect 1368 -2082 1374 -2076
rect 1368 -2088 1374 -2082
rect 1368 -2094 1374 -2088
rect 1368 -2100 1374 -2094
rect 1368 -2106 1374 -2100
rect 1368 -2112 1374 -2106
rect 1368 -2118 1374 -2112
rect 1368 -2124 1374 -2118
rect 1368 -2130 1374 -2124
rect 1368 -2136 1374 -2130
rect 1368 -2142 1374 -2136
rect 1368 -2148 1374 -2142
rect 1368 -2154 1374 -2148
rect 1368 -2160 1374 -2154
rect 1368 -2166 1374 -2160
rect 1368 -2172 1374 -2166
rect 1368 -2178 1374 -2172
rect 1368 -2184 1374 -2178
rect 1368 -2190 1374 -2184
rect 1368 -2196 1374 -2190
rect 1368 -2202 1374 -2196
rect 1368 -2208 1374 -2202
rect 1368 -2214 1374 -2208
rect 1368 -2220 1374 -2214
rect 1368 -2226 1374 -2220
rect 1368 -2232 1374 -2226
rect 1368 -2238 1374 -2232
rect 1368 -2244 1374 -2238
rect 1368 -2250 1374 -2244
rect 1368 -2256 1374 -2250
rect 1368 -2262 1374 -2256
rect 1368 -2268 1374 -2262
rect 1368 -2274 1374 -2268
rect 1368 -2280 1374 -2274
rect 1368 -2286 1374 -2280
rect 1368 -2292 1374 -2286
rect 1368 -2298 1374 -2292
rect 1368 -2304 1374 -2298
rect 1368 -2310 1374 -2304
rect 1368 -2316 1374 -2310
rect 1368 -2322 1374 -2316
rect 1368 -2328 1374 -2322
rect 1368 -2334 1374 -2328
rect 1368 -2340 1374 -2334
rect 1368 -2346 1374 -2340
rect 1368 -2352 1374 -2346
rect 1368 -2358 1374 -2352
rect 1368 -2364 1374 -2358
rect 1368 -2442 1374 -2436
rect 1368 -2448 1374 -2442
rect 1368 -2454 1374 -2448
rect 1368 -2460 1374 -2454
rect 1368 -2466 1374 -2460
rect 1368 -2472 1374 -2466
rect 1368 -2478 1374 -2472
rect 1368 -2484 1374 -2478
rect 1368 -2490 1374 -2484
rect 1368 -2496 1374 -2490
rect 1368 -2502 1374 -2496
rect 1368 -2508 1374 -2502
rect 1368 -2514 1374 -2508
rect 1368 -2520 1374 -2514
rect 1368 -2526 1374 -2520
rect 1368 -2532 1374 -2526
rect 1368 -2538 1374 -2532
rect 1368 -2544 1374 -2538
rect 1368 -2550 1374 -2544
rect 1368 -2556 1374 -2550
rect 1368 -2562 1374 -2556
rect 1368 -2568 1374 -2562
rect 1368 -2574 1374 -2568
rect 1368 -2580 1374 -2574
rect 1368 -2586 1374 -2580
rect 1368 -2592 1374 -2586
rect 1368 -2598 1374 -2592
rect 1368 -2604 1374 -2598
rect 1368 -2610 1374 -2604
rect 1368 -2616 1374 -2610
rect 1368 -2622 1374 -2616
rect 1368 -2628 1374 -2622
rect 1368 -2634 1374 -2628
rect 1368 -2640 1374 -2634
rect 1368 -2646 1374 -2640
rect 1368 -2652 1374 -2646
rect 1368 -2658 1374 -2652
rect 1368 -2664 1374 -2658
rect 1368 -2670 1374 -2664
rect 1368 -2676 1374 -2670
rect 1368 -2682 1374 -2676
rect 1368 -2688 1374 -2682
rect 1368 -2694 1374 -2688
rect 1368 -2700 1374 -2694
rect 1368 -2706 1374 -2700
rect 1368 -2712 1374 -2706
rect 1368 -2718 1374 -2712
rect 1368 -2724 1374 -2718
rect 1368 -2730 1374 -2724
rect 1368 -2736 1374 -2730
rect 1368 -2742 1374 -2736
rect 1368 -2748 1374 -2742
rect 1368 -2754 1374 -2748
rect 1368 -2760 1374 -2754
rect 1368 -2766 1374 -2760
rect 1368 -2772 1374 -2766
rect 1368 -2778 1374 -2772
rect 1368 -2784 1374 -2778
rect 1368 -2790 1374 -2784
rect 1368 -2796 1374 -2790
rect 1368 -2802 1374 -2796
rect 1368 -2808 1374 -2802
rect 1368 -2814 1374 -2808
rect 1368 -2820 1374 -2814
rect 1368 -2826 1374 -2820
rect 1368 -2832 1374 -2826
rect 1368 -2838 1374 -2832
rect 1368 -2844 1374 -2838
rect 1368 -2850 1374 -2844
rect 1368 -2856 1374 -2850
rect 1368 -2862 1374 -2856
rect 1368 -2868 1374 -2862
rect 1368 -2874 1374 -2868
rect 1368 -2880 1374 -2874
rect 1368 -2886 1374 -2880
rect 1368 -2892 1374 -2886
rect 1368 -2898 1374 -2892
rect 1368 -2982 1374 -2976
rect 1368 -2988 1374 -2982
rect 1368 -2994 1374 -2988
rect 1368 -3000 1374 -2994
rect 1368 -3006 1374 -3000
rect 1368 -3012 1374 -3006
rect 1368 -3018 1374 -3012
rect 1368 -3024 1374 -3018
rect 1368 -3030 1374 -3024
rect 1368 -3036 1374 -3030
rect 1368 -3042 1374 -3036
rect 1368 -3048 1374 -3042
rect 1368 -3054 1374 -3048
rect 1368 -3060 1374 -3054
rect 1368 -3066 1374 -3060
rect 1368 -3072 1374 -3066
rect 1368 -3078 1374 -3072
rect 1368 -3084 1374 -3078
rect 1368 -3090 1374 -3084
rect 1368 -3096 1374 -3090
rect 1368 -3102 1374 -3096
rect 1368 -3108 1374 -3102
rect 1368 -3114 1374 -3108
rect 1368 -3120 1374 -3114
rect 1368 -3126 1374 -3120
rect 1368 -3132 1374 -3126
rect 1368 -3138 1374 -3132
rect 1368 -3144 1374 -3138
rect 1368 -3150 1374 -3144
rect 1368 -3156 1374 -3150
rect 1368 -3162 1374 -3156
rect 1368 -3168 1374 -3162
rect 1368 -3174 1374 -3168
rect 1368 -3180 1374 -3174
rect 1368 -3186 1374 -3180
rect 1368 -3192 1374 -3186
rect 1368 -3198 1374 -3192
rect 1368 -3204 1374 -3198
rect 1368 -3210 1374 -3204
rect 1368 -3216 1374 -3210
rect 1368 -3222 1374 -3216
rect 1368 -3228 1374 -3222
rect 1368 -3234 1374 -3228
rect 1368 -3312 1374 -3306
rect 1368 -3318 1374 -3312
rect 1368 -3324 1374 -3318
rect 1368 -3330 1374 -3324
rect 1368 -3336 1374 -3330
rect 1368 -3342 1374 -3336
rect 1368 -3348 1374 -3342
rect 1368 -3354 1374 -3348
rect 1368 -3360 1374 -3354
rect 1368 -3366 1374 -3360
rect 1368 -3372 1374 -3366
rect 1368 -3378 1374 -3372
rect 1368 -3384 1374 -3378
rect 1368 -3390 1374 -3384
rect 1368 -3396 1374 -3390
rect 1368 -3402 1374 -3396
rect 1368 -3408 1374 -3402
rect 1368 -3414 1374 -3408
rect 1368 -3420 1374 -3414
rect 1368 -3426 1374 -3420
rect 1368 -3432 1374 -3426
rect 1368 -3438 1374 -3432
rect 1368 -3444 1374 -3438
rect 1368 -3450 1374 -3444
rect 1368 -3456 1374 -3450
rect 1368 -3462 1374 -3456
rect 1368 -3468 1374 -3462
rect 1368 -3474 1374 -3468
rect 1368 -3480 1374 -3474
rect 1368 -3486 1374 -3480
rect 1368 -3492 1374 -3486
rect 1368 -3498 1374 -3492
rect 1368 -3504 1374 -3498
rect 1368 -3510 1374 -3504
rect 1374 -1116 1380 -1110
rect 1374 -1122 1380 -1116
rect 1374 -1128 1380 -1122
rect 1374 -1134 1380 -1128
rect 1374 -1140 1380 -1134
rect 1374 -1146 1380 -1140
rect 1374 -1152 1380 -1146
rect 1374 -1158 1380 -1152
rect 1374 -1164 1380 -1158
rect 1374 -1170 1380 -1164
rect 1374 -1176 1380 -1170
rect 1374 -1182 1380 -1176
rect 1374 -1188 1380 -1182
rect 1374 -1194 1380 -1188
rect 1374 -1200 1380 -1194
rect 1374 -1206 1380 -1200
rect 1374 -1212 1380 -1206
rect 1374 -1218 1380 -1212
rect 1374 -1224 1380 -1218
rect 1374 -1230 1380 -1224
rect 1374 -1236 1380 -1230
rect 1374 -1242 1380 -1236
rect 1374 -1248 1380 -1242
rect 1374 -1254 1380 -1248
rect 1374 -1260 1380 -1254
rect 1374 -1266 1380 -1260
rect 1374 -1272 1380 -1266
rect 1374 -1278 1380 -1272
rect 1374 -1284 1380 -1278
rect 1374 -1290 1380 -1284
rect 1374 -1296 1380 -1290
rect 1374 -1416 1380 -1410
rect 1374 -1422 1380 -1416
rect 1374 -1428 1380 -1422
rect 1374 -1434 1380 -1428
rect 1374 -1440 1380 -1434
rect 1374 -1446 1380 -1440
rect 1374 -1452 1380 -1446
rect 1374 -1458 1380 -1452
rect 1374 -1464 1380 -1458
rect 1374 -1470 1380 -1464
rect 1374 -1476 1380 -1470
rect 1374 -1482 1380 -1476
rect 1374 -1488 1380 -1482
rect 1374 -1494 1380 -1488
rect 1374 -1500 1380 -1494
rect 1374 -1506 1380 -1500
rect 1374 -1512 1380 -1506
rect 1374 -1518 1380 -1512
rect 1374 -1524 1380 -1518
rect 1374 -1530 1380 -1524
rect 1374 -1536 1380 -1530
rect 1374 -1542 1380 -1536
rect 1374 -1548 1380 -1542
rect 1374 -1554 1380 -1548
rect 1374 -1560 1380 -1554
rect 1374 -1566 1380 -1560
rect 1374 -1572 1380 -1566
rect 1374 -1578 1380 -1572
rect 1374 -1584 1380 -1578
rect 1374 -1590 1380 -1584
rect 1374 -1596 1380 -1590
rect 1374 -1602 1380 -1596
rect 1374 -1608 1380 -1602
rect 1374 -1614 1380 -1608
rect 1374 -1620 1380 -1614
rect 1374 -1626 1380 -1620
rect 1374 -1632 1380 -1626
rect 1374 -1638 1380 -1632
rect 1374 -1644 1380 -1638
rect 1374 -1650 1380 -1644
rect 1374 -1656 1380 -1650
rect 1374 -1662 1380 -1656
rect 1374 -1668 1380 -1662
rect 1374 -1674 1380 -1668
rect 1374 -1680 1380 -1674
rect 1374 -1686 1380 -1680
rect 1374 -1692 1380 -1686
rect 1374 -1698 1380 -1692
rect 1374 -1704 1380 -1698
rect 1374 -1710 1380 -1704
rect 1374 -1716 1380 -1710
rect 1374 -1722 1380 -1716
rect 1374 -1728 1380 -1722
rect 1374 -1734 1380 -1728
rect 1374 -1740 1380 -1734
rect 1374 -1746 1380 -1740
rect 1374 -1752 1380 -1746
rect 1374 -1758 1380 -1752
rect 1374 -1764 1380 -1758
rect 1374 -1770 1380 -1764
rect 1374 -1776 1380 -1770
rect 1374 -1782 1380 -1776
rect 1374 -1788 1380 -1782
rect 1374 -1794 1380 -1788
rect 1374 -1800 1380 -1794
rect 1374 -1806 1380 -1800
rect 1374 -1812 1380 -1806
rect 1374 -1818 1380 -1812
rect 1374 -1824 1380 -1818
rect 1374 -1830 1380 -1824
rect 1374 -1836 1380 -1830
rect 1374 -1842 1380 -1836
rect 1374 -1848 1380 -1842
rect 1374 -1854 1380 -1848
rect 1374 -1860 1380 -1854
rect 1374 -1866 1380 -1860
rect 1374 -1872 1380 -1866
rect 1374 -1878 1380 -1872
rect 1374 -1884 1380 -1878
rect 1374 -1890 1380 -1884
rect 1374 -1896 1380 -1890
rect 1374 -1902 1380 -1896
rect 1374 -1908 1380 -1902
rect 1374 -1914 1380 -1908
rect 1374 -1920 1380 -1914
rect 1374 -1926 1380 -1920
rect 1374 -1932 1380 -1926
rect 1374 -1938 1380 -1932
rect 1374 -1944 1380 -1938
rect 1374 -1950 1380 -1944
rect 1374 -1956 1380 -1950
rect 1374 -1962 1380 -1956
rect 1374 -1968 1380 -1962
rect 1374 -1974 1380 -1968
rect 1374 -1980 1380 -1974
rect 1374 -1986 1380 -1980
rect 1374 -1992 1380 -1986
rect 1374 -1998 1380 -1992
rect 1374 -2004 1380 -1998
rect 1374 -2010 1380 -2004
rect 1374 -2016 1380 -2010
rect 1374 -2022 1380 -2016
rect 1374 -2028 1380 -2022
rect 1374 -2034 1380 -2028
rect 1374 -2040 1380 -2034
rect 1374 -2046 1380 -2040
rect 1374 -2052 1380 -2046
rect 1374 -2058 1380 -2052
rect 1374 -2064 1380 -2058
rect 1374 -2070 1380 -2064
rect 1374 -2076 1380 -2070
rect 1374 -2082 1380 -2076
rect 1374 -2088 1380 -2082
rect 1374 -2094 1380 -2088
rect 1374 -2100 1380 -2094
rect 1374 -2106 1380 -2100
rect 1374 -2112 1380 -2106
rect 1374 -2118 1380 -2112
rect 1374 -2124 1380 -2118
rect 1374 -2130 1380 -2124
rect 1374 -2136 1380 -2130
rect 1374 -2142 1380 -2136
rect 1374 -2148 1380 -2142
rect 1374 -2154 1380 -2148
rect 1374 -2160 1380 -2154
rect 1374 -2166 1380 -2160
rect 1374 -2172 1380 -2166
rect 1374 -2178 1380 -2172
rect 1374 -2184 1380 -2178
rect 1374 -2190 1380 -2184
rect 1374 -2196 1380 -2190
rect 1374 -2202 1380 -2196
rect 1374 -2208 1380 -2202
rect 1374 -2214 1380 -2208
rect 1374 -2220 1380 -2214
rect 1374 -2226 1380 -2220
rect 1374 -2232 1380 -2226
rect 1374 -2238 1380 -2232
rect 1374 -2244 1380 -2238
rect 1374 -2250 1380 -2244
rect 1374 -2256 1380 -2250
rect 1374 -2262 1380 -2256
rect 1374 -2268 1380 -2262
rect 1374 -2274 1380 -2268
rect 1374 -2280 1380 -2274
rect 1374 -2286 1380 -2280
rect 1374 -2292 1380 -2286
rect 1374 -2298 1380 -2292
rect 1374 -2304 1380 -2298
rect 1374 -2310 1380 -2304
rect 1374 -2316 1380 -2310
rect 1374 -2322 1380 -2316
rect 1374 -2328 1380 -2322
rect 1374 -2334 1380 -2328
rect 1374 -2340 1380 -2334
rect 1374 -2346 1380 -2340
rect 1374 -2352 1380 -2346
rect 1374 -2358 1380 -2352
rect 1374 -2436 1380 -2430
rect 1374 -2442 1380 -2436
rect 1374 -2448 1380 -2442
rect 1374 -2454 1380 -2448
rect 1374 -2460 1380 -2454
rect 1374 -2466 1380 -2460
rect 1374 -2472 1380 -2466
rect 1374 -2478 1380 -2472
rect 1374 -2484 1380 -2478
rect 1374 -2490 1380 -2484
rect 1374 -2496 1380 -2490
rect 1374 -2502 1380 -2496
rect 1374 -2508 1380 -2502
rect 1374 -2514 1380 -2508
rect 1374 -2520 1380 -2514
rect 1374 -2526 1380 -2520
rect 1374 -2532 1380 -2526
rect 1374 -2538 1380 -2532
rect 1374 -2544 1380 -2538
rect 1374 -2550 1380 -2544
rect 1374 -2556 1380 -2550
rect 1374 -2562 1380 -2556
rect 1374 -2568 1380 -2562
rect 1374 -2574 1380 -2568
rect 1374 -2580 1380 -2574
rect 1374 -2586 1380 -2580
rect 1374 -2592 1380 -2586
rect 1374 -2598 1380 -2592
rect 1374 -2604 1380 -2598
rect 1374 -2610 1380 -2604
rect 1374 -2616 1380 -2610
rect 1374 -2622 1380 -2616
rect 1374 -2628 1380 -2622
rect 1374 -2634 1380 -2628
rect 1374 -2640 1380 -2634
rect 1374 -2646 1380 -2640
rect 1374 -2652 1380 -2646
rect 1374 -2658 1380 -2652
rect 1374 -2664 1380 -2658
rect 1374 -2670 1380 -2664
rect 1374 -2676 1380 -2670
rect 1374 -2682 1380 -2676
rect 1374 -2688 1380 -2682
rect 1374 -2694 1380 -2688
rect 1374 -2700 1380 -2694
rect 1374 -2706 1380 -2700
rect 1374 -2712 1380 -2706
rect 1374 -2718 1380 -2712
rect 1374 -2724 1380 -2718
rect 1374 -2730 1380 -2724
rect 1374 -2736 1380 -2730
rect 1374 -2742 1380 -2736
rect 1374 -2748 1380 -2742
rect 1374 -2754 1380 -2748
rect 1374 -2760 1380 -2754
rect 1374 -2766 1380 -2760
rect 1374 -2772 1380 -2766
rect 1374 -2778 1380 -2772
rect 1374 -2784 1380 -2778
rect 1374 -2790 1380 -2784
rect 1374 -2796 1380 -2790
rect 1374 -2802 1380 -2796
rect 1374 -2808 1380 -2802
rect 1374 -2814 1380 -2808
rect 1374 -2820 1380 -2814
rect 1374 -2826 1380 -2820
rect 1374 -2832 1380 -2826
rect 1374 -2838 1380 -2832
rect 1374 -2844 1380 -2838
rect 1374 -2850 1380 -2844
rect 1374 -2856 1380 -2850
rect 1374 -2862 1380 -2856
rect 1374 -2868 1380 -2862
rect 1374 -2874 1380 -2868
rect 1374 -2880 1380 -2874
rect 1374 -2886 1380 -2880
rect 1374 -2892 1380 -2886
rect 1374 -2976 1380 -2970
rect 1374 -2982 1380 -2976
rect 1374 -2988 1380 -2982
rect 1374 -2994 1380 -2988
rect 1374 -3000 1380 -2994
rect 1374 -3006 1380 -3000
rect 1374 -3012 1380 -3006
rect 1374 -3018 1380 -3012
rect 1374 -3024 1380 -3018
rect 1374 -3030 1380 -3024
rect 1374 -3036 1380 -3030
rect 1374 -3042 1380 -3036
rect 1374 -3048 1380 -3042
rect 1374 -3054 1380 -3048
rect 1374 -3060 1380 -3054
rect 1374 -3066 1380 -3060
rect 1374 -3072 1380 -3066
rect 1374 -3078 1380 -3072
rect 1374 -3084 1380 -3078
rect 1374 -3090 1380 -3084
rect 1374 -3096 1380 -3090
rect 1374 -3102 1380 -3096
rect 1374 -3108 1380 -3102
rect 1374 -3114 1380 -3108
rect 1374 -3120 1380 -3114
rect 1374 -3126 1380 -3120
rect 1374 -3132 1380 -3126
rect 1374 -3138 1380 -3132
rect 1374 -3144 1380 -3138
rect 1374 -3150 1380 -3144
rect 1374 -3156 1380 -3150
rect 1374 -3162 1380 -3156
rect 1374 -3168 1380 -3162
rect 1374 -3174 1380 -3168
rect 1374 -3180 1380 -3174
rect 1374 -3186 1380 -3180
rect 1374 -3192 1380 -3186
rect 1374 -3198 1380 -3192
rect 1374 -3204 1380 -3198
rect 1374 -3210 1380 -3204
rect 1374 -3216 1380 -3210
rect 1374 -3222 1380 -3216
rect 1374 -3228 1380 -3222
rect 1374 -3234 1380 -3228
rect 1374 -3306 1380 -3300
rect 1374 -3312 1380 -3306
rect 1374 -3318 1380 -3312
rect 1374 -3324 1380 -3318
rect 1374 -3330 1380 -3324
rect 1374 -3336 1380 -3330
rect 1374 -3342 1380 -3336
rect 1374 -3348 1380 -3342
rect 1374 -3354 1380 -3348
rect 1374 -3360 1380 -3354
rect 1374 -3366 1380 -3360
rect 1374 -3372 1380 -3366
rect 1374 -3378 1380 -3372
rect 1374 -3384 1380 -3378
rect 1374 -3390 1380 -3384
rect 1374 -3396 1380 -3390
rect 1374 -3402 1380 -3396
rect 1374 -3408 1380 -3402
rect 1374 -3414 1380 -3408
rect 1374 -3420 1380 -3414
rect 1374 -3426 1380 -3420
rect 1374 -3432 1380 -3426
rect 1374 -3438 1380 -3432
rect 1374 -3444 1380 -3438
rect 1374 -3450 1380 -3444
rect 1374 -3456 1380 -3450
rect 1374 -3462 1380 -3456
rect 1374 -3468 1380 -3462
rect 1374 -3474 1380 -3468
rect 1374 -3480 1380 -3474
rect 1374 -3486 1380 -3480
rect 1374 -3492 1380 -3486
rect 1374 -3498 1380 -3492
rect 1374 -3504 1380 -3498
rect 1374 -3510 1380 -3504
rect 1380 -1116 1386 -1110
rect 1380 -1122 1386 -1116
rect 1380 -1128 1386 -1122
rect 1380 -1134 1386 -1128
rect 1380 -1140 1386 -1134
rect 1380 -1146 1386 -1140
rect 1380 -1152 1386 -1146
rect 1380 -1158 1386 -1152
rect 1380 -1164 1386 -1158
rect 1380 -1170 1386 -1164
rect 1380 -1176 1386 -1170
rect 1380 -1182 1386 -1176
rect 1380 -1188 1386 -1182
rect 1380 -1194 1386 -1188
rect 1380 -1200 1386 -1194
rect 1380 -1206 1386 -1200
rect 1380 -1212 1386 -1206
rect 1380 -1218 1386 -1212
rect 1380 -1224 1386 -1218
rect 1380 -1230 1386 -1224
rect 1380 -1236 1386 -1230
rect 1380 -1242 1386 -1236
rect 1380 -1248 1386 -1242
rect 1380 -1254 1386 -1248
rect 1380 -1260 1386 -1254
rect 1380 -1266 1386 -1260
rect 1380 -1272 1386 -1266
rect 1380 -1278 1386 -1272
rect 1380 -1284 1386 -1278
rect 1380 -1404 1386 -1398
rect 1380 -1410 1386 -1404
rect 1380 -1416 1386 -1410
rect 1380 -1422 1386 -1416
rect 1380 -1428 1386 -1422
rect 1380 -1434 1386 -1428
rect 1380 -1440 1386 -1434
rect 1380 -1446 1386 -1440
rect 1380 -1452 1386 -1446
rect 1380 -1458 1386 -1452
rect 1380 -1464 1386 -1458
rect 1380 -1470 1386 -1464
rect 1380 -1476 1386 -1470
rect 1380 -1482 1386 -1476
rect 1380 -1488 1386 -1482
rect 1380 -1494 1386 -1488
rect 1380 -1500 1386 -1494
rect 1380 -1506 1386 -1500
rect 1380 -1512 1386 -1506
rect 1380 -1518 1386 -1512
rect 1380 -1524 1386 -1518
rect 1380 -1530 1386 -1524
rect 1380 -1536 1386 -1530
rect 1380 -1542 1386 -1536
rect 1380 -1548 1386 -1542
rect 1380 -1554 1386 -1548
rect 1380 -1560 1386 -1554
rect 1380 -1566 1386 -1560
rect 1380 -1572 1386 -1566
rect 1380 -1578 1386 -1572
rect 1380 -1584 1386 -1578
rect 1380 -1590 1386 -1584
rect 1380 -1596 1386 -1590
rect 1380 -1602 1386 -1596
rect 1380 -1608 1386 -1602
rect 1380 -1614 1386 -1608
rect 1380 -1620 1386 -1614
rect 1380 -1626 1386 -1620
rect 1380 -1632 1386 -1626
rect 1380 -1638 1386 -1632
rect 1380 -1644 1386 -1638
rect 1380 -1650 1386 -1644
rect 1380 -1656 1386 -1650
rect 1380 -1662 1386 -1656
rect 1380 -1668 1386 -1662
rect 1380 -1674 1386 -1668
rect 1380 -1680 1386 -1674
rect 1380 -1686 1386 -1680
rect 1380 -1692 1386 -1686
rect 1380 -1698 1386 -1692
rect 1380 -1704 1386 -1698
rect 1380 -1710 1386 -1704
rect 1380 -1716 1386 -1710
rect 1380 -1722 1386 -1716
rect 1380 -1728 1386 -1722
rect 1380 -1734 1386 -1728
rect 1380 -1740 1386 -1734
rect 1380 -1746 1386 -1740
rect 1380 -1752 1386 -1746
rect 1380 -1758 1386 -1752
rect 1380 -1764 1386 -1758
rect 1380 -1770 1386 -1764
rect 1380 -1776 1386 -1770
rect 1380 -1782 1386 -1776
rect 1380 -1788 1386 -1782
rect 1380 -1794 1386 -1788
rect 1380 -1800 1386 -1794
rect 1380 -1806 1386 -1800
rect 1380 -1812 1386 -1806
rect 1380 -1818 1386 -1812
rect 1380 -1824 1386 -1818
rect 1380 -1830 1386 -1824
rect 1380 -1836 1386 -1830
rect 1380 -1842 1386 -1836
rect 1380 -1848 1386 -1842
rect 1380 -1854 1386 -1848
rect 1380 -1860 1386 -1854
rect 1380 -1866 1386 -1860
rect 1380 -1872 1386 -1866
rect 1380 -1878 1386 -1872
rect 1380 -1884 1386 -1878
rect 1380 -1890 1386 -1884
rect 1380 -1896 1386 -1890
rect 1380 -1902 1386 -1896
rect 1380 -1908 1386 -1902
rect 1380 -1914 1386 -1908
rect 1380 -1920 1386 -1914
rect 1380 -1926 1386 -1920
rect 1380 -1932 1386 -1926
rect 1380 -1938 1386 -1932
rect 1380 -1944 1386 -1938
rect 1380 -1950 1386 -1944
rect 1380 -1956 1386 -1950
rect 1380 -1962 1386 -1956
rect 1380 -1968 1386 -1962
rect 1380 -1974 1386 -1968
rect 1380 -1980 1386 -1974
rect 1380 -1986 1386 -1980
rect 1380 -1992 1386 -1986
rect 1380 -1998 1386 -1992
rect 1380 -2004 1386 -1998
rect 1380 -2010 1386 -2004
rect 1380 -2016 1386 -2010
rect 1380 -2022 1386 -2016
rect 1380 -2028 1386 -2022
rect 1380 -2034 1386 -2028
rect 1380 -2040 1386 -2034
rect 1380 -2046 1386 -2040
rect 1380 -2052 1386 -2046
rect 1380 -2058 1386 -2052
rect 1380 -2064 1386 -2058
rect 1380 -2070 1386 -2064
rect 1380 -2076 1386 -2070
rect 1380 -2082 1386 -2076
rect 1380 -2088 1386 -2082
rect 1380 -2094 1386 -2088
rect 1380 -2100 1386 -2094
rect 1380 -2106 1386 -2100
rect 1380 -2112 1386 -2106
rect 1380 -2118 1386 -2112
rect 1380 -2124 1386 -2118
rect 1380 -2130 1386 -2124
rect 1380 -2136 1386 -2130
rect 1380 -2142 1386 -2136
rect 1380 -2148 1386 -2142
rect 1380 -2154 1386 -2148
rect 1380 -2160 1386 -2154
rect 1380 -2166 1386 -2160
rect 1380 -2172 1386 -2166
rect 1380 -2178 1386 -2172
rect 1380 -2184 1386 -2178
rect 1380 -2190 1386 -2184
rect 1380 -2196 1386 -2190
rect 1380 -2202 1386 -2196
rect 1380 -2208 1386 -2202
rect 1380 -2214 1386 -2208
rect 1380 -2220 1386 -2214
rect 1380 -2226 1386 -2220
rect 1380 -2232 1386 -2226
rect 1380 -2238 1386 -2232
rect 1380 -2244 1386 -2238
rect 1380 -2250 1386 -2244
rect 1380 -2256 1386 -2250
rect 1380 -2262 1386 -2256
rect 1380 -2268 1386 -2262
rect 1380 -2274 1386 -2268
rect 1380 -2280 1386 -2274
rect 1380 -2286 1386 -2280
rect 1380 -2292 1386 -2286
rect 1380 -2298 1386 -2292
rect 1380 -2304 1386 -2298
rect 1380 -2310 1386 -2304
rect 1380 -2316 1386 -2310
rect 1380 -2322 1386 -2316
rect 1380 -2328 1386 -2322
rect 1380 -2334 1386 -2328
rect 1380 -2340 1386 -2334
rect 1380 -2346 1386 -2340
rect 1380 -2352 1386 -2346
rect 1380 -2430 1386 -2424
rect 1380 -2436 1386 -2430
rect 1380 -2442 1386 -2436
rect 1380 -2448 1386 -2442
rect 1380 -2454 1386 -2448
rect 1380 -2460 1386 -2454
rect 1380 -2466 1386 -2460
rect 1380 -2472 1386 -2466
rect 1380 -2478 1386 -2472
rect 1380 -2484 1386 -2478
rect 1380 -2490 1386 -2484
rect 1380 -2496 1386 -2490
rect 1380 -2502 1386 -2496
rect 1380 -2508 1386 -2502
rect 1380 -2514 1386 -2508
rect 1380 -2520 1386 -2514
rect 1380 -2526 1386 -2520
rect 1380 -2532 1386 -2526
rect 1380 -2538 1386 -2532
rect 1380 -2544 1386 -2538
rect 1380 -2550 1386 -2544
rect 1380 -2556 1386 -2550
rect 1380 -2562 1386 -2556
rect 1380 -2568 1386 -2562
rect 1380 -2574 1386 -2568
rect 1380 -2580 1386 -2574
rect 1380 -2586 1386 -2580
rect 1380 -2592 1386 -2586
rect 1380 -2598 1386 -2592
rect 1380 -2604 1386 -2598
rect 1380 -2610 1386 -2604
rect 1380 -2616 1386 -2610
rect 1380 -2622 1386 -2616
rect 1380 -2628 1386 -2622
rect 1380 -2634 1386 -2628
rect 1380 -2640 1386 -2634
rect 1380 -2646 1386 -2640
rect 1380 -2652 1386 -2646
rect 1380 -2658 1386 -2652
rect 1380 -2664 1386 -2658
rect 1380 -2670 1386 -2664
rect 1380 -2676 1386 -2670
rect 1380 -2682 1386 -2676
rect 1380 -2688 1386 -2682
rect 1380 -2694 1386 -2688
rect 1380 -2700 1386 -2694
rect 1380 -2706 1386 -2700
rect 1380 -2712 1386 -2706
rect 1380 -2718 1386 -2712
rect 1380 -2724 1386 -2718
rect 1380 -2730 1386 -2724
rect 1380 -2736 1386 -2730
rect 1380 -2742 1386 -2736
rect 1380 -2748 1386 -2742
rect 1380 -2754 1386 -2748
rect 1380 -2760 1386 -2754
rect 1380 -2766 1386 -2760
rect 1380 -2772 1386 -2766
rect 1380 -2778 1386 -2772
rect 1380 -2784 1386 -2778
rect 1380 -2790 1386 -2784
rect 1380 -2796 1386 -2790
rect 1380 -2802 1386 -2796
rect 1380 -2808 1386 -2802
rect 1380 -2814 1386 -2808
rect 1380 -2820 1386 -2814
rect 1380 -2826 1386 -2820
rect 1380 -2832 1386 -2826
rect 1380 -2838 1386 -2832
rect 1380 -2844 1386 -2838
rect 1380 -2850 1386 -2844
rect 1380 -2856 1386 -2850
rect 1380 -2862 1386 -2856
rect 1380 -2868 1386 -2862
rect 1380 -2874 1386 -2868
rect 1380 -2880 1386 -2874
rect 1380 -2886 1386 -2880
rect 1380 -2976 1386 -2970
rect 1380 -2982 1386 -2976
rect 1380 -2988 1386 -2982
rect 1380 -2994 1386 -2988
rect 1380 -3000 1386 -2994
rect 1380 -3006 1386 -3000
rect 1380 -3012 1386 -3006
rect 1380 -3018 1386 -3012
rect 1380 -3024 1386 -3018
rect 1380 -3030 1386 -3024
rect 1380 -3036 1386 -3030
rect 1380 -3042 1386 -3036
rect 1380 -3048 1386 -3042
rect 1380 -3054 1386 -3048
rect 1380 -3060 1386 -3054
rect 1380 -3066 1386 -3060
rect 1380 -3072 1386 -3066
rect 1380 -3078 1386 -3072
rect 1380 -3084 1386 -3078
rect 1380 -3090 1386 -3084
rect 1380 -3096 1386 -3090
rect 1380 -3102 1386 -3096
rect 1380 -3108 1386 -3102
rect 1380 -3114 1386 -3108
rect 1380 -3120 1386 -3114
rect 1380 -3126 1386 -3120
rect 1380 -3132 1386 -3126
rect 1380 -3138 1386 -3132
rect 1380 -3144 1386 -3138
rect 1380 -3150 1386 -3144
rect 1380 -3156 1386 -3150
rect 1380 -3162 1386 -3156
rect 1380 -3168 1386 -3162
rect 1380 -3174 1386 -3168
rect 1380 -3180 1386 -3174
rect 1380 -3186 1386 -3180
rect 1380 -3192 1386 -3186
rect 1380 -3198 1386 -3192
rect 1380 -3204 1386 -3198
rect 1380 -3210 1386 -3204
rect 1380 -3216 1386 -3210
rect 1380 -3222 1386 -3216
rect 1380 -3228 1386 -3222
rect 1380 -3234 1386 -3228
rect 1380 -3306 1386 -3300
rect 1380 -3312 1386 -3306
rect 1380 -3318 1386 -3312
rect 1380 -3324 1386 -3318
rect 1380 -3330 1386 -3324
rect 1380 -3336 1386 -3330
rect 1380 -3342 1386 -3336
rect 1380 -3348 1386 -3342
rect 1380 -3354 1386 -3348
rect 1380 -3360 1386 -3354
rect 1380 -3366 1386 -3360
rect 1380 -3372 1386 -3366
rect 1380 -3378 1386 -3372
rect 1380 -3384 1386 -3378
rect 1380 -3390 1386 -3384
rect 1380 -3396 1386 -3390
rect 1380 -3402 1386 -3396
rect 1380 -3408 1386 -3402
rect 1380 -3414 1386 -3408
rect 1380 -3420 1386 -3414
rect 1380 -3426 1386 -3420
rect 1380 -3432 1386 -3426
rect 1380 -3438 1386 -3432
rect 1380 -3444 1386 -3438
rect 1380 -3450 1386 -3444
rect 1380 -3456 1386 -3450
rect 1380 -3462 1386 -3456
rect 1380 -3468 1386 -3462
rect 1380 -3474 1386 -3468
rect 1380 -3480 1386 -3474
rect 1380 -3486 1386 -3480
rect 1380 -3492 1386 -3486
rect 1380 -3498 1386 -3492
rect 1380 -3504 1386 -3498
rect 1380 -3510 1386 -3504
rect 1386 -1116 1392 -1110
rect 1386 -1122 1392 -1116
rect 1386 -1128 1392 -1122
rect 1386 -1134 1392 -1128
rect 1386 -1140 1392 -1134
rect 1386 -1146 1392 -1140
rect 1386 -1152 1392 -1146
rect 1386 -1158 1392 -1152
rect 1386 -1164 1392 -1158
rect 1386 -1170 1392 -1164
rect 1386 -1176 1392 -1170
rect 1386 -1182 1392 -1176
rect 1386 -1188 1392 -1182
rect 1386 -1194 1392 -1188
rect 1386 -1200 1392 -1194
rect 1386 -1206 1392 -1200
rect 1386 -1212 1392 -1206
rect 1386 -1218 1392 -1212
rect 1386 -1224 1392 -1218
rect 1386 -1230 1392 -1224
rect 1386 -1236 1392 -1230
rect 1386 -1242 1392 -1236
rect 1386 -1248 1392 -1242
rect 1386 -1254 1392 -1248
rect 1386 -1260 1392 -1254
rect 1386 -1266 1392 -1260
rect 1386 -1272 1392 -1266
rect 1386 -1392 1392 -1386
rect 1386 -1398 1392 -1392
rect 1386 -1404 1392 -1398
rect 1386 -1410 1392 -1404
rect 1386 -1416 1392 -1410
rect 1386 -1422 1392 -1416
rect 1386 -1428 1392 -1422
rect 1386 -1434 1392 -1428
rect 1386 -1440 1392 -1434
rect 1386 -1446 1392 -1440
rect 1386 -1452 1392 -1446
rect 1386 -1458 1392 -1452
rect 1386 -1464 1392 -1458
rect 1386 -1470 1392 -1464
rect 1386 -1476 1392 -1470
rect 1386 -1482 1392 -1476
rect 1386 -1488 1392 -1482
rect 1386 -1494 1392 -1488
rect 1386 -1500 1392 -1494
rect 1386 -1506 1392 -1500
rect 1386 -1512 1392 -1506
rect 1386 -1518 1392 -1512
rect 1386 -1524 1392 -1518
rect 1386 -1530 1392 -1524
rect 1386 -1536 1392 -1530
rect 1386 -1542 1392 -1536
rect 1386 -1548 1392 -1542
rect 1386 -1554 1392 -1548
rect 1386 -1560 1392 -1554
rect 1386 -1566 1392 -1560
rect 1386 -1572 1392 -1566
rect 1386 -1578 1392 -1572
rect 1386 -1584 1392 -1578
rect 1386 -1590 1392 -1584
rect 1386 -1596 1392 -1590
rect 1386 -1602 1392 -1596
rect 1386 -1608 1392 -1602
rect 1386 -1614 1392 -1608
rect 1386 -1620 1392 -1614
rect 1386 -1626 1392 -1620
rect 1386 -1632 1392 -1626
rect 1386 -1638 1392 -1632
rect 1386 -1644 1392 -1638
rect 1386 -1650 1392 -1644
rect 1386 -1656 1392 -1650
rect 1386 -1662 1392 -1656
rect 1386 -1668 1392 -1662
rect 1386 -1674 1392 -1668
rect 1386 -1680 1392 -1674
rect 1386 -1686 1392 -1680
rect 1386 -1692 1392 -1686
rect 1386 -1698 1392 -1692
rect 1386 -1704 1392 -1698
rect 1386 -1710 1392 -1704
rect 1386 -1716 1392 -1710
rect 1386 -1722 1392 -1716
rect 1386 -1728 1392 -1722
rect 1386 -1734 1392 -1728
rect 1386 -1740 1392 -1734
rect 1386 -1746 1392 -1740
rect 1386 -1752 1392 -1746
rect 1386 -1758 1392 -1752
rect 1386 -1764 1392 -1758
rect 1386 -1770 1392 -1764
rect 1386 -1776 1392 -1770
rect 1386 -1782 1392 -1776
rect 1386 -1788 1392 -1782
rect 1386 -1794 1392 -1788
rect 1386 -1800 1392 -1794
rect 1386 -1806 1392 -1800
rect 1386 -1812 1392 -1806
rect 1386 -1818 1392 -1812
rect 1386 -1824 1392 -1818
rect 1386 -1830 1392 -1824
rect 1386 -1836 1392 -1830
rect 1386 -1842 1392 -1836
rect 1386 -1848 1392 -1842
rect 1386 -1854 1392 -1848
rect 1386 -1860 1392 -1854
rect 1386 -1866 1392 -1860
rect 1386 -1872 1392 -1866
rect 1386 -1878 1392 -1872
rect 1386 -1884 1392 -1878
rect 1386 -1890 1392 -1884
rect 1386 -1896 1392 -1890
rect 1386 -1902 1392 -1896
rect 1386 -1908 1392 -1902
rect 1386 -1914 1392 -1908
rect 1386 -1920 1392 -1914
rect 1386 -1926 1392 -1920
rect 1386 -1932 1392 -1926
rect 1386 -1938 1392 -1932
rect 1386 -1944 1392 -1938
rect 1386 -1950 1392 -1944
rect 1386 -1956 1392 -1950
rect 1386 -1962 1392 -1956
rect 1386 -1968 1392 -1962
rect 1386 -1974 1392 -1968
rect 1386 -1980 1392 -1974
rect 1386 -1986 1392 -1980
rect 1386 -1992 1392 -1986
rect 1386 -1998 1392 -1992
rect 1386 -2004 1392 -1998
rect 1386 -2010 1392 -2004
rect 1386 -2016 1392 -2010
rect 1386 -2022 1392 -2016
rect 1386 -2028 1392 -2022
rect 1386 -2034 1392 -2028
rect 1386 -2040 1392 -2034
rect 1386 -2046 1392 -2040
rect 1386 -2052 1392 -2046
rect 1386 -2058 1392 -2052
rect 1386 -2064 1392 -2058
rect 1386 -2070 1392 -2064
rect 1386 -2076 1392 -2070
rect 1386 -2082 1392 -2076
rect 1386 -2088 1392 -2082
rect 1386 -2094 1392 -2088
rect 1386 -2100 1392 -2094
rect 1386 -2106 1392 -2100
rect 1386 -2112 1392 -2106
rect 1386 -2118 1392 -2112
rect 1386 -2124 1392 -2118
rect 1386 -2130 1392 -2124
rect 1386 -2136 1392 -2130
rect 1386 -2142 1392 -2136
rect 1386 -2148 1392 -2142
rect 1386 -2154 1392 -2148
rect 1386 -2160 1392 -2154
rect 1386 -2166 1392 -2160
rect 1386 -2172 1392 -2166
rect 1386 -2178 1392 -2172
rect 1386 -2184 1392 -2178
rect 1386 -2190 1392 -2184
rect 1386 -2196 1392 -2190
rect 1386 -2202 1392 -2196
rect 1386 -2208 1392 -2202
rect 1386 -2214 1392 -2208
rect 1386 -2220 1392 -2214
rect 1386 -2226 1392 -2220
rect 1386 -2232 1392 -2226
rect 1386 -2238 1392 -2232
rect 1386 -2244 1392 -2238
rect 1386 -2250 1392 -2244
rect 1386 -2256 1392 -2250
rect 1386 -2262 1392 -2256
rect 1386 -2268 1392 -2262
rect 1386 -2274 1392 -2268
rect 1386 -2280 1392 -2274
rect 1386 -2286 1392 -2280
rect 1386 -2292 1392 -2286
rect 1386 -2298 1392 -2292
rect 1386 -2304 1392 -2298
rect 1386 -2310 1392 -2304
rect 1386 -2316 1392 -2310
rect 1386 -2322 1392 -2316
rect 1386 -2328 1392 -2322
rect 1386 -2334 1392 -2328
rect 1386 -2340 1392 -2334
rect 1386 -2418 1392 -2412
rect 1386 -2424 1392 -2418
rect 1386 -2430 1392 -2424
rect 1386 -2436 1392 -2430
rect 1386 -2442 1392 -2436
rect 1386 -2448 1392 -2442
rect 1386 -2454 1392 -2448
rect 1386 -2460 1392 -2454
rect 1386 -2466 1392 -2460
rect 1386 -2472 1392 -2466
rect 1386 -2478 1392 -2472
rect 1386 -2484 1392 -2478
rect 1386 -2490 1392 -2484
rect 1386 -2496 1392 -2490
rect 1386 -2502 1392 -2496
rect 1386 -2508 1392 -2502
rect 1386 -2514 1392 -2508
rect 1386 -2520 1392 -2514
rect 1386 -2526 1392 -2520
rect 1386 -2532 1392 -2526
rect 1386 -2538 1392 -2532
rect 1386 -2544 1392 -2538
rect 1386 -2550 1392 -2544
rect 1386 -2556 1392 -2550
rect 1386 -2562 1392 -2556
rect 1386 -2568 1392 -2562
rect 1386 -2574 1392 -2568
rect 1386 -2580 1392 -2574
rect 1386 -2586 1392 -2580
rect 1386 -2592 1392 -2586
rect 1386 -2598 1392 -2592
rect 1386 -2604 1392 -2598
rect 1386 -2610 1392 -2604
rect 1386 -2616 1392 -2610
rect 1386 -2622 1392 -2616
rect 1386 -2628 1392 -2622
rect 1386 -2634 1392 -2628
rect 1386 -2640 1392 -2634
rect 1386 -2646 1392 -2640
rect 1386 -2652 1392 -2646
rect 1386 -2658 1392 -2652
rect 1386 -2664 1392 -2658
rect 1386 -2670 1392 -2664
rect 1386 -2676 1392 -2670
rect 1386 -2682 1392 -2676
rect 1386 -2688 1392 -2682
rect 1386 -2694 1392 -2688
rect 1386 -2700 1392 -2694
rect 1386 -2706 1392 -2700
rect 1386 -2712 1392 -2706
rect 1386 -2718 1392 -2712
rect 1386 -2724 1392 -2718
rect 1386 -2730 1392 -2724
rect 1386 -2736 1392 -2730
rect 1386 -2742 1392 -2736
rect 1386 -2748 1392 -2742
rect 1386 -2754 1392 -2748
rect 1386 -2760 1392 -2754
rect 1386 -2766 1392 -2760
rect 1386 -2772 1392 -2766
rect 1386 -2778 1392 -2772
rect 1386 -2784 1392 -2778
rect 1386 -2790 1392 -2784
rect 1386 -2796 1392 -2790
rect 1386 -2802 1392 -2796
rect 1386 -2808 1392 -2802
rect 1386 -2814 1392 -2808
rect 1386 -2820 1392 -2814
rect 1386 -2826 1392 -2820
rect 1386 -2832 1392 -2826
rect 1386 -2838 1392 -2832
rect 1386 -2844 1392 -2838
rect 1386 -2850 1392 -2844
rect 1386 -2856 1392 -2850
rect 1386 -2862 1392 -2856
rect 1386 -2868 1392 -2862
rect 1386 -2874 1392 -2868
rect 1386 -2880 1392 -2874
rect 1386 -2886 1392 -2880
rect 1386 -2970 1392 -2964
rect 1386 -2976 1392 -2970
rect 1386 -2982 1392 -2976
rect 1386 -2988 1392 -2982
rect 1386 -2994 1392 -2988
rect 1386 -3000 1392 -2994
rect 1386 -3006 1392 -3000
rect 1386 -3012 1392 -3006
rect 1386 -3018 1392 -3012
rect 1386 -3024 1392 -3018
rect 1386 -3030 1392 -3024
rect 1386 -3036 1392 -3030
rect 1386 -3042 1392 -3036
rect 1386 -3048 1392 -3042
rect 1386 -3054 1392 -3048
rect 1386 -3060 1392 -3054
rect 1386 -3066 1392 -3060
rect 1386 -3072 1392 -3066
rect 1386 -3078 1392 -3072
rect 1386 -3084 1392 -3078
rect 1386 -3090 1392 -3084
rect 1386 -3096 1392 -3090
rect 1386 -3102 1392 -3096
rect 1386 -3108 1392 -3102
rect 1386 -3114 1392 -3108
rect 1386 -3120 1392 -3114
rect 1386 -3126 1392 -3120
rect 1386 -3132 1392 -3126
rect 1386 -3138 1392 -3132
rect 1386 -3144 1392 -3138
rect 1386 -3150 1392 -3144
rect 1386 -3156 1392 -3150
rect 1386 -3162 1392 -3156
rect 1386 -3168 1392 -3162
rect 1386 -3174 1392 -3168
rect 1386 -3180 1392 -3174
rect 1386 -3186 1392 -3180
rect 1386 -3192 1392 -3186
rect 1386 -3198 1392 -3192
rect 1386 -3204 1392 -3198
rect 1386 -3210 1392 -3204
rect 1386 -3216 1392 -3210
rect 1386 -3222 1392 -3216
rect 1386 -3228 1392 -3222
rect 1386 -3234 1392 -3228
rect 1386 -3306 1392 -3300
rect 1386 -3312 1392 -3306
rect 1386 -3318 1392 -3312
rect 1386 -3324 1392 -3318
rect 1386 -3330 1392 -3324
rect 1386 -3336 1392 -3330
rect 1386 -3342 1392 -3336
rect 1386 -3348 1392 -3342
rect 1386 -3354 1392 -3348
rect 1386 -3360 1392 -3354
rect 1386 -3366 1392 -3360
rect 1386 -3372 1392 -3366
rect 1386 -3378 1392 -3372
rect 1386 -3384 1392 -3378
rect 1386 -3390 1392 -3384
rect 1386 -3396 1392 -3390
rect 1386 -3402 1392 -3396
rect 1386 -3408 1392 -3402
rect 1386 -3414 1392 -3408
rect 1386 -3420 1392 -3414
rect 1386 -3426 1392 -3420
rect 1386 -3432 1392 -3426
rect 1386 -3438 1392 -3432
rect 1386 -3444 1392 -3438
rect 1386 -3450 1392 -3444
rect 1386 -3456 1392 -3450
rect 1386 -3462 1392 -3456
rect 1386 -3468 1392 -3462
rect 1386 -3474 1392 -3468
rect 1386 -3480 1392 -3474
rect 1386 -3486 1392 -3480
rect 1386 -3492 1392 -3486
rect 1386 -3498 1392 -3492
rect 1386 -3504 1392 -3498
rect 1386 -3510 1392 -3504
rect 1392 -1116 1398 -1110
rect 1392 -1122 1398 -1116
rect 1392 -1128 1398 -1122
rect 1392 -1134 1398 -1128
rect 1392 -1140 1398 -1134
rect 1392 -1146 1398 -1140
rect 1392 -1152 1398 -1146
rect 1392 -1158 1398 -1152
rect 1392 -1164 1398 -1158
rect 1392 -1170 1398 -1164
rect 1392 -1176 1398 -1170
rect 1392 -1182 1398 -1176
rect 1392 -1188 1398 -1182
rect 1392 -1194 1398 -1188
rect 1392 -1200 1398 -1194
rect 1392 -1206 1398 -1200
rect 1392 -1212 1398 -1206
rect 1392 -1218 1398 -1212
rect 1392 -1224 1398 -1218
rect 1392 -1230 1398 -1224
rect 1392 -1236 1398 -1230
rect 1392 -1242 1398 -1236
rect 1392 -1248 1398 -1242
rect 1392 -1254 1398 -1248
rect 1392 -1260 1398 -1254
rect 1392 -1380 1398 -1374
rect 1392 -1386 1398 -1380
rect 1392 -1392 1398 -1386
rect 1392 -1398 1398 -1392
rect 1392 -1404 1398 -1398
rect 1392 -1410 1398 -1404
rect 1392 -1416 1398 -1410
rect 1392 -1422 1398 -1416
rect 1392 -1428 1398 -1422
rect 1392 -1434 1398 -1428
rect 1392 -1440 1398 -1434
rect 1392 -1446 1398 -1440
rect 1392 -1452 1398 -1446
rect 1392 -1458 1398 -1452
rect 1392 -1464 1398 -1458
rect 1392 -1470 1398 -1464
rect 1392 -1476 1398 -1470
rect 1392 -1482 1398 -1476
rect 1392 -1488 1398 -1482
rect 1392 -1494 1398 -1488
rect 1392 -1500 1398 -1494
rect 1392 -1506 1398 -1500
rect 1392 -1512 1398 -1506
rect 1392 -1518 1398 -1512
rect 1392 -1524 1398 -1518
rect 1392 -1530 1398 -1524
rect 1392 -1536 1398 -1530
rect 1392 -1542 1398 -1536
rect 1392 -1548 1398 -1542
rect 1392 -1554 1398 -1548
rect 1392 -1560 1398 -1554
rect 1392 -1566 1398 -1560
rect 1392 -1572 1398 -1566
rect 1392 -1578 1398 -1572
rect 1392 -1584 1398 -1578
rect 1392 -1590 1398 -1584
rect 1392 -1596 1398 -1590
rect 1392 -1602 1398 -1596
rect 1392 -1608 1398 -1602
rect 1392 -1614 1398 -1608
rect 1392 -1620 1398 -1614
rect 1392 -1626 1398 -1620
rect 1392 -1632 1398 -1626
rect 1392 -1638 1398 -1632
rect 1392 -1644 1398 -1638
rect 1392 -1650 1398 -1644
rect 1392 -1656 1398 -1650
rect 1392 -1662 1398 -1656
rect 1392 -1668 1398 -1662
rect 1392 -1674 1398 -1668
rect 1392 -1680 1398 -1674
rect 1392 -1686 1398 -1680
rect 1392 -1692 1398 -1686
rect 1392 -1698 1398 -1692
rect 1392 -1704 1398 -1698
rect 1392 -1710 1398 -1704
rect 1392 -1716 1398 -1710
rect 1392 -1722 1398 -1716
rect 1392 -1728 1398 -1722
rect 1392 -1734 1398 -1728
rect 1392 -1740 1398 -1734
rect 1392 -1746 1398 -1740
rect 1392 -1752 1398 -1746
rect 1392 -1758 1398 -1752
rect 1392 -1764 1398 -1758
rect 1392 -1770 1398 -1764
rect 1392 -1776 1398 -1770
rect 1392 -1782 1398 -1776
rect 1392 -1788 1398 -1782
rect 1392 -1794 1398 -1788
rect 1392 -1800 1398 -1794
rect 1392 -1806 1398 -1800
rect 1392 -1812 1398 -1806
rect 1392 -1818 1398 -1812
rect 1392 -1824 1398 -1818
rect 1392 -1830 1398 -1824
rect 1392 -1836 1398 -1830
rect 1392 -1842 1398 -1836
rect 1392 -1848 1398 -1842
rect 1392 -1854 1398 -1848
rect 1392 -1860 1398 -1854
rect 1392 -1866 1398 -1860
rect 1392 -1872 1398 -1866
rect 1392 -1878 1398 -1872
rect 1392 -1884 1398 -1878
rect 1392 -1890 1398 -1884
rect 1392 -1896 1398 -1890
rect 1392 -1902 1398 -1896
rect 1392 -1908 1398 -1902
rect 1392 -1914 1398 -1908
rect 1392 -1920 1398 -1914
rect 1392 -1926 1398 -1920
rect 1392 -1932 1398 -1926
rect 1392 -1938 1398 -1932
rect 1392 -1944 1398 -1938
rect 1392 -1950 1398 -1944
rect 1392 -1956 1398 -1950
rect 1392 -1962 1398 -1956
rect 1392 -1968 1398 -1962
rect 1392 -1974 1398 -1968
rect 1392 -1980 1398 -1974
rect 1392 -1986 1398 -1980
rect 1392 -1992 1398 -1986
rect 1392 -1998 1398 -1992
rect 1392 -2004 1398 -1998
rect 1392 -2010 1398 -2004
rect 1392 -2016 1398 -2010
rect 1392 -2022 1398 -2016
rect 1392 -2028 1398 -2022
rect 1392 -2034 1398 -2028
rect 1392 -2040 1398 -2034
rect 1392 -2046 1398 -2040
rect 1392 -2052 1398 -2046
rect 1392 -2058 1398 -2052
rect 1392 -2064 1398 -2058
rect 1392 -2070 1398 -2064
rect 1392 -2076 1398 -2070
rect 1392 -2082 1398 -2076
rect 1392 -2088 1398 -2082
rect 1392 -2094 1398 -2088
rect 1392 -2100 1398 -2094
rect 1392 -2106 1398 -2100
rect 1392 -2112 1398 -2106
rect 1392 -2118 1398 -2112
rect 1392 -2124 1398 -2118
rect 1392 -2130 1398 -2124
rect 1392 -2136 1398 -2130
rect 1392 -2142 1398 -2136
rect 1392 -2148 1398 -2142
rect 1392 -2154 1398 -2148
rect 1392 -2160 1398 -2154
rect 1392 -2166 1398 -2160
rect 1392 -2172 1398 -2166
rect 1392 -2178 1398 -2172
rect 1392 -2184 1398 -2178
rect 1392 -2190 1398 -2184
rect 1392 -2196 1398 -2190
rect 1392 -2202 1398 -2196
rect 1392 -2208 1398 -2202
rect 1392 -2214 1398 -2208
rect 1392 -2220 1398 -2214
rect 1392 -2226 1398 -2220
rect 1392 -2232 1398 -2226
rect 1392 -2238 1398 -2232
rect 1392 -2244 1398 -2238
rect 1392 -2250 1398 -2244
rect 1392 -2256 1398 -2250
rect 1392 -2262 1398 -2256
rect 1392 -2268 1398 -2262
rect 1392 -2274 1398 -2268
rect 1392 -2280 1398 -2274
rect 1392 -2286 1398 -2280
rect 1392 -2292 1398 -2286
rect 1392 -2298 1398 -2292
rect 1392 -2304 1398 -2298
rect 1392 -2310 1398 -2304
rect 1392 -2316 1398 -2310
rect 1392 -2322 1398 -2316
rect 1392 -2328 1398 -2322
rect 1392 -2334 1398 -2328
rect 1392 -2412 1398 -2406
rect 1392 -2418 1398 -2412
rect 1392 -2424 1398 -2418
rect 1392 -2430 1398 -2424
rect 1392 -2436 1398 -2430
rect 1392 -2442 1398 -2436
rect 1392 -2448 1398 -2442
rect 1392 -2454 1398 -2448
rect 1392 -2460 1398 -2454
rect 1392 -2466 1398 -2460
rect 1392 -2472 1398 -2466
rect 1392 -2478 1398 -2472
rect 1392 -2484 1398 -2478
rect 1392 -2490 1398 -2484
rect 1392 -2496 1398 -2490
rect 1392 -2502 1398 -2496
rect 1392 -2508 1398 -2502
rect 1392 -2514 1398 -2508
rect 1392 -2520 1398 -2514
rect 1392 -2526 1398 -2520
rect 1392 -2532 1398 -2526
rect 1392 -2538 1398 -2532
rect 1392 -2544 1398 -2538
rect 1392 -2550 1398 -2544
rect 1392 -2556 1398 -2550
rect 1392 -2562 1398 -2556
rect 1392 -2568 1398 -2562
rect 1392 -2574 1398 -2568
rect 1392 -2580 1398 -2574
rect 1392 -2586 1398 -2580
rect 1392 -2592 1398 -2586
rect 1392 -2598 1398 -2592
rect 1392 -2604 1398 -2598
rect 1392 -2610 1398 -2604
rect 1392 -2616 1398 -2610
rect 1392 -2622 1398 -2616
rect 1392 -2628 1398 -2622
rect 1392 -2634 1398 -2628
rect 1392 -2640 1398 -2634
rect 1392 -2646 1398 -2640
rect 1392 -2652 1398 -2646
rect 1392 -2658 1398 -2652
rect 1392 -2664 1398 -2658
rect 1392 -2670 1398 -2664
rect 1392 -2676 1398 -2670
rect 1392 -2682 1398 -2676
rect 1392 -2688 1398 -2682
rect 1392 -2694 1398 -2688
rect 1392 -2700 1398 -2694
rect 1392 -2706 1398 -2700
rect 1392 -2712 1398 -2706
rect 1392 -2718 1398 -2712
rect 1392 -2724 1398 -2718
rect 1392 -2730 1398 -2724
rect 1392 -2736 1398 -2730
rect 1392 -2742 1398 -2736
rect 1392 -2748 1398 -2742
rect 1392 -2754 1398 -2748
rect 1392 -2760 1398 -2754
rect 1392 -2766 1398 -2760
rect 1392 -2772 1398 -2766
rect 1392 -2778 1398 -2772
rect 1392 -2784 1398 -2778
rect 1392 -2790 1398 -2784
rect 1392 -2796 1398 -2790
rect 1392 -2802 1398 -2796
rect 1392 -2808 1398 -2802
rect 1392 -2814 1398 -2808
rect 1392 -2820 1398 -2814
rect 1392 -2826 1398 -2820
rect 1392 -2832 1398 -2826
rect 1392 -2838 1398 -2832
rect 1392 -2844 1398 -2838
rect 1392 -2850 1398 -2844
rect 1392 -2856 1398 -2850
rect 1392 -2862 1398 -2856
rect 1392 -2868 1398 -2862
rect 1392 -2874 1398 -2868
rect 1392 -2880 1398 -2874
rect 1392 -2964 1398 -2958
rect 1392 -2970 1398 -2964
rect 1392 -2976 1398 -2970
rect 1392 -2982 1398 -2976
rect 1392 -2988 1398 -2982
rect 1392 -2994 1398 -2988
rect 1392 -3000 1398 -2994
rect 1392 -3006 1398 -3000
rect 1392 -3012 1398 -3006
rect 1392 -3018 1398 -3012
rect 1392 -3024 1398 -3018
rect 1392 -3030 1398 -3024
rect 1392 -3036 1398 -3030
rect 1392 -3042 1398 -3036
rect 1392 -3048 1398 -3042
rect 1392 -3054 1398 -3048
rect 1392 -3060 1398 -3054
rect 1392 -3066 1398 -3060
rect 1392 -3072 1398 -3066
rect 1392 -3078 1398 -3072
rect 1392 -3084 1398 -3078
rect 1392 -3090 1398 -3084
rect 1392 -3096 1398 -3090
rect 1392 -3102 1398 -3096
rect 1392 -3108 1398 -3102
rect 1392 -3114 1398 -3108
rect 1392 -3120 1398 -3114
rect 1392 -3126 1398 -3120
rect 1392 -3132 1398 -3126
rect 1392 -3138 1398 -3132
rect 1392 -3144 1398 -3138
rect 1392 -3150 1398 -3144
rect 1392 -3156 1398 -3150
rect 1392 -3162 1398 -3156
rect 1392 -3168 1398 -3162
rect 1392 -3174 1398 -3168
rect 1392 -3180 1398 -3174
rect 1392 -3186 1398 -3180
rect 1392 -3192 1398 -3186
rect 1392 -3198 1398 -3192
rect 1392 -3204 1398 -3198
rect 1392 -3210 1398 -3204
rect 1392 -3216 1398 -3210
rect 1392 -3222 1398 -3216
rect 1392 -3228 1398 -3222
rect 1392 -3234 1398 -3228
rect 1392 -3306 1398 -3300
rect 1392 -3312 1398 -3306
rect 1392 -3318 1398 -3312
rect 1392 -3324 1398 -3318
rect 1392 -3330 1398 -3324
rect 1392 -3336 1398 -3330
rect 1392 -3342 1398 -3336
rect 1392 -3348 1398 -3342
rect 1392 -3354 1398 -3348
rect 1392 -3360 1398 -3354
rect 1392 -3366 1398 -3360
rect 1392 -3372 1398 -3366
rect 1392 -3378 1398 -3372
rect 1392 -3384 1398 -3378
rect 1392 -3390 1398 -3384
rect 1392 -3396 1398 -3390
rect 1392 -3402 1398 -3396
rect 1392 -3408 1398 -3402
rect 1392 -3414 1398 -3408
rect 1392 -3420 1398 -3414
rect 1392 -3426 1398 -3420
rect 1392 -3432 1398 -3426
rect 1392 -3438 1398 -3432
rect 1392 -3444 1398 -3438
rect 1392 -3450 1398 -3444
rect 1392 -3456 1398 -3450
rect 1392 -3462 1398 -3456
rect 1392 -3468 1398 -3462
rect 1392 -3474 1398 -3468
rect 1392 -3480 1398 -3474
rect 1392 -3486 1398 -3480
rect 1392 -3492 1398 -3486
rect 1392 -3498 1398 -3492
rect 1392 -3504 1398 -3498
rect 1392 -3510 1398 -3504
rect 1398 -1116 1404 -1110
rect 1398 -1122 1404 -1116
rect 1398 -1128 1404 -1122
rect 1398 -1134 1404 -1128
rect 1398 -1140 1404 -1134
rect 1398 -1146 1404 -1140
rect 1398 -1152 1404 -1146
rect 1398 -1158 1404 -1152
rect 1398 -1164 1404 -1158
rect 1398 -1170 1404 -1164
rect 1398 -1176 1404 -1170
rect 1398 -1182 1404 -1176
rect 1398 -1188 1404 -1182
rect 1398 -1194 1404 -1188
rect 1398 -1200 1404 -1194
rect 1398 -1206 1404 -1200
rect 1398 -1212 1404 -1206
rect 1398 -1218 1404 -1212
rect 1398 -1224 1404 -1218
rect 1398 -1230 1404 -1224
rect 1398 -1236 1404 -1230
rect 1398 -1242 1404 -1236
rect 1398 -1248 1404 -1242
rect 1398 -1368 1404 -1362
rect 1398 -1374 1404 -1368
rect 1398 -1380 1404 -1374
rect 1398 -1386 1404 -1380
rect 1398 -1392 1404 -1386
rect 1398 -1398 1404 -1392
rect 1398 -1404 1404 -1398
rect 1398 -1410 1404 -1404
rect 1398 -1416 1404 -1410
rect 1398 -1422 1404 -1416
rect 1398 -1428 1404 -1422
rect 1398 -1434 1404 -1428
rect 1398 -1440 1404 -1434
rect 1398 -1446 1404 -1440
rect 1398 -1452 1404 -1446
rect 1398 -1458 1404 -1452
rect 1398 -1464 1404 -1458
rect 1398 -1470 1404 -1464
rect 1398 -1476 1404 -1470
rect 1398 -1482 1404 -1476
rect 1398 -1488 1404 -1482
rect 1398 -1494 1404 -1488
rect 1398 -1500 1404 -1494
rect 1398 -1506 1404 -1500
rect 1398 -1512 1404 -1506
rect 1398 -1518 1404 -1512
rect 1398 -1524 1404 -1518
rect 1398 -1530 1404 -1524
rect 1398 -1536 1404 -1530
rect 1398 -1542 1404 -1536
rect 1398 -1548 1404 -1542
rect 1398 -1554 1404 -1548
rect 1398 -1560 1404 -1554
rect 1398 -1566 1404 -1560
rect 1398 -1572 1404 -1566
rect 1398 -1578 1404 -1572
rect 1398 -1584 1404 -1578
rect 1398 -1590 1404 -1584
rect 1398 -1596 1404 -1590
rect 1398 -1602 1404 -1596
rect 1398 -1608 1404 -1602
rect 1398 -1614 1404 -1608
rect 1398 -1620 1404 -1614
rect 1398 -1626 1404 -1620
rect 1398 -1632 1404 -1626
rect 1398 -1638 1404 -1632
rect 1398 -1644 1404 -1638
rect 1398 -1650 1404 -1644
rect 1398 -1656 1404 -1650
rect 1398 -1662 1404 -1656
rect 1398 -1668 1404 -1662
rect 1398 -1674 1404 -1668
rect 1398 -1680 1404 -1674
rect 1398 -1686 1404 -1680
rect 1398 -1692 1404 -1686
rect 1398 -1698 1404 -1692
rect 1398 -1704 1404 -1698
rect 1398 -1710 1404 -1704
rect 1398 -1716 1404 -1710
rect 1398 -1722 1404 -1716
rect 1398 -1728 1404 -1722
rect 1398 -1734 1404 -1728
rect 1398 -1740 1404 -1734
rect 1398 -1746 1404 -1740
rect 1398 -1752 1404 -1746
rect 1398 -1758 1404 -1752
rect 1398 -1764 1404 -1758
rect 1398 -1770 1404 -1764
rect 1398 -1776 1404 -1770
rect 1398 -1782 1404 -1776
rect 1398 -1788 1404 -1782
rect 1398 -1794 1404 -1788
rect 1398 -1800 1404 -1794
rect 1398 -1806 1404 -1800
rect 1398 -1812 1404 -1806
rect 1398 -1818 1404 -1812
rect 1398 -1824 1404 -1818
rect 1398 -1830 1404 -1824
rect 1398 -1836 1404 -1830
rect 1398 -1842 1404 -1836
rect 1398 -1848 1404 -1842
rect 1398 -1854 1404 -1848
rect 1398 -1860 1404 -1854
rect 1398 -1866 1404 -1860
rect 1398 -1872 1404 -1866
rect 1398 -1878 1404 -1872
rect 1398 -1884 1404 -1878
rect 1398 -1890 1404 -1884
rect 1398 -1896 1404 -1890
rect 1398 -1902 1404 -1896
rect 1398 -1908 1404 -1902
rect 1398 -1914 1404 -1908
rect 1398 -1920 1404 -1914
rect 1398 -1926 1404 -1920
rect 1398 -1932 1404 -1926
rect 1398 -1938 1404 -1932
rect 1398 -1944 1404 -1938
rect 1398 -1950 1404 -1944
rect 1398 -1956 1404 -1950
rect 1398 -1962 1404 -1956
rect 1398 -1968 1404 -1962
rect 1398 -1974 1404 -1968
rect 1398 -1980 1404 -1974
rect 1398 -1986 1404 -1980
rect 1398 -1992 1404 -1986
rect 1398 -1998 1404 -1992
rect 1398 -2004 1404 -1998
rect 1398 -2010 1404 -2004
rect 1398 -2016 1404 -2010
rect 1398 -2022 1404 -2016
rect 1398 -2028 1404 -2022
rect 1398 -2034 1404 -2028
rect 1398 -2040 1404 -2034
rect 1398 -2046 1404 -2040
rect 1398 -2052 1404 -2046
rect 1398 -2058 1404 -2052
rect 1398 -2064 1404 -2058
rect 1398 -2070 1404 -2064
rect 1398 -2076 1404 -2070
rect 1398 -2082 1404 -2076
rect 1398 -2088 1404 -2082
rect 1398 -2094 1404 -2088
rect 1398 -2100 1404 -2094
rect 1398 -2106 1404 -2100
rect 1398 -2112 1404 -2106
rect 1398 -2118 1404 -2112
rect 1398 -2124 1404 -2118
rect 1398 -2130 1404 -2124
rect 1398 -2136 1404 -2130
rect 1398 -2142 1404 -2136
rect 1398 -2148 1404 -2142
rect 1398 -2154 1404 -2148
rect 1398 -2160 1404 -2154
rect 1398 -2166 1404 -2160
rect 1398 -2172 1404 -2166
rect 1398 -2178 1404 -2172
rect 1398 -2184 1404 -2178
rect 1398 -2190 1404 -2184
rect 1398 -2196 1404 -2190
rect 1398 -2202 1404 -2196
rect 1398 -2208 1404 -2202
rect 1398 -2214 1404 -2208
rect 1398 -2220 1404 -2214
rect 1398 -2226 1404 -2220
rect 1398 -2232 1404 -2226
rect 1398 -2238 1404 -2232
rect 1398 -2244 1404 -2238
rect 1398 -2250 1404 -2244
rect 1398 -2256 1404 -2250
rect 1398 -2262 1404 -2256
rect 1398 -2268 1404 -2262
rect 1398 -2274 1404 -2268
rect 1398 -2280 1404 -2274
rect 1398 -2286 1404 -2280
rect 1398 -2292 1404 -2286
rect 1398 -2298 1404 -2292
rect 1398 -2304 1404 -2298
rect 1398 -2310 1404 -2304
rect 1398 -2316 1404 -2310
rect 1398 -2322 1404 -2316
rect 1398 -2400 1404 -2394
rect 1398 -2406 1404 -2400
rect 1398 -2412 1404 -2406
rect 1398 -2418 1404 -2412
rect 1398 -2424 1404 -2418
rect 1398 -2430 1404 -2424
rect 1398 -2436 1404 -2430
rect 1398 -2442 1404 -2436
rect 1398 -2448 1404 -2442
rect 1398 -2454 1404 -2448
rect 1398 -2460 1404 -2454
rect 1398 -2466 1404 -2460
rect 1398 -2472 1404 -2466
rect 1398 -2478 1404 -2472
rect 1398 -2484 1404 -2478
rect 1398 -2490 1404 -2484
rect 1398 -2496 1404 -2490
rect 1398 -2502 1404 -2496
rect 1398 -2508 1404 -2502
rect 1398 -2514 1404 -2508
rect 1398 -2520 1404 -2514
rect 1398 -2526 1404 -2520
rect 1398 -2532 1404 -2526
rect 1398 -2538 1404 -2532
rect 1398 -2544 1404 -2538
rect 1398 -2550 1404 -2544
rect 1398 -2556 1404 -2550
rect 1398 -2562 1404 -2556
rect 1398 -2568 1404 -2562
rect 1398 -2574 1404 -2568
rect 1398 -2580 1404 -2574
rect 1398 -2586 1404 -2580
rect 1398 -2592 1404 -2586
rect 1398 -2598 1404 -2592
rect 1398 -2604 1404 -2598
rect 1398 -2610 1404 -2604
rect 1398 -2616 1404 -2610
rect 1398 -2622 1404 -2616
rect 1398 -2628 1404 -2622
rect 1398 -2634 1404 -2628
rect 1398 -2640 1404 -2634
rect 1398 -2646 1404 -2640
rect 1398 -2652 1404 -2646
rect 1398 -2658 1404 -2652
rect 1398 -2664 1404 -2658
rect 1398 -2670 1404 -2664
rect 1398 -2676 1404 -2670
rect 1398 -2682 1404 -2676
rect 1398 -2688 1404 -2682
rect 1398 -2694 1404 -2688
rect 1398 -2700 1404 -2694
rect 1398 -2706 1404 -2700
rect 1398 -2712 1404 -2706
rect 1398 -2718 1404 -2712
rect 1398 -2724 1404 -2718
rect 1398 -2730 1404 -2724
rect 1398 -2736 1404 -2730
rect 1398 -2742 1404 -2736
rect 1398 -2748 1404 -2742
rect 1398 -2754 1404 -2748
rect 1398 -2760 1404 -2754
rect 1398 -2766 1404 -2760
rect 1398 -2772 1404 -2766
rect 1398 -2778 1404 -2772
rect 1398 -2784 1404 -2778
rect 1398 -2790 1404 -2784
rect 1398 -2796 1404 -2790
rect 1398 -2802 1404 -2796
rect 1398 -2808 1404 -2802
rect 1398 -2814 1404 -2808
rect 1398 -2820 1404 -2814
rect 1398 -2826 1404 -2820
rect 1398 -2832 1404 -2826
rect 1398 -2838 1404 -2832
rect 1398 -2844 1404 -2838
rect 1398 -2850 1404 -2844
rect 1398 -2856 1404 -2850
rect 1398 -2862 1404 -2856
rect 1398 -2868 1404 -2862
rect 1398 -2874 1404 -2868
rect 1398 -2964 1404 -2958
rect 1398 -2970 1404 -2964
rect 1398 -2976 1404 -2970
rect 1398 -2982 1404 -2976
rect 1398 -2988 1404 -2982
rect 1398 -2994 1404 -2988
rect 1398 -3000 1404 -2994
rect 1398 -3006 1404 -3000
rect 1398 -3012 1404 -3006
rect 1398 -3018 1404 -3012
rect 1398 -3024 1404 -3018
rect 1398 -3030 1404 -3024
rect 1398 -3036 1404 -3030
rect 1398 -3042 1404 -3036
rect 1398 -3048 1404 -3042
rect 1398 -3054 1404 -3048
rect 1398 -3060 1404 -3054
rect 1398 -3066 1404 -3060
rect 1398 -3072 1404 -3066
rect 1398 -3078 1404 -3072
rect 1398 -3084 1404 -3078
rect 1398 -3090 1404 -3084
rect 1398 -3096 1404 -3090
rect 1398 -3102 1404 -3096
rect 1398 -3108 1404 -3102
rect 1398 -3114 1404 -3108
rect 1398 -3120 1404 -3114
rect 1398 -3126 1404 -3120
rect 1398 -3132 1404 -3126
rect 1398 -3138 1404 -3132
rect 1398 -3144 1404 -3138
rect 1398 -3150 1404 -3144
rect 1398 -3156 1404 -3150
rect 1398 -3162 1404 -3156
rect 1398 -3168 1404 -3162
rect 1398 -3174 1404 -3168
rect 1398 -3180 1404 -3174
rect 1398 -3186 1404 -3180
rect 1398 -3192 1404 -3186
rect 1398 -3198 1404 -3192
rect 1398 -3204 1404 -3198
rect 1398 -3210 1404 -3204
rect 1398 -3216 1404 -3210
rect 1398 -3222 1404 -3216
rect 1398 -3228 1404 -3222
rect 1398 -3234 1404 -3228
rect 1398 -3306 1404 -3300
rect 1398 -3312 1404 -3306
rect 1398 -3318 1404 -3312
rect 1398 -3324 1404 -3318
rect 1398 -3330 1404 -3324
rect 1398 -3336 1404 -3330
rect 1398 -3342 1404 -3336
rect 1398 -3348 1404 -3342
rect 1398 -3354 1404 -3348
rect 1398 -3360 1404 -3354
rect 1398 -3366 1404 -3360
rect 1398 -3372 1404 -3366
rect 1398 -3378 1404 -3372
rect 1398 -3384 1404 -3378
rect 1398 -3390 1404 -3384
rect 1398 -3396 1404 -3390
rect 1398 -3402 1404 -3396
rect 1398 -3408 1404 -3402
rect 1398 -3414 1404 -3408
rect 1398 -3420 1404 -3414
rect 1398 -3426 1404 -3420
rect 1398 -3432 1404 -3426
rect 1398 -3438 1404 -3432
rect 1398 -3444 1404 -3438
rect 1398 -3450 1404 -3444
rect 1398 -3456 1404 -3450
rect 1398 -3462 1404 -3456
rect 1398 -3468 1404 -3462
rect 1398 -3474 1404 -3468
rect 1398 -3480 1404 -3474
rect 1398 -3486 1404 -3480
rect 1398 -3492 1404 -3486
rect 1398 -3498 1404 -3492
rect 1398 -3504 1404 -3498
rect 1398 -3510 1404 -3504
rect 1404 -1116 1410 -1110
rect 1404 -1122 1410 -1116
rect 1404 -1128 1410 -1122
rect 1404 -1134 1410 -1128
rect 1404 -1140 1410 -1134
rect 1404 -1146 1410 -1140
rect 1404 -1152 1410 -1146
rect 1404 -1158 1410 -1152
rect 1404 -1164 1410 -1158
rect 1404 -1170 1410 -1164
rect 1404 -1176 1410 -1170
rect 1404 -1182 1410 -1176
rect 1404 -1188 1410 -1182
rect 1404 -1194 1410 -1188
rect 1404 -1200 1410 -1194
rect 1404 -1206 1410 -1200
rect 1404 -1212 1410 -1206
rect 1404 -1218 1410 -1212
rect 1404 -1224 1410 -1218
rect 1404 -1230 1410 -1224
rect 1404 -1236 1410 -1230
rect 1404 -1242 1410 -1236
rect 1404 -1356 1410 -1350
rect 1404 -1362 1410 -1356
rect 1404 -1368 1410 -1362
rect 1404 -1374 1410 -1368
rect 1404 -1380 1410 -1374
rect 1404 -1386 1410 -1380
rect 1404 -1392 1410 -1386
rect 1404 -1398 1410 -1392
rect 1404 -1404 1410 -1398
rect 1404 -1410 1410 -1404
rect 1404 -1416 1410 -1410
rect 1404 -1422 1410 -1416
rect 1404 -1428 1410 -1422
rect 1404 -1434 1410 -1428
rect 1404 -1440 1410 -1434
rect 1404 -1446 1410 -1440
rect 1404 -1452 1410 -1446
rect 1404 -1458 1410 -1452
rect 1404 -1464 1410 -1458
rect 1404 -1470 1410 -1464
rect 1404 -1476 1410 -1470
rect 1404 -1482 1410 -1476
rect 1404 -1488 1410 -1482
rect 1404 -1494 1410 -1488
rect 1404 -1500 1410 -1494
rect 1404 -1506 1410 -1500
rect 1404 -1512 1410 -1506
rect 1404 -1518 1410 -1512
rect 1404 -1524 1410 -1518
rect 1404 -1530 1410 -1524
rect 1404 -1536 1410 -1530
rect 1404 -1542 1410 -1536
rect 1404 -1548 1410 -1542
rect 1404 -1554 1410 -1548
rect 1404 -1560 1410 -1554
rect 1404 -1566 1410 -1560
rect 1404 -1572 1410 -1566
rect 1404 -1578 1410 -1572
rect 1404 -1584 1410 -1578
rect 1404 -1590 1410 -1584
rect 1404 -1596 1410 -1590
rect 1404 -1602 1410 -1596
rect 1404 -1608 1410 -1602
rect 1404 -1614 1410 -1608
rect 1404 -1620 1410 -1614
rect 1404 -1626 1410 -1620
rect 1404 -1632 1410 -1626
rect 1404 -1638 1410 -1632
rect 1404 -1644 1410 -1638
rect 1404 -1650 1410 -1644
rect 1404 -1656 1410 -1650
rect 1404 -1662 1410 -1656
rect 1404 -1668 1410 -1662
rect 1404 -1674 1410 -1668
rect 1404 -1680 1410 -1674
rect 1404 -1686 1410 -1680
rect 1404 -1692 1410 -1686
rect 1404 -1698 1410 -1692
rect 1404 -1704 1410 -1698
rect 1404 -1710 1410 -1704
rect 1404 -1716 1410 -1710
rect 1404 -1722 1410 -1716
rect 1404 -1728 1410 -1722
rect 1404 -1734 1410 -1728
rect 1404 -1740 1410 -1734
rect 1404 -1746 1410 -1740
rect 1404 -1752 1410 -1746
rect 1404 -1758 1410 -1752
rect 1404 -1764 1410 -1758
rect 1404 -1770 1410 -1764
rect 1404 -1776 1410 -1770
rect 1404 -1782 1410 -1776
rect 1404 -1788 1410 -1782
rect 1404 -1794 1410 -1788
rect 1404 -1800 1410 -1794
rect 1404 -1806 1410 -1800
rect 1404 -1812 1410 -1806
rect 1404 -1818 1410 -1812
rect 1404 -1824 1410 -1818
rect 1404 -1830 1410 -1824
rect 1404 -1836 1410 -1830
rect 1404 -1842 1410 -1836
rect 1404 -1848 1410 -1842
rect 1404 -1854 1410 -1848
rect 1404 -1860 1410 -1854
rect 1404 -1866 1410 -1860
rect 1404 -1872 1410 -1866
rect 1404 -1878 1410 -1872
rect 1404 -1884 1410 -1878
rect 1404 -1890 1410 -1884
rect 1404 -1896 1410 -1890
rect 1404 -1902 1410 -1896
rect 1404 -1908 1410 -1902
rect 1404 -1914 1410 -1908
rect 1404 -1920 1410 -1914
rect 1404 -1926 1410 -1920
rect 1404 -1932 1410 -1926
rect 1404 -1938 1410 -1932
rect 1404 -1944 1410 -1938
rect 1404 -1950 1410 -1944
rect 1404 -1956 1410 -1950
rect 1404 -1962 1410 -1956
rect 1404 -1968 1410 -1962
rect 1404 -1974 1410 -1968
rect 1404 -1980 1410 -1974
rect 1404 -1986 1410 -1980
rect 1404 -1992 1410 -1986
rect 1404 -1998 1410 -1992
rect 1404 -2004 1410 -1998
rect 1404 -2010 1410 -2004
rect 1404 -2016 1410 -2010
rect 1404 -2022 1410 -2016
rect 1404 -2028 1410 -2022
rect 1404 -2034 1410 -2028
rect 1404 -2040 1410 -2034
rect 1404 -2046 1410 -2040
rect 1404 -2052 1410 -2046
rect 1404 -2058 1410 -2052
rect 1404 -2064 1410 -2058
rect 1404 -2070 1410 -2064
rect 1404 -2076 1410 -2070
rect 1404 -2082 1410 -2076
rect 1404 -2088 1410 -2082
rect 1404 -2094 1410 -2088
rect 1404 -2100 1410 -2094
rect 1404 -2106 1410 -2100
rect 1404 -2112 1410 -2106
rect 1404 -2118 1410 -2112
rect 1404 -2124 1410 -2118
rect 1404 -2130 1410 -2124
rect 1404 -2136 1410 -2130
rect 1404 -2142 1410 -2136
rect 1404 -2148 1410 -2142
rect 1404 -2154 1410 -2148
rect 1404 -2160 1410 -2154
rect 1404 -2166 1410 -2160
rect 1404 -2172 1410 -2166
rect 1404 -2178 1410 -2172
rect 1404 -2184 1410 -2178
rect 1404 -2190 1410 -2184
rect 1404 -2196 1410 -2190
rect 1404 -2202 1410 -2196
rect 1404 -2208 1410 -2202
rect 1404 -2214 1410 -2208
rect 1404 -2220 1410 -2214
rect 1404 -2226 1410 -2220
rect 1404 -2232 1410 -2226
rect 1404 -2238 1410 -2232
rect 1404 -2244 1410 -2238
rect 1404 -2250 1410 -2244
rect 1404 -2256 1410 -2250
rect 1404 -2262 1410 -2256
rect 1404 -2268 1410 -2262
rect 1404 -2274 1410 -2268
rect 1404 -2280 1410 -2274
rect 1404 -2286 1410 -2280
rect 1404 -2292 1410 -2286
rect 1404 -2298 1410 -2292
rect 1404 -2304 1410 -2298
rect 1404 -2310 1410 -2304
rect 1404 -2316 1410 -2310
rect 1404 -2394 1410 -2388
rect 1404 -2400 1410 -2394
rect 1404 -2406 1410 -2400
rect 1404 -2412 1410 -2406
rect 1404 -2418 1410 -2412
rect 1404 -2424 1410 -2418
rect 1404 -2430 1410 -2424
rect 1404 -2436 1410 -2430
rect 1404 -2442 1410 -2436
rect 1404 -2448 1410 -2442
rect 1404 -2454 1410 -2448
rect 1404 -2460 1410 -2454
rect 1404 -2466 1410 -2460
rect 1404 -2472 1410 -2466
rect 1404 -2478 1410 -2472
rect 1404 -2484 1410 -2478
rect 1404 -2490 1410 -2484
rect 1404 -2496 1410 -2490
rect 1404 -2502 1410 -2496
rect 1404 -2508 1410 -2502
rect 1404 -2514 1410 -2508
rect 1404 -2520 1410 -2514
rect 1404 -2526 1410 -2520
rect 1404 -2532 1410 -2526
rect 1404 -2538 1410 -2532
rect 1404 -2544 1410 -2538
rect 1404 -2550 1410 -2544
rect 1404 -2556 1410 -2550
rect 1404 -2562 1410 -2556
rect 1404 -2568 1410 -2562
rect 1404 -2574 1410 -2568
rect 1404 -2580 1410 -2574
rect 1404 -2586 1410 -2580
rect 1404 -2592 1410 -2586
rect 1404 -2598 1410 -2592
rect 1404 -2604 1410 -2598
rect 1404 -2610 1410 -2604
rect 1404 -2616 1410 -2610
rect 1404 -2622 1410 -2616
rect 1404 -2628 1410 -2622
rect 1404 -2634 1410 -2628
rect 1404 -2640 1410 -2634
rect 1404 -2646 1410 -2640
rect 1404 -2652 1410 -2646
rect 1404 -2658 1410 -2652
rect 1404 -2664 1410 -2658
rect 1404 -2670 1410 -2664
rect 1404 -2676 1410 -2670
rect 1404 -2682 1410 -2676
rect 1404 -2688 1410 -2682
rect 1404 -2694 1410 -2688
rect 1404 -2700 1410 -2694
rect 1404 -2706 1410 -2700
rect 1404 -2712 1410 -2706
rect 1404 -2718 1410 -2712
rect 1404 -2724 1410 -2718
rect 1404 -2730 1410 -2724
rect 1404 -2736 1410 -2730
rect 1404 -2742 1410 -2736
rect 1404 -2748 1410 -2742
rect 1404 -2754 1410 -2748
rect 1404 -2760 1410 -2754
rect 1404 -2766 1410 -2760
rect 1404 -2772 1410 -2766
rect 1404 -2778 1410 -2772
rect 1404 -2784 1410 -2778
rect 1404 -2790 1410 -2784
rect 1404 -2796 1410 -2790
rect 1404 -2802 1410 -2796
rect 1404 -2808 1410 -2802
rect 1404 -2814 1410 -2808
rect 1404 -2820 1410 -2814
rect 1404 -2826 1410 -2820
rect 1404 -2832 1410 -2826
rect 1404 -2838 1410 -2832
rect 1404 -2844 1410 -2838
rect 1404 -2850 1410 -2844
rect 1404 -2856 1410 -2850
rect 1404 -2862 1410 -2856
rect 1404 -2868 1410 -2862
rect 1404 -2874 1410 -2868
rect 1404 -2958 1410 -2952
rect 1404 -2964 1410 -2958
rect 1404 -2970 1410 -2964
rect 1404 -2976 1410 -2970
rect 1404 -2982 1410 -2976
rect 1404 -2988 1410 -2982
rect 1404 -2994 1410 -2988
rect 1404 -3000 1410 -2994
rect 1404 -3006 1410 -3000
rect 1404 -3012 1410 -3006
rect 1404 -3018 1410 -3012
rect 1404 -3024 1410 -3018
rect 1404 -3030 1410 -3024
rect 1404 -3036 1410 -3030
rect 1404 -3042 1410 -3036
rect 1404 -3048 1410 -3042
rect 1404 -3054 1410 -3048
rect 1404 -3060 1410 -3054
rect 1404 -3066 1410 -3060
rect 1404 -3072 1410 -3066
rect 1404 -3078 1410 -3072
rect 1404 -3084 1410 -3078
rect 1404 -3090 1410 -3084
rect 1404 -3096 1410 -3090
rect 1404 -3102 1410 -3096
rect 1404 -3108 1410 -3102
rect 1404 -3114 1410 -3108
rect 1404 -3120 1410 -3114
rect 1404 -3126 1410 -3120
rect 1404 -3132 1410 -3126
rect 1404 -3138 1410 -3132
rect 1404 -3144 1410 -3138
rect 1404 -3150 1410 -3144
rect 1404 -3156 1410 -3150
rect 1404 -3162 1410 -3156
rect 1404 -3168 1410 -3162
rect 1404 -3174 1410 -3168
rect 1404 -3180 1410 -3174
rect 1404 -3186 1410 -3180
rect 1404 -3192 1410 -3186
rect 1404 -3198 1410 -3192
rect 1404 -3204 1410 -3198
rect 1404 -3210 1410 -3204
rect 1404 -3216 1410 -3210
rect 1404 -3222 1410 -3216
rect 1404 -3228 1410 -3222
rect 1404 -3234 1410 -3228
rect 1404 -3306 1410 -3300
rect 1404 -3312 1410 -3306
rect 1404 -3318 1410 -3312
rect 1404 -3324 1410 -3318
rect 1404 -3330 1410 -3324
rect 1404 -3336 1410 -3330
rect 1404 -3342 1410 -3336
rect 1404 -3348 1410 -3342
rect 1404 -3354 1410 -3348
rect 1404 -3360 1410 -3354
rect 1404 -3366 1410 -3360
rect 1404 -3372 1410 -3366
rect 1404 -3378 1410 -3372
rect 1404 -3384 1410 -3378
rect 1404 -3390 1410 -3384
rect 1404 -3396 1410 -3390
rect 1404 -3402 1410 -3396
rect 1404 -3408 1410 -3402
rect 1404 -3414 1410 -3408
rect 1404 -3420 1410 -3414
rect 1404 -3426 1410 -3420
rect 1404 -3432 1410 -3426
rect 1404 -3438 1410 -3432
rect 1404 -3444 1410 -3438
rect 1404 -3450 1410 -3444
rect 1404 -3456 1410 -3450
rect 1404 -3462 1410 -3456
rect 1404 -3468 1410 -3462
rect 1404 -3474 1410 -3468
rect 1404 -3480 1410 -3474
rect 1404 -3486 1410 -3480
rect 1404 -3492 1410 -3486
rect 1404 -3498 1410 -3492
rect 1404 -3504 1410 -3498
rect 1404 -3510 1410 -3504
rect 1410 -1116 1416 -1110
rect 1410 -1122 1416 -1116
rect 1410 -1128 1416 -1122
rect 1410 -1134 1416 -1128
rect 1410 -1140 1416 -1134
rect 1410 -1146 1416 -1140
rect 1410 -1152 1416 -1146
rect 1410 -1158 1416 -1152
rect 1410 -1164 1416 -1158
rect 1410 -1170 1416 -1164
rect 1410 -1176 1416 -1170
rect 1410 -1182 1416 -1176
rect 1410 -1188 1416 -1182
rect 1410 -1194 1416 -1188
rect 1410 -1200 1416 -1194
rect 1410 -1206 1416 -1200
rect 1410 -1212 1416 -1206
rect 1410 -1218 1416 -1212
rect 1410 -1224 1416 -1218
rect 1410 -1230 1416 -1224
rect 1410 -1344 1416 -1338
rect 1410 -1350 1416 -1344
rect 1410 -1356 1416 -1350
rect 1410 -1362 1416 -1356
rect 1410 -1368 1416 -1362
rect 1410 -1374 1416 -1368
rect 1410 -1380 1416 -1374
rect 1410 -1386 1416 -1380
rect 1410 -1392 1416 -1386
rect 1410 -1398 1416 -1392
rect 1410 -1404 1416 -1398
rect 1410 -1410 1416 -1404
rect 1410 -1416 1416 -1410
rect 1410 -1422 1416 -1416
rect 1410 -1428 1416 -1422
rect 1410 -1434 1416 -1428
rect 1410 -1440 1416 -1434
rect 1410 -1446 1416 -1440
rect 1410 -1452 1416 -1446
rect 1410 -1458 1416 -1452
rect 1410 -1464 1416 -1458
rect 1410 -1470 1416 -1464
rect 1410 -1476 1416 -1470
rect 1410 -1482 1416 -1476
rect 1410 -1488 1416 -1482
rect 1410 -1494 1416 -1488
rect 1410 -1500 1416 -1494
rect 1410 -1506 1416 -1500
rect 1410 -1512 1416 -1506
rect 1410 -1518 1416 -1512
rect 1410 -1524 1416 -1518
rect 1410 -1530 1416 -1524
rect 1410 -1536 1416 -1530
rect 1410 -1542 1416 -1536
rect 1410 -1548 1416 -1542
rect 1410 -1554 1416 -1548
rect 1410 -1560 1416 -1554
rect 1410 -1566 1416 -1560
rect 1410 -1572 1416 -1566
rect 1410 -1578 1416 -1572
rect 1410 -1584 1416 -1578
rect 1410 -1590 1416 -1584
rect 1410 -1596 1416 -1590
rect 1410 -1602 1416 -1596
rect 1410 -1608 1416 -1602
rect 1410 -1614 1416 -1608
rect 1410 -1620 1416 -1614
rect 1410 -1626 1416 -1620
rect 1410 -1632 1416 -1626
rect 1410 -1638 1416 -1632
rect 1410 -1644 1416 -1638
rect 1410 -1650 1416 -1644
rect 1410 -1656 1416 -1650
rect 1410 -1662 1416 -1656
rect 1410 -1668 1416 -1662
rect 1410 -1674 1416 -1668
rect 1410 -1680 1416 -1674
rect 1410 -1686 1416 -1680
rect 1410 -1692 1416 -1686
rect 1410 -1698 1416 -1692
rect 1410 -1704 1416 -1698
rect 1410 -1710 1416 -1704
rect 1410 -1716 1416 -1710
rect 1410 -1722 1416 -1716
rect 1410 -1728 1416 -1722
rect 1410 -1734 1416 -1728
rect 1410 -1740 1416 -1734
rect 1410 -1746 1416 -1740
rect 1410 -1752 1416 -1746
rect 1410 -1758 1416 -1752
rect 1410 -1764 1416 -1758
rect 1410 -1770 1416 -1764
rect 1410 -1776 1416 -1770
rect 1410 -1782 1416 -1776
rect 1410 -1788 1416 -1782
rect 1410 -1794 1416 -1788
rect 1410 -1800 1416 -1794
rect 1410 -1806 1416 -1800
rect 1410 -1812 1416 -1806
rect 1410 -1818 1416 -1812
rect 1410 -1824 1416 -1818
rect 1410 -1830 1416 -1824
rect 1410 -1836 1416 -1830
rect 1410 -1842 1416 -1836
rect 1410 -1848 1416 -1842
rect 1410 -1854 1416 -1848
rect 1410 -1860 1416 -1854
rect 1410 -1866 1416 -1860
rect 1410 -1872 1416 -1866
rect 1410 -1878 1416 -1872
rect 1410 -1884 1416 -1878
rect 1410 -1890 1416 -1884
rect 1410 -1896 1416 -1890
rect 1410 -1902 1416 -1896
rect 1410 -1908 1416 -1902
rect 1410 -1914 1416 -1908
rect 1410 -1920 1416 -1914
rect 1410 -1926 1416 -1920
rect 1410 -1932 1416 -1926
rect 1410 -1938 1416 -1932
rect 1410 -1944 1416 -1938
rect 1410 -1950 1416 -1944
rect 1410 -1956 1416 -1950
rect 1410 -1962 1416 -1956
rect 1410 -1968 1416 -1962
rect 1410 -1974 1416 -1968
rect 1410 -1980 1416 -1974
rect 1410 -1986 1416 -1980
rect 1410 -1992 1416 -1986
rect 1410 -1998 1416 -1992
rect 1410 -2004 1416 -1998
rect 1410 -2010 1416 -2004
rect 1410 -2016 1416 -2010
rect 1410 -2022 1416 -2016
rect 1410 -2028 1416 -2022
rect 1410 -2034 1416 -2028
rect 1410 -2040 1416 -2034
rect 1410 -2046 1416 -2040
rect 1410 -2052 1416 -2046
rect 1410 -2058 1416 -2052
rect 1410 -2064 1416 -2058
rect 1410 -2070 1416 -2064
rect 1410 -2076 1416 -2070
rect 1410 -2082 1416 -2076
rect 1410 -2088 1416 -2082
rect 1410 -2094 1416 -2088
rect 1410 -2100 1416 -2094
rect 1410 -2106 1416 -2100
rect 1410 -2112 1416 -2106
rect 1410 -2118 1416 -2112
rect 1410 -2124 1416 -2118
rect 1410 -2130 1416 -2124
rect 1410 -2136 1416 -2130
rect 1410 -2142 1416 -2136
rect 1410 -2148 1416 -2142
rect 1410 -2154 1416 -2148
rect 1410 -2160 1416 -2154
rect 1410 -2166 1416 -2160
rect 1410 -2172 1416 -2166
rect 1410 -2178 1416 -2172
rect 1410 -2184 1416 -2178
rect 1410 -2190 1416 -2184
rect 1410 -2196 1416 -2190
rect 1410 -2202 1416 -2196
rect 1410 -2208 1416 -2202
rect 1410 -2214 1416 -2208
rect 1410 -2220 1416 -2214
rect 1410 -2226 1416 -2220
rect 1410 -2232 1416 -2226
rect 1410 -2238 1416 -2232
rect 1410 -2244 1416 -2238
rect 1410 -2250 1416 -2244
rect 1410 -2256 1416 -2250
rect 1410 -2262 1416 -2256
rect 1410 -2268 1416 -2262
rect 1410 -2274 1416 -2268
rect 1410 -2280 1416 -2274
rect 1410 -2286 1416 -2280
rect 1410 -2292 1416 -2286
rect 1410 -2298 1416 -2292
rect 1410 -2304 1416 -2298
rect 1410 -2310 1416 -2304
rect 1410 -2382 1416 -2376
rect 1410 -2388 1416 -2382
rect 1410 -2394 1416 -2388
rect 1410 -2400 1416 -2394
rect 1410 -2406 1416 -2400
rect 1410 -2412 1416 -2406
rect 1410 -2418 1416 -2412
rect 1410 -2424 1416 -2418
rect 1410 -2430 1416 -2424
rect 1410 -2436 1416 -2430
rect 1410 -2442 1416 -2436
rect 1410 -2448 1416 -2442
rect 1410 -2454 1416 -2448
rect 1410 -2460 1416 -2454
rect 1410 -2466 1416 -2460
rect 1410 -2472 1416 -2466
rect 1410 -2478 1416 -2472
rect 1410 -2484 1416 -2478
rect 1410 -2490 1416 -2484
rect 1410 -2496 1416 -2490
rect 1410 -2502 1416 -2496
rect 1410 -2508 1416 -2502
rect 1410 -2514 1416 -2508
rect 1410 -2520 1416 -2514
rect 1410 -2526 1416 -2520
rect 1410 -2532 1416 -2526
rect 1410 -2538 1416 -2532
rect 1410 -2544 1416 -2538
rect 1410 -2550 1416 -2544
rect 1410 -2556 1416 -2550
rect 1410 -2562 1416 -2556
rect 1410 -2568 1416 -2562
rect 1410 -2574 1416 -2568
rect 1410 -2580 1416 -2574
rect 1410 -2586 1416 -2580
rect 1410 -2592 1416 -2586
rect 1410 -2598 1416 -2592
rect 1410 -2604 1416 -2598
rect 1410 -2610 1416 -2604
rect 1410 -2616 1416 -2610
rect 1410 -2622 1416 -2616
rect 1410 -2628 1416 -2622
rect 1410 -2634 1416 -2628
rect 1410 -2640 1416 -2634
rect 1410 -2646 1416 -2640
rect 1410 -2652 1416 -2646
rect 1410 -2658 1416 -2652
rect 1410 -2664 1416 -2658
rect 1410 -2670 1416 -2664
rect 1410 -2676 1416 -2670
rect 1410 -2682 1416 -2676
rect 1410 -2688 1416 -2682
rect 1410 -2694 1416 -2688
rect 1410 -2700 1416 -2694
rect 1410 -2706 1416 -2700
rect 1410 -2712 1416 -2706
rect 1410 -2718 1416 -2712
rect 1410 -2724 1416 -2718
rect 1410 -2730 1416 -2724
rect 1410 -2736 1416 -2730
rect 1410 -2742 1416 -2736
rect 1410 -2748 1416 -2742
rect 1410 -2754 1416 -2748
rect 1410 -2760 1416 -2754
rect 1410 -2766 1416 -2760
rect 1410 -2772 1416 -2766
rect 1410 -2778 1416 -2772
rect 1410 -2784 1416 -2778
rect 1410 -2790 1416 -2784
rect 1410 -2796 1416 -2790
rect 1410 -2802 1416 -2796
rect 1410 -2808 1416 -2802
rect 1410 -2814 1416 -2808
rect 1410 -2820 1416 -2814
rect 1410 -2826 1416 -2820
rect 1410 -2832 1416 -2826
rect 1410 -2838 1416 -2832
rect 1410 -2844 1416 -2838
rect 1410 -2850 1416 -2844
rect 1410 -2856 1416 -2850
rect 1410 -2862 1416 -2856
rect 1410 -2868 1416 -2862
rect 1410 -2952 1416 -2946
rect 1410 -2958 1416 -2952
rect 1410 -2964 1416 -2958
rect 1410 -2970 1416 -2964
rect 1410 -2976 1416 -2970
rect 1410 -2982 1416 -2976
rect 1410 -2988 1416 -2982
rect 1410 -2994 1416 -2988
rect 1410 -3000 1416 -2994
rect 1410 -3006 1416 -3000
rect 1410 -3012 1416 -3006
rect 1410 -3018 1416 -3012
rect 1410 -3024 1416 -3018
rect 1410 -3030 1416 -3024
rect 1410 -3036 1416 -3030
rect 1410 -3042 1416 -3036
rect 1410 -3048 1416 -3042
rect 1410 -3054 1416 -3048
rect 1410 -3060 1416 -3054
rect 1410 -3066 1416 -3060
rect 1410 -3072 1416 -3066
rect 1410 -3078 1416 -3072
rect 1410 -3084 1416 -3078
rect 1410 -3090 1416 -3084
rect 1410 -3096 1416 -3090
rect 1410 -3102 1416 -3096
rect 1410 -3108 1416 -3102
rect 1410 -3114 1416 -3108
rect 1410 -3120 1416 -3114
rect 1410 -3126 1416 -3120
rect 1410 -3132 1416 -3126
rect 1410 -3138 1416 -3132
rect 1410 -3144 1416 -3138
rect 1410 -3150 1416 -3144
rect 1410 -3156 1416 -3150
rect 1410 -3162 1416 -3156
rect 1410 -3168 1416 -3162
rect 1410 -3174 1416 -3168
rect 1410 -3180 1416 -3174
rect 1410 -3186 1416 -3180
rect 1410 -3192 1416 -3186
rect 1410 -3198 1416 -3192
rect 1410 -3204 1416 -3198
rect 1410 -3210 1416 -3204
rect 1410 -3216 1416 -3210
rect 1410 -3222 1416 -3216
rect 1410 -3228 1416 -3222
rect 1410 -3234 1416 -3228
rect 1410 -3300 1416 -3294
rect 1410 -3306 1416 -3300
rect 1410 -3312 1416 -3306
rect 1410 -3318 1416 -3312
rect 1410 -3324 1416 -3318
rect 1410 -3330 1416 -3324
rect 1410 -3336 1416 -3330
rect 1410 -3342 1416 -3336
rect 1410 -3348 1416 -3342
rect 1410 -3354 1416 -3348
rect 1410 -3360 1416 -3354
rect 1410 -3366 1416 -3360
rect 1410 -3372 1416 -3366
rect 1410 -3378 1416 -3372
rect 1410 -3384 1416 -3378
rect 1410 -3390 1416 -3384
rect 1410 -3396 1416 -3390
rect 1410 -3402 1416 -3396
rect 1410 -3408 1416 -3402
rect 1410 -3414 1416 -3408
rect 1410 -3420 1416 -3414
rect 1410 -3426 1416 -3420
rect 1410 -3432 1416 -3426
rect 1410 -3438 1416 -3432
rect 1410 -3444 1416 -3438
rect 1410 -3450 1416 -3444
rect 1410 -3456 1416 -3450
rect 1410 -3462 1416 -3456
rect 1410 -3468 1416 -3462
rect 1410 -3474 1416 -3468
rect 1410 -3480 1416 -3474
rect 1410 -3486 1416 -3480
rect 1410 -3492 1416 -3486
rect 1410 -3498 1416 -3492
rect 1410 -3504 1416 -3498
rect 1416 -1116 1422 -1110
rect 1416 -1122 1422 -1116
rect 1416 -1128 1422 -1122
rect 1416 -1134 1422 -1128
rect 1416 -1140 1422 -1134
rect 1416 -1146 1422 -1140
rect 1416 -1152 1422 -1146
rect 1416 -1158 1422 -1152
rect 1416 -1164 1422 -1158
rect 1416 -1170 1422 -1164
rect 1416 -1176 1422 -1170
rect 1416 -1182 1422 -1176
rect 1416 -1188 1422 -1182
rect 1416 -1194 1422 -1188
rect 1416 -1200 1422 -1194
rect 1416 -1206 1422 -1200
rect 1416 -1212 1422 -1206
rect 1416 -1218 1422 -1212
rect 1416 -1332 1422 -1326
rect 1416 -1338 1422 -1332
rect 1416 -1344 1422 -1338
rect 1416 -1350 1422 -1344
rect 1416 -1356 1422 -1350
rect 1416 -1362 1422 -1356
rect 1416 -1368 1422 -1362
rect 1416 -1374 1422 -1368
rect 1416 -1380 1422 -1374
rect 1416 -1386 1422 -1380
rect 1416 -1392 1422 -1386
rect 1416 -1398 1422 -1392
rect 1416 -1404 1422 -1398
rect 1416 -1410 1422 -1404
rect 1416 -1416 1422 -1410
rect 1416 -1422 1422 -1416
rect 1416 -1428 1422 -1422
rect 1416 -1434 1422 -1428
rect 1416 -1440 1422 -1434
rect 1416 -1446 1422 -1440
rect 1416 -1452 1422 -1446
rect 1416 -1458 1422 -1452
rect 1416 -1464 1422 -1458
rect 1416 -1470 1422 -1464
rect 1416 -1476 1422 -1470
rect 1416 -1482 1422 -1476
rect 1416 -1488 1422 -1482
rect 1416 -1494 1422 -1488
rect 1416 -1500 1422 -1494
rect 1416 -1506 1422 -1500
rect 1416 -1512 1422 -1506
rect 1416 -1518 1422 -1512
rect 1416 -1524 1422 -1518
rect 1416 -1530 1422 -1524
rect 1416 -1536 1422 -1530
rect 1416 -1542 1422 -1536
rect 1416 -1548 1422 -1542
rect 1416 -1554 1422 -1548
rect 1416 -1560 1422 -1554
rect 1416 -1566 1422 -1560
rect 1416 -1572 1422 -1566
rect 1416 -1578 1422 -1572
rect 1416 -1584 1422 -1578
rect 1416 -1590 1422 -1584
rect 1416 -1596 1422 -1590
rect 1416 -1602 1422 -1596
rect 1416 -1608 1422 -1602
rect 1416 -1614 1422 -1608
rect 1416 -1620 1422 -1614
rect 1416 -1626 1422 -1620
rect 1416 -1632 1422 -1626
rect 1416 -1638 1422 -1632
rect 1416 -1644 1422 -1638
rect 1416 -1650 1422 -1644
rect 1416 -1656 1422 -1650
rect 1416 -1662 1422 -1656
rect 1416 -1668 1422 -1662
rect 1416 -1674 1422 -1668
rect 1416 -1680 1422 -1674
rect 1416 -1686 1422 -1680
rect 1416 -1692 1422 -1686
rect 1416 -1698 1422 -1692
rect 1416 -1704 1422 -1698
rect 1416 -1710 1422 -1704
rect 1416 -1716 1422 -1710
rect 1416 -1722 1422 -1716
rect 1416 -1728 1422 -1722
rect 1416 -1734 1422 -1728
rect 1416 -1740 1422 -1734
rect 1416 -1746 1422 -1740
rect 1416 -1752 1422 -1746
rect 1416 -1758 1422 -1752
rect 1416 -1764 1422 -1758
rect 1416 -1770 1422 -1764
rect 1416 -1776 1422 -1770
rect 1416 -1782 1422 -1776
rect 1416 -1788 1422 -1782
rect 1416 -1794 1422 -1788
rect 1416 -1800 1422 -1794
rect 1416 -1806 1422 -1800
rect 1416 -1812 1422 -1806
rect 1416 -1818 1422 -1812
rect 1416 -1824 1422 -1818
rect 1416 -1830 1422 -1824
rect 1416 -1836 1422 -1830
rect 1416 -1842 1422 -1836
rect 1416 -1848 1422 -1842
rect 1416 -1854 1422 -1848
rect 1416 -1860 1422 -1854
rect 1416 -1866 1422 -1860
rect 1416 -1872 1422 -1866
rect 1416 -1878 1422 -1872
rect 1416 -1884 1422 -1878
rect 1416 -1890 1422 -1884
rect 1416 -1896 1422 -1890
rect 1416 -1902 1422 -1896
rect 1416 -1908 1422 -1902
rect 1416 -1914 1422 -1908
rect 1416 -1920 1422 -1914
rect 1416 -1926 1422 -1920
rect 1416 -1932 1422 -1926
rect 1416 -1938 1422 -1932
rect 1416 -1944 1422 -1938
rect 1416 -1950 1422 -1944
rect 1416 -1956 1422 -1950
rect 1416 -1962 1422 -1956
rect 1416 -1968 1422 -1962
rect 1416 -1974 1422 -1968
rect 1416 -1980 1422 -1974
rect 1416 -1986 1422 -1980
rect 1416 -1992 1422 -1986
rect 1416 -1998 1422 -1992
rect 1416 -2004 1422 -1998
rect 1416 -2010 1422 -2004
rect 1416 -2016 1422 -2010
rect 1416 -2022 1422 -2016
rect 1416 -2028 1422 -2022
rect 1416 -2034 1422 -2028
rect 1416 -2040 1422 -2034
rect 1416 -2046 1422 -2040
rect 1416 -2052 1422 -2046
rect 1416 -2058 1422 -2052
rect 1416 -2064 1422 -2058
rect 1416 -2070 1422 -2064
rect 1416 -2076 1422 -2070
rect 1416 -2082 1422 -2076
rect 1416 -2088 1422 -2082
rect 1416 -2094 1422 -2088
rect 1416 -2100 1422 -2094
rect 1416 -2106 1422 -2100
rect 1416 -2112 1422 -2106
rect 1416 -2118 1422 -2112
rect 1416 -2124 1422 -2118
rect 1416 -2130 1422 -2124
rect 1416 -2136 1422 -2130
rect 1416 -2142 1422 -2136
rect 1416 -2148 1422 -2142
rect 1416 -2154 1422 -2148
rect 1416 -2160 1422 -2154
rect 1416 -2166 1422 -2160
rect 1416 -2172 1422 -2166
rect 1416 -2178 1422 -2172
rect 1416 -2184 1422 -2178
rect 1416 -2190 1422 -2184
rect 1416 -2196 1422 -2190
rect 1416 -2202 1422 -2196
rect 1416 -2208 1422 -2202
rect 1416 -2214 1422 -2208
rect 1416 -2220 1422 -2214
rect 1416 -2226 1422 -2220
rect 1416 -2232 1422 -2226
rect 1416 -2238 1422 -2232
rect 1416 -2244 1422 -2238
rect 1416 -2250 1422 -2244
rect 1416 -2256 1422 -2250
rect 1416 -2262 1422 -2256
rect 1416 -2268 1422 -2262
rect 1416 -2274 1422 -2268
rect 1416 -2280 1422 -2274
rect 1416 -2286 1422 -2280
rect 1416 -2292 1422 -2286
rect 1416 -2298 1422 -2292
rect 1416 -2376 1422 -2370
rect 1416 -2382 1422 -2376
rect 1416 -2388 1422 -2382
rect 1416 -2394 1422 -2388
rect 1416 -2400 1422 -2394
rect 1416 -2406 1422 -2400
rect 1416 -2412 1422 -2406
rect 1416 -2418 1422 -2412
rect 1416 -2424 1422 -2418
rect 1416 -2430 1422 -2424
rect 1416 -2436 1422 -2430
rect 1416 -2442 1422 -2436
rect 1416 -2448 1422 -2442
rect 1416 -2454 1422 -2448
rect 1416 -2460 1422 -2454
rect 1416 -2466 1422 -2460
rect 1416 -2472 1422 -2466
rect 1416 -2478 1422 -2472
rect 1416 -2484 1422 -2478
rect 1416 -2490 1422 -2484
rect 1416 -2496 1422 -2490
rect 1416 -2502 1422 -2496
rect 1416 -2508 1422 -2502
rect 1416 -2514 1422 -2508
rect 1416 -2520 1422 -2514
rect 1416 -2526 1422 -2520
rect 1416 -2532 1422 -2526
rect 1416 -2538 1422 -2532
rect 1416 -2544 1422 -2538
rect 1416 -2550 1422 -2544
rect 1416 -2556 1422 -2550
rect 1416 -2562 1422 -2556
rect 1416 -2568 1422 -2562
rect 1416 -2574 1422 -2568
rect 1416 -2580 1422 -2574
rect 1416 -2586 1422 -2580
rect 1416 -2592 1422 -2586
rect 1416 -2598 1422 -2592
rect 1416 -2604 1422 -2598
rect 1416 -2610 1422 -2604
rect 1416 -2616 1422 -2610
rect 1416 -2622 1422 -2616
rect 1416 -2628 1422 -2622
rect 1416 -2634 1422 -2628
rect 1416 -2640 1422 -2634
rect 1416 -2646 1422 -2640
rect 1416 -2652 1422 -2646
rect 1416 -2658 1422 -2652
rect 1416 -2664 1422 -2658
rect 1416 -2670 1422 -2664
rect 1416 -2676 1422 -2670
rect 1416 -2682 1422 -2676
rect 1416 -2688 1422 -2682
rect 1416 -2694 1422 -2688
rect 1416 -2700 1422 -2694
rect 1416 -2706 1422 -2700
rect 1416 -2712 1422 -2706
rect 1416 -2718 1422 -2712
rect 1416 -2724 1422 -2718
rect 1416 -2730 1422 -2724
rect 1416 -2736 1422 -2730
rect 1416 -2742 1422 -2736
rect 1416 -2748 1422 -2742
rect 1416 -2754 1422 -2748
rect 1416 -2760 1422 -2754
rect 1416 -2766 1422 -2760
rect 1416 -2772 1422 -2766
rect 1416 -2778 1422 -2772
rect 1416 -2784 1422 -2778
rect 1416 -2790 1422 -2784
rect 1416 -2796 1422 -2790
rect 1416 -2802 1422 -2796
rect 1416 -2808 1422 -2802
rect 1416 -2814 1422 -2808
rect 1416 -2820 1422 -2814
rect 1416 -2826 1422 -2820
rect 1416 -2832 1422 -2826
rect 1416 -2838 1422 -2832
rect 1416 -2844 1422 -2838
rect 1416 -2850 1422 -2844
rect 1416 -2856 1422 -2850
rect 1416 -2862 1422 -2856
rect 1416 -2952 1422 -2946
rect 1416 -2958 1422 -2952
rect 1416 -2964 1422 -2958
rect 1416 -2970 1422 -2964
rect 1416 -2976 1422 -2970
rect 1416 -2982 1422 -2976
rect 1416 -2988 1422 -2982
rect 1416 -2994 1422 -2988
rect 1416 -3000 1422 -2994
rect 1416 -3006 1422 -3000
rect 1416 -3012 1422 -3006
rect 1416 -3018 1422 -3012
rect 1416 -3024 1422 -3018
rect 1416 -3030 1422 -3024
rect 1416 -3036 1422 -3030
rect 1416 -3042 1422 -3036
rect 1416 -3048 1422 -3042
rect 1416 -3054 1422 -3048
rect 1416 -3060 1422 -3054
rect 1416 -3066 1422 -3060
rect 1416 -3072 1422 -3066
rect 1416 -3078 1422 -3072
rect 1416 -3084 1422 -3078
rect 1416 -3090 1422 -3084
rect 1416 -3096 1422 -3090
rect 1416 -3102 1422 -3096
rect 1416 -3108 1422 -3102
rect 1416 -3114 1422 -3108
rect 1416 -3120 1422 -3114
rect 1416 -3126 1422 -3120
rect 1416 -3132 1422 -3126
rect 1416 -3138 1422 -3132
rect 1416 -3144 1422 -3138
rect 1416 -3150 1422 -3144
rect 1416 -3156 1422 -3150
rect 1416 -3162 1422 -3156
rect 1416 -3168 1422 -3162
rect 1416 -3174 1422 -3168
rect 1416 -3180 1422 -3174
rect 1416 -3186 1422 -3180
rect 1416 -3192 1422 -3186
rect 1416 -3198 1422 -3192
rect 1416 -3204 1422 -3198
rect 1416 -3210 1422 -3204
rect 1416 -3216 1422 -3210
rect 1416 -3222 1422 -3216
rect 1416 -3228 1422 -3222
rect 1416 -3234 1422 -3228
rect 1416 -3300 1422 -3294
rect 1416 -3306 1422 -3300
rect 1416 -3312 1422 -3306
rect 1416 -3318 1422 -3312
rect 1416 -3324 1422 -3318
rect 1416 -3330 1422 -3324
rect 1416 -3336 1422 -3330
rect 1416 -3342 1422 -3336
rect 1416 -3348 1422 -3342
rect 1416 -3354 1422 -3348
rect 1416 -3360 1422 -3354
rect 1416 -3366 1422 -3360
rect 1416 -3372 1422 -3366
rect 1416 -3378 1422 -3372
rect 1416 -3384 1422 -3378
rect 1416 -3390 1422 -3384
rect 1416 -3396 1422 -3390
rect 1416 -3402 1422 -3396
rect 1416 -3408 1422 -3402
rect 1416 -3414 1422 -3408
rect 1416 -3420 1422 -3414
rect 1416 -3426 1422 -3420
rect 1416 -3432 1422 -3426
rect 1416 -3438 1422 -3432
rect 1416 -3444 1422 -3438
rect 1416 -3450 1422 -3444
rect 1416 -3456 1422 -3450
rect 1416 -3462 1422 -3456
rect 1416 -3468 1422 -3462
rect 1416 -3474 1422 -3468
rect 1416 -3480 1422 -3474
rect 1416 -3486 1422 -3480
rect 1416 -3492 1422 -3486
rect 1416 -3498 1422 -3492
rect 1416 -3504 1422 -3498
rect 1422 -1116 1428 -1110
rect 1422 -1122 1428 -1116
rect 1422 -1128 1428 -1122
rect 1422 -1134 1428 -1128
rect 1422 -1140 1428 -1134
rect 1422 -1146 1428 -1140
rect 1422 -1152 1428 -1146
rect 1422 -1158 1428 -1152
rect 1422 -1164 1428 -1158
rect 1422 -1170 1428 -1164
rect 1422 -1176 1428 -1170
rect 1422 -1182 1428 -1176
rect 1422 -1188 1428 -1182
rect 1422 -1194 1428 -1188
rect 1422 -1200 1428 -1194
rect 1422 -1206 1428 -1200
rect 1422 -1320 1428 -1314
rect 1422 -1326 1428 -1320
rect 1422 -1332 1428 -1326
rect 1422 -1338 1428 -1332
rect 1422 -1344 1428 -1338
rect 1422 -1350 1428 -1344
rect 1422 -1356 1428 -1350
rect 1422 -1362 1428 -1356
rect 1422 -1368 1428 -1362
rect 1422 -1374 1428 -1368
rect 1422 -1380 1428 -1374
rect 1422 -1386 1428 -1380
rect 1422 -1392 1428 -1386
rect 1422 -1398 1428 -1392
rect 1422 -1404 1428 -1398
rect 1422 -1410 1428 -1404
rect 1422 -1416 1428 -1410
rect 1422 -1422 1428 -1416
rect 1422 -1428 1428 -1422
rect 1422 -1434 1428 -1428
rect 1422 -1440 1428 -1434
rect 1422 -1446 1428 -1440
rect 1422 -1452 1428 -1446
rect 1422 -1458 1428 -1452
rect 1422 -1464 1428 -1458
rect 1422 -1470 1428 -1464
rect 1422 -1476 1428 -1470
rect 1422 -1482 1428 -1476
rect 1422 -1488 1428 -1482
rect 1422 -1494 1428 -1488
rect 1422 -1500 1428 -1494
rect 1422 -1506 1428 -1500
rect 1422 -1512 1428 -1506
rect 1422 -1518 1428 -1512
rect 1422 -1524 1428 -1518
rect 1422 -1530 1428 -1524
rect 1422 -1536 1428 -1530
rect 1422 -1542 1428 -1536
rect 1422 -1548 1428 -1542
rect 1422 -1554 1428 -1548
rect 1422 -1560 1428 -1554
rect 1422 -1566 1428 -1560
rect 1422 -1572 1428 -1566
rect 1422 -1578 1428 -1572
rect 1422 -1584 1428 -1578
rect 1422 -1590 1428 -1584
rect 1422 -1596 1428 -1590
rect 1422 -1602 1428 -1596
rect 1422 -1608 1428 -1602
rect 1422 -1614 1428 -1608
rect 1422 -1620 1428 -1614
rect 1422 -1626 1428 -1620
rect 1422 -1632 1428 -1626
rect 1422 -1638 1428 -1632
rect 1422 -1644 1428 -1638
rect 1422 -1650 1428 -1644
rect 1422 -1656 1428 -1650
rect 1422 -1662 1428 -1656
rect 1422 -1668 1428 -1662
rect 1422 -1674 1428 -1668
rect 1422 -1680 1428 -1674
rect 1422 -1686 1428 -1680
rect 1422 -1692 1428 -1686
rect 1422 -1698 1428 -1692
rect 1422 -1704 1428 -1698
rect 1422 -1710 1428 -1704
rect 1422 -1716 1428 -1710
rect 1422 -1722 1428 -1716
rect 1422 -1728 1428 -1722
rect 1422 -1734 1428 -1728
rect 1422 -1740 1428 -1734
rect 1422 -1746 1428 -1740
rect 1422 -1752 1428 -1746
rect 1422 -1758 1428 -1752
rect 1422 -1764 1428 -1758
rect 1422 -1770 1428 -1764
rect 1422 -1776 1428 -1770
rect 1422 -1782 1428 -1776
rect 1422 -1788 1428 -1782
rect 1422 -1794 1428 -1788
rect 1422 -1800 1428 -1794
rect 1422 -1806 1428 -1800
rect 1422 -1812 1428 -1806
rect 1422 -1818 1428 -1812
rect 1422 -1824 1428 -1818
rect 1422 -1830 1428 -1824
rect 1422 -1836 1428 -1830
rect 1422 -1842 1428 -1836
rect 1422 -1848 1428 -1842
rect 1422 -1854 1428 -1848
rect 1422 -1860 1428 -1854
rect 1422 -1866 1428 -1860
rect 1422 -1872 1428 -1866
rect 1422 -1878 1428 -1872
rect 1422 -1884 1428 -1878
rect 1422 -1890 1428 -1884
rect 1422 -1896 1428 -1890
rect 1422 -1902 1428 -1896
rect 1422 -1908 1428 -1902
rect 1422 -1914 1428 -1908
rect 1422 -1920 1428 -1914
rect 1422 -1926 1428 -1920
rect 1422 -1932 1428 -1926
rect 1422 -1938 1428 -1932
rect 1422 -1944 1428 -1938
rect 1422 -1950 1428 -1944
rect 1422 -1956 1428 -1950
rect 1422 -1962 1428 -1956
rect 1422 -1968 1428 -1962
rect 1422 -1974 1428 -1968
rect 1422 -1980 1428 -1974
rect 1422 -1986 1428 -1980
rect 1422 -1992 1428 -1986
rect 1422 -1998 1428 -1992
rect 1422 -2004 1428 -1998
rect 1422 -2010 1428 -2004
rect 1422 -2016 1428 -2010
rect 1422 -2022 1428 -2016
rect 1422 -2028 1428 -2022
rect 1422 -2034 1428 -2028
rect 1422 -2040 1428 -2034
rect 1422 -2046 1428 -2040
rect 1422 -2052 1428 -2046
rect 1422 -2058 1428 -2052
rect 1422 -2064 1428 -2058
rect 1422 -2070 1428 -2064
rect 1422 -2076 1428 -2070
rect 1422 -2082 1428 -2076
rect 1422 -2088 1428 -2082
rect 1422 -2094 1428 -2088
rect 1422 -2100 1428 -2094
rect 1422 -2106 1428 -2100
rect 1422 -2112 1428 -2106
rect 1422 -2118 1428 -2112
rect 1422 -2124 1428 -2118
rect 1422 -2130 1428 -2124
rect 1422 -2136 1428 -2130
rect 1422 -2142 1428 -2136
rect 1422 -2148 1428 -2142
rect 1422 -2154 1428 -2148
rect 1422 -2160 1428 -2154
rect 1422 -2166 1428 -2160
rect 1422 -2172 1428 -2166
rect 1422 -2178 1428 -2172
rect 1422 -2184 1428 -2178
rect 1422 -2190 1428 -2184
rect 1422 -2196 1428 -2190
rect 1422 -2202 1428 -2196
rect 1422 -2208 1428 -2202
rect 1422 -2214 1428 -2208
rect 1422 -2220 1428 -2214
rect 1422 -2226 1428 -2220
rect 1422 -2232 1428 -2226
rect 1422 -2238 1428 -2232
rect 1422 -2244 1428 -2238
rect 1422 -2250 1428 -2244
rect 1422 -2256 1428 -2250
rect 1422 -2262 1428 -2256
rect 1422 -2268 1428 -2262
rect 1422 -2274 1428 -2268
rect 1422 -2280 1428 -2274
rect 1422 -2286 1428 -2280
rect 1422 -2292 1428 -2286
rect 1422 -2370 1428 -2364
rect 1422 -2376 1428 -2370
rect 1422 -2382 1428 -2376
rect 1422 -2388 1428 -2382
rect 1422 -2394 1428 -2388
rect 1422 -2400 1428 -2394
rect 1422 -2406 1428 -2400
rect 1422 -2412 1428 -2406
rect 1422 -2418 1428 -2412
rect 1422 -2424 1428 -2418
rect 1422 -2430 1428 -2424
rect 1422 -2436 1428 -2430
rect 1422 -2442 1428 -2436
rect 1422 -2448 1428 -2442
rect 1422 -2454 1428 -2448
rect 1422 -2460 1428 -2454
rect 1422 -2466 1428 -2460
rect 1422 -2472 1428 -2466
rect 1422 -2478 1428 -2472
rect 1422 -2484 1428 -2478
rect 1422 -2490 1428 -2484
rect 1422 -2496 1428 -2490
rect 1422 -2502 1428 -2496
rect 1422 -2508 1428 -2502
rect 1422 -2514 1428 -2508
rect 1422 -2520 1428 -2514
rect 1422 -2526 1428 -2520
rect 1422 -2532 1428 -2526
rect 1422 -2538 1428 -2532
rect 1422 -2544 1428 -2538
rect 1422 -2550 1428 -2544
rect 1422 -2556 1428 -2550
rect 1422 -2562 1428 -2556
rect 1422 -2568 1428 -2562
rect 1422 -2574 1428 -2568
rect 1422 -2580 1428 -2574
rect 1422 -2586 1428 -2580
rect 1422 -2592 1428 -2586
rect 1422 -2598 1428 -2592
rect 1422 -2604 1428 -2598
rect 1422 -2610 1428 -2604
rect 1422 -2616 1428 -2610
rect 1422 -2622 1428 -2616
rect 1422 -2628 1428 -2622
rect 1422 -2634 1428 -2628
rect 1422 -2640 1428 -2634
rect 1422 -2646 1428 -2640
rect 1422 -2652 1428 -2646
rect 1422 -2658 1428 -2652
rect 1422 -2664 1428 -2658
rect 1422 -2670 1428 -2664
rect 1422 -2676 1428 -2670
rect 1422 -2682 1428 -2676
rect 1422 -2688 1428 -2682
rect 1422 -2694 1428 -2688
rect 1422 -2700 1428 -2694
rect 1422 -2706 1428 -2700
rect 1422 -2712 1428 -2706
rect 1422 -2718 1428 -2712
rect 1422 -2724 1428 -2718
rect 1422 -2730 1428 -2724
rect 1422 -2736 1428 -2730
rect 1422 -2742 1428 -2736
rect 1422 -2748 1428 -2742
rect 1422 -2754 1428 -2748
rect 1422 -2760 1428 -2754
rect 1422 -2766 1428 -2760
rect 1422 -2772 1428 -2766
rect 1422 -2778 1428 -2772
rect 1422 -2784 1428 -2778
rect 1422 -2790 1428 -2784
rect 1422 -2796 1428 -2790
rect 1422 -2802 1428 -2796
rect 1422 -2808 1428 -2802
rect 1422 -2814 1428 -2808
rect 1422 -2820 1428 -2814
rect 1422 -2826 1428 -2820
rect 1422 -2832 1428 -2826
rect 1422 -2838 1428 -2832
rect 1422 -2844 1428 -2838
rect 1422 -2850 1428 -2844
rect 1422 -2856 1428 -2850
rect 1422 -2862 1428 -2856
rect 1422 -2946 1428 -2940
rect 1422 -2952 1428 -2946
rect 1422 -2958 1428 -2952
rect 1422 -2964 1428 -2958
rect 1422 -2970 1428 -2964
rect 1422 -2976 1428 -2970
rect 1422 -2982 1428 -2976
rect 1422 -2988 1428 -2982
rect 1422 -2994 1428 -2988
rect 1422 -3000 1428 -2994
rect 1422 -3006 1428 -3000
rect 1422 -3012 1428 -3006
rect 1422 -3018 1428 -3012
rect 1422 -3024 1428 -3018
rect 1422 -3030 1428 -3024
rect 1422 -3036 1428 -3030
rect 1422 -3042 1428 -3036
rect 1422 -3048 1428 -3042
rect 1422 -3054 1428 -3048
rect 1422 -3060 1428 -3054
rect 1422 -3066 1428 -3060
rect 1422 -3072 1428 -3066
rect 1422 -3078 1428 -3072
rect 1422 -3084 1428 -3078
rect 1422 -3090 1428 -3084
rect 1422 -3096 1428 -3090
rect 1422 -3102 1428 -3096
rect 1422 -3108 1428 -3102
rect 1422 -3114 1428 -3108
rect 1422 -3120 1428 -3114
rect 1422 -3126 1428 -3120
rect 1422 -3132 1428 -3126
rect 1422 -3138 1428 -3132
rect 1422 -3144 1428 -3138
rect 1422 -3150 1428 -3144
rect 1422 -3156 1428 -3150
rect 1422 -3162 1428 -3156
rect 1422 -3168 1428 -3162
rect 1422 -3174 1428 -3168
rect 1422 -3180 1428 -3174
rect 1422 -3186 1428 -3180
rect 1422 -3192 1428 -3186
rect 1422 -3198 1428 -3192
rect 1422 -3204 1428 -3198
rect 1422 -3210 1428 -3204
rect 1422 -3216 1428 -3210
rect 1422 -3222 1428 -3216
rect 1422 -3228 1428 -3222
rect 1422 -3234 1428 -3228
rect 1422 -3300 1428 -3294
rect 1422 -3306 1428 -3300
rect 1422 -3312 1428 -3306
rect 1422 -3318 1428 -3312
rect 1422 -3324 1428 -3318
rect 1422 -3330 1428 -3324
rect 1422 -3336 1428 -3330
rect 1422 -3342 1428 -3336
rect 1422 -3348 1428 -3342
rect 1422 -3354 1428 -3348
rect 1422 -3360 1428 -3354
rect 1422 -3366 1428 -3360
rect 1422 -3372 1428 -3366
rect 1422 -3378 1428 -3372
rect 1422 -3384 1428 -3378
rect 1422 -3390 1428 -3384
rect 1422 -3396 1428 -3390
rect 1422 -3402 1428 -3396
rect 1422 -3408 1428 -3402
rect 1422 -3414 1428 -3408
rect 1422 -3420 1428 -3414
rect 1422 -3426 1428 -3420
rect 1422 -3432 1428 -3426
rect 1422 -3438 1428 -3432
rect 1422 -3444 1428 -3438
rect 1422 -3450 1428 -3444
rect 1422 -3456 1428 -3450
rect 1422 -3462 1428 -3456
rect 1422 -3468 1428 -3462
rect 1422 -3474 1428 -3468
rect 1422 -3480 1428 -3474
rect 1422 -3486 1428 -3480
rect 1422 -3492 1428 -3486
rect 1422 -3498 1428 -3492
rect 1422 -3504 1428 -3498
rect 1428 -1122 1434 -1116
rect 1428 -1128 1434 -1122
rect 1428 -1134 1434 -1128
rect 1428 -1140 1434 -1134
rect 1428 -1146 1434 -1140
rect 1428 -1152 1434 -1146
rect 1428 -1158 1434 -1152
rect 1428 -1164 1434 -1158
rect 1428 -1170 1434 -1164
rect 1428 -1176 1434 -1170
rect 1428 -1182 1434 -1176
rect 1428 -1188 1434 -1182
rect 1428 -1194 1434 -1188
rect 1428 -1308 1434 -1302
rect 1428 -1314 1434 -1308
rect 1428 -1320 1434 -1314
rect 1428 -1326 1434 -1320
rect 1428 -1332 1434 -1326
rect 1428 -1338 1434 -1332
rect 1428 -1344 1434 -1338
rect 1428 -1350 1434 -1344
rect 1428 -1356 1434 -1350
rect 1428 -1362 1434 -1356
rect 1428 -1368 1434 -1362
rect 1428 -1374 1434 -1368
rect 1428 -1380 1434 -1374
rect 1428 -1386 1434 -1380
rect 1428 -1392 1434 -1386
rect 1428 -1398 1434 -1392
rect 1428 -1404 1434 -1398
rect 1428 -1410 1434 -1404
rect 1428 -1416 1434 -1410
rect 1428 -1422 1434 -1416
rect 1428 -1428 1434 -1422
rect 1428 -1434 1434 -1428
rect 1428 -1440 1434 -1434
rect 1428 -1446 1434 -1440
rect 1428 -1452 1434 -1446
rect 1428 -1458 1434 -1452
rect 1428 -1464 1434 -1458
rect 1428 -1470 1434 -1464
rect 1428 -1476 1434 -1470
rect 1428 -1482 1434 -1476
rect 1428 -1488 1434 -1482
rect 1428 -1494 1434 -1488
rect 1428 -1500 1434 -1494
rect 1428 -1506 1434 -1500
rect 1428 -1512 1434 -1506
rect 1428 -1518 1434 -1512
rect 1428 -1524 1434 -1518
rect 1428 -1530 1434 -1524
rect 1428 -1536 1434 -1530
rect 1428 -1542 1434 -1536
rect 1428 -1548 1434 -1542
rect 1428 -1554 1434 -1548
rect 1428 -1560 1434 -1554
rect 1428 -1566 1434 -1560
rect 1428 -1572 1434 -1566
rect 1428 -1578 1434 -1572
rect 1428 -1584 1434 -1578
rect 1428 -1590 1434 -1584
rect 1428 -1596 1434 -1590
rect 1428 -1602 1434 -1596
rect 1428 -1608 1434 -1602
rect 1428 -1614 1434 -1608
rect 1428 -1620 1434 -1614
rect 1428 -1626 1434 -1620
rect 1428 -1632 1434 -1626
rect 1428 -1638 1434 -1632
rect 1428 -1644 1434 -1638
rect 1428 -1650 1434 -1644
rect 1428 -1656 1434 -1650
rect 1428 -1662 1434 -1656
rect 1428 -1668 1434 -1662
rect 1428 -1674 1434 -1668
rect 1428 -1680 1434 -1674
rect 1428 -1686 1434 -1680
rect 1428 -1692 1434 -1686
rect 1428 -1698 1434 -1692
rect 1428 -1704 1434 -1698
rect 1428 -1710 1434 -1704
rect 1428 -1716 1434 -1710
rect 1428 -1722 1434 -1716
rect 1428 -1728 1434 -1722
rect 1428 -1734 1434 -1728
rect 1428 -1740 1434 -1734
rect 1428 -1746 1434 -1740
rect 1428 -1752 1434 -1746
rect 1428 -1758 1434 -1752
rect 1428 -1764 1434 -1758
rect 1428 -1770 1434 -1764
rect 1428 -1776 1434 -1770
rect 1428 -1782 1434 -1776
rect 1428 -1788 1434 -1782
rect 1428 -1794 1434 -1788
rect 1428 -1800 1434 -1794
rect 1428 -1806 1434 -1800
rect 1428 -1812 1434 -1806
rect 1428 -1818 1434 -1812
rect 1428 -1824 1434 -1818
rect 1428 -1830 1434 -1824
rect 1428 -1836 1434 -1830
rect 1428 -1842 1434 -1836
rect 1428 -1848 1434 -1842
rect 1428 -1854 1434 -1848
rect 1428 -1860 1434 -1854
rect 1428 -1866 1434 -1860
rect 1428 -1872 1434 -1866
rect 1428 -1878 1434 -1872
rect 1428 -1884 1434 -1878
rect 1428 -1890 1434 -1884
rect 1428 -1896 1434 -1890
rect 1428 -1902 1434 -1896
rect 1428 -1908 1434 -1902
rect 1428 -1914 1434 -1908
rect 1428 -1920 1434 -1914
rect 1428 -1926 1434 -1920
rect 1428 -1932 1434 -1926
rect 1428 -1938 1434 -1932
rect 1428 -1944 1434 -1938
rect 1428 -1950 1434 -1944
rect 1428 -1956 1434 -1950
rect 1428 -1962 1434 -1956
rect 1428 -1968 1434 -1962
rect 1428 -1974 1434 -1968
rect 1428 -1980 1434 -1974
rect 1428 -1986 1434 -1980
rect 1428 -1992 1434 -1986
rect 1428 -1998 1434 -1992
rect 1428 -2004 1434 -1998
rect 1428 -2010 1434 -2004
rect 1428 -2016 1434 -2010
rect 1428 -2022 1434 -2016
rect 1428 -2028 1434 -2022
rect 1428 -2034 1434 -2028
rect 1428 -2040 1434 -2034
rect 1428 -2046 1434 -2040
rect 1428 -2052 1434 -2046
rect 1428 -2058 1434 -2052
rect 1428 -2064 1434 -2058
rect 1428 -2070 1434 -2064
rect 1428 -2076 1434 -2070
rect 1428 -2082 1434 -2076
rect 1428 -2088 1434 -2082
rect 1428 -2094 1434 -2088
rect 1428 -2100 1434 -2094
rect 1428 -2106 1434 -2100
rect 1428 -2112 1434 -2106
rect 1428 -2118 1434 -2112
rect 1428 -2124 1434 -2118
rect 1428 -2130 1434 -2124
rect 1428 -2136 1434 -2130
rect 1428 -2142 1434 -2136
rect 1428 -2148 1434 -2142
rect 1428 -2154 1434 -2148
rect 1428 -2160 1434 -2154
rect 1428 -2166 1434 -2160
rect 1428 -2172 1434 -2166
rect 1428 -2178 1434 -2172
rect 1428 -2184 1434 -2178
rect 1428 -2190 1434 -2184
rect 1428 -2196 1434 -2190
rect 1428 -2202 1434 -2196
rect 1428 -2208 1434 -2202
rect 1428 -2214 1434 -2208
rect 1428 -2220 1434 -2214
rect 1428 -2226 1434 -2220
rect 1428 -2232 1434 -2226
rect 1428 -2238 1434 -2232
rect 1428 -2244 1434 -2238
rect 1428 -2250 1434 -2244
rect 1428 -2256 1434 -2250
rect 1428 -2262 1434 -2256
rect 1428 -2268 1434 -2262
rect 1428 -2274 1434 -2268
rect 1428 -2280 1434 -2274
rect 1428 -2286 1434 -2280
rect 1428 -2358 1434 -2352
rect 1428 -2364 1434 -2358
rect 1428 -2370 1434 -2364
rect 1428 -2376 1434 -2370
rect 1428 -2382 1434 -2376
rect 1428 -2388 1434 -2382
rect 1428 -2394 1434 -2388
rect 1428 -2400 1434 -2394
rect 1428 -2406 1434 -2400
rect 1428 -2412 1434 -2406
rect 1428 -2418 1434 -2412
rect 1428 -2424 1434 -2418
rect 1428 -2430 1434 -2424
rect 1428 -2436 1434 -2430
rect 1428 -2442 1434 -2436
rect 1428 -2448 1434 -2442
rect 1428 -2454 1434 -2448
rect 1428 -2460 1434 -2454
rect 1428 -2466 1434 -2460
rect 1428 -2472 1434 -2466
rect 1428 -2478 1434 -2472
rect 1428 -2484 1434 -2478
rect 1428 -2490 1434 -2484
rect 1428 -2496 1434 -2490
rect 1428 -2502 1434 -2496
rect 1428 -2508 1434 -2502
rect 1428 -2514 1434 -2508
rect 1428 -2520 1434 -2514
rect 1428 -2526 1434 -2520
rect 1428 -2532 1434 -2526
rect 1428 -2538 1434 -2532
rect 1428 -2544 1434 -2538
rect 1428 -2550 1434 -2544
rect 1428 -2556 1434 -2550
rect 1428 -2562 1434 -2556
rect 1428 -2568 1434 -2562
rect 1428 -2574 1434 -2568
rect 1428 -2580 1434 -2574
rect 1428 -2586 1434 -2580
rect 1428 -2592 1434 -2586
rect 1428 -2598 1434 -2592
rect 1428 -2604 1434 -2598
rect 1428 -2610 1434 -2604
rect 1428 -2616 1434 -2610
rect 1428 -2622 1434 -2616
rect 1428 -2628 1434 -2622
rect 1428 -2634 1434 -2628
rect 1428 -2640 1434 -2634
rect 1428 -2646 1434 -2640
rect 1428 -2652 1434 -2646
rect 1428 -2658 1434 -2652
rect 1428 -2664 1434 -2658
rect 1428 -2670 1434 -2664
rect 1428 -2676 1434 -2670
rect 1428 -2682 1434 -2676
rect 1428 -2688 1434 -2682
rect 1428 -2694 1434 -2688
rect 1428 -2700 1434 -2694
rect 1428 -2706 1434 -2700
rect 1428 -2712 1434 -2706
rect 1428 -2718 1434 -2712
rect 1428 -2724 1434 -2718
rect 1428 -2730 1434 -2724
rect 1428 -2736 1434 -2730
rect 1428 -2742 1434 -2736
rect 1428 -2748 1434 -2742
rect 1428 -2754 1434 -2748
rect 1428 -2760 1434 -2754
rect 1428 -2766 1434 -2760
rect 1428 -2772 1434 -2766
rect 1428 -2778 1434 -2772
rect 1428 -2784 1434 -2778
rect 1428 -2790 1434 -2784
rect 1428 -2796 1434 -2790
rect 1428 -2802 1434 -2796
rect 1428 -2808 1434 -2802
rect 1428 -2814 1434 -2808
rect 1428 -2820 1434 -2814
rect 1428 -2826 1434 -2820
rect 1428 -2832 1434 -2826
rect 1428 -2838 1434 -2832
rect 1428 -2844 1434 -2838
rect 1428 -2850 1434 -2844
rect 1428 -2856 1434 -2850
rect 1428 -2940 1434 -2934
rect 1428 -2946 1434 -2940
rect 1428 -2952 1434 -2946
rect 1428 -2958 1434 -2952
rect 1428 -2964 1434 -2958
rect 1428 -2970 1434 -2964
rect 1428 -2976 1434 -2970
rect 1428 -2982 1434 -2976
rect 1428 -2988 1434 -2982
rect 1428 -2994 1434 -2988
rect 1428 -3000 1434 -2994
rect 1428 -3006 1434 -3000
rect 1428 -3012 1434 -3006
rect 1428 -3018 1434 -3012
rect 1428 -3024 1434 -3018
rect 1428 -3030 1434 -3024
rect 1428 -3036 1434 -3030
rect 1428 -3042 1434 -3036
rect 1428 -3048 1434 -3042
rect 1428 -3054 1434 -3048
rect 1428 -3060 1434 -3054
rect 1428 -3066 1434 -3060
rect 1428 -3072 1434 -3066
rect 1428 -3078 1434 -3072
rect 1428 -3084 1434 -3078
rect 1428 -3090 1434 -3084
rect 1428 -3096 1434 -3090
rect 1428 -3102 1434 -3096
rect 1428 -3108 1434 -3102
rect 1428 -3114 1434 -3108
rect 1428 -3120 1434 -3114
rect 1428 -3126 1434 -3120
rect 1428 -3132 1434 -3126
rect 1428 -3138 1434 -3132
rect 1428 -3144 1434 -3138
rect 1428 -3150 1434 -3144
rect 1428 -3156 1434 -3150
rect 1428 -3162 1434 -3156
rect 1428 -3168 1434 -3162
rect 1428 -3174 1434 -3168
rect 1428 -3180 1434 -3174
rect 1428 -3186 1434 -3180
rect 1428 -3192 1434 -3186
rect 1428 -3198 1434 -3192
rect 1428 -3204 1434 -3198
rect 1428 -3210 1434 -3204
rect 1428 -3216 1434 -3210
rect 1428 -3222 1434 -3216
rect 1428 -3228 1434 -3222
rect 1428 -3234 1434 -3228
rect 1428 -3300 1434 -3294
rect 1428 -3306 1434 -3300
rect 1428 -3312 1434 -3306
rect 1428 -3318 1434 -3312
rect 1428 -3324 1434 -3318
rect 1428 -3330 1434 -3324
rect 1428 -3336 1434 -3330
rect 1428 -3342 1434 -3336
rect 1428 -3348 1434 -3342
rect 1428 -3354 1434 -3348
rect 1428 -3360 1434 -3354
rect 1428 -3366 1434 -3360
rect 1428 -3372 1434 -3366
rect 1428 -3378 1434 -3372
rect 1428 -3384 1434 -3378
rect 1428 -3390 1434 -3384
rect 1428 -3396 1434 -3390
rect 1428 -3402 1434 -3396
rect 1428 -3408 1434 -3402
rect 1428 -3414 1434 -3408
rect 1428 -3420 1434 -3414
rect 1428 -3426 1434 -3420
rect 1428 -3432 1434 -3426
rect 1428 -3438 1434 -3432
rect 1428 -3444 1434 -3438
rect 1428 -3450 1434 -3444
rect 1428 -3456 1434 -3450
rect 1428 -3462 1434 -3456
rect 1428 -3468 1434 -3462
rect 1428 -3474 1434 -3468
rect 1428 -3480 1434 -3474
rect 1428 -3486 1434 -3480
rect 1428 -3492 1434 -3486
rect 1428 -3498 1434 -3492
rect 1428 -3504 1434 -3498
rect 1434 -1122 1440 -1116
rect 1434 -1128 1440 -1122
rect 1434 -1134 1440 -1128
rect 1434 -1140 1440 -1134
rect 1434 -1146 1440 -1140
rect 1434 -1152 1440 -1146
rect 1434 -1158 1440 -1152
rect 1434 -1164 1440 -1158
rect 1434 -1170 1440 -1164
rect 1434 -1176 1440 -1170
rect 1434 -1182 1440 -1176
rect 1434 -1296 1440 -1290
rect 1434 -1302 1440 -1296
rect 1434 -1308 1440 -1302
rect 1434 -1314 1440 -1308
rect 1434 -1320 1440 -1314
rect 1434 -1326 1440 -1320
rect 1434 -1332 1440 -1326
rect 1434 -1338 1440 -1332
rect 1434 -1344 1440 -1338
rect 1434 -1350 1440 -1344
rect 1434 -1356 1440 -1350
rect 1434 -1362 1440 -1356
rect 1434 -1368 1440 -1362
rect 1434 -1374 1440 -1368
rect 1434 -1380 1440 -1374
rect 1434 -1386 1440 -1380
rect 1434 -1392 1440 -1386
rect 1434 -1398 1440 -1392
rect 1434 -1404 1440 -1398
rect 1434 -1410 1440 -1404
rect 1434 -1416 1440 -1410
rect 1434 -1422 1440 -1416
rect 1434 -1428 1440 -1422
rect 1434 -1434 1440 -1428
rect 1434 -1440 1440 -1434
rect 1434 -1446 1440 -1440
rect 1434 -1452 1440 -1446
rect 1434 -1458 1440 -1452
rect 1434 -1464 1440 -1458
rect 1434 -1470 1440 -1464
rect 1434 -1476 1440 -1470
rect 1434 -1482 1440 -1476
rect 1434 -1488 1440 -1482
rect 1434 -1494 1440 -1488
rect 1434 -1500 1440 -1494
rect 1434 -1506 1440 -1500
rect 1434 -1512 1440 -1506
rect 1434 -1518 1440 -1512
rect 1434 -1524 1440 -1518
rect 1434 -1530 1440 -1524
rect 1434 -1536 1440 -1530
rect 1434 -1542 1440 -1536
rect 1434 -1548 1440 -1542
rect 1434 -1554 1440 -1548
rect 1434 -1560 1440 -1554
rect 1434 -1566 1440 -1560
rect 1434 -1572 1440 -1566
rect 1434 -1578 1440 -1572
rect 1434 -1584 1440 -1578
rect 1434 -1590 1440 -1584
rect 1434 -1596 1440 -1590
rect 1434 -1602 1440 -1596
rect 1434 -1608 1440 -1602
rect 1434 -1614 1440 -1608
rect 1434 -1620 1440 -1614
rect 1434 -1626 1440 -1620
rect 1434 -1632 1440 -1626
rect 1434 -1638 1440 -1632
rect 1434 -1644 1440 -1638
rect 1434 -1650 1440 -1644
rect 1434 -1656 1440 -1650
rect 1434 -1662 1440 -1656
rect 1434 -1668 1440 -1662
rect 1434 -1674 1440 -1668
rect 1434 -1680 1440 -1674
rect 1434 -1686 1440 -1680
rect 1434 -1692 1440 -1686
rect 1434 -1698 1440 -1692
rect 1434 -1704 1440 -1698
rect 1434 -1710 1440 -1704
rect 1434 -1716 1440 -1710
rect 1434 -1722 1440 -1716
rect 1434 -1728 1440 -1722
rect 1434 -1734 1440 -1728
rect 1434 -1740 1440 -1734
rect 1434 -1746 1440 -1740
rect 1434 -1752 1440 -1746
rect 1434 -1758 1440 -1752
rect 1434 -1764 1440 -1758
rect 1434 -1770 1440 -1764
rect 1434 -1776 1440 -1770
rect 1434 -1782 1440 -1776
rect 1434 -1788 1440 -1782
rect 1434 -1794 1440 -1788
rect 1434 -1800 1440 -1794
rect 1434 -1806 1440 -1800
rect 1434 -1812 1440 -1806
rect 1434 -1818 1440 -1812
rect 1434 -1824 1440 -1818
rect 1434 -1830 1440 -1824
rect 1434 -1836 1440 -1830
rect 1434 -1842 1440 -1836
rect 1434 -1848 1440 -1842
rect 1434 -1854 1440 -1848
rect 1434 -1860 1440 -1854
rect 1434 -1866 1440 -1860
rect 1434 -1872 1440 -1866
rect 1434 -1878 1440 -1872
rect 1434 -1884 1440 -1878
rect 1434 -1890 1440 -1884
rect 1434 -1896 1440 -1890
rect 1434 -1902 1440 -1896
rect 1434 -1908 1440 -1902
rect 1434 -1914 1440 -1908
rect 1434 -1920 1440 -1914
rect 1434 -1926 1440 -1920
rect 1434 -1932 1440 -1926
rect 1434 -1938 1440 -1932
rect 1434 -1944 1440 -1938
rect 1434 -1950 1440 -1944
rect 1434 -1956 1440 -1950
rect 1434 -1962 1440 -1956
rect 1434 -1968 1440 -1962
rect 1434 -1974 1440 -1968
rect 1434 -1980 1440 -1974
rect 1434 -1986 1440 -1980
rect 1434 -1992 1440 -1986
rect 1434 -1998 1440 -1992
rect 1434 -2004 1440 -1998
rect 1434 -2010 1440 -2004
rect 1434 -2016 1440 -2010
rect 1434 -2022 1440 -2016
rect 1434 -2028 1440 -2022
rect 1434 -2034 1440 -2028
rect 1434 -2040 1440 -2034
rect 1434 -2046 1440 -2040
rect 1434 -2052 1440 -2046
rect 1434 -2058 1440 -2052
rect 1434 -2064 1440 -2058
rect 1434 -2070 1440 -2064
rect 1434 -2076 1440 -2070
rect 1434 -2082 1440 -2076
rect 1434 -2088 1440 -2082
rect 1434 -2094 1440 -2088
rect 1434 -2100 1440 -2094
rect 1434 -2106 1440 -2100
rect 1434 -2112 1440 -2106
rect 1434 -2118 1440 -2112
rect 1434 -2124 1440 -2118
rect 1434 -2130 1440 -2124
rect 1434 -2136 1440 -2130
rect 1434 -2142 1440 -2136
rect 1434 -2148 1440 -2142
rect 1434 -2154 1440 -2148
rect 1434 -2160 1440 -2154
rect 1434 -2166 1440 -2160
rect 1434 -2172 1440 -2166
rect 1434 -2178 1440 -2172
rect 1434 -2184 1440 -2178
rect 1434 -2190 1440 -2184
rect 1434 -2196 1440 -2190
rect 1434 -2202 1440 -2196
rect 1434 -2208 1440 -2202
rect 1434 -2214 1440 -2208
rect 1434 -2220 1440 -2214
rect 1434 -2226 1440 -2220
rect 1434 -2232 1440 -2226
rect 1434 -2238 1440 -2232
rect 1434 -2244 1440 -2238
rect 1434 -2250 1440 -2244
rect 1434 -2256 1440 -2250
rect 1434 -2262 1440 -2256
rect 1434 -2268 1440 -2262
rect 1434 -2274 1440 -2268
rect 1434 -2352 1440 -2346
rect 1434 -2358 1440 -2352
rect 1434 -2364 1440 -2358
rect 1434 -2370 1440 -2364
rect 1434 -2376 1440 -2370
rect 1434 -2382 1440 -2376
rect 1434 -2388 1440 -2382
rect 1434 -2394 1440 -2388
rect 1434 -2400 1440 -2394
rect 1434 -2406 1440 -2400
rect 1434 -2412 1440 -2406
rect 1434 -2418 1440 -2412
rect 1434 -2424 1440 -2418
rect 1434 -2430 1440 -2424
rect 1434 -2436 1440 -2430
rect 1434 -2442 1440 -2436
rect 1434 -2448 1440 -2442
rect 1434 -2454 1440 -2448
rect 1434 -2460 1440 -2454
rect 1434 -2466 1440 -2460
rect 1434 -2472 1440 -2466
rect 1434 -2478 1440 -2472
rect 1434 -2484 1440 -2478
rect 1434 -2490 1440 -2484
rect 1434 -2496 1440 -2490
rect 1434 -2502 1440 -2496
rect 1434 -2508 1440 -2502
rect 1434 -2514 1440 -2508
rect 1434 -2520 1440 -2514
rect 1434 -2526 1440 -2520
rect 1434 -2532 1440 -2526
rect 1434 -2538 1440 -2532
rect 1434 -2544 1440 -2538
rect 1434 -2550 1440 -2544
rect 1434 -2556 1440 -2550
rect 1434 -2562 1440 -2556
rect 1434 -2568 1440 -2562
rect 1434 -2574 1440 -2568
rect 1434 -2580 1440 -2574
rect 1434 -2586 1440 -2580
rect 1434 -2592 1440 -2586
rect 1434 -2598 1440 -2592
rect 1434 -2604 1440 -2598
rect 1434 -2610 1440 -2604
rect 1434 -2616 1440 -2610
rect 1434 -2622 1440 -2616
rect 1434 -2628 1440 -2622
rect 1434 -2634 1440 -2628
rect 1434 -2640 1440 -2634
rect 1434 -2646 1440 -2640
rect 1434 -2652 1440 -2646
rect 1434 -2658 1440 -2652
rect 1434 -2664 1440 -2658
rect 1434 -2670 1440 -2664
rect 1434 -2676 1440 -2670
rect 1434 -2682 1440 -2676
rect 1434 -2688 1440 -2682
rect 1434 -2694 1440 -2688
rect 1434 -2700 1440 -2694
rect 1434 -2706 1440 -2700
rect 1434 -2712 1440 -2706
rect 1434 -2718 1440 -2712
rect 1434 -2724 1440 -2718
rect 1434 -2730 1440 -2724
rect 1434 -2736 1440 -2730
rect 1434 -2742 1440 -2736
rect 1434 -2748 1440 -2742
rect 1434 -2754 1440 -2748
rect 1434 -2760 1440 -2754
rect 1434 -2766 1440 -2760
rect 1434 -2772 1440 -2766
rect 1434 -2778 1440 -2772
rect 1434 -2784 1440 -2778
rect 1434 -2790 1440 -2784
rect 1434 -2796 1440 -2790
rect 1434 -2802 1440 -2796
rect 1434 -2808 1440 -2802
rect 1434 -2814 1440 -2808
rect 1434 -2820 1440 -2814
rect 1434 -2826 1440 -2820
rect 1434 -2832 1440 -2826
rect 1434 -2838 1440 -2832
rect 1434 -2844 1440 -2838
rect 1434 -2850 1440 -2844
rect 1434 -2940 1440 -2934
rect 1434 -2946 1440 -2940
rect 1434 -2952 1440 -2946
rect 1434 -2958 1440 -2952
rect 1434 -2964 1440 -2958
rect 1434 -2970 1440 -2964
rect 1434 -2976 1440 -2970
rect 1434 -2982 1440 -2976
rect 1434 -2988 1440 -2982
rect 1434 -2994 1440 -2988
rect 1434 -3000 1440 -2994
rect 1434 -3006 1440 -3000
rect 1434 -3012 1440 -3006
rect 1434 -3018 1440 -3012
rect 1434 -3024 1440 -3018
rect 1434 -3030 1440 -3024
rect 1434 -3036 1440 -3030
rect 1434 -3042 1440 -3036
rect 1434 -3048 1440 -3042
rect 1434 -3054 1440 -3048
rect 1434 -3060 1440 -3054
rect 1434 -3066 1440 -3060
rect 1434 -3072 1440 -3066
rect 1434 -3078 1440 -3072
rect 1434 -3084 1440 -3078
rect 1434 -3090 1440 -3084
rect 1434 -3096 1440 -3090
rect 1434 -3102 1440 -3096
rect 1434 -3108 1440 -3102
rect 1434 -3114 1440 -3108
rect 1434 -3120 1440 -3114
rect 1434 -3126 1440 -3120
rect 1434 -3132 1440 -3126
rect 1434 -3138 1440 -3132
rect 1434 -3144 1440 -3138
rect 1434 -3150 1440 -3144
rect 1434 -3156 1440 -3150
rect 1434 -3162 1440 -3156
rect 1434 -3168 1440 -3162
rect 1434 -3174 1440 -3168
rect 1434 -3180 1440 -3174
rect 1434 -3186 1440 -3180
rect 1434 -3192 1440 -3186
rect 1434 -3198 1440 -3192
rect 1434 -3204 1440 -3198
rect 1434 -3210 1440 -3204
rect 1434 -3216 1440 -3210
rect 1434 -3222 1440 -3216
rect 1434 -3228 1440 -3222
rect 1434 -3234 1440 -3228
rect 1434 -3300 1440 -3294
rect 1434 -3306 1440 -3300
rect 1434 -3312 1440 -3306
rect 1434 -3318 1440 -3312
rect 1434 -3324 1440 -3318
rect 1434 -3330 1440 -3324
rect 1434 -3336 1440 -3330
rect 1434 -3342 1440 -3336
rect 1434 -3348 1440 -3342
rect 1434 -3354 1440 -3348
rect 1434 -3360 1440 -3354
rect 1434 -3366 1440 -3360
rect 1434 -3372 1440 -3366
rect 1434 -3378 1440 -3372
rect 1434 -3384 1440 -3378
rect 1434 -3390 1440 -3384
rect 1434 -3396 1440 -3390
rect 1434 -3402 1440 -3396
rect 1434 -3408 1440 -3402
rect 1434 -3414 1440 -3408
rect 1434 -3420 1440 -3414
rect 1434 -3426 1440 -3420
rect 1434 -3432 1440 -3426
rect 1434 -3438 1440 -3432
rect 1434 -3444 1440 -3438
rect 1434 -3450 1440 -3444
rect 1434 -3456 1440 -3450
rect 1434 -3462 1440 -3456
rect 1434 -3468 1440 -3462
rect 1434 -3474 1440 -3468
rect 1434 -3480 1440 -3474
rect 1434 -3486 1440 -3480
rect 1434 -3492 1440 -3486
rect 1434 -3498 1440 -3492
rect 1434 -3504 1440 -3498
rect 1440 -1122 1446 -1116
rect 1440 -1128 1446 -1122
rect 1440 -1134 1446 -1128
rect 1440 -1140 1446 -1134
rect 1440 -1146 1446 -1140
rect 1440 -1152 1446 -1146
rect 1440 -1158 1446 -1152
rect 1440 -1164 1446 -1158
rect 1440 -1170 1446 -1164
rect 1440 -1290 1446 -1284
rect 1440 -1296 1446 -1290
rect 1440 -1302 1446 -1296
rect 1440 -1308 1446 -1302
rect 1440 -1314 1446 -1308
rect 1440 -1320 1446 -1314
rect 1440 -1326 1446 -1320
rect 1440 -1332 1446 -1326
rect 1440 -1338 1446 -1332
rect 1440 -1344 1446 -1338
rect 1440 -1350 1446 -1344
rect 1440 -1356 1446 -1350
rect 1440 -1362 1446 -1356
rect 1440 -1368 1446 -1362
rect 1440 -1374 1446 -1368
rect 1440 -1380 1446 -1374
rect 1440 -1386 1446 -1380
rect 1440 -1392 1446 -1386
rect 1440 -1398 1446 -1392
rect 1440 -1404 1446 -1398
rect 1440 -1410 1446 -1404
rect 1440 -1416 1446 -1410
rect 1440 -1422 1446 -1416
rect 1440 -1428 1446 -1422
rect 1440 -1434 1446 -1428
rect 1440 -1440 1446 -1434
rect 1440 -1446 1446 -1440
rect 1440 -1452 1446 -1446
rect 1440 -1458 1446 -1452
rect 1440 -1464 1446 -1458
rect 1440 -1470 1446 -1464
rect 1440 -1476 1446 -1470
rect 1440 -1482 1446 -1476
rect 1440 -1488 1446 -1482
rect 1440 -1494 1446 -1488
rect 1440 -1500 1446 -1494
rect 1440 -1506 1446 -1500
rect 1440 -1512 1446 -1506
rect 1440 -1518 1446 -1512
rect 1440 -1524 1446 -1518
rect 1440 -1530 1446 -1524
rect 1440 -1536 1446 -1530
rect 1440 -1542 1446 -1536
rect 1440 -1548 1446 -1542
rect 1440 -1554 1446 -1548
rect 1440 -1560 1446 -1554
rect 1440 -1566 1446 -1560
rect 1440 -1572 1446 -1566
rect 1440 -1578 1446 -1572
rect 1440 -1584 1446 -1578
rect 1440 -1590 1446 -1584
rect 1440 -1596 1446 -1590
rect 1440 -1602 1446 -1596
rect 1440 -1608 1446 -1602
rect 1440 -1614 1446 -1608
rect 1440 -1620 1446 -1614
rect 1440 -1626 1446 -1620
rect 1440 -1632 1446 -1626
rect 1440 -1638 1446 -1632
rect 1440 -1644 1446 -1638
rect 1440 -1650 1446 -1644
rect 1440 -1656 1446 -1650
rect 1440 -1662 1446 -1656
rect 1440 -1668 1446 -1662
rect 1440 -1674 1446 -1668
rect 1440 -1680 1446 -1674
rect 1440 -1686 1446 -1680
rect 1440 -1692 1446 -1686
rect 1440 -1698 1446 -1692
rect 1440 -1704 1446 -1698
rect 1440 -1710 1446 -1704
rect 1440 -1716 1446 -1710
rect 1440 -1722 1446 -1716
rect 1440 -1728 1446 -1722
rect 1440 -1734 1446 -1728
rect 1440 -1740 1446 -1734
rect 1440 -1746 1446 -1740
rect 1440 -1752 1446 -1746
rect 1440 -1758 1446 -1752
rect 1440 -1764 1446 -1758
rect 1440 -1770 1446 -1764
rect 1440 -1776 1446 -1770
rect 1440 -1782 1446 -1776
rect 1440 -1788 1446 -1782
rect 1440 -1794 1446 -1788
rect 1440 -1800 1446 -1794
rect 1440 -1806 1446 -1800
rect 1440 -1812 1446 -1806
rect 1440 -1818 1446 -1812
rect 1440 -1824 1446 -1818
rect 1440 -1830 1446 -1824
rect 1440 -1836 1446 -1830
rect 1440 -1842 1446 -1836
rect 1440 -1848 1446 -1842
rect 1440 -1854 1446 -1848
rect 1440 -1860 1446 -1854
rect 1440 -1866 1446 -1860
rect 1440 -1872 1446 -1866
rect 1440 -1878 1446 -1872
rect 1440 -1884 1446 -1878
rect 1440 -1890 1446 -1884
rect 1440 -1896 1446 -1890
rect 1440 -1902 1446 -1896
rect 1440 -1908 1446 -1902
rect 1440 -1914 1446 -1908
rect 1440 -1920 1446 -1914
rect 1440 -1926 1446 -1920
rect 1440 -1932 1446 -1926
rect 1440 -1938 1446 -1932
rect 1440 -1944 1446 -1938
rect 1440 -1950 1446 -1944
rect 1440 -1956 1446 -1950
rect 1440 -1962 1446 -1956
rect 1440 -1968 1446 -1962
rect 1440 -1974 1446 -1968
rect 1440 -1980 1446 -1974
rect 1440 -1986 1446 -1980
rect 1440 -1992 1446 -1986
rect 1440 -1998 1446 -1992
rect 1440 -2004 1446 -1998
rect 1440 -2010 1446 -2004
rect 1440 -2016 1446 -2010
rect 1440 -2022 1446 -2016
rect 1440 -2028 1446 -2022
rect 1440 -2034 1446 -2028
rect 1440 -2040 1446 -2034
rect 1440 -2046 1446 -2040
rect 1440 -2052 1446 -2046
rect 1440 -2058 1446 -2052
rect 1440 -2064 1446 -2058
rect 1440 -2070 1446 -2064
rect 1440 -2076 1446 -2070
rect 1440 -2082 1446 -2076
rect 1440 -2088 1446 -2082
rect 1440 -2094 1446 -2088
rect 1440 -2100 1446 -2094
rect 1440 -2106 1446 -2100
rect 1440 -2112 1446 -2106
rect 1440 -2118 1446 -2112
rect 1440 -2124 1446 -2118
rect 1440 -2130 1446 -2124
rect 1440 -2136 1446 -2130
rect 1440 -2142 1446 -2136
rect 1440 -2148 1446 -2142
rect 1440 -2154 1446 -2148
rect 1440 -2160 1446 -2154
rect 1440 -2166 1446 -2160
rect 1440 -2172 1446 -2166
rect 1440 -2178 1446 -2172
rect 1440 -2184 1446 -2178
rect 1440 -2190 1446 -2184
rect 1440 -2196 1446 -2190
rect 1440 -2202 1446 -2196
rect 1440 -2208 1446 -2202
rect 1440 -2214 1446 -2208
rect 1440 -2220 1446 -2214
rect 1440 -2226 1446 -2220
rect 1440 -2232 1446 -2226
rect 1440 -2238 1446 -2232
rect 1440 -2244 1446 -2238
rect 1440 -2250 1446 -2244
rect 1440 -2256 1446 -2250
rect 1440 -2262 1446 -2256
rect 1440 -2268 1446 -2262
rect 1440 -2346 1446 -2340
rect 1440 -2352 1446 -2346
rect 1440 -2358 1446 -2352
rect 1440 -2364 1446 -2358
rect 1440 -2370 1446 -2364
rect 1440 -2376 1446 -2370
rect 1440 -2382 1446 -2376
rect 1440 -2388 1446 -2382
rect 1440 -2394 1446 -2388
rect 1440 -2400 1446 -2394
rect 1440 -2406 1446 -2400
rect 1440 -2412 1446 -2406
rect 1440 -2418 1446 -2412
rect 1440 -2424 1446 -2418
rect 1440 -2430 1446 -2424
rect 1440 -2436 1446 -2430
rect 1440 -2442 1446 -2436
rect 1440 -2448 1446 -2442
rect 1440 -2454 1446 -2448
rect 1440 -2460 1446 -2454
rect 1440 -2466 1446 -2460
rect 1440 -2472 1446 -2466
rect 1440 -2478 1446 -2472
rect 1440 -2484 1446 -2478
rect 1440 -2490 1446 -2484
rect 1440 -2496 1446 -2490
rect 1440 -2502 1446 -2496
rect 1440 -2508 1446 -2502
rect 1440 -2514 1446 -2508
rect 1440 -2520 1446 -2514
rect 1440 -2526 1446 -2520
rect 1440 -2532 1446 -2526
rect 1440 -2538 1446 -2532
rect 1440 -2544 1446 -2538
rect 1440 -2550 1446 -2544
rect 1440 -2556 1446 -2550
rect 1440 -2562 1446 -2556
rect 1440 -2568 1446 -2562
rect 1440 -2574 1446 -2568
rect 1440 -2580 1446 -2574
rect 1440 -2586 1446 -2580
rect 1440 -2592 1446 -2586
rect 1440 -2598 1446 -2592
rect 1440 -2604 1446 -2598
rect 1440 -2610 1446 -2604
rect 1440 -2616 1446 -2610
rect 1440 -2622 1446 -2616
rect 1440 -2628 1446 -2622
rect 1440 -2634 1446 -2628
rect 1440 -2640 1446 -2634
rect 1440 -2646 1446 -2640
rect 1440 -2652 1446 -2646
rect 1440 -2658 1446 -2652
rect 1440 -2664 1446 -2658
rect 1440 -2670 1446 -2664
rect 1440 -2676 1446 -2670
rect 1440 -2682 1446 -2676
rect 1440 -2688 1446 -2682
rect 1440 -2694 1446 -2688
rect 1440 -2700 1446 -2694
rect 1440 -2706 1446 -2700
rect 1440 -2712 1446 -2706
rect 1440 -2718 1446 -2712
rect 1440 -2724 1446 -2718
rect 1440 -2730 1446 -2724
rect 1440 -2736 1446 -2730
rect 1440 -2742 1446 -2736
rect 1440 -2748 1446 -2742
rect 1440 -2754 1446 -2748
rect 1440 -2760 1446 -2754
rect 1440 -2766 1446 -2760
rect 1440 -2772 1446 -2766
rect 1440 -2778 1446 -2772
rect 1440 -2784 1446 -2778
rect 1440 -2790 1446 -2784
rect 1440 -2796 1446 -2790
rect 1440 -2802 1446 -2796
rect 1440 -2808 1446 -2802
rect 1440 -2814 1446 -2808
rect 1440 -2820 1446 -2814
rect 1440 -2826 1446 -2820
rect 1440 -2832 1446 -2826
rect 1440 -2838 1446 -2832
rect 1440 -2844 1446 -2838
rect 1440 -2850 1446 -2844
rect 1440 -2934 1446 -2928
rect 1440 -2940 1446 -2934
rect 1440 -2946 1446 -2940
rect 1440 -2952 1446 -2946
rect 1440 -2958 1446 -2952
rect 1440 -2964 1446 -2958
rect 1440 -2970 1446 -2964
rect 1440 -2976 1446 -2970
rect 1440 -2982 1446 -2976
rect 1440 -2988 1446 -2982
rect 1440 -2994 1446 -2988
rect 1440 -3000 1446 -2994
rect 1440 -3006 1446 -3000
rect 1440 -3012 1446 -3006
rect 1440 -3018 1446 -3012
rect 1440 -3024 1446 -3018
rect 1440 -3030 1446 -3024
rect 1440 -3036 1446 -3030
rect 1440 -3042 1446 -3036
rect 1440 -3048 1446 -3042
rect 1440 -3054 1446 -3048
rect 1440 -3060 1446 -3054
rect 1440 -3066 1446 -3060
rect 1440 -3072 1446 -3066
rect 1440 -3078 1446 -3072
rect 1440 -3084 1446 -3078
rect 1440 -3090 1446 -3084
rect 1440 -3096 1446 -3090
rect 1440 -3102 1446 -3096
rect 1440 -3108 1446 -3102
rect 1440 -3114 1446 -3108
rect 1440 -3120 1446 -3114
rect 1440 -3126 1446 -3120
rect 1440 -3132 1446 -3126
rect 1440 -3138 1446 -3132
rect 1440 -3144 1446 -3138
rect 1440 -3150 1446 -3144
rect 1440 -3156 1446 -3150
rect 1440 -3162 1446 -3156
rect 1440 -3168 1446 -3162
rect 1440 -3174 1446 -3168
rect 1440 -3180 1446 -3174
rect 1440 -3186 1446 -3180
rect 1440 -3192 1446 -3186
rect 1440 -3198 1446 -3192
rect 1440 -3204 1446 -3198
rect 1440 -3210 1446 -3204
rect 1440 -3216 1446 -3210
rect 1440 -3222 1446 -3216
rect 1440 -3228 1446 -3222
rect 1440 -3234 1446 -3228
rect 1440 -3294 1446 -3288
rect 1440 -3300 1446 -3294
rect 1440 -3306 1446 -3300
rect 1440 -3312 1446 -3306
rect 1440 -3318 1446 -3312
rect 1440 -3324 1446 -3318
rect 1440 -3330 1446 -3324
rect 1440 -3336 1446 -3330
rect 1440 -3342 1446 -3336
rect 1440 -3348 1446 -3342
rect 1440 -3354 1446 -3348
rect 1440 -3360 1446 -3354
rect 1440 -3366 1446 -3360
rect 1440 -3372 1446 -3366
rect 1440 -3378 1446 -3372
rect 1440 -3384 1446 -3378
rect 1440 -3390 1446 -3384
rect 1440 -3396 1446 -3390
rect 1440 -3402 1446 -3396
rect 1440 -3408 1446 -3402
rect 1440 -3414 1446 -3408
rect 1440 -3420 1446 -3414
rect 1440 -3426 1446 -3420
rect 1440 -3432 1446 -3426
rect 1440 -3438 1446 -3432
rect 1440 -3444 1446 -3438
rect 1440 -3450 1446 -3444
rect 1440 -3456 1446 -3450
rect 1440 -3462 1446 -3456
rect 1440 -3468 1446 -3462
rect 1440 -3474 1446 -3468
rect 1440 -3480 1446 -3474
rect 1440 -3486 1446 -3480
rect 1440 -3492 1446 -3486
rect 1440 -3498 1446 -3492
rect 1440 -3504 1446 -3498
rect 1446 -1122 1452 -1116
rect 1446 -1128 1452 -1122
rect 1446 -1134 1452 -1128
rect 1446 -1140 1452 -1134
rect 1446 -1146 1452 -1140
rect 1446 -1152 1452 -1146
rect 1446 -1158 1452 -1152
rect 1446 -1164 1452 -1158
rect 1446 -1278 1452 -1272
rect 1446 -1284 1452 -1278
rect 1446 -1290 1452 -1284
rect 1446 -1296 1452 -1290
rect 1446 -1302 1452 -1296
rect 1446 -1308 1452 -1302
rect 1446 -1314 1452 -1308
rect 1446 -1320 1452 -1314
rect 1446 -1326 1452 -1320
rect 1446 -1332 1452 -1326
rect 1446 -1338 1452 -1332
rect 1446 -1344 1452 -1338
rect 1446 -1350 1452 -1344
rect 1446 -1356 1452 -1350
rect 1446 -1362 1452 -1356
rect 1446 -1368 1452 -1362
rect 1446 -1374 1452 -1368
rect 1446 -1380 1452 -1374
rect 1446 -1386 1452 -1380
rect 1446 -1392 1452 -1386
rect 1446 -1398 1452 -1392
rect 1446 -1404 1452 -1398
rect 1446 -1410 1452 -1404
rect 1446 -1416 1452 -1410
rect 1446 -1422 1452 -1416
rect 1446 -1428 1452 -1422
rect 1446 -1434 1452 -1428
rect 1446 -1440 1452 -1434
rect 1446 -1446 1452 -1440
rect 1446 -1452 1452 -1446
rect 1446 -1458 1452 -1452
rect 1446 -1464 1452 -1458
rect 1446 -1470 1452 -1464
rect 1446 -1476 1452 -1470
rect 1446 -1482 1452 -1476
rect 1446 -1488 1452 -1482
rect 1446 -1494 1452 -1488
rect 1446 -1500 1452 -1494
rect 1446 -1506 1452 -1500
rect 1446 -1512 1452 -1506
rect 1446 -1518 1452 -1512
rect 1446 -1524 1452 -1518
rect 1446 -1530 1452 -1524
rect 1446 -1536 1452 -1530
rect 1446 -1542 1452 -1536
rect 1446 -1548 1452 -1542
rect 1446 -1554 1452 -1548
rect 1446 -1560 1452 -1554
rect 1446 -1566 1452 -1560
rect 1446 -1572 1452 -1566
rect 1446 -1578 1452 -1572
rect 1446 -1584 1452 -1578
rect 1446 -1590 1452 -1584
rect 1446 -1596 1452 -1590
rect 1446 -1602 1452 -1596
rect 1446 -1608 1452 -1602
rect 1446 -1614 1452 -1608
rect 1446 -1620 1452 -1614
rect 1446 -1626 1452 -1620
rect 1446 -1632 1452 -1626
rect 1446 -1638 1452 -1632
rect 1446 -1644 1452 -1638
rect 1446 -1650 1452 -1644
rect 1446 -1656 1452 -1650
rect 1446 -1662 1452 -1656
rect 1446 -1668 1452 -1662
rect 1446 -1674 1452 -1668
rect 1446 -1680 1452 -1674
rect 1446 -1686 1452 -1680
rect 1446 -1692 1452 -1686
rect 1446 -1698 1452 -1692
rect 1446 -1704 1452 -1698
rect 1446 -1710 1452 -1704
rect 1446 -1716 1452 -1710
rect 1446 -1722 1452 -1716
rect 1446 -1728 1452 -1722
rect 1446 -1734 1452 -1728
rect 1446 -1740 1452 -1734
rect 1446 -1746 1452 -1740
rect 1446 -1752 1452 -1746
rect 1446 -1758 1452 -1752
rect 1446 -1764 1452 -1758
rect 1446 -1770 1452 -1764
rect 1446 -1776 1452 -1770
rect 1446 -1782 1452 -1776
rect 1446 -1788 1452 -1782
rect 1446 -1794 1452 -1788
rect 1446 -1800 1452 -1794
rect 1446 -1806 1452 -1800
rect 1446 -1812 1452 -1806
rect 1446 -1818 1452 -1812
rect 1446 -1824 1452 -1818
rect 1446 -1830 1452 -1824
rect 1446 -1836 1452 -1830
rect 1446 -1842 1452 -1836
rect 1446 -1848 1452 -1842
rect 1446 -1854 1452 -1848
rect 1446 -1860 1452 -1854
rect 1446 -1866 1452 -1860
rect 1446 -1872 1452 -1866
rect 1446 -1878 1452 -1872
rect 1446 -1884 1452 -1878
rect 1446 -1890 1452 -1884
rect 1446 -1896 1452 -1890
rect 1446 -1902 1452 -1896
rect 1446 -1908 1452 -1902
rect 1446 -1914 1452 -1908
rect 1446 -1920 1452 -1914
rect 1446 -1926 1452 -1920
rect 1446 -1932 1452 -1926
rect 1446 -1938 1452 -1932
rect 1446 -1944 1452 -1938
rect 1446 -1950 1452 -1944
rect 1446 -1956 1452 -1950
rect 1446 -1962 1452 -1956
rect 1446 -1968 1452 -1962
rect 1446 -1974 1452 -1968
rect 1446 -1980 1452 -1974
rect 1446 -1986 1452 -1980
rect 1446 -1992 1452 -1986
rect 1446 -1998 1452 -1992
rect 1446 -2004 1452 -1998
rect 1446 -2010 1452 -2004
rect 1446 -2016 1452 -2010
rect 1446 -2022 1452 -2016
rect 1446 -2028 1452 -2022
rect 1446 -2034 1452 -2028
rect 1446 -2040 1452 -2034
rect 1446 -2046 1452 -2040
rect 1446 -2052 1452 -2046
rect 1446 -2058 1452 -2052
rect 1446 -2064 1452 -2058
rect 1446 -2070 1452 -2064
rect 1446 -2076 1452 -2070
rect 1446 -2082 1452 -2076
rect 1446 -2088 1452 -2082
rect 1446 -2094 1452 -2088
rect 1446 -2100 1452 -2094
rect 1446 -2106 1452 -2100
rect 1446 -2112 1452 -2106
rect 1446 -2118 1452 -2112
rect 1446 -2124 1452 -2118
rect 1446 -2130 1452 -2124
rect 1446 -2136 1452 -2130
rect 1446 -2142 1452 -2136
rect 1446 -2148 1452 -2142
rect 1446 -2154 1452 -2148
rect 1446 -2160 1452 -2154
rect 1446 -2166 1452 -2160
rect 1446 -2172 1452 -2166
rect 1446 -2178 1452 -2172
rect 1446 -2184 1452 -2178
rect 1446 -2190 1452 -2184
rect 1446 -2196 1452 -2190
rect 1446 -2202 1452 -2196
rect 1446 -2208 1452 -2202
rect 1446 -2214 1452 -2208
rect 1446 -2220 1452 -2214
rect 1446 -2226 1452 -2220
rect 1446 -2232 1452 -2226
rect 1446 -2238 1452 -2232
rect 1446 -2244 1452 -2238
rect 1446 -2250 1452 -2244
rect 1446 -2256 1452 -2250
rect 1446 -2262 1452 -2256
rect 1446 -2334 1452 -2328
rect 1446 -2340 1452 -2334
rect 1446 -2346 1452 -2340
rect 1446 -2352 1452 -2346
rect 1446 -2358 1452 -2352
rect 1446 -2364 1452 -2358
rect 1446 -2370 1452 -2364
rect 1446 -2376 1452 -2370
rect 1446 -2382 1452 -2376
rect 1446 -2388 1452 -2382
rect 1446 -2394 1452 -2388
rect 1446 -2400 1452 -2394
rect 1446 -2406 1452 -2400
rect 1446 -2412 1452 -2406
rect 1446 -2418 1452 -2412
rect 1446 -2424 1452 -2418
rect 1446 -2430 1452 -2424
rect 1446 -2436 1452 -2430
rect 1446 -2442 1452 -2436
rect 1446 -2448 1452 -2442
rect 1446 -2454 1452 -2448
rect 1446 -2460 1452 -2454
rect 1446 -2466 1452 -2460
rect 1446 -2472 1452 -2466
rect 1446 -2478 1452 -2472
rect 1446 -2484 1452 -2478
rect 1446 -2490 1452 -2484
rect 1446 -2496 1452 -2490
rect 1446 -2502 1452 -2496
rect 1446 -2508 1452 -2502
rect 1446 -2514 1452 -2508
rect 1446 -2520 1452 -2514
rect 1446 -2526 1452 -2520
rect 1446 -2532 1452 -2526
rect 1446 -2538 1452 -2532
rect 1446 -2544 1452 -2538
rect 1446 -2550 1452 -2544
rect 1446 -2556 1452 -2550
rect 1446 -2562 1452 -2556
rect 1446 -2568 1452 -2562
rect 1446 -2574 1452 -2568
rect 1446 -2580 1452 -2574
rect 1446 -2586 1452 -2580
rect 1446 -2592 1452 -2586
rect 1446 -2598 1452 -2592
rect 1446 -2604 1452 -2598
rect 1446 -2610 1452 -2604
rect 1446 -2616 1452 -2610
rect 1446 -2622 1452 -2616
rect 1446 -2628 1452 -2622
rect 1446 -2634 1452 -2628
rect 1446 -2640 1452 -2634
rect 1446 -2646 1452 -2640
rect 1446 -2652 1452 -2646
rect 1446 -2658 1452 -2652
rect 1446 -2664 1452 -2658
rect 1446 -2670 1452 -2664
rect 1446 -2676 1452 -2670
rect 1446 -2682 1452 -2676
rect 1446 -2688 1452 -2682
rect 1446 -2694 1452 -2688
rect 1446 -2700 1452 -2694
rect 1446 -2706 1452 -2700
rect 1446 -2712 1452 -2706
rect 1446 -2718 1452 -2712
rect 1446 -2724 1452 -2718
rect 1446 -2730 1452 -2724
rect 1446 -2736 1452 -2730
rect 1446 -2742 1452 -2736
rect 1446 -2748 1452 -2742
rect 1446 -2754 1452 -2748
rect 1446 -2760 1452 -2754
rect 1446 -2766 1452 -2760
rect 1446 -2772 1452 -2766
rect 1446 -2778 1452 -2772
rect 1446 -2784 1452 -2778
rect 1446 -2790 1452 -2784
rect 1446 -2796 1452 -2790
rect 1446 -2802 1452 -2796
rect 1446 -2808 1452 -2802
rect 1446 -2814 1452 -2808
rect 1446 -2820 1452 -2814
rect 1446 -2826 1452 -2820
rect 1446 -2832 1452 -2826
rect 1446 -2838 1452 -2832
rect 1446 -2844 1452 -2838
rect 1446 -2928 1452 -2922
rect 1446 -2934 1452 -2928
rect 1446 -2940 1452 -2934
rect 1446 -2946 1452 -2940
rect 1446 -2952 1452 -2946
rect 1446 -2958 1452 -2952
rect 1446 -2964 1452 -2958
rect 1446 -2970 1452 -2964
rect 1446 -2976 1452 -2970
rect 1446 -2982 1452 -2976
rect 1446 -2988 1452 -2982
rect 1446 -2994 1452 -2988
rect 1446 -3000 1452 -2994
rect 1446 -3006 1452 -3000
rect 1446 -3012 1452 -3006
rect 1446 -3018 1452 -3012
rect 1446 -3024 1452 -3018
rect 1446 -3030 1452 -3024
rect 1446 -3036 1452 -3030
rect 1446 -3042 1452 -3036
rect 1446 -3048 1452 -3042
rect 1446 -3054 1452 -3048
rect 1446 -3060 1452 -3054
rect 1446 -3066 1452 -3060
rect 1446 -3072 1452 -3066
rect 1446 -3078 1452 -3072
rect 1446 -3084 1452 -3078
rect 1446 -3090 1452 -3084
rect 1446 -3096 1452 -3090
rect 1446 -3102 1452 -3096
rect 1446 -3108 1452 -3102
rect 1446 -3114 1452 -3108
rect 1446 -3120 1452 -3114
rect 1446 -3126 1452 -3120
rect 1446 -3132 1452 -3126
rect 1446 -3138 1452 -3132
rect 1446 -3144 1452 -3138
rect 1446 -3150 1452 -3144
rect 1446 -3156 1452 -3150
rect 1446 -3162 1452 -3156
rect 1446 -3168 1452 -3162
rect 1446 -3174 1452 -3168
rect 1446 -3180 1452 -3174
rect 1446 -3186 1452 -3180
rect 1446 -3192 1452 -3186
rect 1446 -3198 1452 -3192
rect 1446 -3204 1452 -3198
rect 1446 -3210 1452 -3204
rect 1446 -3216 1452 -3210
rect 1446 -3222 1452 -3216
rect 1446 -3228 1452 -3222
rect 1446 -3234 1452 -3228
rect 1446 -3294 1452 -3288
rect 1446 -3300 1452 -3294
rect 1446 -3306 1452 -3300
rect 1446 -3312 1452 -3306
rect 1446 -3318 1452 -3312
rect 1446 -3324 1452 -3318
rect 1446 -3330 1452 -3324
rect 1446 -3336 1452 -3330
rect 1446 -3342 1452 -3336
rect 1446 -3348 1452 -3342
rect 1446 -3354 1452 -3348
rect 1446 -3360 1452 -3354
rect 1446 -3366 1452 -3360
rect 1446 -3372 1452 -3366
rect 1446 -3378 1452 -3372
rect 1446 -3384 1452 -3378
rect 1446 -3390 1452 -3384
rect 1446 -3396 1452 -3390
rect 1446 -3402 1452 -3396
rect 1446 -3408 1452 -3402
rect 1446 -3414 1452 -3408
rect 1446 -3420 1452 -3414
rect 1446 -3426 1452 -3420
rect 1446 -3432 1452 -3426
rect 1446 -3438 1452 -3432
rect 1446 -3444 1452 -3438
rect 1446 -3450 1452 -3444
rect 1446 -3456 1452 -3450
rect 1446 -3462 1452 -3456
rect 1446 -3468 1452 -3462
rect 1446 -3474 1452 -3468
rect 1446 -3480 1452 -3474
rect 1446 -3486 1452 -3480
rect 1446 -3492 1452 -3486
rect 1446 -3498 1452 -3492
rect 1452 -1122 1458 -1116
rect 1452 -1128 1458 -1122
rect 1452 -1134 1458 -1128
rect 1452 -1140 1458 -1134
rect 1452 -1146 1458 -1140
rect 1452 -1152 1458 -1146
rect 1452 -1266 1458 -1260
rect 1452 -1272 1458 -1266
rect 1452 -1278 1458 -1272
rect 1452 -1284 1458 -1278
rect 1452 -1290 1458 -1284
rect 1452 -1296 1458 -1290
rect 1452 -1302 1458 -1296
rect 1452 -1308 1458 -1302
rect 1452 -1314 1458 -1308
rect 1452 -1320 1458 -1314
rect 1452 -1326 1458 -1320
rect 1452 -1332 1458 -1326
rect 1452 -1338 1458 -1332
rect 1452 -1344 1458 -1338
rect 1452 -1350 1458 -1344
rect 1452 -1356 1458 -1350
rect 1452 -1362 1458 -1356
rect 1452 -1368 1458 -1362
rect 1452 -1374 1458 -1368
rect 1452 -1380 1458 -1374
rect 1452 -1386 1458 -1380
rect 1452 -1392 1458 -1386
rect 1452 -1398 1458 -1392
rect 1452 -1404 1458 -1398
rect 1452 -1410 1458 -1404
rect 1452 -1416 1458 -1410
rect 1452 -1422 1458 -1416
rect 1452 -1428 1458 -1422
rect 1452 -1434 1458 -1428
rect 1452 -1440 1458 -1434
rect 1452 -1446 1458 -1440
rect 1452 -1452 1458 -1446
rect 1452 -1458 1458 -1452
rect 1452 -1464 1458 -1458
rect 1452 -1470 1458 -1464
rect 1452 -1476 1458 -1470
rect 1452 -1482 1458 -1476
rect 1452 -1488 1458 -1482
rect 1452 -1494 1458 -1488
rect 1452 -1500 1458 -1494
rect 1452 -1506 1458 -1500
rect 1452 -1512 1458 -1506
rect 1452 -1518 1458 -1512
rect 1452 -1524 1458 -1518
rect 1452 -1530 1458 -1524
rect 1452 -1536 1458 -1530
rect 1452 -1542 1458 -1536
rect 1452 -1548 1458 -1542
rect 1452 -1554 1458 -1548
rect 1452 -1560 1458 -1554
rect 1452 -1566 1458 -1560
rect 1452 -1572 1458 -1566
rect 1452 -1578 1458 -1572
rect 1452 -1584 1458 -1578
rect 1452 -1590 1458 -1584
rect 1452 -1596 1458 -1590
rect 1452 -1602 1458 -1596
rect 1452 -1608 1458 -1602
rect 1452 -1614 1458 -1608
rect 1452 -1620 1458 -1614
rect 1452 -1626 1458 -1620
rect 1452 -1632 1458 -1626
rect 1452 -1638 1458 -1632
rect 1452 -1644 1458 -1638
rect 1452 -1650 1458 -1644
rect 1452 -1656 1458 -1650
rect 1452 -1662 1458 -1656
rect 1452 -1668 1458 -1662
rect 1452 -1674 1458 -1668
rect 1452 -1680 1458 -1674
rect 1452 -1686 1458 -1680
rect 1452 -1692 1458 -1686
rect 1452 -1698 1458 -1692
rect 1452 -1704 1458 -1698
rect 1452 -1710 1458 -1704
rect 1452 -1716 1458 -1710
rect 1452 -1722 1458 -1716
rect 1452 -1728 1458 -1722
rect 1452 -1734 1458 -1728
rect 1452 -1740 1458 -1734
rect 1452 -1746 1458 -1740
rect 1452 -1752 1458 -1746
rect 1452 -1758 1458 -1752
rect 1452 -1764 1458 -1758
rect 1452 -1770 1458 -1764
rect 1452 -1776 1458 -1770
rect 1452 -1782 1458 -1776
rect 1452 -1788 1458 -1782
rect 1452 -1794 1458 -1788
rect 1452 -1800 1458 -1794
rect 1452 -1806 1458 -1800
rect 1452 -1812 1458 -1806
rect 1452 -1818 1458 -1812
rect 1452 -1824 1458 -1818
rect 1452 -1830 1458 -1824
rect 1452 -1836 1458 -1830
rect 1452 -1842 1458 -1836
rect 1452 -1848 1458 -1842
rect 1452 -1854 1458 -1848
rect 1452 -1860 1458 -1854
rect 1452 -1866 1458 -1860
rect 1452 -1872 1458 -1866
rect 1452 -1878 1458 -1872
rect 1452 -1884 1458 -1878
rect 1452 -1890 1458 -1884
rect 1452 -1896 1458 -1890
rect 1452 -1902 1458 -1896
rect 1452 -1908 1458 -1902
rect 1452 -1914 1458 -1908
rect 1452 -1920 1458 -1914
rect 1452 -1926 1458 -1920
rect 1452 -1932 1458 -1926
rect 1452 -1938 1458 -1932
rect 1452 -1944 1458 -1938
rect 1452 -1950 1458 -1944
rect 1452 -1956 1458 -1950
rect 1452 -1962 1458 -1956
rect 1452 -1968 1458 -1962
rect 1452 -1974 1458 -1968
rect 1452 -1980 1458 -1974
rect 1452 -1986 1458 -1980
rect 1452 -1992 1458 -1986
rect 1452 -1998 1458 -1992
rect 1452 -2004 1458 -1998
rect 1452 -2010 1458 -2004
rect 1452 -2016 1458 -2010
rect 1452 -2022 1458 -2016
rect 1452 -2028 1458 -2022
rect 1452 -2034 1458 -2028
rect 1452 -2040 1458 -2034
rect 1452 -2046 1458 -2040
rect 1452 -2052 1458 -2046
rect 1452 -2058 1458 -2052
rect 1452 -2064 1458 -2058
rect 1452 -2070 1458 -2064
rect 1452 -2076 1458 -2070
rect 1452 -2082 1458 -2076
rect 1452 -2088 1458 -2082
rect 1452 -2094 1458 -2088
rect 1452 -2100 1458 -2094
rect 1452 -2106 1458 -2100
rect 1452 -2112 1458 -2106
rect 1452 -2118 1458 -2112
rect 1452 -2124 1458 -2118
rect 1452 -2130 1458 -2124
rect 1452 -2136 1458 -2130
rect 1452 -2142 1458 -2136
rect 1452 -2148 1458 -2142
rect 1452 -2154 1458 -2148
rect 1452 -2160 1458 -2154
rect 1452 -2166 1458 -2160
rect 1452 -2172 1458 -2166
rect 1452 -2178 1458 -2172
rect 1452 -2184 1458 -2178
rect 1452 -2190 1458 -2184
rect 1452 -2196 1458 -2190
rect 1452 -2202 1458 -2196
rect 1452 -2208 1458 -2202
rect 1452 -2214 1458 -2208
rect 1452 -2220 1458 -2214
rect 1452 -2226 1458 -2220
rect 1452 -2232 1458 -2226
rect 1452 -2238 1458 -2232
rect 1452 -2244 1458 -2238
rect 1452 -2250 1458 -2244
rect 1452 -2328 1458 -2322
rect 1452 -2334 1458 -2328
rect 1452 -2340 1458 -2334
rect 1452 -2346 1458 -2340
rect 1452 -2352 1458 -2346
rect 1452 -2358 1458 -2352
rect 1452 -2364 1458 -2358
rect 1452 -2370 1458 -2364
rect 1452 -2376 1458 -2370
rect 1452 -2382 1458 -2376
rect 1452 -2388 1458 -2382
rect 1452 -2394 1458 -2388
rect 1452 -2400 1458 -2394
rect 1452 -2406 1458 -2400
rect 1452 -2412 1458 -2406
rect 1452 -2418 1458 -2412
rect 1452 -2424 1458 -2418
rect 1452 -2430 1458 -2424
rect 1452 -2436 1458 -2430
rect 1452 -2442 1458 -2436
rect 1452 -2448 1458 -2442
rect 1452 -2454 1458 -2448
rect 1452 -2460 1458 -2454
rect 1452 -2466 1458 -2460
rect 1452 -2472 1458 -2466
rect 1452 -2478 1458 -2472
rect 1452 -2484 1458 -2478
rect 1452 -2490 1458 -2484
rect 1452 -2496 1458 -2490
rect 1452 -2502 1458 -2496
rect 1452 -2508 1458 -2502
rect 1452 -2514 1458 -2508
rect 1452 -2520 1458 -2514
rect 1452 -2526 1458 -2520
rect 1452 -2532 1458 -2526
rect 1452 -2538 1458 -2532
rect 1452 -2544 1458 -2538
rect 1452 -2550 1458 -2544
rect 1452 -2556 1458 -2550
rect 1452 -2562 1458 -2556
rect 1452 -2568 1458 -2562
rect 1452 -2574 1458 -2568
rect 1452 -2580 1458 -2574
rect 1452 -2586 1458 -2580
rect 1452 -2592 1458 -2586
rect 1452 -2598 1458 -2592
rect 1452 -2604 1458 -2598
rect 1452 -2610 1458 -2604
rect 1452 -2616 1458 -2610
rect 1452 -2622 1458 -2616
rect 1452 -2628 1458 -2622
rect 1452 -2634 1458 -2628
rect 1452 -2640 1458 -2634
rect 1452 -2646 1458 -2640
rect 1452 -2652 1458 -2646
rect 1452 -2658 1458 -2652
rect 1452 -2664 1458 -2658
rect 1452 -2670 1458 -2664
rect 1452 -2676 1458 -2670
rect 1452 -2682 1458 -2676
rect 1452 -2688 1458 -2682
rect 1452 -2694 1458 -2688
rect 1452 -2700 1458 -2694
rect 1452 -2706 1458 -2700
rect 1452 -2712 1458 -2706
rect 1452 -2718 1458 -2712
rect 1452 -2724 1458 -2718
rect 1452 -2730 1458 -2724
rect 1452 -2736 1458 -2730
rect 1452 -2742 1458 -2736
rect 1452 -2748 1458 -2742
rect 1452 -2754 1458 -2748
rect 1452 -2760 1458 -2754
rect 1452 -2766 1458 -2760
rect 1452 -2772 1458 -2766
rect 1452 -2778 1458 -2772
rect 1452 -2784 1458 -2778
rect 1452 -2790 1458 -2784
rect 1452 -2796 1458 -2790
rect 1452 -2802 1458 -2796
rect 1452 -2808 1458 -2802
rect 1452 -2814 1458 -2808
rect 1452 -2820 1458 -2814
rect 1452 -2826 1458 -2820
rect 1452 -2832 1458 -2826
rect 1452 -2838 1458 -2832
rect 1452 -2928 1458 -2922
rect 1452 -2934 1458 -2928
rect 1452 -2940 1458 -2934
rect 1452 -2946 1458 -2940
rect 1452 -2952 1458 -2946
rect 1452 -2958 1458 -2952
rect 1452 -2964 1458 -2958
rect 1452 -2970 1458 -2964
rect 1452 -2976 1458 -2970
rect 1452 -2982 1458 -2976
rect 1452 -2988 1458 -2982
rect 1452 -2994 1458 -2988
rect 1452 -3000 1458 -2994
rect 1452 -3006 1458 -3000
rect 1452 -3012 1458 -3006
rect 1452 -3018 1458 -3012
rect 1452 -3024 1458 -3018
rect 1452 -3030 1458 -3024
rect 1452 -3036 1458 -3030
rect 1452 -3042 1458 -3036
rect 1452 -3048 1458 -3042
rect 1452 -3054 1458 -3048
rect 1452 -3060 1458 -3054
rect 1452 -3066 1458 -3060
rect 1452 -3072 1458 -3066
rect 1452 -3078 1458 -3072
rect 1452 -3084 1458 -3078
rect 1452 -3090 1458 -3084
rect 1452 -3096 1458 -3090
rect 1452 -3102 1458 -3096
rect 1452 -3108 1458 -3102
rect 1452 -3114 1458 -3108
rect 1452 -3120 1458 -3114
rect 1452 -3126 1458 -3120
rect 1452 -3132 1458 -3126
rect 1452 -3138 1458 -3132
rect 1452 -3144 1458 -3138
rect 1452 -3150 1458 -3144
rect 1452 -3156 1458 -3150
rect 1452 -3162 1458 -3156
rect 1452 -3168 1458 -3162
rect 1452 -3174 1458 -3168
rect 1452 -3180 1458 -3174
rect 1452 -3186 1458 -3180
rect 1452 -3192 1458 -3186
rect 1452 -3198 1458 -3192
rect 1452 -3204 1458 -3198
rect 1452 -3210 1458 -3204
rect 1452 -3216 1458 -3210
rect 1452 -3222 1458 -3216
rect 1452 -3228 1458 -3222
rect 1452 -3234 1458 -3228
rect 1452 -3294 1458 -3288
rect 1452 -3300 1458 -3294
rect 1452 -3306 1458 -3300
rect 1452 -3312 1458 -3306
rect 1452 -3318 1458 -3312
rect 1452 -3324 1458 -3318
rect 1452 -3330 1458 -3324
rect 1452 -3336 1458 -3330
rect 1452 -3342 1458 -3336
rect 1452 -3348 1458 -3342
rect 1452 -3354 1458 -3348
rect 1452 -3360 1458 -3354
rect 1452 -3366 1458 -3360
rect 1452 -3372 1458 -3366
rect 1452 -3378 1458 -3372
rect 1452 -3384 1458 -3378
rect 1452 -3390 1458 -3384
rect 1452 -3396 1458 -3390
rect 1452 -3402 1458 -3396
rect 1452 -3408 1458 -3402
rect 1452 -3414 1458 -3408
rect 1452 -3420 1458 -3414
rect 1452 -3426 1458 -3420
rect 1452 -3432 1458 -3426
rect 1452 -3438 1458 -3432
rect 1452 -3444 1458 -3438
rect 1452 -3450 1458 -3444
rect 1452 -3456 1458 -3450
rect 1452 -3462 1458 -3456
rect 1452 -3468 1458 -3462
rect 1452 -3474 1458 -3468
rect 1452 -3480 1458 -3474
rect 1452 -3486 1458 -3480
rect 1452 -3492 1458 -3486
rect 1452 -3498 1458 -3492
rect 1458 -1122 1464 -1116
rect 1458 -1128 1464 -1122
rect 1458 -1134 1464 -1128
rect 1458 -1140 1464 -1134
rect 1458 -1254 1464 -1248
rect 1458 -1260 1464 -1254
rect 1458 -1266 1464 -1260
rect 1458 -1272 1464 -1266
rect 1458 -1278 1464 -1272
rect 1458 -1284 1464 -1278
rect 1458 -1290 1464 -1284
rect 1458 -1296 1464 -1290
rect 1458 -1302 1464 -1296
rect 1458 -1308 1464 -1302
rect 1458 -1314 1464 -1308
rect 1458 -1320 1464 -1314
rect 1458 -1326 1464 -1320
rect 1458 -1332 1464 -1326
rect 1458 -1338 1464 -1332
rect 1458 -1344 1464 -1338
rect 1458 -1350 1464 -1344
rect 1458 -1356 1464 -1350
rect 1458 -1362 1464 -1356
rect 1458 -1368 1464 -1362
rect 1458 -1374 1464 -1368
rect 1458 -1380 1464 -1374
rect 1458 -1386 1464 -1380
rect 1458 -1392 1464 -1386
rect 1458 -1398 1464 -1392
rect 1458 -1404 1464 -1398
rect 1458 -1410 1464 -1404
rect 1458 -1416 1464 -1410
rect 1458 -1422 1464 -1416
rect 1458 -1428 1464 -1422
rect 1458 -1434 1464 -1428
rect 1458 -1440 1464 -1434
rect 1458 -1446 1464 -1440
rect 1458 -1452 1464 -1446
rect 1458 -1458 1464 -1452
rect 1458 -1464 1464 -1458
rect 1458 -1470 1464 -1464
rect 1458 -1476 1464 -1470
rect 1458 -1482 1464 -1476
rect 1458 -1488 1464 -1482
rect 1458 -1494 1464 -1488
rect 1458 -1500 1464 -1494
rect 1458 -1506 1464 -1500
rect 1458 -1512 1464 -1506
rect 1458 -1518 1464 -1512
rect 1458 -1524 1464 -1518
rect 1458 -1530 1464 -1524
rect 1458 -1536 1464 -1530
rect 1458 -1542 1464 -1536
rect 1458 -1548 1464 -1542
rect 1458 -1554 1464 -1548
rect 1458 -1560 1464 -1554
rect 1458 -1566 1464 -1560
rect 1458 -1572 1464 -1566
rect 1458 -1578 1464 -1572
rect 1458 -1584 1464 -1578
rect 1458 -1590 1464 -1584
rect 1458 -1596 1464 -1590
rect 1458 -1602 1464 -1596
rect 1458 -1608 1464 -1602
rect 1458 -1614 1464 -1608
rect 1458 -1620 1464 -1614
rect 1458 -1626 1464 -1620
rect 1458 -1632 1464 -1626
rect 1458 -1638 1464 -1632
rect 1458 -1644 1464 -1638
rect 1458 -1650 1464 -1644
rect 1458 -1656 1464 -1650
rect 1458 -1662 1464 -1656
rect 1458 -1668 1464 -1662
rect 1458 -1674 1464 -1668
rect 1458 -1680 1464 -1674
rect 1458 -1686 1464 -1680
rect 1458 -1692 1464 -1686
rect 1458 -1698 1464 -1692
rect 1458 -1704 1464 -1698
rect 1458 -1710 1464 -1704
rect 1458 -1716 1464 -1710
rect 1458 -1722 1464 -1716
rect 1458 -1728 1464 -1722
rect 1458 -1734 1464 -1728
rect 1458 -1740 1464 -1734
rect 1458 -1746 1464 -1740
rect 1458 -1752 1464 -1746
rect 1458 -1758 1464 -1752
rect 1458 -1764 1464 -1758
rect 1458 -1770 1464 -1764
rect 1458 -1776 1464 -1770
rect 1458 -1782 1464 -1776
rect 1458 -1788 1464 -1782
rect 1458 -1794 1464 -1788
rect 1458 -1800 1464 -1794
rect 1458 -1806 1464 -1800
rect 1458 -1812 1464 -1806
rect 1458 -1818 1464 -1812
rect 1458 -1824 1464 -1818
rect 1458 -1830 1464 -1824
rect 1458 -1836 1464 -1830
rect 1458 -1842 1464 -1836
rect 1458 -1848 1464 -1842
rect 1458 -1854 1464 -1848
rect 1458 -1860 1464 -1854
rect 1458 -1866 1464 -1860
rect 1458 -1872 1464 -1866
rect 1458 -1878 1464 -1872
rect 1458 -1884 1464 -1878
rect 1458 -1890 1464 -1884
rect 1458 -1896 1464 -1890
rect 1458 -1902 1464 -1896
rect 1458 -1908 1464 -1902
rect 1458 -1914 1464 -1908
rect 1458 -1920 1464 -1914
rect 1458 -1926 1464 -1920
rect 1458 -1932 1464 -1926
rect 1458 -1938 1464 -1932
rect 1458 -1944 1464 -1938
rect 1458 -1950 1464 -1944
rect 1458 -1956 1464 -1950
rect 1458 -1962 1464 -1956
rect 1458 -1968 1464 -1962
rect 1458 -1974 1464 -1968
rect 1458 -1980 1464 -1974
rect 1458 -1986 1464 -1980
rect 1458 -1992 1464 -1986
rect 1458 -1998 1464 -1992
rect 1458 -2004 1464 -1998
rect 1458 -2010 1464 -2004
rect 1458 -2016 1464 -2010
rect 1458 -2022 1464 -2016
rect 1458 -2028 1464 -2022
rect 1458 -2034 1464 -2028
rect 1458 -2040 1464 -2034
rect 1458 -2046 1464 -2040
rect 1458 -2052 1464 -2046
rect 1458 -2058 1464 -2052
rect 1458 -2064 1464 -2058
rect 1458 -2070 1464 -2064
rect 1458 -2076 1464 -2070
rect 1458 -2082 1464 -2076
rect 1458 -2088 1464 -2082
rect 1458 -2094 1464 -2088
rect 1458 -2100 1464 -2094
rect 1458 -2106 1464 -2100
rect 1458 -2112 1464 -2106
rect 1458 -2118 1464 -2112
rect 1458 -2124 1464 -2118
rect 1458 -2130 1464 -2124
rect 1458 -2136 1464 -2130
rect 1458 -2142 1464 -2136
rect 1458 -2148 1464 -2142
rect 1458 -2154 1464 -2148
rect 1458 -2160 1464 -2154
rect 1458 -2166 1464 -2160
rect 1458 -2172 1464 -2166
rect 1458 -2178 1464 -2172
rect 1458 -2184 1464 -2178
rect 1458 -2190 1464 -2184
rect 1458 -2196 1464 -2190
rect 1458 -2202 1464 -2196
rect 1458 -2208 1464 -2202
rect 1458 -2214 1464 -2208
rect 1458 -2220 1464 -2214
rect 1458 -2226 1464 -2220
rect 1458 -2232 1464 -2226
rect 1458 -2238 1464 -2232
rect 1458 -2244 1464 -2238
rect 1458 -2316 1464 -2310
rect 1458 -2322 1464 -2316
rect 1458 -2328 1464 -2322
rect 1458 -2334 1464 -2328
rect 1458 -2340 1464 -2334
rect 1458 -2346 1464 -2340
rect 1458 -2352 1464 -2346
rect 1458 -2358 1464 -2352
rect 1458 -2364 1464 -2358
rect 1458 -2370 1464 -2364
rect 1458 -2376 1464 -2370
rect 1458 -2382 1464 -2376
rect 1458 -2388 1464 -2382
rect 1458 -2394 1464 -2388
rect 1458 -2400 1464 -2394
rect 1458 -2406 1464 -2400
rect 1458 -2412 1464 -2406
rect 1458 -2418 1464 -2412
rect 1458 -2424 1464 -2418
rect 1458 -2430 1464 -2424
rect 1458 -2436 1464 -2430
rect 1458 -2442 1464 -2436
rect 1458 -2448 1464 -2442
rect 1458 -2454 1464 -2448
rect 1458 -2460 1464 -2454
rect 1458 -2466 1464 -2460
rect 1458 -2472 1464 -2466
rect 1458 -2478 1464 -2472
rect 1458 -2484 1464 -2478
rect 1458 -2490 1464 -2484
rect 1458 -2496 1464 -2490
rect 1458 -2502 1464 -2496
rect 1458 -2508 1464 -2502
rect 1458 -2514 1464 -2508
rect 1458 -2520 1464 -2514
rect 1458 -2526 1464 -2520
rect 1458 -2532 1464 -2526
rect 1458 -2538 1464 -2532
rect 1458 -2544 1464 -2538
rect 1458 -2550 1464 -2544
rect 1458 -2556 1464 -2550
rect 1458 -2562 1464 -2556
rect 1458 -2568 1464 -2562
rect 1458 -2574 1464 -2568
rect 1458 -2580 1464 -2574
rect 1458 -2586 1464 -2580
rect 1458 -2592 1464 -2586
rect 1458 -2598 1464 -2592
rect 1458 -2604 1464 -2598
rect 1458 -2610 1464 -2604
rect 1458 -2616 1464 -2610
rect 1458 -2622 1464 -2616
rect 1458 -2628 1464 -2622
rect 1458 -2634 1464 -2628
rect 1458 -2640 1464 -2634
rect 1458 -2646 1464 -2640
rect 1458 -2652 1464 -2646
rect 1458 -2658 1464 -2652
rect 1458 -2664 1464 -2658
rect 1458 -2670 1464 -2664
rect 1458 -2676 1464 -2670
rect 1458 -2682 1464 -2676
rect 1458 -2688 1464 -2682
rect 1458 -2694 1464 -2688
rect 1458 -2700 1464 -2694
rect 1458 -2706 1464 -2700
rect 1458 -2712 1464 -2706
rect 1458 -2718 1464 -2712
rect 1458 -2724 1464 -2718
rect 1458 -2730 1464 -2724
rect 1458 -2736 1464 -2730
rect 1458 -2742 1464 -2736
rect 1458 -2748 1464 -2742
rect 1458 -2754 1464 -2748
rect 1458 -2760 1464 -2754
rect 1458 -2766 1464 -2760
rect 1458 -2772 1464 -2766
rect 1458 -2778 1464 -2772
rect 1458 -2784 1464 -2778
rect 1458 -2790 1464 -2784
rect 1458 -2796 1464 -2790
rect 1458 -2802 1464 -2796
rect 1458 -2808 1464 -2802
rect 1458 -2814 1464 -2808
rect 1458 -2820 1464 -2814
rect 1458 -2826 1464 -2820
rect 1458 -2832 1464 -2826
rect 1458 -2838 1464 -2832
rect 1458 -2922 1464 -2916
rect 1458 -2928 1464 -2922
rect 1458 -2934 1464 -2928
rect 1458 -2940 1464 -2934
rect 1458 -2946 1464 -2940
rect 1458 -2952 1464 -2946
rect 1458 -2958 1464 -2952
rect 1458 -2964 1464 -2958
rect 1458 -2970 1464 -2964
rect 1458 -2976 1464 -2970
rect 1458 -2982 1464 -2976
rect 1458 -2988 1464 -2982
rect 1458 -2994 1464 -2988
rect 1458 -3000 1464 -2994
rect 1458 -3006 1464 -3000
rect 1458 -3012 1464 -3006
rect 1458 -3018 1464 -3012
rect 1458 -3024 1464 -3018
rect 1458 -3030 1464 -3024
rect 1458 -3036 1464 -3030
rect 1458 -3042 1464 -3036
rect 1458 -3048 1464 -3042
rect 1458 -3054 1464 -3048
rect 1458 -3060 1464 -3054
rect 1458 -3066 1464 -3060
rect 1458 -3072 1464 -3066
rect 1458 -3078 1464 -3072
rect 1458 -3084 1464 -3078
rect 1458 -3090 1464 -3084
rect 1458 -3096 1464 -3090
rect 1458 -3102 1464 -3096
rect 1458 -3108 1464 -3102
rect 1458 -3114 1464 -3108
rect 1458 -3120 1464 -3114
rect 1458 -3126 1464 -3120
rect 1458 -3132 1464 -3126
rect 1458 -3138 1464 -3132
rect 1458 -3144 1464 -3138
rect 1458 -3150 1464 -3144
rect 1458 -3156 1464 -3150
rect 1458 -3162 1464 -3156
rect 1458 -3168 1464 -3162
rect 1458 -3174 1464 -3168
rect 1458 -3180 1464 -3174
rect 1458 -3186 1464 -3180
rect 1458 -3192 1464 -3186
rect 1458 -3198 1464 -3192
rect 1458 -3204 1464 -3198
rect 1458 -3210 1464 -3204
rect 1458 -3216 1464 -3210
rect 1458 -3222 1464 -3216
rect 1458 -3228 1464 -3222
rect 1458 -3234 1464 -3228
rect 1458 -3294 1464 -3288
rect 1458 -3300 1464 -3294
rect 1458 -3306 1464 -3300
rect 1458 -3312 1464 -3306
rect 1458 -3318 1464 -3312
rect 1458 -3324 1464 -3318
rect 1458 -3330 1464 -3324
rect 1458 -3336 1464 -3330
rect 1458 -3342 1464 -3336
rect 1458 -3348 1464 -3342
rect 1458 -3354 1464 -3348
rect 1458 -3360 1464 -3354
rect 1458 -3366 1464 -3360
rect 1458 -3372 1464 -3366
rect 1458 -3378 1464 -3372
rect 1458 -3384 1464 -3378
rect 1458 -3390 1464 -3384
rect 1458 -3396 1464 -3390
rect 1458 -3402 1464 -3396
rect 1458 -3408 1464 -3402
rect 1458 -3414 1464 -3408
rect 1458 -3420 1464 -3414
rect 1458 -3426 1464 -3420
rect 1458 -3432 1464 -3426
rect 1458 -3438 1464 -3432
rect 1458 -3444 1464 -3438
rect 1458 -3450 1464 -3444
rect 1458 -3456 1464 -3450
rect 1458 -3462 1464 -3456
rect 1458 -3468 1464 -3462
rect 1458 -3474 1464 -3468
rect 1458 -3480 1464 -3474
rect 1458 -3486 1464 -3480
rect 1458 -3492 1464 -3486
rect 1458 -3498 1464 -3492
rect 1464 -1122 1470 -1116
rect 1464 -1128 1470 -1122
rect 1464 -1242 1470 -1236
rect 1464 -1248 1470 -1242
rect 1464 -1254 1470 -1248
rect 1464 -1260 1470 -1254
rect 1464 -1266 1470 -1260
rect 1464 -1272 1470 -1266
rect 1464 -1278 1470 -1272
rect 1464 -1284 1470 -1278
rect 1464 -1290 1470 -1284
rect 1464 -1296 1470 -1290
rect 1464 -1302 1470 -1296
rect 1464 -1308 1470 -1302
rect 1464 -1314 1470 -1308
rect 1464 -1320 1470 -1314
rect 1464 -1326 1470 -1320
rect 1464 -1332 1470 -1326
rect 1464 -1338 1470 -1332
rect 1464 -1344 1470 -1338
rect 1464 -1350 1470 -1344
rect 1464 -1356 1470 -1350
rect 1464 -1362 1470 -1356
rect 1464 -1368 1470 -1362
rect 1464 -1374 1470 -1368
rect 1464 -1380 1470 -1374
rect 1464 -1386 1470 -1380
rect 1464 -1392 1470 -1386
rect 1464 -1398 1470 -1392
rect 1464 -1404 1470 -1398
rect 1464 -1410 1470 -1404
rect 1464 -1416 1470 -1410
rect 1464 -1422 1470 -1416
rect 1464 -1428 1470 -1422
rect 1464 -1434 1470 -1428
rect 1464 -1440 1470 -1434
rect 1464 -1446 1470 -1440
rect 1464 -1452 1470 -1446
rect 1464 -1458 1470 -1452
rect 1464 -1464 1470 -1458
rect 1464 -1470 1470 -1464
rect 1464 -1476 1470 -1470
rect 1464 -1482 1470 -1476
rect 1464 -1488 1470 -1482
rect 1464 -1494 1470 -1488
rect 1464 -1500 1470 -1494
rect 1464 -1506 1470 -1500
rect 1464 -1512 1470 -1506
rect 1464 -1518 1470 -1512
rect 1464 -1524 1470 -1518
rect 1464 -1530 1470 -1524
rect 1464 -1536 1470 -1530
rect 1464 -1542 1470 -1536
rect 1464 -1548 1470 -1542
rect 1464 -1554 1470 -1548
rect 1464 -1560 1470 -1554
rect 1464 -1566 1470 -1560
rect 1464 -1572 1470 -1566
rect 1464 -1578 1470 -1572
rect 1464 -1584 1470 -1578
rect 1464 -1590 1470 -1584
rect 1464 -1596 1470 -1590
rect 1464 -1602 1470 -1596
rect 1464 -1608 1470 -1602
rect 1464 -1614 1470 -1608
rect 1464 -1620 1470 -1614
rect 1464 -1626 1470 -1620
rect 1464 -1632 1470 -1626
rect 1464 -1638 1470 -1632
rect 1464 -1644 1470 -1638
rect 1464 -1650 1470 -1644
rect 1464 -1656 1470 -1650
rect 1464 -1662 1470 -1656
rect 1464 -1668 1470 -1662
rect 1464 -1674 1470 -1668
rect 1464 -1680 1470 -1674
rect 1464 -1686 1470 -1680
rect 1464 -1692 1470 -1686
rect 1464 -1698 1470 -1692
rect 1464 -1704 1470 -1698
rect 1464 -1710 1470 -1704
rect 1464 -1716 1470 -1710
rect 1464 -1722 1470 -1716
rect 1464 -1728 1470 -1722
rect 1464 -1734 1470 -1728
rect 1464 -1740 1470 -1734
rect 1464 -1746 1470 -1740
rect 1464 -1752 1470 -1746
rect 1464 -1758 1470 -1752
rect 1464 -1764 1470 -1758
rect 1464 -1770 1470 -1764
rect 1464 -1776 1470 -1770
rect 1464 -1782 1470 -1776
rect 1464 -1788 1470 -1782
rect 1464 -1794 1470 -1788
rect 1464 -1800 1470 -1794
rect 1464 -1806 1470 -1800
rect 1464 -1812 1470 -1806
rect 1464 -1818 1470 -1812
rect 1464 -1824 1470 -1818
rect 1464 -1830 1470 -1824
rect 1464 -1836 1470 -1830
rect 1464 -1842 1470 -1836
rect 1464 -1848 1470 -1842
rect 1464 -1854 1470 -1848
rect 1464 -1860 1470 -1854
rect 1464 -1866 1470 -1860
rect 1464 -1872 1470 -1866
rect 1464 -1878 1470 -1872
rect 1464 -1884 1470 -1878
rect 1464 -1890 1470 -1884
rect 1464 -1896 1470 -1890
rect 1464 -1902 1470 -1896
rect 1464 -1908 1470 -1902
rect 1464 -1914 1470 -1908
rect 1464 -1920 1470 -1914
rect 1464 -1926 1470 -1920
rect 1464 -1932 1470 -1926
rect 1464 -1938 1470 -1932
rect 1464 -1944 1470 -1938
rect 1464 -1950 1470 -1944
rect 1464 -1956 1470 -1950
rect 1464 -1962 1470 -1956
rect 1464 -1968 1470 -1962
rect 1464 -1974 1470 -1968
rect 1464 -1980 1470 -1974
rect 1464 -1986 1470 -1980
rect 1464 -1992 1470 -1986
rect 1464 -1998 1470 -1992
rect 1464 -2004 1470 -1998
rect 1464 -2010 1470 -2004
rect 1464 -2016 1470 -2010
rect 1464 -2022 1470 -2016
rect 1464 -2028 1470 -2022
rect 1464 -2034 1470 -2028
rect 1464 -2040 1470 -2034
rect 1464 -2046 1470 -2040
rect 1464 -2052 1470 -2046
rect 1464 -2058 1470 -2052
rect 1464 -2064 1470 -2058
rect 1464 -2070 1470 -2064
rect 1464 -2076 1470 -2070
rect 1464 -2082 1470 -2076
rect 1464 -2088 1470 -2082
rect 1464 -2094 1470 -2088
rect 1464 -2100 1470 -2094
rect 1464 -2106 1470 -2100
rect 1464 -2112 1470 -2106
rect 1464 -2118 1470 -2112
rect 1464 -2124 1470 -2118
rect 1464 -2130 1470 -2124
rect 1464 -2136 1470 -2130
rect 1464 -2142 1470 -2136
rect 1464 -2148 1470 -2142
rect 1464 -2154 1470 -2148
rect 1464 -2160 1470 -2154
rect 1464 -2166 1470 -2160
rect 1464 -2172 1470 -2166
rect 1464 -2178 1470 -2172
rect 1464 -2184 1470 -2178
rect 1464 -2190 1470 -2184
rect 1464 -2196 1470 -2190
rect 1464 -2202 1470 -2196
rect 1464 -2208 1470 -2202
rect 1464 -2214 1470 -2208
rect 1464 -2220 1470 -2214
rect 1464 -2226 1470 -2220
rect 1464 -2232 1470 -2226
rect 1464 -2238 1470 -2232
rect 1464 -2310 1470 -2304
rect 1464 -2316 1470 -2310
rect 1464 -2322 1470 -2316
rect 1464 -2328 1470 -2322
rect 1464 -2334 1470 -2328
rect 1464 -2340 1470 -2334
rect 1464 -2346 1470 -2340
rect 1464 -2352 1470 -2346
rect 1464 -2358 1470 -2352
rect 1464 -2364 1470 -2358
rect 1464 -2370 1470 -2364
rect 1464 -2376 1470 -2370
rect 1464 -2382 1470 -2376
rect 1464 -2388 1470 -2382
rect 1464 -2394 1470 -2388
rect 1464 -2400 1470 -2394
rect 1464 -2406 1470 -2400
rect 1464 -2412 1470 -2406
rect 1464 -2418 1470 -2412
rect 1464 -2424 1470 -2418
rect 1464 -2430 1470 -2424
rect 1464 -2436 1470 -2430
rect 1464 -2442 1470 -2436
rect 1464 -2448 1470 -2442
rect 1464 -2454 1470 -2448
rect 1464 -2460 1470 -2454
rect 1464 -2466 1470 -2460
rect 1464 -2472 1470 -2466
rect 1464 -2478 1470 -2472
rect 1464 -2484 1470 -2478
rect 1464 -2490 1470 -2484
rect 1464 -2496 1470 -2490
rect 1464 -2502 1470 -2496
rect 1464 -2508 1470 -2502
rect 1464 -2514 1470 -2508
rect 1464 -2520 1470 -2514
rect 1464 -2526 1470 -2520
rect 1464 -2532 1470 -2526
rect 1464 -2538 1470 -2532
rect 1464 -2544 1470 -2538
rect 1464 -2550 1470 -2544
rect 1464 -2556 1470 -2550
rect 1464 -2562 1470 -2556
rect 1464 -2568 1470 -2562
rect 1464 -2574 1470 -2568
rect 1464 -2580 1470 -2574
rect 1464 -2586 1470 -2580
rect 1464 -2592 1470 -2586
rect 1464 -2598 1470 -2592
rect 1464 -2604 1470 -2598
rect 1464 -2610 1470 -2604
rect 1464 -2616 1470 -2610
rect 1464 -2622 1470 -2616
rect 1464 -2628 1470 -2622
rect 1464 -2634 1470 -2628
rect 1464 -2640 1470 -2634
rect 1464 -2646 1470 -2640
rect 1464 -2652 1470 -2646
rect 1464 -2658 1470 -2652
rect 1464 -2664 1470 -2658
rect 1464 -2670 1470 -2664
rect 1464 -2676 1470 -2670
rect 1464 -2682 1470 -2676
rect 1464 -2688 1470 -2682
rect 1464 -2694 1470 -2688
rect 1464 -2700 1470 -2694
rect 1464 -2706 1470 -2700
rect 1464 -2712 1470 -2706
rect 1464 -2718 1470 -2712
rect 1464 -2724 1470 -2718
rect 1464 -2730 1470 -2724
rect 1464 -2736 1470 -2730
rect 1464 -2742 1470 -2736
rect 1464 -2748 1470 -2742
rect 1464 -2754 1470 -2748
rect 1464 -2760 1470 -2754
rect 1464 -2766 1470 -2760
rect 1464 -2772 1470 -2766
rect 1464 -2778 1470 -2772
rect 1464 -2784 1470 -2778
rect 1464 -2790 1470 -2784
rect 1464 -2796 1470 -2790
rect 1464 -2802 1470 -2796
rect 1464 -2808 1470 -2802
rect 1464 -2814 1470 -2808
rect 1464 -2820 1470 -2814
rect 1464 -2826 1470 -2820
rect 1464 -2832 1470 -2826
rect 1464 -2916 1470 -2910
rect 1464 -2922 1470 -2916
rect 1464 -2928 1470 -2922
rect 1464 -2934 1470 -2928
rect 1464 -2940 1470 -2934
rect 1464 -2946 1470 -2940
rect 1464 -2952 1470 -2946
rect 1464 -2958 1470 -2952
rect 1464 -2964 1470 -2958
rect 1464 -2970 1470 -2964
rect 1464 -2976 1470 -2970
rect 1464 -2982 1470 -2976
rect 1464 -2988 1470 -2982
rect 1464 -2994 1470 -2988
rect 1464 -3000 1470 -2994
rect 1464 -3006 1470 -3000
rect 1464 -3012 1470 -3006
rect 1464 -3018 1470 -3012
rect 1464 -3024 1470 -3018
rect 1464 -3030 1470 -3024
rect 1464 -3036 1470 -3030
rect 1464 -3042 1470 -3036
rect 1464 -3048 1470 -3042
rect 1464 -3054 1470 -3048
rect 1464 -3060 1470 -3054
rect 1464 -3066 1470 -3060
rect 1464 -3072 1470 -3066
rect 1464 -3078 1470 -3072
rect 1464 -3084 1470 -3078
rect 1464 -3090 1470 -3084
rect 1464 -3096 1470 -3090
rect 1464 -3102 1470 -3096
rect 1464 -3108 1470 -3102
rect 1464 -3114 1470 -3108
rect 1464 -3120 1470 -3114
rect 1464 -3126 1470 -3120
rect 1464 -3132 1470 -3126
rect 1464 -3138 1470 -3132
rect 1464 -3144 1470 -3138
rect 1464 -3150 1470 -3144
rect 1464 -3156 1470 -3150
rect 1464 -3162 1470 -3156
rect 1464 -3168 1470 -3162
rect 1464 -3174 1470 -3168
rect 1464 -3180 1470 -3174
rect 1464 -3186 1470 -3180
rect 1464 -3192 1470 -3186
rect 1464 -3198 1470 -3192
rect 1464 -3204 1470 -3198
rect 1464 -3210 1470 -3204
rect 1464 -3216 1470 -3210
rect 1464 -3222 1470 -3216
rect 1464 -3228 1470 -3222
rect 1464 -3234 1470 -3228
rect 1464 -3288 1470 -3282
rect 1464 -3294 1470 -3288
rect 1464 -3300 1470 -3294
rect 1464 -3306 1470 -3300
rect 1464 -3312 1470 -3306
rect 1464 -3318 1470 -3312
rect 1464 -3324 1470 -3318
rect 1464 -3330 1470 -3324
rect 1464 -3336 1470 -3330
rect 1464 -3342 1470 -3336
rect 1464 -3348 1470 -3342
rect 1464 -3354 1470 -3348
rect 1464 -3360 1470 -3354
rect 1464 -3366 1470 -3360
rect 1464 -3372 1470 -3366
rect 1464 -3378 1470 -3372
rect 1464 -3384 1470 -3378
rect 1464 -3390 1470 -3384
rect 1464 -3396 1470 -3390
rect 1464 -3402 1470 -3396
rect 1464 -3408 1470 -3402
rect 1464 -3414 1470 -3408
rect 1464 -3420 1470 -3414
rect 1464 -3426 1470 -3420
rect 1464 -3432 1470 -3426
rect 1464 -3438 1470 -3432
rect 1464 -3444 1470 -3438
rect 1464 -3450 1470 -3444
rect 1464 -3456 1470 -3450
rect 1464 -3462 1470 -3456
rect 1464 -3468 1470 -3462
rect 1464 -3474 1470 -3468
rect 1464 -3480 1470 -3474
rect 1464 -3486 1470 -3480
rect 1464 -3492 1470 -3486
rect 1464 -3498 1470 -3492
rect 1470 -1236 1476 -1230
rect 1470 -1242 1476 -1236
rect 1470 -1248 1476 -1242
rect 1470 -1254 1476 -1248
rect 1470 -1260 1476 -1254
rect 1470 -1266 1476 -1260
rect 1470 -1272 1476 -1266
rect 1470 -1278 1476 -1272
rect 1470 -1284 1476 -1278
rect 1470 -1290 1476 -1284
rect 1470 -1296 1476 -1290
rect 1470 -1302 1476 -1296
rect 1470 -1308 1476 -1302
rect 1470 -1314 1476 -1308
rect 1470 -1320 1476 -1314
rect 1470 -1326 1476 -1320
rect 1470 -1332 1476 -1326
rect 1470 -1338 1476 -1332
rect 1470 -1344 1476 -1338
rect 1470 -1350 1476 -1344
rect 1470 -1356 1476 -1350
rect 1470 -1362 1476 -1356
rect 1470 -1368 1476 -1362
rect 1470 -1374 1476 -1368
rect 1470 -1380 1476 -1374
rect 1470 -1386 1476 -1380
rect 1470 -1392 1476 -1386
rect 1470 -1398 1476 -1392
rect 1470 -1404 1476 -1398
rect 1470 -1410 1476 -1404
rect 1470 -1416 1476 -1410
rect 1470 -1422 1476 -1416
rect 1470 -1428 1476 -1422
rect 1470 -1434 1476 -1428
rect 1470 -1440 1476 -1434
rect 1470 -1446 1476 -1440
rect 1470 -1452 1476 -1446
rect 1470 -1458 1476 -1452
rect 1470 -1464 1476 -1458
rect 1470 -1470 1476 -1464
rect 1470 -1476 1476 -1470
rect 1470 -1482 1476 -1476
rect 1470 -1488 1476 -1482
rect 1470 -1494 1476 -1488
rect 1470 -1500 1476 -1494
rect 1470 -1506 1476 -1500
rect 1470 -1512 1476 -1506
rect 1470 -1518 1476 -1512
rect 1470 -1524 1476 -1518
rect 1470 -1530 1476 -1524
rect 1470 -1536 1476 -1530
rect 1470 -1542 1476 -1536
rect 1470 -1548 1476 -1542
rect 1470 -1554 1476 -1548
rect 1470 -1560 1476 -1554
rect 1470 -1566 1476 -1560
rect 1470 -1572 1476 -1566
rect 1470 -1578 1476 -1572
rect 1470 -1584 1476 -1578
rect 1470 -1590 1476 -1584
rect 1470 -1596 1476 -1590
rect 1470 -1602 1476 -1596
rect 1470 -1608 1476 -1602
rect 1470 -1614 1476 -1608
rect 1470 -1620 1476 -1614
rect 1470 -1626 1476 -1620
rect 1470 -1632 1476 -1626
rect 1470 -1638 1476 -1632
rect 1470 -1644 1476 -1638
rect 1470 -1650 1476 -1644
rect 1470 -1656 1476 -1650
rect 1470 -1662 1476 -1656
rect 1470 -1668 1476 -1662
rect 1470 -1674 1476 -1668
rect 1470 -1680 1476 -1674
rect 1470 -1686 1476 -1680
rect 1470 -1692 1476 -1686
rect 1470 -1698 1476 -1692
rect 1470 -1704 1476 -1698
rect 1470 -1710 1476 -1704
rect 1470 -1716 1476 -1710
rect 1470 -1722 1476 -1716
rect 1470 -1728 1476 -1722
rect 1470 -1734 1476 -1728
rect 1470 -1740 1476 -1734
rect 1470 -1746 1476 -1740
rect 1470 -1752 1476 -1746
rect 1470 -1758 1476 -1752
rect 1470 -1764 1476 -1758
rect 1470 -1770 1476 -1764
rect 1470 -1776 1476 -1770
rect 1470 -1782 1476 -1776
rect 1470 -1788 1476 -1782
rect 1470 -1794 1476 -1788
rect 1470 -1800 1476 -1794
rect 1470 -1806 1476 -1800
rect 1470 -1812 1476 -1806
rect 1470 -1818 1476 -1812
rect 1470 -1824 1476 -1818
rect 1470 -1830 1476 -1824
rect 1470 -1836 1476 -1830
rect 1470 -1842 1476 -1836
rect 1470 -1848 1476 -1842
rect 1470 -1854 1476 -1848
rect 1470 -1860 1476 -1854
rect 1470 -1866 1476 -1860
rect 1470 -1872 1476 -1866
rect 1470 -1878 1476 -1872
rect 1470 -1884 1476 -1878
rect 1470 -1890 1476 -1884
rect 1470 -1896 1476 -1890
rect 1470 -1902 1476 -1896
rect 1470 -1908 1476 -1902
rect 1470 -1914 1476 -1908
rect 1470 -1920 1476 -1914
rect 1470 -1926 1476 -1920
rect 1470 -1932 1476 -1926
rect 1470 -1938 1476 -1932
rect 1470 -1944 1476 -1938
rect 1470 -1950 1476 -1944
rect 1470 -1956 1476 -1950
rect 1470 -1962 1476 -1956
rect 1470 -1968 1476 -1962
rect 1470 -1974 1476 -1968
rect 1470 -1980 1476 -1974
rect 1470 -1986 1476 -1980
rect 1470 -1992 1476 -1986
rect 1470 -1998 1476 -1992
rect 1470 -2004 1476 -1998
rect 1470 -2010 1476 -2004
rect 1470 -2016 1476 -2010
rect 1470 -2022 1476 -2016
rect 1470 -2028 1476 -2022
rect 1470 -2034 1476 -2028
rect 1470 -2040 1476 -2034
rect 1470 -2046 1476 -2040
rect 1470 -2052 1476 -2046
rect 1470 -2058 1476 -2052
rect 1470 -2064 1476 -2058
rect 1470 -2070 1476 -2064
rect 1470 -2076 1476 -2070
rect 1470 -2082 1476 -2076
rect 1470 -2088 1476 -2082
rect 1470 -2094 1476 -2088
rect 1470 -2100 1476 -2094
rect 1470 -2106 1476 -2100
rect 1470 -2112 1476 -2106
rect 1470 -2118 1476 -2112
rect 1470 -2124 1476 -2118
rect 1470 -2130 1476 -2124
rect 1470 -2136 1476 -2130
rect 1470 -2142 1476 -2136
rect 1470 -2148 1476 -2142
rect 1470 -2154 1476 -2148
rect 1470 -2160 1476 -2154
rect 1470 -2166 1476 -2160
rect 1470 -2172 1476 -2166
rect 1470 -2178 1476 -2172
rect 1470 -2184 1476 -2178
rect 1470 -2190 1476 -2184
rect 1470 -2196 1476 -2190
rect 1470 -2202 1476 -2196
rect 1470 -2208 1476 -2202
rect 1470 -2214 1476 -2208
rect 1470 -2220 1476 -2214
rect 1470 -2226 1476 -2220
rect 1470 -2304 1476 -2298
rect 1470 -2310 1476 -2304
rect 1470 -2316 1476 -2310
rect 1470 -2322 1476 -2316
rect 1470 -2328 1476 -2322
rect 1470 -2334 1476 -2328
rect 1470 -2340 1476 -2334
rect 1470 -2346 1476 -2340
rect 1470 -2352 1476 -2346
rect 1470 -2358 1476 -2352
rect 1470 -2364 1476 -2358
rect 1470 -2370 1476 -2364
rect 1470 -2376 1476 -2370
rect 1470 -2382 1476 -2376
rect 1470 -2388 1476 -2382
rect 1470 -2394 1476 -2388
rect 1470 -2400 1476 -2394
rect 1470 -2406 1476 -2400
rect 1470 -2412 1476 -2406
rect 1470 -2418 1476 -2412
rect 1470 -2424 1476 -2418
rect 1470 -2430 1476 -2424
rect 1470 -2436 1476 -2430
rect 1470 -2442 1476 -2436
rect 1470 -2448 1476 -2442
rect 1470 -2454 1476 -2448
rect 1470 -2460 1476 -2454
rect 1470 -2466 1476 -2460
rect 1470 -2472 1476 -2466
rect 1470 -2478 1476 -2472
rect 1470 -2484 1476 -2478
rect 1470 -2490 1476 -2484
rect 1470 -2496 1476 -2490
rect 1470 -2502 1476 -2496
rect 1470 -2508 1476 -2502
rect 1470 -2514 1476 -2508
rect 1470 -2520 1476 -2514
rect 1470 -2526 1476 -2520
rect 1470 -2532 1476 -2526
rect 1470 -2538 1476 -2532
rect 1470 -2544 1476 -2538
rect 1470 -2550 1476 -2544
rect 1470 -2556 1476 -2550
rect 1470 -2562 1476 -2556
rect 1470 -2568 1476 -2562
rect 1470 -2574 1476 -2568
rect 1470 -2580 1476 -2574
rect 1470 -2586 1476 -2580
rect 1470 -2592 1476 -2586
rect 1470 -2598 1476 -2592
rect 1470 -2604 1476 -2598
rect 1470 -2610 1476 -2604
rect 1470 -2616 1476 -2610
rect 1470 -2622 1476 -2616
rect 1470 -2628 1476 -2622
rect 1470 -2634 1476 -2628
rect 1470 -2640 1476 -2634
rect 1470 -2646 1476 -2640
rect 1470 -2652 1476 -2646
rect 1470 -2658 1476 -2652
rect 1470 -2664 1476 -2658
rect 1470 -2670 1476 -2664
rect 1470 -2676 1476 -2670
rect 1470 -2682 1476 -2676
rect 1470 -2688 1476 -2682
rect 1470 -2694 1476 -2688
rect 1470 -2700 1476 -2694
rect 1470 -2706 1476 -2700
rect 1470 -2712 1476 -2706
rect 1470 -2718 1476 -2712
rect 1470 -2724 1476 -2718
rect 1470 -2730 1476 -2724
rect 1470 -2736 1476 -2730
rect 1470 -2742 1476 -2736
rect 1470 -2748 1476 -2742
rect 1470 -2754 1476 -2748
rect 1470 -2760 1476 -2754
rect 1470 -2766 1476 -2760
rect 1470 -2772 1476 -2766
rect 1470 -2778 1476 -2772
rect 1470 -2784 1476 -2778
rect 1470 -2790 1476 -2784
rect 1470 -2796 1476 -2790
rect 1470 -2802 1476 -2796
rect 1470 -2808 1476 -2802
rect 1470 -2814 1476 -2808
rect 1470 -2820 1476 -2814
rect 1470 -2826 1476 -2820
rect 1470 -2916 1476 -2910
rect 1470 -2922 1476 -2916
rect 1470 -2928 1476 -2922
rect 1470 -2934 1476 -2928
rect 1470 -2940 1476 -2934
rect 1470 -2946 1476 -2940
rect 1470 -2952 1476 -2946
rect 1470 -2958 1476 -2952
rect 1470 -2964 1476 -2958
rect 1470 -2970 1476 -2964
rect 1470 -2976 1476 -2970
rect 1470 -2982 1476 -2976
rect 1470 -2988 1476 -2982
rect 1470 -2994 1476 -2988
rect 1470 -3000 1476 -2994
rect 1470 -3006 1476 -3000
rect 1470 -3012 1476 -3006
rect 1470 -3018 1476 -3012
rect 1470 -3024 1476 -3018
rect 1470 -3030 1476 -3024
rect 1470 -3036 1476 -3030
rect 1470 -3042 1476 -3036
rect 1470 -3048 1476 -3042
rect 1470 -3054 1476 -3048
rect 1470 -3060 1476 -3054
rect 1470 -3066 1476 -3060
rect 1470 -3072 1476 -3066
rect 1470 -3078 1476 -3072
rect 1470 -3084 1476 -3078
rect 1470 -3090 1476 -3084
rect 1470 -3096 1476 -3090
rect 1470 -3102 1476 -3096
rect 1470 -3108 1476 -3102
rect 1470 -3114 1476 -3108
rect 1470 -3120 1476 -3114
rect 1470 -3126 1476 -3120
rect 1470 -3132 1476 -3126
rect 1470 -3138 1476 -3132
rect 1470 -3144 1476 -3138
rect 1470 -3150 1476 -3144
rect 1470 -3156 1476 -3150
rect 1470 -3162 1476 -3156
rect 1470 -3168 1476 -3162
rect 1470 -3174 1476 -3168
rect 1470 -3180 1476 -3174
rect 1470 -3186 1476 -3180
rect 1470 -3192 1476 -3186
rect 1470 -3198 1476 -3192
rect 1470 -3204 1476 -3198
rect 1470 -3210 1476 -3204
rect 1470 -3216 1476 -3210
rect 1470 -3222 1476 -3216
rect 1470 -3228 1476 -3222
rect 1470 -3234 1476 -3228
rect 1470 -3288 1476 -3282
rect 1470 -3294 1476 -3288
rect 1470 -3300 1476 -3294
rect 1470 -3306 1476 -3300
rect 1470 -3312 1476 -3306
rect 1470 -3318 1476 -3312
rect 1470 -3324 1476 -3318
rect 1470 -3330 1476 -3324
rect 1470 -3336 1476 -3330
rect 1470 -3342 1476 -3336
rect 1470 -3348 1476 -3342
rect 1470 -3354 1476 -3348
rect 1470 -3360 1476 -3354
rect 1470 -3366 1476 -3360
rect 1470 -3372 1476 -3366
rect 1470 -3378 1476 -3372
rect 1470 -3384 1476 -3378
rect 1470 -3390 1476 -3384
rect 1470 -3396 1476 -3390
rect 1470 -3402 1476 -3396
rect 1470 -3408 1476 -3402
rect 1470 -3414 1476 -3408
rect 1470 -3420 1476 -3414
rect 1470 -3426 1476 -3420
rect 1470 -3432 1476 -3426
rect 1470 -3438 1476 -3432
rect 1470 -3444 1476 -3438
rect 1470 -3450 1476 -3444
rect 1470 -3456 1476 -3450
rect 1470 -3462 1476 -3456
rect 1470 -3468 1476 -3462
rect 1470 -3474 1476 -3468
rect 1470 -3480 1476 -3474
rect 1470 -3486 1476 -3480
rect 1470 -3492 1476 -3486
rect 1476 -1224 1482 -1218
rect 1476 -1230 1482 -1224
rect 1476 -1236 1482 -1230
rect 1476 -1242 1482 -1236
rect 1476 -1248 1482 -1242
rect 1476 -1254 1482 -1248
rect 1476 -1260 1482 -1254
rect 1476 -1266 1482 -1260
rect 1476 -1272 1482 -1266
rect 1476 -1278 1482 -1272
rect 1476 -1284 1482 -1278
rect 1476 -1290 1482 -1284
rect 1476 -1296 1482 -1290
rect 1476 -1302 1482 -1296
rect 1476 -1308 1482 -1302
rect 1476 -1314 1482 -1308
rect 1476 -1320 1482 -1314
rect 1476 -1326 1482 -1320
rect 1476 -1332 1482 -1326
rect 1476 -1338 1482 -1332
rect 1476 -1344 1482 -1338
rect 1476 -1350 1482 -1344
rect 1476 -1356 1482 -1350
rect 1476 -1362 1482 -1356
rect 1476 -1368 1482 -1362
rect 1476 -1374 1482 -1368
rect 1476 -1380 1482 -1374
rect 1476 -1386 1482 -1380
rect 1476 -1392 1482 -1386
rect 1476 -1398 1482 -1392
rect 1476 -1404 1482 -1398
rect 1476 -1410 1482 -1404
rect 1476 -1416 1482 -1410
rect 1476 -1422 1482 -1416
rect 1476 -1428 1482 -1422
rect 1476 -1434 1482 -1428
rect 1476 -1440 1482 -1434
rect 1476 -1446 1482 -1440
rect 1476 -1452 1482 -1446
rect 1476 -1458 1482 -1452
rect 1476 -1464 1482 -1458
rect 1476 -1470 1482 -1464
rect 1476 -1476 1482 -1470
rect 1476 -1482 1482 -1476
rect 1476 -1488 1482 -1482
rect 1476 -1494 1482 -1488
rect 1476 -1500 1482 -1494
rect 1476 -1506 1482 -1500
rect 1476 -1512 1482 -1506
rect 1476 -1518 1482 -1512
rect 1476 -1524 1482 -1518
rect 1476 -1530 1482 -1524
rect 1476 -1536 1482 -1530
rect 1476 -1542 1482 -1536
rect 1476 -1548 1482 -1542
rect 1476 -1554 1482 -1548
rect 1476 -1560 1482 -1554
rect 1476 -1566 1482 -1560
rect 1476 -1572 1482 -1566
rect 1476 -1578 1482 -1572
rect 1476 -1584 1482 -1578
rect 1476 -1590 1482 -1584
rect 1476 -1596 1482 -1590
rect 1476 -1602 1482 -1596
rect 1476 -1608 1482 -1602
rect 1476 -1614 1482 -1608
rect 1476 -1620 1482 -1614
rect 1476 -1626 1482 -1620
rect 1476 -1632 1482 -1626
rect 1476 -1638 1482 -1632
rect 1476 -1644 1482 -1638
rect 1476 -1650 1482 -1644
rect 1476 -1656 1482 -1650
rect 1476 -1662 1482 -1656
rect 1476 -1668 1482 -1662
rect 1476 -1674 1482 -1668
rect 1476 -1680 1482 -1674
rect 1476 -1686 1482 -1680
rect 1476 -1692 1482 -1686
rect 1476 -1698 1482 -1692
rect 1476 -1704 1482 -1698
rect 1476 -1710 1482 -1704
rect 1476 -1716 1482 -1710
rect 1476 -1722 1482 -1716
rect 1476 -1728 1482 -1722
rect 1476 -1734 1482 -1728
rect 1476 -1740 1482 -1734
rect 1476 -1746 1482 -1740
rect 1476 -1752 1482 -1746
rect 1476 -1758 1482 -1752
rect 1476 -1764 1482 -1758
rect 1476 -1770 1482 -1764
rect 1476 -1776 1482 -1770
rect 1476 -1782 1482 -1776
rect 1476 -1788 1482 -1782
rect 1476 -1794 1482 -1788
rect 1476 -1800 1482 -1794
rect 1476 -1806 1482 -1800
rect 1476 -1812 1482 -1806
rect 1476 -1818 1482 -1812
rect 1476 -1824 1482 -1818
rect 1476 -1830 1482 -1824
rect 1476 -1836 1482 -1830
rect 1476 -1842 1482 -1836
rect 1476 -1848 1482 -1842
rect 1476 -1854 1482 -1848
rect 1476 -1860 1482 -1854
rect 1476 -1866 1482 -1860
rect 1476 -1872 1482 -1866
rect 1476 -1878 1482 -1872
rect 1476 -1884 1482 -1878
rect 1476 -1890 1482 -1884
rect 1476 -1896 1482 -1890
rect 1476 -1902 1482 -1896
rect 1476 -1908 1482 -1902
rect 1476 -1914 1482 -1908
rect 1476 -1920 1482 -1914
rect 1476 -1926 1482 -1920
rect 1476 -1932 1482 -1926
rect 1476 -1938 1482 -1932
rect 1476 -1944 1482 -1938
rect 1476 -1950 1482 -1944
rect 1476 -1956 1482 -1950
rect 1476 -1962 1482 -1956
rect 1476 -1968 1482 -1962
rect 1476 -1974 1482 -1968
rect 1476 -1980 1482 -1974
rect 1476 -1986 1482 -1980
rect 1476 -1992 1482 -1986
rect 1476 -1998 1482 -1992
rect 1476 -2004 1482 -1998
rect 1476 -2010 1482 -2004
rect 1476 -2016 1482 -2010
rect 1476 -2022 1482 -2016
rect 1476 -2028 1482 -2022
rect 1476 -2034 1482 -2028
rect 1476 -2040 1482 -2034
rect 1476 -2046 1482 -2040
rect 1476 -2052 1482 -2046
rect 1476 -2058 1482 -2052
rect 1476 -2064 1482 -2058
rect 1476 -2070 1482 -2064
rect 1476 -2076 1482 -2070
rect 1476 -2082 1482 -2076
rect 1476 -2088 1482 -2082
rect 1476 -2094 1482 -2088
rect 1476 -2100 1482 -2094
rect 1476 -2106 1482 -2100
rect 1476 -2112 1482 -2106
rect 1476 -2118 1482 -2112
rect 1476 -2124 1482 -2118
rect 1476 -2130 1482 -2124
rect 1476 -2136 1482 -2130
rect 1476 -2142 1482 -2136
rect 1476 -2148 1482 -2142
rect 1476 -2154 1482 -2148
rect 1476 -2160 1482 -2154
rect 1476 -2166 1482 -2160
rect 1476 -2172 1482 -2166
rect 1476 -2178 1482 -2172
rect 1476 -2184 1482 -2178
rect 1476 -2190 1482 -2184
rect 1476 -2196 1482 -2190
rect 1476 -2202 1482 -2196
rect 1476 -2208 1482 -2202
rect 1476 -2214 1482 -2208
rect 1476 -2220 1482 -2214
rect 1476 -2292 1482 -2286
rect 1476 -2298 1482 -2292
rect 1476 -2304 1482 -2298
rect 1476 -2310 1482 -2304
rect 1476 -2316 1482 -2310
rect 1476 -2322 1482 -2316
rect 1476 -2328 1482 -2322
rect 1476 -2334 1482 -2328
rect 1476 -2340 1482 -2334
rect 1476 -2346 1482 -2340
rect 1476 -2352 1482 -2346
rect 1476 -2358 1482 -2352
rect 1476 -2364 1482 -2358
rect 1476 -2370 1482 -2364
rect 1476 -2376 1482 -2370
rect 1476 -2382 1482 -2376
rect 1476 -2388 1482 -2382
rect 1476 -2394 1482 -2388
rect 1476 -2400 1482 -2394
rect 1476 -2406 1482 -2400
rect 1476 -2412 1482 -2406
rect 1476 -2418 1482 -2412
rect 1476 -2424 1482 -2418
rect 1476 -2430 1482 -2424
rect 1476 -2436 1482 -2430
rect 1476 -2442 1482 -2436
rect 1476 -2448 1482 -2442
rect 1476 -2454 1482 -2448
rect 1476 -2460 1482 -2454
rect 1476 -2466 1482 -2460
rect 1476 -2472 1482 -2466
rect 1476 -2478 1482 -2472
rect 1476 -2484 1482 -2478
rect 1476 -2490 1482 -2484
rect 1476 -2496 1482 -2490
rect 1476 -2502 1482 -2496
rect 1476 -2508 1482 -2502
rect 1476 -2514 1482 -2508
rect 1476 -2520 1482 -2514
rect 1476 -2526 1482 -2520
rect 1476 -2532 1482 -2526
rect 1476 -2538 1482 -2532
rect 1476 -2544 1482 -2538
rect 1476 -2550 1482 -2544
rect 1476 -2556 1482 -2550
rect 1476 -2562 1482 -2556
rect 1476 -2568 1482 -2562
rect 1476 -2574 1482 -2568
rect 1476 -2580 1482 -2574
rect 1476 -2586 1482 -2580
rect 1476 -2592 1482 -2586
rect 1476 -2598 1482 -2592
rect 1476 -2604 1482 -2598
rect 1476 -2610 1482 -2604
rect 1476 -2616 1482 -2610
rect 1476 -2622 1482 -2616
rect 1476 -2628 1482 -2622
rect 1476 -2634 1482 -2628
rect 1476 -2640 1482 -2634
rect 1476 -2646 1482 -2640
rect 1476 -2652 1482 -2646
rect 1476 -2658 1482 -2652
rect 1476 -2664 1482 -2658
rect 1476 -2670 1482 -2664
rect 1476 -2676 1482 -2670
rect 1476 -2682 1482 -2676
rect 1476 -2688 1482 -2682
rect 1476 -2694 1482 -2688
rect 1476 -2700 1482 -2694
rect 1476 -2706 1482 -2700
rect 1476 -2712 1482 -2706
rect 1476 -2718 1482 -2712
rect 1476 -2724 1482 -2718
rect 1476 -2730 1482 -2724
rect 1476 -2736 1482 -2730
rect 1476 -2742 1482 -2736
rect 1476 -2748 1482 -2742
rect 1476 -2754 1482 -2748
rect 1476 -2760 1482 -2754
rect 1476 -2766 1482 -2760
rect 1476 -2772 1482 -2766
rect 1476 -2778 1482 -2772
rect 1476 -2784 1482 -2778
rect 1476 -2790 1482 -2784
rect 1476 -2796 1482 -2790
rect 1476 -2802 1482 -2796
rect 1476 -2808 1482 -2802
rect 1476 -2814 1482 -2808
rect 1476 -2820 1482 -2814
rect 1476 -2826 1482 -2820
rect 1476 -2910 1482 -2904
rect 1476 -2916 1482 -2910
rect 1476 -2922 1482 -2916
rect 1476 -2928 1482 -2922
rect 1476 -2934 1482 -2928
rect 1476 -2940 1482 -2934
rect 1476 -2946 1482 -2940
rect 1476 -2952 1482 -2946
rect 1476 -2958 1482 -2952
rect 1476 -2964 1482 -2958
rect 1476 -2970 1482 -2964
rect 1476 -2976 1482 -2970
rect 1476 -2982 1482 -2976
rect 1476 -2988 1482 -2982
rect 1476 -2994 1482 -2988
rect 1476 -3000 1482 -2994
rect 1476 -3006 1482 -3000
rect 1476 -3012 1482 -3006
rect 1476 -3018 1482 -3012
rect 1476 -3024 1482 -3018
rect 1476 -3030 1482 -3024
rect 1476 -3036 1482 -3030
rect 1476 -3042 1482 -3036
rect 1476 -3048 1482 -3042
rect 1476 -3054 1482 -3048
rect 1476 -3060 1482 -3054
rect 1476 -3066 1482 -3060
rect 1476 -3072 1482 -3066
rect 1476 -3078 1482 -3072
rect 1476 -3084 1482 -3078
rect 1476 -3090 1482 -3084
rect 1476 -3096 1482 -3090
rect 1476 -3102 1482 -3096
rect 1476 -3108 1482 -3102
rect 1476 -3114 1482 -3108
rect 1476 -3120 1482 -3114
rect 1476 -3126 1482 -3120
rect 1476 -3132 1482 -3126
rect 1476 -3138 1482 -3132
rect 1476 -3144 1482 -3138
rect 1476 -3150 1482 -3144
rect 1476 -3156 1482 -3150
rect 1476 -3162 1482 -3156
rect 1476 -3168 1482 -3162
rect 1476 -3174 1482 -3168
rect 1476 -3180 1482 -3174
rect 1476 -3186 1482 -3180
rect 1476 -3192 1482 -3186
rect 1476 -3198 1482 -3192
rect 1476 -3204 1482 -3198
rect 1476 -3210 1482 -3204
rect 1476 -3216 1482 -3210
rect 1476 -3222 1482 -3216
rect 1476 -3228 1482 -3222
rect 1476 -3234 1482 -3228
rect 1476 -3288 1482 -3282
rect 1476 -3294 1482 -3288
rect 1476 -3300 1482 -3294
rect 1476 -3306 1482 -3300
rect 1476 -3312 1482 -3306
rect 1476 -3318 1482 -3312
rect 1476 -3324 1482 -3318
rect 1476 -3330 1482 -3324
rect 1476 -3336 1482 -3330
rect 1476 -3342 1482 -3336
rect 1476 -3348 1482 -3342
rect 1476 -3354 1482 -3348
rect 1476 -3360 1482 -3354
rect 1476 -3366 1482 -3360
rect 1476 -3372 1482 -3366
rect 1476 -3378 1482 -3372
rect 1476 -3384 1482 -3378
rect 1476 -3390 1482 -3384
rect 1476 -3396 1482 -3390
rect 1476 -3402 1482 -3396
rect 1476 -3408 1482 -3402
rect 1476 -3414 1482 -3408
rect 1476 -3420 1482 -3414
rect 1476 -3426 1482 -3420
rect 1476 -3432 1482 -3426
rect 1476 -3438 1482 -3432
rect 1476 -3444 1482 -3438
rect 1476 -3450 1482 -3444
rect 1476 -3456 1482 -3450
rect 1476 -3462 1482 -3456
rect 1476 -3468 1482 -3462
rect 1476 -3474 1482 -3468
rect 1476 -3480 1482 -3474
rect 1476 -3486 1482 -3480
rect 1476 -3492 1482 -3486
rect 1482 -1212 1488 -1206
rect 1482 -1218 1488 -1212
rect 1482 -1224 1488 -1218
rect 1482 -1230 1488 -1224
rect 1482 -1236 1488 -1230
rect 1482 -1242 1488 -1236
rect 1482 -1248 1488 -1242
rect 1482 -1254 1488 -1248
rect 1482 -1260 1488 -1254
rect 1482 -1266 1488 -1260
rect 1482 -1272 1488 -1266
rect 1482 -1278 1488 -1272
rect 1482 -1284 1488 -1278
rect 1482 -1290 1488 -1284
rect 1482 -1296 1488 -1290
rect 1482 -1302 1488 -1296
rect 1482 -1308 1488 -1302
rect 1482 -1314 1488 -1308
rect 1482 -1320 1488 -1314
rect 1482 -1326 1488 -1320
rect 1482 -1332 1488 -1326
rect 1482 -1338 1488 -1332
rect 1482 -1344 1488 -1338
rect 1482 -1350 1488 -1344
rect 1482 -1356 1488 -1350
rect 1482 -1362 1488 -1356
rect 1482 -1368 1488 -1362
rect 1482 -1374 1488 -1368
rect 1482 -1380 1488 -1374
rect 1482 -1386 1488 -1380
rect 1482 -1392 1488 -1386
rect 1482 -1398 1488 -1392
rect 1482 -1404 1488 -1398
rect 1482 -1410 1488 -1404
rect 1482 -1416 1488 -1410
rect 1482 -1422 1488 -1416
rect 1482 -1428 1488 -1422
rect 1482 -1434 1488 -1428
rect 1482 -1440 1488 -1434
rect 1482 -1446 1488 -1440
rect 1482 -1452 1488 -1446
rect 1482 -1458 1488 -1452
rect 1482 -1464 1488 -1458
rect 1482 -1470 1488 -1464
rect 1482 -1476 1488 -1470
rect 1482 -1482 1488 -1476
rect 1482 -1488 1488 -1482
rect 1482 -1494 1488 -1488
rect 1482 -1500 1488 -1494
rect 1482 -1506 1488 -1500
rect 1482 -1512 1488 -1506
rect 1482 -1518 1488 -1512
rect 1482 -1524 1488 -1518
rect 1482 -1530 1488 -1524
rect 1482 -1536 1488 -1530
rect 1482 -1542 1488 -1536
rect 1482 -1548 1488 -1542
rect 1482 -1554 1488 -1548
rect 1482 -1560 1488 -1554
rect 1482 -1566 1488 -1560
rect 1482 -1572 1488 -1566
rect 1482 -1578 1488 -1572
rect 1482 -1584 1488 -1578
rect 1482 -1590 1488 -1584
rect 1482 -1596 1488 -1590
rect 1482 -1602 1488 -1596
rect 1482 -1608 1488 -1602
rect 1482 -1614 1488 -1608
rect 1482 -1620 1488 -1614
rect 1482 -1626 1488 -1620
rect 1482 -1632 1488 -1626
rect 1482 -1638 1488 -1632
rect 1482 -1644 1488 -1638
rect 1482 -1650 1488 -1644
rect 1482 -1656 1488 -1650
rect 1482 -1662 1488 -1656
rect 1482 -1668 1488 -1662
rect 1482 -1674 1488 -1668
rect 1482 -1680 1488 -1674
rect 1482 -1686 1488 -1680
rect 1482 -1692 1488 -1686
rect 1482 -1698 1488 -1692
rect 1482 -1704 1488 -1698
rect 1482 -1710 1488 -1704
rect 1482 -1716 1488 -1710
rect 1482 -1722 1488 -1716
rect 1482 -1728 1488 -1722
rect 1482 -1734 1488 -1728
rect 1482 -1740 1488 -1734
rect 1482 -1746 1488 -1740
rect 1482 -1752 1488 -1746
rect 1482 -1758 1488 -1752
rect 1482 -1764 1488 -1758
rect 1482 -1770 1488 -1764
rect 1482 -1776 1488 -1770
rect 1482 -1782 1488 -1776
rect 1482 -1788 1488 -1782
rect 1482 -1794 1488 -1788
rect 1482 -1800 1488 -1794
rect 1482 -1806 1488 -1800
rect 1482 -1812 1488 -1806
rect 1482 -1818 1488 -1812
rect 1482 -1824 1488 -1818
rect 1482 -1830 1488 -1824
rect 1482 -1836 1488 -1830
rect 1482 -1842 1488 -1836
rect 1482 -1848 1488 -1842
rect 1482 -1854 1488 -1848
rect 1482 -1860 1488 -1854
rect 1482 -1866 1488 -1860
rect 1482 -1872 1488 -1866
rect 1482 -1878 1488 -1872
rect 1482 -1884 1488 -1878
rect 1482 -1890 1488 -1884
rect 1482 -1896 1488 -1890
rect 1482 -1902 1488 -1896
rect 1482 -1908 1488 -1902
rect 1482 -1914 1488 -1908
rect 1482 -1920 1488 -1914
rect 1482 -1926 1488 -1920
rect 1482 -1932 1488 -1926
rect 1482 -1938 1488 -1932
rect 1482 -1944 1488 -1938
rect 1482 -1950 1488 -1944
rect 1482 -1956 1488 -1950
rect 1482 -1962 1488 -1956
rect 1482 -1968 1488 -1962
rect 1482 -1974 1488 -1968
rect 1482 -1980 1488 -1974
rect 1482 -1986 1488 -1980
rect 1482 -1992 1488 -1986
rect 1482 -1998 1488 -1992
rect 1482 -2004 1488 -1998
rect 1482 -2010 1488 -2004
rect 1482 -2016 1488 -2010
rect 1482 -2022 1488 -2016
rect 1482 -2028 1488 -2022
rect 1482 -2034 1488 -2028
rect 1482 -2040 1488 -2034
rect 1482 -2046 1488 -2040
rect 1482 -2052 1488 -2046
rect 1482 -2058 1488 -2052
rect 1482 -2064 1488 -2058
rect 1482 -2070 1488 -2064
rect 1482 -2076 1488 -2070
rect 1482 -2082 1488 -2076
rect 1482 -2088 1488 -2082
rect 1482 -2094 1488 -2088
rect 1482 -2100 1488 -2094
rect 1482 -2106 1488 -2100
rect 1482 -2112 1488 -2106
rect 1482 -2118 1488 -2112
rect 1482 -2124 1488 -2118
rect 1482 -2130 1488 -2124
rect 1482 -2136 1488 -2130
rect 1482 -2142 1488 -2136
rect 1482 -2148 1488 -2142
rect 1482 -2154 1488 -2148
rect 1482 -2160 1488 -2154
rect 1482 -2166 1488 -2160
rect 1482 -2172 1488 -2166
rect 1482 -2178 1488 -2172
rect 1482 -2184 1488 -2178
rect 1482 -2190 1488 -2184
rect 1482 -2196 1488 -2190
rect 1482 -2202 1488 -2196
rect 1482 -2208 1488 -2202
rect 1482 -2214 1488 -2208
rect 1482 -2286 1488 -2280
rect 1482 -2292 1488 -2286
rect 1482 -2298 1488 -2292
rect 1482 -2304 1488 -2298
rect 1482 -2310 1488 -2304
rect 1482 -2316 1488 -2310
rect 1482 -2322 1488 -2316
rect 1482 -2328 1488 -2322
rect 1482 -2334 1488 -2328
rect 1482 -2340 1488 -2334
rect 1482 -2346 1488 -2340
rect 1482 -2352 1488 -2346
rect 1482 -2358 1488 -2352
rect 1482 -2364 1488 -2358
rect 1482 -2370 1488 -2364
rect 1482 -2376 1488 -2370
rect 1482 -2382 1488 -2376
rect 1482 -2388 1488 -2382
rect 1482 -2394 1488 -2388
rect 1482 -2400 1488 -2394
rect 1482 -2406 1488 -2400
rect 1482 -2412 1488 -2406
rect 1482 -2418 1488 -2412
rect 1482 -2424 1488 -2418
rect 1482 -2430 1488 -2424
rect 1482 -2436 1488 -2430
rect 1482 -2442 1488 -2436
rect 1482 -2448 1488 -2442
rect 1482 -2454 1488 -2448
rect 1482 -2460 1488 -2454
rect 1482 -2466 1488 -2460
rect 1482 -2472 1488 -2466
rect 1482 -2478 1488 -2472
rect 1482 -2484 1488 -2478
rect 1482 -2490 1488 -2484
rect 1482 -2496 1488 -2490
rect 1482 -2502 1488 -2496
rect 1482 -2508 1488 -2502
rect 1482 -2514 1488 -2508
rect 1482 -2520 1488 -2514
rect 1482 -2526 1488 -2520
rect 1482 -2532 1488 -2526
rect 1482 -2538 1488 -2532
rect 1482 -2544 1488 -2538
rect 1482 -2550 1488 -2544
rect 1482 -2556 1488 -2550
rect 1482 -2562 1488 -2556
rect 1482 -2568 1488 -2562
rect 1482 -2574 1488 -2568
rect 1482 -2580 1488 -2574
rect 1482 -2586 1488 -2580
rect 1482 -2592 1488 -2586
rect 1482 -2598 1488 -2592
rect 1482 -2604 1488 -2598
rect 1482 -2610 1488 -2604
rect 1482 -2616 1488 -2610
rect 1482 -2622 1488 -2616
rect 1482 -2628 1488 -2622
rect 1482 -2634 1488 -2628
rect 1482 -2640 1488 -2634
rect 1482 -2646 1488 -2640
rect 1482 -2652 1488 -2646
rect 1482 -2658 1488 -2652
rect 1482 -2664 1488 -2658
rect 1482 -2670 1488 -2664
rect 1482 -2676 1488 -2670
rect 1482 -2682 1488 -2676
rect 1482 -2688 1488 -2682
rect 1482 -2694 1488 -2688
rect 1482 -2700 1488 -2694
rect 1482 -2706 1488 -2700
rect 1482 -2712 1488 -2706
rect 1482 -2718 1488 -2712
rect 1482 -2724 1488 -2718
rect 1482 -2730 1488 -2724
rect 1482 -2736 1488 -2730
rect 1482 -2742 1488 -2736
rect 1482 -2748 1488 -2742
rect 1482 -2754 1488 -2748
rect 1482 -2760 1488 -2754
rect 1482 -2766 1488 -2760
rect 1482 -2772 1488 -2766
rect 1482 -2778 1488 -2772
rect 1482 -2784 1488 -2778
rect 1482 -2790 1488 -2784
rect 1482 -2796 1488 -2790
rect 1482 -2802 1488 -2796
rect 1482 -2808 1488 -2802
rect 1482 -2814 1488 -2808
rect 1482 -2820 1488 -2814
rect 1482 -2904 1488 -2898
rect 1482 -2910 1488 -2904
rect 1482 -2916 1488 -2910
rect 1482 -2922 1488 -2916
rect 1482 -2928 1488 -2922
rect 1482 -2934 1488 -2928
rect 1482 -2940 1488 -2934
rect 1482 -2946 1488 -2940
rect 1482 -2952 1488 -2946
rect 1482 -2958 1488 -2952
rect 1482 -2964 1488 -2958
rect 1482 -2970 1488 -2964
rect 1482 -2976 1488 -2970
rect 1482 -2982 1488 -2976
rect 1482 -2988 1488 -2982
rect 1482 -2994 1488 -2988
rect 1482 -3000 1488 -2994
rect 1482 -3006 1488 -3000
rect 1482 -3012 1488 -3006
rect 1482 -3018 1488 -3012
rect 1482 -3024 1488 -3018
rect 1482 -3030 1488 -3024
rect 1482 -3036 1488 -3030
rect 1482 -3042 1488 -3036
rect 1482 -3048 1488 -3042
rect 1482 -3054 1488 -3048
rect 1482 -3060 1488 -3054
rect 1482 -3066 1488 -3060
rect 1482 -3072 1488 -3066
rect 1482 -3078 1488 -3072
rect 1482 -3084 1488 -3078
rect 1482 -3090 1488 -3084
rect 1482 -3096 1488 -3090
rect 1482 -3102 1488 -3096
rect 1482 -3108 1488 -3102
rect 1482 -3114 1488 -3108
rect 1482 -3120 1488 -3114
rect 1482 -3126 1488 -3120
rect 1482 -3132 1488 -3126
rect 1482 -3138 1488 -3132
rect 1482 -3144 1488 -3138
rect 1482 -3150 1488 -3144
rect 1482 -3156 1488 -3150
rect 1482 -3162 1488 -3156
rect 1482 -3168 1488 -3162
rect 1482 -3174 1488 -3168
rect 1482 -3180 1488 -3174
rect 1482 -3186 1488 -3180
rect 1482 -3192 1488 -3186
rect 1482 -3198 1488 -3192
rect 1482 -3204 1488 -3198
rect 1482 -3210 1488 -3204
rect 1482 -3216 1488 -3210
rect 1482 -3222 1488 -3216
rect 1482 -3228 1488 -3222
rect 1482 -3234 1488 -3228
rect 1482 -3282 1488 -3276
rect 1482 -3288 1488 -3282
rect 1482 -3294 1488 -3288
rect 1482 -3300 1488 -3294
rect 1482 -3306 1488 -3300
rect 1482 -3312 1488 -3306
rect 1482 -3318 1488 -3312
rect 1482 -3324 1488 -3318
rect 1482 -3330 1488 -3324
rect 1482 -3336 1488 -3330
rect 1482 -3342 1488 -3336
rect 1482 -3348 1488 -3342
rect 1482 -3354 1488 -3348
rect 1482 -3360 1488 -3354
rect 1482 -3366 1488 -3360
rect 1482 -3372 1488 -3366
rect 1482 -3378 1488 -3372
rect 1482 -3384 1488 -3378
rect 1482 -3390 1488 -3384
rect 1482 -3396 1488 -3390
rect 1482 -3402 1488 -3396
rect 1482 -3408 1488 -3402
rect 1482 -3414 1488 -3408
rect 1482 -3420 1488 -3414
rect 1482 -3426 1488 -3420
rect 1482 -3432 1488 -3426
rect 1482 -3438 1488 -3432
rect 1482 -3444 1488 -3438
rect 1482 -3450 1488 -3444
rect 1482 -3456 1488 -3450
rect 1482 -3462 1488 -3456
rect 1482 -3468 1488 -3462
rect 1482 -3474 1488 -3468
rect 1482 -3480 1488 -3474
rect 1482 -3486 1488 -3480
rect 1482 -3492 1488 -3486
rect 1488 -1200 1494 -1194
rect 1488 -1206 1494 -1200
rect 1488 -1212 1494 -1206
rect 1488 -1218 1494 -1212
rect 1488 -1224 1494 -1218
rect 1488 -1230 1494 -1224
rect 1488 -1236 1494 -1230
rect 1488 -1242 1494 -1236
rect 1488 -1248 1494 -1242
rect 1488 -1254 1494 -1248
rect 1488 -1260 1494 -1254
rect 1488 -1266 1494 -1260
rect 1488 -1272 1494 -1266
rect 1488 -1278 1494 -1272
rect 1488 -1284 1494 -1278
rect 1488 -1290 1494 -1284
rect 1488 -1296 1494 -1290
rect 1488 -1302 1494 -1296
rect 1488 -1308 1494 -1302
rect 1488 -1314 1494 -1308
rect 1488 -1320 1494 -1314
rect 1488 -1326 1494 -1320
rect 1488 -1332 1494 -1326
rect 1488 -1338 1494 -1332
rect 1488 -1344 1494 -1338
rect 1488 -1350 1494 -1344
rect 1488 -1356 1494 -1350
rect 1488 -1362 1494 -1356
rect 1488 -1368 1494 -1362
rect 1488 -1374 1494 -1368
rect 1488 -1380 1494 -1374
rect 1488 -1386 1494 -1380
rect 1488 -1392 1494 -1386
rect 1488 -1398 1494 -1392
rect 1488 -1404 1494 -1398
rect 1488 -1410 1494 -1404
rect 1488 -1416 1494 -1410
rect 1488 -1422 1494 -1416
rect 1488 -1428 1494 -1422
rect 1488 -1434 1494 -1428
rect 1488 -1440 1494 -1434
rect 1488 -1446 1494 -1440
rect 1488 -1452 1494 -1446
rect 1488 -1458 1494 -1452
rect 1488 -1464 1494 -1458
rect 1488 -1470 1494 -1464
rect 1488 -1476 1494 -1470
rect 1488 -1482 1494 -1476
rect 1488 -1488 1494 -1482
rect 1488 -1494 1494 -1488
rect 1488 -1500 1494 -1494
rect 1488 -1506 1494 -1500
rect 1488 -1512 1494 -1506
rect 1488 -1518 1494 -1512
rect 1488 -1524 1494 -1518
rect 1488 -1530 1494 -1524
rect 1488 -1536 1494 -1530
rect 1488 -1542 1494 -1536
rect 1488 -1548 1494 -1542
rect 1488 -1554 1494 -1548
rect 1488 -1560 1494 -1554
rect 1488 -1566 1494 -1560
rect 1488 -1572 1494 -1566
rect 1488 -1578 1494 -1572
rect 1488 -1584 1494 -1578
rect 1488 -1590 1494 -1584
rect 1488 -1596 1494 -1590
rect 1488 -1602 1494 -1596
rect 1488 -1608 1494 -1602
rect 1488 -1614 1494 -1608
rect 1488 -1620 1494 -1614
rect 1488 -1626 1494 -1620
rect 1488 -1632 1494 -1626
rect 1488 -1638 1494 -1632
rect 1488 -1644 1494 -1638
rect 1488 -1650 1494 -1644
rect 1488 -1656 1494 -1650
rect 1488 -1662 1494 -1656
rect 1488 -1668 1494 -1662
rect 1488 -1674 1494 -1668
rect 1488 -1680 1494 -1674
rect 1488 -1686 1494 -1680
rect 1488 -1692 1494 -1686
rect 1488 -1698 1494 -1692
rect 1488 -1704 1494 -1698
rect 1488 -1710 1494 -1704
rect 1488 -1716 1494 -1710
rect 1488 -1722 1494 -1716
rect 1488 -1728 1494 -1722
rect 1488 -1734 1494 -1728
rect 1488 -1740 1494 -1734
rect 1488 -1746 1494 -1740
rect 1488 -1752 1494 -1746
rect 1488 -1758 1494 -1752
rect 1488 -1764 1494 -1758
rect 1488 -1770 1494 -1764
rect 1488 -1776 1494 -1770
rect 1488 -1782 1494 -1776
rect 1488 -1788 1494 -1782
rect 1488 -1794 1494 -1788
rect 1488 -1800 1494 -1794
rect 1488 -1806 1494 -1800
rect 1488 -1812 1494 -1806
rect 1488 -1818 1494 -1812
rect 1488 -1824 1494 -1818
rect 1488 -1830 1494 -1824
rect 1488 -1836 1494 -1830
rect 1488 -1842 1494 -1836
rect 1488 -1848 1494 -1842
rect 1488 -1854 1494 -1848
rect 1488 -1860 1494 -1854
rect 1488 -1866 1494 -1860
rect 1488 -1872 1494 -1866
rect 1488 -1878 1494 -1872
rect 1488 -1884 1494 -1878
rect 1488 -1890 1494 -1884
rect 1488 -1896 1494 -1890
rect 1488 -1902 1494 -1896
rect 1488 -1908 1494 -1902
rect 1488 -1914 1494 -1908
rect 1488 -1920 1494 -1914
rect 1488 -1926 1494 -1920
rect 1488 -1932 1494 -1926
rect 1488 -1938 1494 -1932
rect 1488 -1944 1494 -1938
rect 1488 -1950 1494 -1944
rect 1488 -1956 1494 -1950
rect 1488 -1962 1494 -1956
rect 1488 -1968 1494 -1962
rect 1488 -1974 1494 -1968
rect 1488 -1980 1494 -1974
rect 1488 -1986 1494 -1980
rect 1488 -1992 1494 -1986
rect 1488 -1998 1494 -1992
rect 1488 -2004 1494 -1998
rect 1488 -2010 1494 -2004
rect 1488 -2016 1494 -2010
rect 1488 -2022 1494 -2016
rect 1488 -2028 1494 -2022
rect 1488 -2034 1494 -2028
rect 1488 -2040 1494 -2034
rect 1488 -2046 1494 -2040
rect 1488 -2052 1494 -2046
rect 1488 -2058 1494 -2052
rect 1488 -2064 1494 -2058
rect 1488 -2070 1494 -2064
rect 1488 -2076 1494 -2070
rect 1488 -2082 1494 -2076
rect 1488 -2088 1494 -2082
rect 1488 -2094 1494 -2088
rect 1488 -2100 1494 -2094
rect 1488 -2106 1494 -2100
rect 1488 -2112 1494 -2106
rect 1488 -2118 1494 -2112
rect 1488 -2124 1494 -2118
rect 1488 -2130 1494 -2124
rect 1488 -2136 1494 -2130
rect 1488 -2142 1494 -2136
rect 1488 -2148 1494 -2142
rect 1488 -2154 1494 -2148
rect 1488 -2160 1494 -2154
rect 1488 -2166 1494 -2160
rect 1488 -2172 1494 -2166
rect 1488 -2178 1494 -2172
rect 1488 -2184 1494 -2178
rect 1488 -2190 1494 -2184
rect 1488 -2196 1494 -2190
rect 1488 -2202 1494 -2196
rect 1488 -2208 1494 -2202
rect 1488 -2280 1494 -2274
rect 1488 -2286 1494 -2280
rect 1488 -2292 1494 -2286
rect 1488 -2298 1494 -2292
rect 1488 -2304 1494 -2298
rect 1488 -2310 1494 -2304
rect 1488 -2316 1494 -2310
rect 1488 -2322 1494 -2316
rect 1488 -2328 1494 -2322
rect 1488 -2334 1494 -2328
rect 1488 -2340 1494 -2334
rect 1488 -2346 1494 -2340
rect 1488 -2352 1494 -2346
rect 1488 -2358 1494 -2352
rect 1488 -2364 1494 -2358
rect 1488 -2370 1494 -2364
rect 1488 -2376 1494 -2370
rect 1488 -2382 1494 -2376
rect 1488 -2388 1494 -2382
rect 1488 -2394 1494 -2388
rect 1488 -2400 1494 -2394
rect 1488 -2406 1494 -2400
rect 1488 -2412 1494 -2406
rect 1488 -2418 1494 -2412
rect 1488 -2424 1494 -2418
rect 1488 -2430 1494 -2424
rect 1488 -2436 1494 -2430
rect 1488 -2442 1494 -2436
rect 1488 -2448 1494 -2442
rect 1488 -2454 1494 -2448
rect 1488 -2460 1494 -2454
rect 1488 -2466 1494 -2460
rect 1488 -2472 1494 -2466
rect 1488 -2478 1494 -2472
rect 1488 -2484 1494 -2478
rect 1488 -2490 1494 -2484
rect 1488 -2496 1494 -2490
rect 1488 -2502 1494 -2496
rect 1488 -2508 1494 -2502
rect 1488 -2514 1494 -2508
rect 1488 -2520 1494 -2514
rect 1488 -2526 1494 -2520
rect 1488 -2532 1494 -2526
rect 1488 -2538 1494 -2532
rect 1488 -2544 1494 -2538
rect 1488 -2550 1494 -2544
rect 1488 -2556 1494 -2550
rect 1488 -2562 1494 -2556
rect 1488 -2568 1494 -2562
rect 1488 -2574 1494 -2568
rect 1488 -2580 1494 -2574
rect 1488 -2586 1494 -2580
rect 1488 -2592 1494 -2586
rect 1488 -2598 1494 -2592
rect 1488 -2604 1494 -2598
rect 1488 -2610 1494 -2604
rect 1488 -2616 1494 -2610
rect 1488 -2622 1494 -2616
rect 1488 -2628 1494 -2622
rect 1488 -2634 1494 -2628
rect 1488 -2640 1494 -2634
rect 1488 -2646 1494 -2640
rect 1488 -2652 1494 -2646
rect 1488 -2658 1494 -2652
rect 1488 -2664 1494 -2658
rect 1488 -2670 1494 -2664
rect 1488 -2676 1494 -2670
rect 1488 -2682 1494 -2676
rect 1488 -2688 1494 -2682
rect 1488 -2694 1494 -2688
rect 1488 -2700 1494 -2694
rect 1488 -2706 1494 -2700
rect 1488 -2712 1494 -2706
rect 1488 -2718 1494 -2712
rect 1488 -2724 1494 -2718
rect 1488 -2730 1494 -2724
rect 1488 -2736 1494 -2730
rect 1488 -2742 1494 -2736
rect 1488 -2748 1494 -2742
rect 1488 -2754 1494 -2748
rect 1488 -2760 1494 -2754
rect 1488 -2766 1494 -2760
rect 1488 -2772 1494 -2766
rect 1488 -2778 1494 -2772
rect 1488 -2784 1494 -2778
rect 1488 -2790 1494 -2784
rect 1488 -2796 1494 -2790
rect 1488 -2802 1494 -2796
rect 1488 -2808 1494 -2802
rect 1488 -2814 1494 -2808
rect 1488 -2904 1494 -2898
rect 1488 -2910 1494 -2904
rect 1488 -2916 1494 -2910
rect 1488 -2922 1494 -2916
rect 1488 -2928 1494 -2922
rect 1488 -2934 1494 -2928
rect 1488 -2940 1494 -2934
rect 1488 -2946 1494 -2940
rect 1488 -2952 1494 -2946
rect 1488 -2958 1494 -2952
rect 1488 -2964 1494 -2958
rect 1488 -2970 1494 -2964
rect 1488 -2976 1494 -2970
rect 1488 -2982 1494 -2976
rect 1488 -2988 1494 -2982
rect 1488 -2994 1494 -2988
rect 1488 -3000 1494 -2994
rect 1488 -3006 1494 -3000
rect 1488 -3012 1494 -3006
rect 1488 -3018 1494 -3012
rect 1488 -3024 1494 -3018
rect 1488 -3030 1494 -3024
rect 1488 -3036 1494 -3030
rect 1488 -3042 1494 -3036
rect 1488 -3048 1494 -3042
rect 1488 -3054 1494 -3048
rect 1488 -3060 1494 -3054
rect 1488 -3066 1494 -3060
rect 1488 -3072 1494 -3066
rect 1488 -3078 1494 -3072
rect 1488 -3084 1494 -3078
rect 1488 -3090 1494 -3084
rect 1488 -3096 1494 -3090
rect 1488 -3102 1494 -3096
rect 1488 -3108 1494 -3102
rect 1488 -3114 1494 -3108
rect 1488 -3120 1494 -3114
rect 1488 -3126 1494 -3120
rect 1488 -3132 1494 -3126
rect 1488 -3138 1494 -3132
rect 1488 -3144 1494 -3138
rect 1488 -3150 1494 -3144
rect 1488 -3156 1494 -3150
rect 1488 -3162 1494 -3156
rect 1488 -3168 1494 -3162
rect 1488 -3174 1494 -3168
rect 1488 -3180 1494 -3174
rect 1488 -3186 1494 -3180
rect 1488 -3192 1494 -3186
rect 1488 -3198 1494 -3192
rect 1488 -3204 1494 -3198
rect 1488 -3210 1494 -3204
rect 1488 -3216 1494 -3210
rect 1488 -3222 1494 -3216
rect 1488 -3228 1494 -3222
rect 1488 -3234 1494 -3228
rect 1488 -3282 1494 -3276
rect 1488 -3288 1494 -3282
rect 1488 -3294 1494 -3288
rect 1488 -3300 1494 -3294
rect 1488 -3306 1494 -3300
rect 1488 -3312 1494 -3306
rect 1488 -3318 1494 -3312
rect 1488 -3324 1494 -3318
rect 1488 -3330 1494 -3324
rect 1488 -3336 1494 -3330
rect 1488 -3342 1494 -3336
rect 1488 -3348 1494 -3342
rect 1488 -3354 1494 -3348
rect 1488 -3360 1494 -3354
rect 1488 -3366 1494 -3360
rect 1488 -3372 1494 -3366
rect 1488 -3378 1494 -3372
rect 1488 -3384 1494 -3378
rect 1488 -3390 1494 -3384
rect 1488 -3396 1494 -3390
rect 1488 -3402 1494 -3396
rect 1488 -3408 1494 -3402
rect 1488 -3414 1494 -3408
rect 1488 -3420 1494 -3414
rect 1488 -3426 1494 -3420
rect 1488 -3432 1494 -3426
rect 1488 -3438 1494 -3432
rect 1488 -3444 1494 -3438
rect 1488 -3450 1494 -3444
rect 1488 -3456 1494 -3450
rect 1488 -3462 1494 -3456
rect 1488 -3468 1494 -3462
rect 1488 -3474 1494 -3468
rect 1488 -3480 1494 -3474
rect 1488 -3486 1494 -3480
rect 1488 -3492 1494 -3486
rect 1494 -1188 1500 -1182
rect 1494 -1194 1500 -1188
rect 1494 -1200 1500 -1194
rect 1494 -1206 1500 -1200
rect 1494 -1212 1500 -1206
rect 1494 -1218 1500 -1212
rect 1494 -1224 1500 -1218
rect 1494 -1230 1500 -1224
rect 1494 -1236 1500 -1230
rect 1494 -1242 1500 -1236
rect 1494 -1248 1500 -1242
rect 1494 -1254 1500 -1248
rect 1494 -1260 1500 -1254
rect 1494 -1266 1500 -1260
rect 1494 -1272 1500 -1266
rect 1494 -1278 1500 -1272
rect 1494 -1284 1500 -1278
rect 1494 -1290 1500 -1284
rect 1494 -1296 1500 -1290
rect 1494 -1302 1500 -1296
rect 1494 -1308 1500 -1302
rect 1494 -1314 1500 -1308
rect 1494 -1320 1500 -1314
rect 1494 -1326 1500 -1320
rect 1494 -1332 1500 -1326
rect 1494 -1338 1500 -1332
rect 1494 -1344 1500 -1338
rect 1494 -1350 1500 -1344
rect 1494 -1356 1500 -1350
rect 1494 -1362 1500 -1356
rect 1494 -1368 1500 -1362
rect 1494 -1374 1500 -1368
rect 1494 -1380 1500 -1374
rect 1494 -1386 1500 -1380
rect 1494 -1392 1500 -1386
rect 1494 -1398 1500 -1392
rect 1494 -1404 1500 -1398
rect 1494 -1410 1500 -1404
rect 1494 -1416 1500 -1410
rect 1494 -1422 1500 -1416
rect 1494 -1428 1500 -1422
rect 1494 -1434 1500 -1428
rect 1494 -1440 1500 -1434
rect 1494 -1446 1500 -1440
rect 1494 -1452 1500 -1446
rect 1494 -1458 1500 -1452
rect 1494 -1464 1500 -1458
rect 1494 -1470 1500 -1464
rect 1494 -1476 1500 -1470
rect 1494 -1482 1500 -1476
rect 1494 -1488 1500 -1482
rect 1494 -1494 1500 -1488
rect 1494 -1500 1500 -1494
rect 1494 -1506 1500 -1500
rect 1494 -1512 1500 -1506
rect 1494 -1518 1500 -1512
rect 1494 -1524 1500 -1518
rect 1494 -1530 1500 -1524
rect 1494 -1536 1500 -1530
rect 1494 -1542 1500 -1536
rect 1494 -1548 1500 -1542
rect 1494 -1554 1500 -1548
rect 1494 -1560 1500 -1554
rect 1494 -1566 1500 -1560
rect 1494 -1572 1500 -1566
rect 1494 -1578 1500 -1572
rect 1494 -1584 1500 -1578
rect 1494 -1590 1500 -1584
rect 1494 -1596 1500 -1590
rect 1494 -1602 1500 -1596
rect 1494 -1608 1500 -1602
rect 1494 -1614 1500 -1608
rect 1494 -1620 1500 -1614
rect 1494 -1626 1500 -1620
rect 1494 -1632 1500 -1626
rect 1494 -1638 1500 -1632
rect 1494 -1644 1500 -1638
rect 1494 -1650 1500 -1644
rect 1494 -1656 1500 -1650
rect 1494 -1662 1500 -1656
rect 1494 -1668 1500 -1662
rect 1494 -1674 1500 -1668
rect 1494 -1680 1500 -1674
rect 1494 -1686 1500 -1680
rect 1494 -1692 1500 -1686
rect 1494 -1698 1500 -1692
rect 1494 -1704 1500 -1698
rect 1494 -1710 1500 -1704
rect 1494 -1716 1500 -1710
rect 1494 -1722 1500 -1716
rect 1494 -1728 1500 -1722
rect 1494 -1734 1500 -1728
rect 1494 -1740 1500 -1734
rect 1494 -1746 1500 -1740
rect 1494 -1752 1500 -1746
rect 1494 -1758 1500 -1752
rect 1494 -1764 1500 -1758
rect 1494 -1770 1500 -1764
rect 1494 -1776 1500 -1770
rect 1494 -1782 1500 -1776
rect 1494 -1788 1500 -1782
rect 1494 -1794 1500 -1788
rect 1494 -1800 1500 -1794
rect 1494 -1806 1500 -1800
rect 1494 -1812 1500 -1806
rect 1494 -1818 1500 -1812
rect 1494 -1824 1500 -1818
rect 1494 -1830 1500 -1824
rect 1494 -1836 1500 -1830
rect 1494 -1842 1500 -1836
rect 1494 -1848 1500 -1842
rect 1494 -1854 1500 -1848
rect 1494 -1860 1500 -1854
rect 1494 -1866 1500 -1860
rect 1494 -1872 1500 -1866
rect 1494 -1878 1500 -1872
rect 1494 -1884 1500 -1878
rect 1494 -1890 1500 -1884
rect 1494 -1896 1500 -1890
rect 1494 -1902 1500 -1896
rect 1494 -1908 1500 -1902
rect 1494 -1914 1500 -1908
rect 1494 -1920 1500 -1914
rect 1494 -1926 1500 -1920
rect 1494 -1932 1500 -1926
rect 1494 -1938 1500 -1932
rect 1494 -1944 1500 -1938
rect 1494 -1950 1500 -1944
rect 1494 -1956 1500 -1950
rect 1494 -1962 1500 -1956
rect 1494 -1968 1500 -1962
rect 1494 -1974 1500 -1968
rect 1494 -1980 1500 -1974
rect 1494 -1986 1500 -1980
rect 1494 -1992 1500 -1986
rect 1494 -1998 1500 -1992
rect 1494 -2004 1500 -1998
rect 1494 -2010 1500 -2004
rect 1494 -2016 1500 -2010
rect 1494 -2022 1500 -2016
rect 1494 -2028 1500 -2022
rect 1494 -2034 1500 -2028
rect 1494 -2040 1500 -2034
rect 1494 -2046 1500 -2040
rect 1494 -2052 1500 -2046
rect 1494 -2058 1500 -2052
rect 1494 -2064 1500 -2058
rect 1494 -2070 1500 -2064
rect 1494 -2076 1500 -2070
rect 1494 -2082 1500 -2076
rect 1494 -2088 1500 -2082
rect 1494 -2094 1500 -2088
rect 1494 -2100 1500 -2094
rect 1494 -2106 1500 -2100
rect 1494 -2112 1500 -2106
rect 1494 -2118 1500 -2112
rect 1494 -2124 1500 -2118
rect 1494 -2130 1500 -2124
rect 1494 -2136 1500 -2130
rect 1494 -2142 1500 -2136
rect 1494 -2148 1500 -2142
rect 1494 -2154 1500 -2148
rect 1494 -2160 1500 -2154
rect 1494 -2166 1500 -2160
rect 1494 -2172 1500 -2166
rect 1494 -2178 1500 -2172
rect 1494 -2184 1500 -2178
rect 1494 -2190 1500 -2184
rect 1494 -2196 1500 -2190
rect 1494 -2274 1500 -2268
rect 1494 -2280 1500 -2274
rect 1494 -2286 1500 -2280
rect 1494 -2292 1500 -2286
rect 1494 -2298 1500 -2292
rect 1494 -2304 1500 -2298
rect 1494 -2310 1500 -2304
rect 1494 -2316 1500 -2310
rect 1494 -2322 1500 -2316
rect 1494 -2328 1500 -2322
rect 1494 -2334 1500 -2328
rect 1494 -2340 1500 -2334
rect 1494 -2346 1500 -2340
rect 1494 -2352 1500 -2346
rect 1494 -2358 1500 -2352
rect 1494 -2364 1500 -2358
rect 1494 -2370 1500 -2364
rect 1494 -2376 1500 -2370
rect 1494 -2382 1500 -2376
rect 1494 -2388 1500 -2382
rect 1494 -2394 1500 -2388
rect 1494 -2400 1500 -2394
rect 1494 -2406 1500 -2400
rect 1494 -2412 1500 -2406
rect 1494 -2418 1500 -2412
rect 1494 -2424 1500 -2418
rect 1494 -2430 1500 -2424
rect 1494 -2436 1500 -2430
rect 1494 -2442 1500 -2436
rect 1494 -2448 1500 -2442
rect 1494 -2454 1500 -2448
rect 1494 -2460 1500 -2454
rect 1494 -2466 1500 -2460
rect 1494 -2472 1500 -2466
rect 1494 -2478 1500 -2472
rect 1494 -2484 1500 -2478
rect 1494 -2490 1500 -2484
rect 1494 -2496 1500 -2490
rect 1494 -2502 1500 -2496
rect 1494 -2508 1500 -2502
rect 1494 -2514 1500 -2508
rect 1494 -2520 1500 -2514
rect 1494 -2526 1500 -2520
rect 1494 -2532 1500 -2526
rect 1494 -2538 1500 -2532
rect 1494 -2544 1500 -2538
rect 1494 -2550 1500 -2544
rect 1494 -2556 1500 -2550
rect 1494 -2562 1500 -2556
rect 1494 -2568 1500 -2562
rect 1494 -2574 1500 -2568
rect 1494 -2580 1500 -2574
rect 1494 -2586 1500 -2580
rect 1494 -2592 1500 -2586
rect 1494 -2598 1500 -2592
rect 1494 -2604 1500 -2598
rect 1494 -2610 1500 -2604
rect 1494 -2616 1500 -2610
rect 1494 -2622 1500 -2616
rect 1494 -2628 1500 -2622
rect 1494 -2634 1500 -2628
rect 1494 -2640 1500 -2634
rect 1494 -2646 1500 -2640
rect 1494 -2652 1500 -2646
rect 1494 -2658 1500 -2652
rect 1494 -2664 1500 -2658
rect 1494 -2670 1500 -2664
rect 1494 -2676 1500 -2670
rect 1494 -2682 1500 -2676
rect 1494 -2688 1500 -2682
rect 1494 -2694 1500 -2688
rect 1494 -2700 1500 -2694
rect 1494 -2706 1500 -2700
rect 1494 -2712 1500 -2706
rect 1494 -2718 1500 -2712
rect 1494 -2724 1500 -2718
rect 1494 -2730 1500 -2724
rect 1494 -2736 1500 -2730
rect 1494 -2742 1500 -2736
rect 1494 -2748 1500 -2742
rect 1494 -2754 1500 -2748
rect 1494 -2760 1500 -2754
rect 1494 -2766 1500 -2760
rect 1494 -2772 1500 -2766
rect 1494 -2778 1500 -2772
rect 1494 -2784 1500 -2778
rect 1494 -2790 1500 -2784
rect 1494 -2796 1500 -2790
rect 1494 -2802 1500 -2796
rect 1494 -2808 1500 -2802
rect 1494 -2814 1500 -2808
rect 1494 -2898 1500 -2892
rect 1494 -2904 1500 -2898
rect 1494 -2910 1500 -2904
rect 1494 -2916 1500 -2910
rect 1494 -2922 1500 -2916
rect 1494 -2928 1500 -2922
rect 1494 -2934 1500 -2928
rect 1494 -2940 1500 -2934
rect 1494 -2946 1500 -2940
rect 1494 -2952 1500 -2946
rect 1494 -2958 1500 -2952
rect 1494 -2964 1500 -2958
rect 1494 -2970 1500 -2964
rect 1494 -2976 1500 -2970
rect 1494 -2982 1500 -2976
rect 1494 -2988 1500 -2982
rect 1494 -2994 1500 -2988
rect 1494 -3000 1500 -2994
rect 1494 -3006 1500 -3000
rect 1494 -3012 1500 -3006
rect 1494 -3018 1500 -3012
rect 1494 -3024 1500 -3018
rect 1494 -3030 1500 -3024
rect 1494 -3036 1500 -3030
rect 1494 -3042 1500 -3036
rect 1494 -3048 1500 -3042
rect 1494 -3054 1500 -3048
rect 1494 -3060 1500 -3054
rect 1494 -3066 1500 -3060
rect 1494 -3072 1500 -3066
rect 1494 -3078 1500 -3072
rect 1494 -3084 1500 -3078
rect 1494 -3090 1500 -3084
rect 1494 -3096 1500 -3090
rect 1494 -3102 1500 -3096
rect 1494 -3108 1500 -3102
rect 1494 -3114 1500 -3108
rect 1494 -3120 1500 -3114
rect 1494 -3126 1500 -3120
rect 1494 -3132 1500 -3126
rect 1494 -3138 1500 -3132
rect 1494 -3144 1500 -3138
rect 1494 -3150 1500 -3144
rect 1494 -3156 1500 -3150
rect 1494 -3162 1500 -3156
rect 1494 -3168 1500 -3162
rect 1494 -3174 1500 -3168
rect 1494 -3180 1500 -3174
rect 1494 -3186 1500 -3180
rect 1494 -3192 1500 -3186
rect 1494 -3198 1500 -3192
rect 1494 -3204 1500 -3198
rect 1494 -3210 1500 -3204
rect 1494 -3216 1500 -3210
rect 1494 -3222 1500 -3216
rect 1494 -3228 1500 -3222
rect 1494 -3234 1500 -3228
rect 1494 -3282 1500 -3276
rect 1494 -3288 1500 -3282
rect 1494 -3294 1500 -3288
rect 1494 -3300 1500 -3294
rect 1494 -3306 1500 -3300
rect 1494 -3312 1500 -3306
rect 1494 -3318 1500 -3312
rect 1494 -3324 1500 -3318
rect 1494 -3330 1500 -3324
rect 1494 -3336 1500 -3330
rect 1494 -3342 1500 -3336
rect 1494 -3348 1500 -3342
rect 1494 -3354 1500 -3348
rect 1494 -3360 1500 -3354
rect 1494 -3366 1500 -3360
rect 1494 -3372 1500 -3366
rect 1494 -3378 1500 -3372
rect 1494 -3384 1500 -3378
rect 1494 -3390 1500 -3384
rect 1494 -3396 1500 -3390
rect 1494 -3402 1500 -3396
rect 1494 -3408 1500 -3402
rect 1494 -3414 1500 -3408
rect 1494 -3420 1500 -3414
rect 1494 -3426 1500 -3420
rect 1494 -3432 1500 -3426
rect 1494 -3438 1500 -3432
rect 1494 -3444 1500 -3438
rect 1494 -3450 1500 -3444
rect 1494 -3456 1500 -3450
rect 1494 -3462 1500 -3456
rect 1494 -3468 1500 -3462
rect 1494 -3474 1500 -3468
rect 1494 -3480 1500 -3474
rect 1494 -3486 1500 -3480
rect 1494 -3492 1500 -3486
rect 1500 -1182 1506 -1176
rect 1500 -1188 1506 -1182
rect 1500 -1194 1506 -1188
rect 1500 -1200 1506 -1194
rect 1500 -1206 1506 -1200
rect 1500 -1212 1506 -1206
rect 1500 -1218 1506 -1212
rect 1500 -1224 1506 -1218
rect 1500 -1230 1506 -1224
rect 1500 -1236 1506 -1230
rect 1500 -1242 1506 -1236
rect 1500 -1248 1506 -1242
rect 1500 -1254 1506 -1248
rect 1500 -1260 1506 -1254
rect 1500 -1266 1506 -1260
rect 1500 -1272 1506 -1266
rect 1500 -1278 1506 -1272
rect 1500 -1284 1506 -1278
rect 1500 -1290 1506 -1284
rect 1500 -1296 1506 -1290
rect 1500 -1302 1506 -1296
rect 1500 -1308 1506 -1302
rect 1500 -1314 1506 -1308
rect 1500 -1320 1506 -1314
rect 1500 -1326 1506 -1320
rect 1500 -1332 1506 -1326
rect 1500 -1338 1506 -1332
rect 1500 -1344 1506 -1338
rect 1500 -1350 1506 -1344
rect 1500 -1356 1506 -1350
rect 1500 -1362 1506 -1356
rect 1500 -1368 1506 -1362
rect 1500 -1374 1506 -1368
rect 1500 -1380 1506 -1374
rect 1500 -1386 1506 -1380
rect 1500 -1392 1506 -1386
rect 1500 -1398 1506 -1392
rect 1500 -1404 1506 -1398
rect 1500 -1410 1506 -1404
rect 1500 -1416 1506 -1410
rect 1500 -1422 1506 -1416
rect 1500 -1428 1506 -1422
rect 1500 -1434 1506 -1428
rect 1500 -1440 1506 -1434
rect 1500 -1446 1506 -1440
rect 1500 -1452 1506 -1446
rect 1500 -1458 1506 -1452
rect 1500 -1464 1506 -1458
rect 1500 -1470 1506 -1464
rect 1500 -1476 1506 -1470
rect 1500 -1482 1506 -1476
rect 1500 -1488 1506 -1482
rect 1500 -1494 1506 -1488
rect 1500 -1500 1506 -1494
rect 1500 -1506 1506 -1500
rect 1500 -1512 1506 -1506
rect 1500 -1518 1506 -1512
rect 1500 -1524 1506 -1518
rect 1500 -1530 1506 -1524
rect 1500 -1536 1506 -1530
rect 1500 -1542 1506 -1536
rect 1500 -1548 1506 -1542
rect 1500 -1554 1506 -1548
rect 1500 -1560 1506 -1554
rect 1500 -1566 1506 -1560
rect 1500 -1572 1506 -1566
rect 1500 -1578 1506 -1572
rect 1500 -1584 1506 -1578
rect 1500 -1590 1506 -1584
rect 1500 -1596 1506 -1590
rect 1500 -1602 1506 -1596
rect 1500 -1608 1506 -1602
rect 1500 -1614 1506 -1608
rect 1500 -1620 1506 -1614
rect 1500 -1626 1506 -1620
rect 1500 -1632 1506 -1626
rect 1500 -1638 1506 -1632
rect 1500 -1644 1506 -1638
rect 1500 -1650 1506 -1644
rect 1500 -1656 1506 -1650
rect 1500 -1662 1506 -1656
rect 1500 -1668 1506 -1662
rect 1500 -1674 1506 -1668
rect 1500 -1680 1506 -1674
rect 1500 -1686 1506 -1680
rect 1500 -1692 1506 -1686
rect 1500 -1698 1506 -1692
rect 1500 -1704 1506 -1698
rect 1500 -1710 1506 -1704
rect 1500 -1716 1506 -1710
rect 1500 -1722 1506 -1716
rect 1500 -1728 1506 -1722
rect 1500 -1734 1506 -1728
rect 1500 -1740 1506 -1734
rect 1500 -1746 1506 -1740
rect 1500 -1752 1506 -1746
rect 1500 -1758 1506 -1752
rect 1500 -1764 1506 -1758
rect 1500 -1770 1506 -1764
rect 1500 -1776 1506 -1770
rect 1500 -1782 1506 -1776
rect 1500 -1788 1506 -1782
rect 1500 -1794 1506 -1788
rect 1500 -1800 1506 -1794
rect 1500 -1806 1506 -1800
rect 1500 -1812 1506 -1806
rect 1500 -1818 1506 -1812
rect 1500 -1824 1506 -1818
rect 1500 -1830 1506 -1824
rect 1500 -1836 1506 -1830
rect 1500 -1842 1506 -1836
rect 1500 -1848 1506 -1842
rect 1500 -1854 1506 -1848
rect 1500 -1860 1506 -1854
rect 1500 -1866 1506 -1860
rect 1500 -1872 1506 -1866
rect 1500 -1878 1506 -1872
rect 1500 -1884 1506 -1878
rect 1500 -1890 1506 -1884
rect 1500 -1896 1506 -1890
rect 1500 -1902 1506 -1896
rect 1500 -1908 1506 -1902
rect 1500 -1914 1506 -1908
rect 1500 -1920 1506 -1914
rect 1500 -1926 1506 -1920
rect 1500 -1932 1506 -1926
rect 1500 -1938 1506 -1932
rect 1500 -1944 1506 -1938
rect 1500 -1950 1506 -1944
rect 1500 -1956 1506 -1950
rect 1500 -1962 1506 -1956
rect 1500 -1968 1506 -1962
rect 1500 -1974 1506 -1968
rect 1500 -1980 1506 -1974
rect 1500 -1986 1506 -1980
rect 1500 -1992 1506 -1986
rect 1500 -1998 1506 -1992
rect 1500 -2004 1506 -1998
rect 1500 -2010 1506 -2004
rect 1500 -2016 1506 -2010
rect 1500 -2022 1506 -2016
rect 1500 -2028 1506 -2022
rect 1500 -2034 1506 -2028
rect 1500 -2040 1506 -2034
rect 1500 -2046 1506 -2040
rect 1500 -2052 1506 -2046
rect 1500 -2058 1506 -2052
rect 1500 -2064 1506 -2058
rect 1500 -2070 1506 -2064
rect 1500 -2076 1506 -2070
rect 1500 -2082 1506 -2076
rect 1500 -2088 1506 -2082
rect 1500 -2094 1506 -2088
rect 1500 -2100 1506 -2094
rect 1500 -2106 1506 -2100
rect 1500 -2112 1506 -2106
rect 1500 -2118 1506 -2112
rect 1500 -2124 1506 -2118
rect 1500 -2130 1506 -2124
rect 1500 -2136 1506 -2130
rect 1500 -2142 1506 -2136
rect 1500 -2148 1506 -2142
rect 1500 -2154 1506 -2148
rect 1500 -2160 1506 -2154
rect 1500 -2166 1506 -2160
rect 1500 -2172 1506 -2166
rect 1500 -2178 1506 -2172
rect 1500 -2184 1506 -2178
rect 1500 -2190 1506 -2184
rect 1500 -2262 1506 -2256
rect 1500 -2268 1506 -2262
rect 1500 -2274 1506 -2268
rect 1500 -2280 1506 -2274
rect 1500 -2286 1506 -2280
rect 1500 -2292 1506 -2286
rect 1500 -2298 1506 -2292
rect 1500 -2304 1506 -2298
rect 1500 -2310 1506 -2304
rect 1500 -2316 1506 -2310
rect 1500 -2322 1506 -2316
rect 1500 -2328 1506 -2322
rect 1500 -2334 1506 -2328
rect 1500 -2340 1506 -2334
rect 1500 -2346 1506 -2340
rect 1500 -2352 1506 -2346
rect 1500 -2358 1506 -2352
rect 1500 -2364 1506 -2358
rect 1500 -2370 1506 -2364
rect 1500 -2376 1506 -2370
rect 1500 -2382 1506 -2376
rect 1500 -2388 1506 -2382
rect 1500 -2394 1506 -2388
rect 1500 -2400 1506 -2394
rect 1500 -2406 1506 -2400
rect 1500 -2412 1506 -2406
rect 1500 -2418 1506 -2412
rect 1500 -2424 1506 -2418
rect 1500 -2430 1506 -2424
rect 1500 -2436 1506 -2430
rect 1500 -2442 1506 -2436
rect 1500 -2448 1506 -2442
rect 1500 -2454 1506 -2448
rect 1500 -2460 1506 -2454
rect 1500 -2466 1506 -2460
rect 1500 -2472 1506 -2466
rect 1500 -2478 1506 -2472
rect 1500 -2484 1506 -2478
rect 1500 -2490 1506 -2484
rect 1500 -2496 1506 -2490
rect 1500 -2502 1506 -2496
rect 1500 -2508 1506 -2502
rect 1500 -2514 1506 -2508
rect 1500 -2520 1506 -2514
rect 1500 -2526 1506 -2520
rect 1500 -2532 1506 -2526
rect 1500 -2538 1506 -2532
rect 1500 -2544 1506 -2538
rect 1500 -2550 1506 -2544
rect 1500 -2556 1506 -2550
rect 1500 -2562 1506 -2556
rect 1500 -2568 1506 -2562
rect 1500 -2574 1506 -2568
rect 1500 -2580 1506 -2574
rect 1500 -2586 1506 -2580
rect 1500 -2592 1506 -2586
rect 1500 -2598 1506 -2592
rect 1500 -2604 1506 -2598
rect 1500 -2610 1506 -2604
rect 1500 -2616 1506 -2610
rect 1500 -2622 1506 -2616
rect 1500 -2628 1506 -2622
rect 1500 -2634 1506 -2628
rect 1500 -2640 1506 -2634
rect 1500 -2646 1506 -2640
rect 1500 -2652 1506 -2646
rect 1500 -2658 1506 -2652
rect 1500 -2664 1506 -2658
rect 1500 -2670 1506 -2664
rect 1500 -2676 1506 -2670
rect 1500 -2682 1506 -2676
rect 1500 -2688 1506 -2682
rect 1500 -2694 1506 -2688
rect 1500 -2700 1506 -2694
rect 1500 -2706 1506 -2700
rect 1500 -2712 1506 -2706
rect 1500 -2718 1506 -2712
rect 1500 -2724 1506 -2718
rect 1500 -2730 1506 -2724
rect 1500 -2736 1506 -2730
rect 1500 -2742 1506 -2736
rect 1500 -2748 1506 -2742
rect 1500 -2754 1506 -2748
rect 1500 -2760 1506 -2754
rect 1500 -2766 1506 -2760
rect 1500 -2772 1506 -2766
rect 1500 -2778 1506 -2772
rect 1500 -2784 1506 -2778
rect 1500 -2790 1506 -2784
rect 1500 -2796 1506 -2790
rect 1500 -2802 1506 -2796
rect 1500 -2808 1506 -2802
rect 1500 -2892 1506 -2886
rect 1500 -2898 1506 -2892
rect 1500 -2904 1506 -2898
rect 1500 -2910 1506 -2904
rect 1500 -2916 1506 -2910
rect 1500 -2922 1506 -2916
rect 1500 -2928 1506 -2922
rect 1500 -2934 1506 -2928
rect 1500 -2940 1506 -2934
rect 1500 -2946 1506 -2940
rect 1500 -2952 1506 -2946
rect 1500 -2958 1506 -2952
rect 1500 -2964 1506 -2958
rect 1500 -2970 1506 -2964
rect 1500 -2976 1506 -2970
rect 1500 -2982 1506 -2976
rect 1500 -2988 1506 -2982
rect 1500 -2994 1506 -2988
rect 1500 -3000 1506 -2994
rect 1500 -3006 1506 -3000
rect 1500 -3012 1506 -3006
rect 1500 -3018 1506 -3012
rect 1500 -3024 1506 -3018
rect 1500 -3030 1506 -3024
rect 1500 -3036 1506 -3030
rect 1500 -3042 1506 -3036
rect 1500 -3048 1506 -3042
rect 1500 -3054 1506 -3048
rect 1500 -3060 1506 -3054
rect 1500 -3066 1506 -3060
rect 1500 -3072 1506 -3066
rect 1500 -3078 1506 -3072
rect 1500 -3084 1506 -3078
rect 1500 -3090 1506 -3084
rect 1500 -3096 1506 -3090
rect 1500 -3102 1506 -3096
rect 1500 -3108 1506 -3102
rect 1500 -3114 1506 -3108
rect 1500 -3120 1506 -3114
rect 1500 -3126 1506 -3120
rect 1500 -3132 1506 -3126
rect 1500 -3138 1506 -3132
rect 1500 -3144 1506 -3138
rect 1500 -3150 1506 -3144
rect 1500 -3156 1506 -3150
rect 1500 -3162 1506 -3156
rect 1500 -3168 1506 -3162
rect 1500 -3174 1506 -3168
rect 1500 -3180 1506 -3174
rect 1500 -3186 1506 -3180
rect 1500 -3192 1506 -3186
rect 1500 -3198 1506 -3192
rect 1500 -3204 1506 -3198
rect 1500 -3210 1506 -3204
rect 1500 -3216 1506 -3210
rect 1500 -3222 1506 -3216
rect 1500 -3228 1506 -3222
rect 1500 -3234 1506 -3228
rect 1500 -3282 1506 -3276
rect 1500 -3288 1506 -3282
rect 1500 -3294 1506 -3288
rect 1500 -3300 1506 -3294
rect 1500 -3306 1506 -3300
rect 1500 -3312 1506 -3306
rect 1500 -3318 1506 -3312
rect 1500 -3324 1506 -3318
rect 1500 -3330 1506 -3324
rect 1500 -3336 1506 -3330
rect 1500 -3342 1506 -3336
rect 1500 -3348 1506 -3342
rect 1500 -3354 1506 -3348
rect 1500 -3360 1506 -3354
rect 1500 -3366 1506 -3360
rect 1500 -3372 1506 -3366
rect 1500 -3378 1506 -3372
rect 1500 -3384 1506 -3378
rect 1500 -3390 1506 -3384
rect 1500 -3396 1506 -3390
rect 1500 -3402 1506 -3396
rect 1500 -3408 1506 -3402
rect 1500 -3414 1506 -3408
rect 1500 -3420 1506 -3414
rect 1500 -3426 1506 -3420
rect 1500 -3432 1506 -3426
rect 1500 -3438 1506 -3432
rect 1500 -3444 1506 -3438
rect 1500 -3450 1506 -3444
rect 1500 -3456 1506 -3450
rect 1500 -3462 1506 -3456
rect 1500 -3468 1506 -3462
rect 1500 -3474 1506 -3468
rect 1500 -3480 1506 -3474
rect 1500 -3486 1506 -3480
rect 1506 -1170 1512 -1164
rect 1506 -1176 1512 -1170
rect 1506 -1182 1512 -1176
rect 1506 -1188 1512 -1182
rect 1506 -1194 1512 -1188
rect 1506 -1200 1512 -1194
rect 1506 -1206 1512 -1200
rect 1506 -1212 1512 -1206
rect 1506 -1218 1512 -1212
rect 1506 -1224 1512 -1218
rect 1506 -1230 1512 -1224
rect 1506 -1236 1512 -1230
rect 1506 -1242 1512 -1236
rect 1506 -1248 1512 -1242
rect 1506 -1254 1512 -1248
rect 1506 -1260 1512 -1254
rect 1506 -1266 1512 -1260
rect 1506 -1272 1512 -1266
rect 1506 -1278 1512 -1272
rect 1506 -1284 1512 -1278
rect 1506 -1290 1512 -1284
rect 1506 -1296 1512 -1290
rect 1506 -1302 1512 -1296
rect 1506 -1308 1512 -1302
rect 1506 -1314 1512 -1308
rect 1506 -1320 1512 -1314
rect 1506 -1326 1512 -1320
rect 1506 -1332 1512 -1326
rect 1506 -1338 1512 -1332
rect 1506 -1344 1512 -1338
rect 1506 -1350 1512 -1344
rect 1506 -1356 1512 -1350
rect 1506 -1362 1512 -1356
rect 1506 -1368 1512 -1362
rect 1506 -1374 1512 -1368
rect 1506 -1380 1512 -1374
rect 1506 -1386 1512 -1380
rect 1506 -1392 1512 -1386
rect 1506 -1398 1512 -1392
rect 1506 -1404 1512 -1398
rect 1506 -1410 1512 -1404
rect 1506 -1416 1512 -1410
rect 1506 -1422 1512 -1416
rect 1506 -1428 1512 -1422
rect 1506 -1434 1512 -1428
rect 1506 -1440 1512 -1434
rect 1506 -1446 1512 -1440
rect 1506 -1452 1512 -1446
rect 1506 -1458 1512 -1452
rect 1506 -1464 1512 -1458
rect 1506 -1470 1512 -1464
rect 1506 -1476 1512 -1470
rect 1506 -1482 1512 -1476
rect 1506 -1488 1512 -1482
rect 1506 -1494 1512 -1488
rect 1506 -1500 1512 -1494
rect 1506 -1506 1512 -1500
rect 1506 -1512 1512 -1506
rect 1506 -1518 1512 -1512
rect 1506 -1524 1512 -1518
rect 1506 -1530 1512 -1524
rect 1506 -1536 1512 -1530
rect 1506 -1542 1512 -1536
rect 1506 -1548 1512 -1542
rect 1506 -1554 1512 -1548
rect 1506 -1560 1512 -1554
rect 1506 -1566 1512 -1560
rect 1506 -1572 1512 -1566
rect 1506 -1578 1512 -1572
rect 1506 -1584 1512 -1578
rect 1506 -1590 1512 -1584
rect 1506 -1596 1512 -1590
rect 1506 -1602 1512 -1596
rect 1506 -1608 1512 -1602
rect 1506 -1614 1512 -1608
rect 1506 -1620 1512 -1614
rect 1506 -1626 1512 -1620
rect 1506 -1632 1512 -1626
rect 1506 -1638 1512 -1632
rect 1506 -1644 1512 -1638
rect 1506 -1650 1512 -1644
rect 1506 -1656 1512 -1650
rect 1506 -1662 1512 -1656
rect 1506 -1668 1512 -1662
rect 1506 -1674 1512 -1668
rect 1506 -1680 1512 -1674
rect 1506 -1686 1512 -1680
rect 1506 -1692 1512 -1686
rect 1506 -1698 1512 -1692
rect 1506 -1704 1512 -1698
rect 1506 -1710 1512 -1704
rect 1506 -1716 1512 -1710
rect 1506 -1722 1512 -1716
rect 1506 -1728 1512 -1722
rect 1506 -1734 1512 -1728
rect 1506 -1740 1512 -1734
rect 1506 -1746 1512 -1740
rect 1506 -1752 1512 -1746
rect 1506 -1758 1512 -1752
rect 1506 -1764 1512 -1758
rect 1506 -1770 1512 -1764
rect 1506 -1776 1512 -1770
rect 1506 -1782 1512 -1776
rect 1506 -1788 1512 -1782
rect 1506 -1794 1512 -1788
rect 1506 -1800 1512 -1794
rect 1506 -1806 1512 -1800
rect 1506 -1812 1512 -1806
rect 1506 -1818 1512 -1812
rect 1506 -1824 1512 -1818
rect 1506 -1830 1512 -1824
rect 1506 -1836 1512 -1830
rect 1506 -1842 1512 -1836
rect 1506 -1848 1512 -1842
rect 1506 -1854 1512 -1848
rect 1506 -1860 1512 -1854
rect 1506 -1866 1512 -1860
rect 1506 -1872 1512 -1866
rect 1506 -1878 1512 -1872
rect 1506 -1884 1512 -1878
rect 1506 -1890 1512 -1884
rect 1506 -1896 1512 -1890
rect 1506 -1902 1512 -1896
rect 1506 -1908 1512 -1902
rect 1506 -1914 1512 -1908
rect 1506 -1920 1512 -1914
rect 1506 -1926 1512 -1920
rect 1506 -1932 1512 -1926
rect 1506 -1938 1512 -1932
rect 1506 -1944 1512 -1938
rect 1506 -1950 1512 -1944
rect 1506 -1956 1512 -1950
rect 1506 -1962 1512 -1956
rect 1506 -1968 1512 -1962
rect 1506 -1974 1512 -1968
rect 1506 -1980 1512 -1974
rect 1506 -1986 1512 -1980
rect 1506 -1992 1512 -1986
rect 1506 -1998 1512 -1992
rect 1506 -2004 1512 -1998
rect 1506 -2010 1512 -2004
rect 1506 -2016 1512 -2010
rect 1506 -2022 1512 -2016
rect 1506 -2028 1512 -2022
rect 1506 -2034 1512 -2028
rect 1506 -2040 1512 -2034
rect 1506 -2046 1512 -2040
rect 1506 -2052 1512 -2046
rect 1506 -2058 1512 -2052
rect 1506 -2064 1512 -2058
rect 1506 -2070 1512 -2064
rect 1506 -2076 1512 -2070
rect 1506 -2082 1512 -2076
rect 1506 -2088 1512 -2082
rect 1506 -2094 1512 -2088
rect 1506 -2100 1512 -2094
rect 1506 -2106 1512 -2100
rect 1506 -2112 1512 -2106
rect 1506 -2118 1512 -2112
rect 1506 -2124 1512 -2118
rect 1506 -2130 1512 -2124
rect 1506 -2136 1512 -2130
rect 1506 -2142 1512 -2136
rect 1506 -2148 1512 -2142
rect 1506 -2154 1512 -2148
rect 1506 -2160 1512 -2154
rect 1506 -2166 1512 -2160
rect 1506 -2172 1512 -2166
rect 1506 -2178 1512 -2172
rect 1506 -2184 1512 -2178
rect 1506 -2256 1512 -2250
rect 1506 -2262 1512 -2256
rect 1506 -2268 1512 -2262
rect 1506 -2274 1512 -2268
rect 1506 -2280 1512 -2274
rect 1506 -2286 1512 -2280
rect 1506 -2292 1512 -2286
rect 1506 -2298 1512 -2292
rect 1506 -2304 1512 -2298
rect 1506 -2310 1512 -2304
rect 1506 -2316 1512 -2310
rect 1506 -2322 1512 -2316
rect 1506 -2328 1512 -2322
rect 1506 -2334 1512 -2328
rect 1506 -2340 1512 -2334
rect 1506 -2346 1512 -2340
rect 1506 -2352 1512 -2346
rect 1506 -2358 1512 -2352
rect 1506 -2364 1512 -2358
rect 1506 -2370 1512 -2364
rect 1506 -2376 1512 -2370
rect 1506 -2382 1512 -2376
rect 1506 -2388 1512 -2382
rect 1506 -2394 1512 -2388
rect 1506 -2400 1512 -2394
rect 1506 -2406 1512 -2400
rect 1506 -2412 1512 -2406
rect 1506 -2418 1512 -2412
rect 1506 -2424 1512 -2418
rect 1506 -2430 1512 -2424
rect 1506 -2436 1512 -2430
rect 1506 -2442 1512 -2436
rect 1506 -2448 1512 -2442
rect 1506 -2454 1512 -2448
rect 1506 -2460 1512 -2454
rect 1506 -2466 1512 -2460
rect 1506 -2472 1512 -2466
rect 1506 -2478 1512 -2472
rect 1506 -2484 1512 -2478
rect 1506 -2490 1512 -2484
rect 1506 -2496 1512 -2490
rect 1506 -2502 1512 -2496
rect 1506 -2508 1512 -2502
rect 1506 -2514 1512 -2508
rect 1506 -2520 1512 -2514
rect 1506 -2526 1512 -2520
rect 1506 -2532 1512 -2526
rect 1506 -2538 1512 -2532
rect 1506 -2544 1512 -2538
rect 1506 -2550 1512 -2544
rect 1506 -2556 1512 -2550
rect 1506 -2562 1512 -2556
rect 1506 -2568 1512 -2562
rect 1506 -2574 1512 -2568
rect 1506 -2580 1512 -2574
rect 1506 -2586 1512 -2580
rect 1506 -2592 1512 -2586
rect 1506 -2598 1512 -2592
rect 1506 -2604 1512 -2598
rect 1506 -2610 1512 -2604
rect 1506 -2616 1512 -2610
rect 1506 -2622 1512 -2616
rect 1506 -2628 1512 -2622
rect 1506 -2634 1512 -2628
rect 1506 -2640 1512 -2634
rect 1506 -2646 1512 -2640
rect 1506 -2652 1512 -2646
rect 1506 -2658 1512 -2652
rect 1506 -2664 1512 -2658
rect 1506 -2670 1512 -2664
rect 1506 -2676 1512 -2670
rect 1506 -2682 1512 -2676
rect 1506 -2688 1512 -2682
rect 1506 -2694 1512 -2688
rect 1506 -2700 1512 -2694
rect 1506 -2706 1512 -2700
rect 1506 -2712 1512 -2706
rect 1506 -2718 1512 -2712
rect 1506 -2724 1512 -2718
rect 1506 -2730 1512 -2724
rect 1506 -2736 1512 -2730
rect 1506 -2742 1512 -2736
rect 1506 -2748 1512 -2742
rect 1506 -2754 1512 -2748
rect 1506 -2760 1512 -2754
rect 1506 -2766 1512 -2760
rect 1506 -2772 1512 -2766
rect 1506 -2778 1512 -2772
rect 1506 -2784 1512 -2778
rect 1506 -2790 1512 -2784
rect 1506 -2796 1512 -2790
rect 1506 -2802 1512 -2796
rect 1506 -2808 1512 -2802
rect 1506 -2892 1512 -2886
rect 1506 -2898 1512 -2892
rect 1506 -2904 1512 -2898
rect 1506 -2910 1512 -2904
rect 1506 -2916 1512 -2910
rect 1506 -2922 1512 -2916
rect 1506 -2928 1512 -2922
rect 1506 -2934 1512 -2928
rect 1506 -2940 1512 -2934
rect 1506 -2946 1512 -2940
rect 1506 -2952 1512 -2946
rect 1506 -2958 1512 -2952
rect 1506 -2964 1512 -2958
rect 1506 -2970 1512 -2964
rect 1506 -2976 1512 -2970
rect 1506 -2982 1512 -2976
rect 1506 -2988 1512 -2982
rect 1506 -2994 1512 -2988
rect 1506 -3000 1512 -2994
rect 1506 -3006 1512 -3000
rect 1506 -3012 1512 -3006
rect 1506 -3018 1512 -3012
rect 1506 -3024 1512 -3018
rect 1506 -3030 1512 -3024
rect 1506 -3036 1512 -3030
rect 1506 -3042 1512 -3036
rect 1506 -3048 1512 -3042
rect 1506 -3054 1512 -3048
rect 1506 -3060 1512 -3054
rect 1506 -3066 1512 -3060
rect 1506 -3072 1512 -3066
rect 1506 -3078 1512 -3072
rect 1506 -3084 1512 -3078
rect 1506 -3090 1512 -3084
rect 1506 -3096 1512 -3090
rect 1506 -3102 1512 -3096
rect 1506 -3108 1512 -3102
rect 1506 -3114 1512 -3108
rect 1506 -3120 1512 -3114
rect 1506 -3126 1512 -3120
rect 1506 -3132 1512 -3126
rect 1506 -3138 1512 -3132
rect 1506 -3144 1512 -3138
rect 1506 -3150 1512 -3144
rect 1506 -3156 1512 -3150
rect 1506 -3162 1512 -3156
rect 1506 -3168 1512 -3162
rect 1506 -3174 1512 -3168
rect 1506 -3180 1512 -3174
rect 1506 -3186 1512 -3180
rect 1506 -3192 1512 -3186
rect 1506 -3198 1512 -3192
rect 1506 -3204 1512 -3198
rect 1506 -3210 1512 -3204
rect 1506 -3216 1512 -3210
rect 1506 -3222 1512 -3216
rect 1506 -3228 1512 -3222
rect 1506 -3234 1512 -3228
rect 1506 -3276 1512 -3270
rect 1506 -3282 1512 -3276
rect 1506 -3288 1512 -3282
rect 1506 -3294 1512 -3288
rect 1506 -3300 1512 -3294
rect 1506 -3306 1512 -3300
rect 1506 -3312 1512 -3306
rect 1506 -3318 1512 -3312
rect 1506 -3324 1512 -3318
rect 1506 -3330 1512 -3324
rect 1506 -3336 1512 -3330
rect 1506 -3342 1512 -3336
rect 1506 -3348 1512 -3342
rect 1506 -3354 1512 -3348
rect 1506 -3360 1512 -3354
rect 1506 -3366 1512 -3360
rect 1506 -3372 1512 -3366
rect 1506 -3378 1512 -3372
rect 1506 -3384 1512 -3378
rect 1506 -3390 1512 -3384
rect 1506 -3396 1512 -3390
rect 1506 -3402 1512 -3396
rect 1506 -3408 1512 -3402
rect 1506 -3414 1512 -3408
rect 1506 -3420 1512 -3414
rect 1506 -3426 1512 -3420
rect 1506 -3432 1512 -3426
rect 1506 -3438 1512 -3432
rect 1506 -3444 1512 -3438
rect 1506 -3450 1512 -3444
rect 1506 -3456 1512 -3450
rect 1506 -3462 1512 -3456
rect 1506 -3468 1512 -3462
rect 1506 -3474 1512 -3468
rect 1506 -3480 1512 -3474
rect 1506 -3486 1512 -3480
rect 1512 -1158 1518 -1152
rect 1512 -1164 1518 -1158
rect 1512 -1170 1518 -1164
rect 1512 -1176 1518 -1170
rect 1512 -1182 1518 -1176
rect 1512 -1188 1518 -1182
rect 1512 -1194 1518 -1188
rect 1512 -1200 1518 -1194
rect 1512 -1206 1518 -1200
rect 1512 -1212 1518 -1206
rect 1512 -1218 1518 -1212
rect 1512 -1224 1518 -1218
rect 1512 -1230 1518 -1224
rect 1512 -1236 1518 -1230
rect 1512 -1242 1518 -1236
rect 1512 -1248 1518 -1242
rect 1512 -1254 1518 -1248
rect 1512 -1260 1518 -1254
rect 1512 -1266 1518 -1260
rect 1512 -1272 1518 -1266
rect 1512 -1278 1518 -1272
rect 1512 -1284 1518 -1278
rect 1512 -1290 1518 -1284
rect 1512 -1296 1518 -1290
rect 1512 -1302 1518 -1296
rect 1512 -1308 1518 -1302
rect 1512 -1314 1518 -1308
rect 1512 -1320 1518 -1314
rect 1512 -1326 1518 -1320
rect 1512 -1332 1518 -1326
rect 1512 -1338 1518 -1332
rect 1512 -1344 1518 -1338
rect 1512 -1350 1518 -1344
rect 1512 -1356 1518 -1350
rect 1512 -1362 1518 -1356
rect 1512 -1368 1518 -1362
rect 1512 -1374 1518 -1368
rect 1512 -1380 1518 -1374
rect 1512 -1386 1518 -1380
rect 1512 -1392 1518 -1386
rect 1512 -1398 1518 -1392
rect 1512 -1404 1518 -1398
rect 1512 -1410 1518 -1404
rect 1512 -1416 1518 -1410
rect 1512 -1422 1518 -1416
rect 1512 -1428 1518 -1422
rect 1512 -1434 1518 -1428
rect 1512 -1440 1518 -1434
rect 1512 -1446 1518 -1440
rect 1512 -1452 1518 -1446
rect 1512 -1458 1518 -1452
rect 1512 -1464 1518 -1458
rect 1512 -1470 1518 -1464
rect 1512 -1476 1518 -1470
rect 1512 -1482 1518 -1476
rect 1512 -1488 1518 -1482
rect 1512 -1494 1518 -1488
rect 1512 -1500 1518 -1494
rect 1512 -1506 1518 -1500
rect 1512 -1512 1518 -1506
rect 1512 -1518 1518 -1512
rect 1512 -1524 1518 -1518
rect 1512 -1530 1518 -1524
rect 1512 -1536 1518 -1530
rect 1512 -1542 1518 -1536
rect 1512 -1548 1518 -1542
rect 1512 -1554 1518 -1548
rect 1512 -1560 1518 -1554
rect 1512 -1566 1518 -1560
rect 1512 -1572 1518 -1566
rect 1512 -1578 1518 -1572
rect 1512 -1584 1518 -1578
rect 1512 -1590 1518 -1584
rect 1512 -1596 1518 -1590
rect 1512 -1602 1518 -1596
rect 1512 -1608 1518 -1602
rect 1512 -1614 1518 -1608
rect 1512 -1620 1518 -1614
rect 1512 -1626 1518 -1620
rect 1512 -1632 1518 -1626
rect 1512 -1638 1518 -1632
rect 1512 -1644 1518 -1638
rect 1512 -1650 1518 -1644
rect 1512 -1656 1518 -1650
rect 1512 -1662 1518 -1656
rect 1512 -1668 1518 -1662
rect 1512 -1674 1518 -1668
rect 1512 -1680 1518 -1674
rect 1512 -1686 1518 -1680
rect 1512 -1692 1518 -1686
rect 1512 -1698 1518 -1692
rect 1512 -1704 1518 -1698
rect 1512 -1710 1518 -1704
rect 1512 -1716 1518 -1710
rect 1512 -1722 1518 -1716
rect 1512 -1728 1518 -1722
rect 1512 -1734 1518 -1728
rect 1512 -1740 1518 -1734
rect 1512 -1746 1518 -1740
rect 1512 -1752 1518 -1746
rect 1512 -1758 1518 -1752
rect 1512 -1764 1518 -1758
rect 1512 -1770 1518 -1764
rect 1512 -1776 1518 -1770
rect 1512 -1782 1518 -1776
rect 1512 -1788 1518 -1782
rect 1512 -1794 1518 -1788
rect 1512 -1800 1518 -1794
rect 1512 -1806 1518 -1800
rect 1512 -1812 1518 -1806
rect 1512 -1818 1518 -1812
rect 1512 -1824 1518 -1818
rect 1512 -1830 1518 -1824
rect 1512 -1836 1518 -1830
rect 1512 -1842 1518 -1836
rect 1512 -1848 1518 -1842
rect 1512 -1854 1518 -1848
rect 1512 -1860 1518 -1854
rect 1512 -1866 1518 -1860
rect 1512 -1872 1518 -1866
rect 1512 -1878 1518 -1872
rect 1512 -1884 1518 -1878
rect 1512 -1890 1518 -1884
rect 1512 -1896 1518 -1890
rect 1512 -1902 1518 -1896
rect 1512 -1908 1518 -1902
rect 1512 -1914 1518 -1908
rect 1512 -1920 1518 -1914
rect 1512 -1926 1518 -1920
rect 1512 -1932 1518 -1926
rect 1512 -1938 1518 -1932
rect 1512 -1944 1518 -1938
rect 1512 -1950 1518 -1944
rect 1512 -1956 1518 -1950
rect 1512 -1962 1518 -1956
rect 1512 -1968 1518 -1962
rect 1512 -1974 1518 -1968
rect 1512 -1980 1518 -1974
rect 1512 -1986 1518 -1980
rect 1512 -1992 1518 -1986
rect 1512 -1998 1518 -1992
rect 1512 -2004 1518 -1998
rect 1512 -2010 1518 -2004
rect 1512 -2016 1518 -2010
rect 1512 -2022 1518 -2016
rect 1512 -2028 1518 -2022
rect 1512 -2034 1518 -2028
rect 1512 -2040 1518 -2034
rect 1512 -2046 1518 -2040
rect 1512 -2052 1518 -2046
rect 1512 -2058 1518 -2052
rect 1512 -2064 1518 -2058
rect 1512 -2070 1518 -2064
rect 1512 -2076 1518 -2070
rect 1512 -2082 1518 -2076
rect 1512 -2088 1518 -2082
rect 1512 -2094 1518 -2088
rect 1512 -2100 1518 -2094
rect 1512 -2106 1518 -2100
rect 1512 -2112 1518 -2106
rect 1512 -2118 1518 -2112
rect 1512 -2124 1518 -2118
rect 1512 -2130 1518 -2124
rect 1512 -2136 1518 -2130
rect 1512 -2142 1518 -2136
rect 1512 -2148 1518 -2142
rect 1512 -2154 1518 -2148
rect 1512 -2160 1518 -2154
rect 1512 -2166 1518 -2160
rect 1512 -2172 1518 -2166
rect 1512 -2250 1518 -2244
rect 1512 -2256 1518 -2250
rect 1512 -2262 1518 -2256
rect 1512 -2268 1518 -2262
rect 1512 -2274 1518 -2268
rect 1512 -2280 1518 -2274
rect 1512 -2286 1518 -2280
rect 1512 -2292 1518 -2286
rect 1512 -2298 1518 -2292
rect 1512 -2304 1518 -2298
rect 1512 -2310 1518 -2304
rect 1512 -2316 1518 -2310
rect 1512 -2322 1518 -2316
rect 1512 -2328 1518 -2322
rect 1512 -2334 1518 -2328
rect 1512 -2340 1518 -2334
rect 1512 -2346 1518 -2340
rect 1512 -2352 1518 -2346
rect 1512 -2358 1518 -2352
rect 1512 -2364 1518 -2358
rect 1512 -2370 1518 -2364
rect 1512 -2376 1518 -2370
rect 1512 -2382 1518 -2376
rect 1512 -2388 1518 -2382
rect 1512 -2394 1518 -2388
rect 1512 -2400 1518 -2394
rect 1512 -2406 1518 -2400
rect 1512 -2412 1518 -2406
rect 1512 -2418 1518 -2412
rect 1512 -2424 1518 -2418
rect 1512 -2430 1518 -2424
rect 1512 -2436 1518 -2430
rect 1512 -2442 1518 -2436
rect 1512 -2448 1518 -2442
rect 1512 -2454 1518 -2448
rect 1512 -2460 1518 -2454
rect 1512 -2466 1518 -2460
rect 1512 -2472 1518 -2466
rect 1512 -2478 1518 -2472
rect 1512 -2484 1518 -2478
rect 1512 -2490 1518 -2484
rect 1512 -2496 1518 -2490
rect 1512 -2502 1518 -2496
rect 1512 -2508 1518 -2502
rect 1512 -2514 1518 -2508
rect 1512 -2520 1518 -2514
rect 1512 -2526 1518 -2520
rect 1512 -2532 1518 -2526
rect 1512 -2538 1518 -2532
rect 1512 -2544 1518 -2538
rect 1512 -2550 1518 -2544
rect 1512 -2556 1518 -2550
rect 1512 -2562 1518 -2556
rect 1512 -2568 1518 -2562
rect 1512 -2574 1518 -2568
rect 1512 -2580 1518 -2574
rect 1512 -2586 1518 -2580
rect 1512 -2592 1518 -2586
rect 1512 -2598 1518 -2592
rect 1512 -2604 1518 -2598
rect 1512 -2610 1518 -2604
rect 1512 -2616 1518 -2610
rect 1512 -2622 1518 -2616
rect 1512 -2628 1518 -2622
rect 1512 -2634 1518 -2628
rect 1512 -2640 1518 -2634
rect 1512 -2646 1518 -2640
rect 1512 -2652 1518 -2646
rect 1512 -2658 1518 -2652
rect 1512 -2664 1518 -2658
rect 1512 -2670 1518 -2664
rect 1512 -2676 1518 -2670
rect 1512 -2682 1518 -2676
rect 1512 -2688 1518 -2682
rect 1512 -2694 1518 -2688
rect 1512 -2700 1518 -2694
rect 1512 -2706 1518 -2700
rect 1512 -2712 1518 -2706
rect 1512 -2718 1518 -2712
rect 1512 -2724 1518 -2718
rect 1512 -2730 1518 -2724
rect 1512 -2736 1518 -2730
rect 1512 -2742 1518 -2736
rect 1512 -2748 1518 -2742
rect 1512 -2754 1518 -2748
rect 1512 -2760 1518 -2754
rect 1512 -2766 1518 -2760
rect 1512 -2772 1518 -2766
rect 1512 -2778 1518 -2772
rect 1512 -2784 1518 -2778
rect 1512 -2790 1518 -2784
rect 1512 -2796 1518 -2790
rect 1512 -2802 1518 -2796
rect 1512 -2886 1518 -2880
rect 1512 -2892 1518 -2886
rect 1512 -2898 1518 -2892
rect 1512 -2904 1518 -2898
rect 1512 -2910 1518 -2904
rect 1512 -2916 1518 -2910
rect 1512 -2922 1518 -2916
rect 1512 -2928 1518 -2922
rect 1512 -2934 1518 -2928
rect 1512 -2940 1518 -2934
rect 1512 -2946 1518 -2940
rect 1512 -2952 1518 -2946
rect 1512 -2958 1518 -2952
rect 1512 -2964 1518 -2958
rect 1512 -2970 1518 -2964
rect 1512 -2976 1518 -2970
rect 1512 -2982 1518 -2976
rect 1512 -2988 1518 -2982
rect 1512 -2994 1518 -2988
rect 1512 -3000 1518 -2994
rect 1512 -3006 1518 -3000
rect 1512 -3012 1518 -3006
rect 1512 -3018 1518 -3012
rect 1512 -3024 1518 -3018
rect 1512 -3030 1518 -3024
rect 1512 -3036 1518 -3030
rect 1512 -3042 1518 -3036
rect 1512 -3048 1518 -3042
rect 1512 -3054 1518 -3048
rect 1512 -3060 1518 -3054
rect 1512 -3066 1518 -3060
rect 1512 -3072 1518 -3066
rect 1512 -3078 1518 -3072
rect 1512 -3084 1518 -3078
rect 1512 -3090 1518 -3084
rect 1512 -3096 1518 -3090
rect 1512 -3102 1518 -3096
rect 1512 -3108 1518 -3102
rect 1512 -3114 1518 -3108
rect 1512 -3120 1518 -3114
rect 1512 -3126 1518 -3120
rect 1512 -3132 1518 -3126
rect 1512 -3138 1518 -3132
rect 1512 -3144 1518 -3138
rect 1512 -3150 1518 -3144
rect 1512 -3156 1518 -3150
rect 1512 -3162 1518 -3156
rect 1512 -3168 1518 -3162
rect 1512 -3174 1518 -3168
rect 1512 -3180 1518 -3174
rect 1512 -3186 1518 -3180
rect 1512 -3192 1518 -3186
rect 1512 -3198 1518 -3192
rect 1512 -3204 1518 -3198
rect 1512 -3210 1518 -3204
rect 1512 -3216 1518 -3210
rect 1512 -3222 1518 -3216
rect 1512 -3228 1518 -3222
rect 1512 -3234 1518 -3228
rect 1512 -3276 1518 -3270
rect 1512 -3282 1518 -3276
rect 1512 -3288 1518 -3282
rect 1512 -3294 1518 -3288
rect 1512 -3300 1518 -3294
rect 1512 -3306 1518 -3300
rect 1512 -3312 1518 -3306
rect 1512 -3318 1518 -3312
rect 1512 -3324 1518 -3318
rect 1512 -3330 1518 -3324
rect 1512 -3336 1518 -3330
rect 1512 -3342 1518 -3336
rect 1512 -3348 1518 -3342
rect 1512 -3354 1518 -3348
rect 1512 -3360 1518 -3354
rect 1512 -3366 1518 -3360
rect 1512 -3372 1518 -3366
rect 1512 -3378 1518 -3372
rect 1512 -3384 1518 -3378
rect 1512 -3390 1518 -3384
rect 1512 -3396 1518 -3390
rect 1512 -3402 1518 -3396
rect 1512 -3408 1518 -3402
rect 1512 -3414 1518 -3408
rect 1512 -3420 1518 -3414
rect 1512 -3426 1518 -3420
rect 1512 -3432 1518 -3426
rect 1512 -3438 1518 -3432
rect 1512 -3444 1518 -3438
rect 1512 -3450 1518 -3444
rect 1512 -3456 1518 -3450
rect 1512 -3462 1518 -3456
rect 1512 -3468 1518 -3462
rect 1512 -3474 1518 -3468
rect 1512 -3480 1518 -3474
rect 1512 -3486 1518 -3480
rect 1518 -1152 1524 -1146
rect 1518 -1158 1524 -1152
rect 1518 -1164 1524 -1158
rect 1518 -1170 1524 -1164
rect 1518 -1176 1524 -1170
rect 1518 -1182 1524 -1176
rect 1518 -1188 1524 -1182
rect 1518 -1194 1524 -1188
rect 1518 -1200 1524 -1194
rect 1518 -1206 1524 -1200
rect 1518 -1212 1524 -1206
rect 1518 -1218 1524 -1212
rect 1518 -1224 1524 -1218
rect 1518 -1230 1524 -1224
rect 1518 -1236 1524 -1230
rect 1518 -1242 1524 -1236
rect 1518 -1248 1524 -1242
rect 1518 -1254 1524 -1248
rect 1518 -1260 1524 -1254
rect 1518 -1266 1524 -1260
rect 1518 -1272 1524 -1266
rect 1518 -1278 1524 -1272
rect 1518 -1284 1524 -1278
rect 1518 -1290 1524 -1284
rect 1518 -1296 1524 -1290
rect 1518 -1302 1524 -1296
rect 1518 -1308 1524 -1302
rect 1518 -1314 1524 -1308
rect 1518 -1320 1524 -1314
rect 1518 -1326 1524 -1320
rect 1518 -1332 1524 -1326
rect 1518 -1338 1524 -1332
rect 1518 -1344 1524 -1338
rect 1518 -1350 1524 -1344
rect 1518 -1356 1524 -1350
rect 1518 -1362 1524 -1356
rect 1518 -1368 1524 -1362
rect 1518 -1374 1524 -1368
rect 1518 -1380 1524 -1374
rect 1518 -1386 1524 -1380
rect 1518 -1392 1524 -1386
rect 1518 -1398 1524 -1392
rect 1518 -1404 1524 -1398
rect 1518 -1410 1524 -1404
rect 1518 -1416 1524 -1410
rect 1518 -1422 1524 -1416
rect 1518 -1428 1524 -1422
rect 1518 -1434 1524 -1428
rect 1518 -1440 1524 -1434
rect 1518 -1446 1524 -1440
rect 1518 -1452 1524 -1446
rect 1518 -1458 1524 -1452
rect 1518 -1464 1524 -1458
rect 1518 -1470 1524 -1464
rect 1518 -1476 1524 -1470
rect 1518 -1482 1524 -1476
rect 1518 -1488 1524 -1482
rect 1518 -1494 1524 -1488
rect 1518 -1500 1524 -1494
rect 1518 -1506 1524 -1500
rect 1518 -1512 1524 -1506
rect 1518 -1518 1524 -1512
rect 1518 -1524 1524 -1518
rect 1518 -1530 1524 -1524
rect 1518 -1536 1524 -1530
rect 1518 -1542 1524 -1536
rect 1518 -1548 1524 -1542
rect 1518 -1554 1524 -1548
rect 1518 -1560 1524 -1554
rect 1518 -1566 1524 -1560
rect 1518 -1572 1524 -1566
rect 1518 -1578 1524 -1572
rect 1518 -1584 1524 -1578
rect 1518 -1590 1524 -1584
rect 1518 -1596 1524 -1590
rect 1518 -1602 1524 -1596
rect 1518 -1608 1524 -1602
rect 1518 -1614 1524 -1608
rect 1518 -1620 1524 -1614
rect 1518 -1626 1524 -1620
rect 1518 -1632 1524 -1626
rect 1518 -1638 1524 -1632
rect 1518 -1644 1524 -1638
rect 1518 -1650 1524 -1644
rect 1518 -1656 1524 -1650
rect 1518 -1662 1524 -1656
rect 1518 -1668 1524 -1662
rect 1518 -1674 1524 -1668
rect 1518 -1680 1524 -1674
rect 1518 -1686 1524 -1680
rect 1518 -1692 1524 -1686
rect 1518 -1698 1524 -1692
rect 1518 -1704 1524 -1698
rect 1518 -1710 1524 -1704
rect 1518 -1716 1524 -1710
rect 1518 -1722 1524 -1716
rect 1518 -1728 1524 -1722
rect 1518 -1734 1524 -1728
rect 1518 -1740 1524 -1734
rect 1518 -1746 1524 -1740
rect 1518 -1752 1524 -1746
rect 1518 -1758 1524 -1752
rect 1518 -1764 1524 -1758
rect 1518 -1770 1524 -1764
rect 1518 -1776 1524 -1770
rect 1518 -1782 1524 -1776
rect 1518 -1788 1524 -1782
rect 1518 -1794 1524 -1788
rect 1518 -1800 1524 -1794
rect 1518 -1806 1524 -1800
rect 1518 -1812 1524 -1806
rect 1518 -1818 1524 -1812
rect 1518 -1824 1524 -1818
rect 1518 -1830 1524 -1824
rect 1518 -1836 1524 -1830
rect 1518 -1842 1524 -1836
rect 1518 -1848 1524 -1842
rect 1518 -1854 1524 -1848
rect 1518 -1860 1524 -1854
rect 1518 -1866 1524 -1860
rect 1518 -1872 1524 -1866
rect 1518 -1878 1524 -1872
rect 1518 -1884 1524 -1878
rect 1518 -1890 1524 -1884
rect 1518 -1896 1524 -1890
rect 1518 -1902 1524 -1896
rect 1518 -1908 1524 -1902
rect 1518 -1914 1524 -1908
rect 1518 -1920 1524 -1914
rect 1518 -1926 1524 -1920
rect 1518 -1932 1524 -1926
rect 1518 -1938 1524 -1932
rect 1518 -1944 1524 -1938
rect 1518 -1950 1524 -1944
rect 1518 -1956 1524 -1950
rect 1518 -1962 1524 -1956
rect 1518 -1968 1524 -1962
rect 1518 -1974 1524 -1968
rect 1518 -1980 1524 -1974
rect 1518 -1986 1524 -1980
rect 1518 -1992 1524 -1986
rect 1518 -1998 1524 -1992
rect 1518 -2004 1524 -1998
rect 1518 -2010 1524 -2004
rect 1518 -2016 1524 -2010
rect 1518 -2022 1524 -2016
rect 1518 -2028 1524 -2022
rect 1518 -2034 1524 -2028
rect 1518 -2040 1524 -2034
rect 1518 -2046 1524 -2040
rect 1518 -2052 1524 -2046
rect 1518 -2058 1524 -2052
rect 1518 -2064 1524 -2058
rect 1518 -2070 1524 -2064
rect 1518 -2076 1524 -2070
rect 1518 -2082 1524 -2076
rect 1518 -2088 1524 -2082
rect 1518 -2094 1524 -2088
rect 1518 -2100 1524 -2094
rect 1518 -2106 1524 -2100
rect 1518 -2112 1524 -2106
rect 1518 -2118 1524 -2112
rect 1518 -2124 1524 -2118
rect 1518 -2130 1524 -2124
rect 1518 -2136 1524 -2130
rect 1518 -2142 1524 -2136
rect 1518 -2148 1524 -2142
rect 1518 -2154 1524 -2148
rect 1518 -2160 1524 -2154
rect 1518 -2166 1524 -2160
rect 1518 -2238 1524 -2232
rect 1518 -2244 1524 -2238
rect 1518 -2250 1524 -2244
rect 1518 -2256 1524 -2250
rect 1518 -2262 1524 -2256
rect 1518 -2268 1524 -2262
rect 1518 -2274 1524 -2268
rect 1518 -2280 1524 -2274
rect 1518 -2286 1524 -2280
rect 1518 -2292 1524 -2286
rect 1518 -2298 1524 -2292
rect 1518 -2304 1524 -2298
rect 1518 -2310 1524 -2304
rect 1518 -2316 1524 -2310
rect 1518 -2322 1524 -2316
rect 1518 -2328 1524 -2322
rect 1518 -2334 1524 -2328
rect 1518 -2340 1524 -2334
rect 1518 -2346 1524 -2340
rect 1518 -2352 1524 -2346
rect 1518 -2358 1524 -2352
rect 1518 -2364 1524 -2358
rect 1518 -2370 1524 -2364
rect 1518 -2376 1524 -2370
rect 1518 -2382 1524 -2376
rect 1518 -2388 1524 -2382
rect 1518 -2394 1524 -2388
rect 1518 -2400 1524 -2394
rect 1518 -2406 1524 -2400
rect 1518 -2412 1524 -2406
rect 1518 -2418 1524 -2412
rect 1518 -2424 1524 -2418
rect 1518 -2430 1524 -2424
rect 1518 -2436 1524 -2430
rect 1518 -2442 1524 -2436
rect 1518 -2448 1524 -2442
rect 1518 -2454 1524 -2448
rect 1518 -2460 1524 -2454
rect 1518 -2466 1524 -2460
rect 1518 -2472 1524 -2466
rect 1518 -2478 1524 -2472
rect 1518 -2484 1524 -2478
rect 1518 -2490 1524 -2484
rect 1518 -2496 1524 -2490
rect 1518 -2502 1524 -2496
rect 1518 -2508 1524 -2502
rect 1518 -2514 1524 -2508
rect 1518 -2520 1524 -2514
rect 1518 -2526 1524 -2520
rect 1518 -2532 1524 -2526
rect 1518 -2538 1524 -2532
rect 1518 -2544 1524 -2538
rect 1518 -2550 1524 -2544
rect 1518 -2556 1524 -2550
rect 1518 -2562 1524 -2556
rect 1518 -2568 1524 -2562
rect 1518 -2574 1524 -2568
rect 1518 -2580 1524 -2574
rect 1518 -2586 1524 -2580
rect 1518 -2592 1524 -2586
rect 1518 -2598 1524 -2592
rect 1518 -2604 1524 -2598
rect 1518 -2610 1524 -2604
rect 1518 -2616 1524 -2610
rect 1518 -2622 1524 -2616
rect 1518 -2628 1524 -2622
rect 1518 -2634 1524 -2628
rect 1518 -2640 1524 -2634
rect 1518 -2646 1524 -2640
rect 1518 -2652 1524 -2646
rect 1518 -2658 1524 -2652
rect 1518 -2664 1524 -2658
rect 1518 -2670 1524 -2664
rect 1518 -2676 1524 -2670
rect 1518 -2682 1524 -2676
rect 1518 -2688 1524 -2682
rect 1518 -2694 1524 -2688
rect 1518 -2700 1524 -2694
rect 1518 -2706 1524 -2700
rect 1518 -2712 1524 -2706
rect 1518 -2718 1524 -2712
rect 1518 -2724 1524 -2718
rect 1518 -2730 1524 -2724
rect 1518 -2736 1524 -2730
rect 1518 -2742 1524 -2736
rect 1518 -2748 1524 -2742
rect 1518 -2754 1524 -2748
rect 1518 -2760 1524 -2754
rect 1518 -2766 1524 -2760
rect 1518 -2772 1524 -2766
rect 1518 -2778 1524 -2772
rect 1518 -2784 1524 -2778
rect 1518 -2790 1524 -2784
rect 1518 -2796 1524 -2790
rect 1518 -2880 1524 -2874
rect 1518 -2886 1524 -2880
rect 1518 -2892 1524 -2886
rect 1518 -2898 1524 -2892
rect 1518 -2904 1524 -2898
rect 1518 -2910 1524 -2904
rect 1518 -2916 1524 -2910
rect 1518 -2922 1524 -2916
rect 1518 -2928 1524 -2922
rect 1518 -2934 1524 -2928
rect 1518 -2940 1524 -2934
rect 1518 -2946 1524 -2940
rect 1518 -2952 1524 -2946
rect 1518 -2958 1524 -2952
rect 1518 -2964 1524 -2958
rect 1518 -2970 1524 -2964
rect 1518 -2976 1524 -2970
rect 1518 -2982 1524 -2976
rect 1518 -2988 1524 -2982
rect 1518 -2994 1524 -2988
rect 1518 -3000 1524 -2994
rect 1518 -3006 1524 -3000
rect 1518 -3012 1524 -3006
rect 1518 -3018 1524 -3012
rect 1518 -3024 1524 -3018
rect 1518 -3030 1524 -3024
rect 1518 -3036 1524 -3030
rect 1518 -3042 1524 -3036
rect 1518 -3048 1524 -3042
rect 1518 -3054 1524 -3048
rect 1518 -3060 1524 -3054
rect 1518 -3066 1524 -3060
rect 1518 -3072 1524 -3066
rect 1518 -3078 1524 -3072
rect 1518 -3084 1524 -3078
rect 1518 -3090 1524 -3084
rect 1518 -3096 1524 -3090
rect 1518 -3102 1524 -3096
rect 1518 -3108 1524 -3102
rect 1518 -3114 1524 -3108
rect 1518 -3120 1524 -3114
rect 1518 -3126 1524 -3120
rect 1518 -3132 1524 -3126
rect 1518 -3138 1524 -3132
rect 1518 -3144 1524 -3138
rect 1518 -3150 1524 -3144
rect 1518 -3156 1524 -3150
rect 1518 -3162 1524 -3156
rect 1518 -3168 1524 -3162
rect 1518 -3174 1524 -3168
rect 1518 -3180 1524 -3174
rect 1518 -3186 1524 -3180
rect 1518 -3192 1524 -3186
rect 1518 -3198 1524 -3192
rect 1518 -3204 1524 -3198
rect 1518 -3210 1524 -3204
rect 1518 -3216 1524 -3210
rect 1518 -3222 1524 -3216
rect 1518 -3228 1524 -3222
rect 1518 -3234 1524 -3228
rect 1518 -3276 1524 -3270
rect 1518 -3282 1524 -3276
rect 1518 -3288 1524 -3282
rect 1518 -3294 1524 -3288
rect 1518 -3300 1524 -3294
rect 1518 -3306 1524 -3300
rect 1518 -3312 1524 -3306
rect 1518 -3318 1524 -3312
rect 1518 -3324 1524 -3318
rect 1518 -3330 1524 -3324
rect 1518 -3336 1524 -3330
rect 1518 -3342 1524 -3336
rect 1518 -3348 1524 -3342
rect 1518 -3354 1524 -3348
rect 1518 -3360 1524 -3354
rect 1518 -3366 1524 -3360
rect 1518 -3372 1524 -3366
rect 1518 -3378 1524 -3372
rect 1518 -3384 1524 -3378
rect 1518 -3390 1524 -3384
rect 1518 -3396 1524 -3390
rect 1518 -3402 1524 -3396
rect 1518 -3408 1524 -3402
rect 1518 -3414 1524 -3408
rect 1518 -3420 1524 -3414
rect 1518 -3426 1524 -3420
rect 1518 -3432 1524 -3426
rect 1518 -3438 1524 -3432
rect 1518 -3444 1524 -3438
rect 1518 -3450 1524 -3444
rect 1518 -3456 1524 -3450
rect 1518 -3462 1524 -3456
rect 1518 -3468 1524 -3462
rect 1518 -3474 1524 -3468
rect 1518 -3480 1524 -3474
rect 1518 -3486 1524 -3480
rect 1524 -1140 1530 -1134
rect 1524 -1146 1530 -1140
rect 1524 -1152 1530 -1146
rect 1524 -1158 1530 -1152
rect 1524 -1164 1530 -1158
rect 1524 -1170 1530 -1164
rect 1524 -1176 1530 -1170
rect 1524 -1182 1530 -1176
rect 1524 -1188 1530 -1182
rect 1524 -1194 1530 -1188
rect 1524 -1200 1530 -1194
rect 1524 -1206 1530 -1200
rect 1524 -1212 1530 -1206
rect 1524 -1218 1530 -1212
rect 1524 -1224 1530 -1218
rect 1524 -1230 1530 -1224
rect 1524 -1236 1530 -1230
rect 1524 -1242 1530 -1236
rect 1524 -1248 1530 -1242
rect 1524 -1254 1530 -1248
rect 1524 -1260 1530 -1254
rect 1524 -1266 1530 -1260
rect 1524 -1272 1530 -1266
rect 1524 -1278 1530 -1272
rect 1524 -1284 1530 -1278
rect 1524 -1290 1530 -1284
rect 1524 -1296 1530 -1290
rect 1524 -1302 1530 -1296
rect 1524 -1308 1530 -1302
rect 1524 -1314 1530 -1308
rect 1524 -1320 1530 -1314
rect 1524 -1326 1530 -1320
rect 1524 -1332 1530 -1326
rect 1524 -1338 1530 -1332
rect 1524 -1344 1530 -1338
rect 1524 -1350 1530 -1344
rect 1524 -1356 1530 -1350
rect 1524 -1362 1530 -1356
rect 1524 -1368 1530 -1362
rect 1524 -1374 1530 -1368
rect 1524 -1380 1530 -1374
rect 1524 -1386 1530 -1380
rect 1524 -1392 1530 -1386
rect 1524 -1398 1530 -1392
rect 1524 -1404 1530 -1398
rect 1524 -1410 1530 -1404
rect 1524 -1416 1530 -1410
rect 1524 -1422 1530 -1416
rect 1524 -1428 1530 -1422
rect 1524 -1434 1530 -1428
rect 1524 -1440 1530 -1434
rect 1524 -1446 1530 -1440
rect 1524 -1452 1530 -1446
rect 1524 -1458 1530 -1452
rect 1524 -1464 1530 -1458
rect 1524 -1470 1530 -1464
rect 1524 -1476 1530 -1470
rect 1524 -1482 1530 -1476
rect 1524 -1488 1530 -1482
rect 1524 -1494 1530 -1488
rect 1524 -1500 1530 -1494
rect 1524 -1506 1530 -1500
rect 1524 -1512 1530 -1506
rect 1524 -1518 1530 -1512
rect 1524 -1524 1530 -1518
rect 1524 -1530 1530 -1524
rect 1524 -1536 1530 -1530
rect 1524 -1542 1530 -1536
rect 1524 -1548 1530 -1542
rect 1524 -1554 1530 -1548
rect 1524 -1560 1530 -1554
rect 1524 -1566 1530 -1560
rect 1524 -1572 1530 -1566
rect 1524 -1578 1530 -1572
rect 1524 -1584 1530 -1578
rect 1524 -1590 1530 -1584
rect 1524 -1596 1530 -1590
rect 1524 -1602 1530 -1596
rect 1524 -1608 1530 -1602
rect 1524 -1614 1530 -1608
rect 1524 -1620 1530 -1614
rect 1524 -1626 1530 -1620
rect 1524 -1632 1530 -1626
rect 1524 -1638 1530 -1632
rect 1524 -1644 1530 -1638
rect 1524 -1650 1530 -1644
rect 1524 -1656 1530 -1650
rect 1524 -1662 1530 -1656
rect 1524 -1668 1530 -1662
rect 1524 -1674 1530 -1668
rect 1524 -1680 1530 -1674
rect 1524 -1686 1530 -1680
rect 1524 -1692 1530 -1686
rect 1524 -1698 1530 -1692
rect 1524 -1704 1530 -1698
rect 1524 -1710 1530 -1704
rect 1524 -1716 1530 -1710
rect 1524 -1722 1530 -1716
rect 1524 -1728 1530 -1722
rect 1524 -1734 1530 -1728
rect 1524 -1740 1530 -1734
rect 1524 -1746 1530 -1740
rect 1524 -1752 1530 -1746
rect 1524 -1758 1530 -1752
rect 1524 -1764 1530 -1758
rect 1524 -1770 1530 -1764
rect 1524 -1776 1530 -1770
rect 1524 -1782 1530 -1776
rect 1524 -1788 1530 -1782
rect 1524 -1794 1530 -1788
rect 1524 -1800 1530 -1794
rect 1524 -1806 1530 -1800
rect 1524 -1812 1530 -1806
rect 1524 -1818 1530 -1812
rect 1524 -1824 1530 -1818
rect 1524 -1830 1530 -1824
rect 1524 -1836 1530 -1830
rect 1524 -1842 1530 -1836
rect 1524 -1848 1530 -1842
rect 1524 -1854 1530 -1848
rect 1524 -1860 1530 -1854
rect 1524 -1866 1530 -1860
rect 1524 -1872 1530 -1866
rect 1524 -1878 1530 -1872
rect 1524 -1884 1530 -1878
rect 1524 -1890 1530 -1884
rect 1524 -1896 1530 -1890
rect 1524 -1902 1530 -1896
rect 1524 -1908 1530 -1902
rect 1524 -1914 1530 -1908
rect 1524 -1920 1530 -1914
rect 1524 -1926 1530 -1920
rect 1524 -1932 1530 -1926
rect 1524 -1938 1530 -1932
rect 1524 -1944 1530 -1938
rect 1524 -1950 1530 -1944
rect 1524 -1956 1530 -1950
rect 1524 -1962 1530 -1956
rect 1524 -1968 1530 -1962
rect 1524 -1974 1530 -1968
rect 1524 -1980 1530 -1974
rect 1524 -1986 1530 -1980
rect 1524 -1992 1530 -1986
rect 1524 -1998 1530 -1992
rect 1524 -2004 1530 -1998
rect 1524 -2010 1530 -2004
rect 1524 -2016 1530 -2010
rect 1524 -2022 1530 -2016
rect 1524 -2028 1530 -2022
rect 1524 -2034 1530 -2028
rect 1524 -2040 1530 -2034
rect 1524 -2046 1530 -2040
rect 1524 -2052 1530 -2046
rect 1524 -2058 1530 -2052
rect 1524 -2064 1530 -2058
rect 1524 -2070 1530 -2064
rect 1524 -2076 1530 -2070
rect 1524 -2082 1530 -2076
rect 1524 -2088 1530 -2082
rect 1524 -2094 1530 -2088
rect 1524 -2100 1530 -2094
rect 1524 -2106 1530 -2100
rect 1524 -2112 1530 -2106
rect 1524 -2118 1530 -2112
rect 1524 -2124 1530 -2118
rect 1524 -2130 1530 -2124
rect 1524 -2136 1530 -2130
rect 1524 -2142 1530 -2136
rect 1524 -2148 1530 -2142
rect 1524 -2154 1530 -2148
rect 1524 -2160 1530 -2154
rect 1524 -2232 1530 -2226
rect 1524 -2238 1530 -2232
rect 1524 -2244 1530 -2238
rect 1524 -2250 1530 -2244
rect 1524 -2256 1530 -2250
rect 1524 -2262 1530 -2256
rect 1524 -2268 1530 -2262
rect 1524 -2274 1530 -2268
rect 1524 -2280 1530 -2274
rect 1524 -2286 1530 -2280
rect 1524 -2292 1530 -2286
rect 1524 -2298 1530 -2292
rect 1524 -2304 1530 -2298
rect 1524 -2310 1530 -2304
rect 1524 -2316 1530 -2310
rect 1524 -2322 1530 -2316
rect 1524 -2328 1530 -2322
rect 1524 -2334 1530 -2328
rect 1524 -2340 1530 -2334
rect 1524 -2346 1530 -2340
rect 1524 -2352 1530 -2346
rect 1524 -2358 1530 -2352
rect 1524 -2364 1530 -2358
rect 1524 -2370 1530 -2364
rect 1524 -2376 1530 -2370
rect 1524 -2382 1530 -2376
rect 1524 -2388 1530 -2382
rect 1524 -2394 1530 -2388
rect 1524 -2400 1530 -2394
rect 1524 -2406 1530 -2400
rect 1524 -2412 1530 -2406
rect 1524 -2418 1530 -2412
rect 1524 -2424 1530 -2418
rect 1524 -2430 1530 -2424
rect 1524 -2436 1530 -2430
rect 1524 -2442 1530 -2436
rect 1524 -2448 1530 -2442
rect 1524 -2454 1530 -2448
rect 1524 -2460 1530 -2454
rect 1524 -2466 1530 -2460
rect 1524 -2472 1530 -2466
rect 1524 -2478 1530 -2472
rect 1524 -2484 1530 -2478
rect 1524 -2490 1530 -2484
rect 1524 -2496 1530 -2490
rect 1524 -2502 1530 -2496
rect 1524 -2508 1530 -2502
rect 1524 -2514 1530 -2508
rect 1524 -2520 1530 -2514
rect 1524 -2526 1530 -2520
rect 1524 -2532 1530 -2526
rect 1524 -2538 1530 -2532
rect 1524 -2544 1530 -2538
rect 1524 -2550 1530 -2544
rect 1524 -2556 1530 -2550
rect 1524 -2562 1530 -2556
rect 1524 -2568 1530 -2562
rect 1524 -2574 1530 -2568
rect 1524 -2580 1530 -2574
rect 1524 -2586 1530 -2580
rect 1524 -2592 1530 -2586
rect 1524 -2598 1530 -2592
rect 1524 -2604 1530 -2598
rect 1524 -2610 1530 -2604
rect 1524 -2616 1530 -2610
rect 1524 -2622 1530 -2616
rect 1524 -2628 1530 -2622
rect 1524 -2634 1530 -2628
rect 1524 -2640 1530 -2634
rect 1524 -2646 1530 -2640
rect 1524 -2652 1530 -2646
rect 1524 -2658 1530 -2652
rect 1524 -2664 1530 -2658
rect 1524 -2670 1530 -2664
rect 1524 -2676 1530 -2670
rect 1524 -2682 1530 -2676
rect 1524 -2688 1530 -2682
rect 1524 -2694 1530 -2688
rect 1524 -2700 1530 -2694
rect 1524 -2706 1530 -2700
rect 1524 -2712 1530 -2706
rect 1524 -2718 1530 -2712
rect 1524 -2724 1530 -2718
rect 1524 -2730 1530 -2724
rect 1524 -2736 1530 -2730
rect 1524 -2742 1530 -2736
rect 1524 -2748 1530 -2742
rect 1524 -2754 1530 -2748
rect 1524 -2760 1530 -2754
rect 1524 -2766 1530 -2760
rect 1524 -2772 1530 -2766
rect 1524 -2778 1530 -2772
rect 1524 -2784 1530 -2778
rect 1524 -2790 1530 -2784
rect 1524 -2796 1530 -2790
rect 1524 -2880 1530 -2874
rect 1524 -2886 1530 -2880
rect 1524 -2892 1530 -2886
rect 1524 -2898 1530 -2892
rect 1524 -2904 1530 -2898
rect 1524 -2910 1530 -2904
rect 1524 -2916 1530 -2910
rect 1524 -2922 1530 -2916
rect 1524 -2928 1530 -2922
rect 1524 -2934 1530 -2928
rect 1524 -2940 1530 -2934
rect 1524 -2946 1530 -2940
rect 1524 -2952 1530 -2946
rect 1524 -2958 1530 -2952
rect 1524 -2964 1530 -2958
rect 1524 -2970 1530 -2964
rect 1524 -2976 1530 -2970
rect 1524 -2982 1530 -2976
rect 1524 -2988 1530 -2982
rect 1524 -2994 1530 -2988
rect 1524 -3000 1530 -2994
rect 1524 -3006 1530 -3000
rect 1524 -3012 1530 -3006
rect 1524 -3018 1530 -3012
rect 1524 -3024 1530 -3018
rect 1524 -3030 1530 -3024
rect 1524 -3036 1530 -3030
rect 1524 -3042 1530 -3036
rect 1524 -3048 1530 -3042
rect 1524 -3054 1530 -3048
rect 1524 -3060 1530 -3054
rect 1524 -3066 1530 -3060
rect 1524 -3072 1530 -3066
rect 1524 -3078 1530 -3072
rect 1524 -3084 1530 -3078
rect 1524 -3090 1530 -3084
rect 1524 -3096 1530 -3090
rect 1524 -3102 1530 -3096
rect 1524 -3108 1530 -3102
rect 1524 -3114 1530 -3108
rect 1524 -3120 1530 -3114
rect 1524 -3126 1530 -3120
rect 1524 -3132 1530 -3126
rect 1524 -3138 1530 -3132
rect 1524 -3144 1530 -3138
rect 1524 -3150 1530 -3144
rect 1524 -3156 1530 -3150
rect 1524 -3162 1530 -3156
rect 1524 -3168 1530 -3162
rect 1524 -3174 1530 -3168
rect 1524 -3180 1530 -3174
rect 1524 -3186 1530 -3180
rect 1524 -3192 1530 -3186
rect 1524 -3198 1530 -3192
rect 1524 -3204 1530 -3198
rect 1524 -3210 1530 -3204
rect 1524 -3216 1530 -3210
rect 1524 -3222 1530 -3216
rect 1524 -3228 1530 -3222
rect 1524 -3234 1530 -3228
rect 1524 -3276 1530 -3270
rect 1524 -3282 1530 -3276
rect 1524 -3288 1530 -3282
rect 1524 -3294 1530 -3288
rect 1524 -3300 1530 -3294
rect 1524 -3306 1530 -3300
rect 1524 -3312 1530 -3306
rect 1524 -3318 1530 -3312
rect 1524 -3324 1530 -3318
rect 1524 -3330 1530 -3324
rect 1524 -3336 1530 -3330
rect 1524 -3342 1530 -3336
rect 1524 -3348 1530 -3342
rect 1524 -3354 1530 -3348
rect 1524 -3360 1530 -3354
rect 1524 -3366 1530 -3360
rect 1524 -3372 1530 -3366
rect 1524 -3378 1530 -3372
rect 1524 -3384 1530 -3378
rect 1524 -3390 1530 -3384
rect 1524 -3396 1530 -3390
rect 1524 -3402 1530 -3396
rect 1524 -3408 1530 -3402
rect 1524 -3414 1530 -3408
rect 1524 -3420 1530 -3414
rect 1524 -3426 1530 -3420
rect 1524 -3432 1530 -3426
rect 1524 -3438 1530 -3432
rect 1524 -3444 1530 -3438
rect 1524 -3450 1530 -3444
rect 1524 -3456 1530 -3450
rect 1524 -3462 1530 -3456
rect 1524 -3468 1530 -3462
rect 1524 -3474 1530 -3468
rect 1524 -3480 1530 -3474
rect 1530 -1128 1536 -1122
rect 1530 -1134 1536 -1128
rect 1530 -1140 1536 -1134
rect 1530 -1146 1536 -1140
rect 1530 -1152 1536 -1146
rect 1530 -1158 1536 -1152
rect 1530 -1164 1536 -1158
rect 1530 -1170 1536 -1164
rect 1530 -1176 1536 -1170
rect 1530 -1182 1536 -1176
rect 1530 -1188 1536 -1182
rect 1530 -1194 1536 -1188
rect 1530 -1200 1536 -1194
rect 1530 -1206 1536 -1200
rect 1530 -1212 1536 -1206
rect 1530 -1218 1536 -1212
rect 1530 -1224 1536 -1218
rect 1530 -1230 1536 -1224
rect 1530 -1236 1536 -1230
rect 1530 -1242 1536 -1236
rect 1530 -1248 1536 -1242
rect 1530 -1254 1536 -1248
rect 1530 -1260 1536 -1254
rect 1530 -1266 1536 -1260
rect 1530 -1272 1536 -1266
rect 1530 -1278 1536 -1272
rect 1530 -1284 1536 -1278
rect 1530 -1290 1536 -1284
rect 1530 -1296 1536 -1290
rect 1530 -1302 1536 -1296
rect 1530 -1308 1536 -1302
rect 1530 -1314 1536 -1308
rect 1530 -1320 1536 -1314
rect 1530 -1326 1536 -1320
rect 1530 -1332 1536 -1326
rect 1530 -1338 1536 -1332
rect 1530 -1344 1536 -1338
rect 1530 -1350 1536 -1344
rect 1530 -1356 1536 -1350
rect 1530 -1362 1536 -1356
rect 1530 -1368 1536 -1362
rect 1530 -1374 1536 -1368
rect 1530 -1380 1536 -1374
rect 1530 -1386 1536 -1380
rect 1530 -1392 1536 -1386
rect 1530 -1398 1536 -1392
rect 1530 -1404 1536 -1398
rect 1530 -1410 1536 -1404
rect 1530 -1416 1536 -1410
rect 1530 -1422 1536 -1416
rect 1530 -1428 1536 -1422
rect 1530 -1434 1536 -1428
rect 1530 -1440 1536 -1434
rect 1530 -1446 1536 -1440
rect 1530 -1452 1536 -1446
rect 1530 -1458 1536 -1452
rect 1530 -1464 1536 -1458
rect 1530 -1470 1536 -1464
rect 1530 -1476 1536 -1470
rect 1530 -1482 1536 -1476
rect 1530 -1488 1536 -1482
rect 1530 -1494 1536 -1488
rect 1530 -1500 1536 -1494
rect 1530 -1506 1536 -1500
rect 1530 -1512 1536 -1506
rect 1530 -1518 1536 -1512
rect 1530 -1524 1536 -1518
rect 1530 -1530 1536 -1524
rect 1530 -1536 1536 -1530
rect 1530 -1542 1536 -1536
rect 1530 -1548 1536 -1542
rect 1530 -1554 1536 -1548
rect 1530 -1560 1536 -1554
rect 1530 -1566 1536 -1560
rect 1530 -1572 1536 -1566
rect 1530 -1578 1536 -1572
rect 1530 -1584 1536 -1578
rect 1530 -1590 1536 -1584
rect 1530 -1596 1536 -1590
rect 1530 -1602 1536 -1596
rect 1530 -1608 1536 -1602
rect 1530 -1614 1536 -1608
rect 1530 -1620 1536 -1614
rect 1530 -1626 1536 -1620
rect 1530 -1632 1536 -1626
rect 1530 -1638 1536 -1632
rect 1530 -1644 1536 -1638
rect 1530 -1650 1536 -1644
rect 1530 -1656 1536 -1650
rect 1530 -1662 1536 -1656
rect 1530 -1668 1536 -1662
rect 1530 -1674 1536 -1668
rect 1530 -1680 1536 -1674
rect 1530 -1686 1536 -1680
rect 1530 -1692 1536 -1686
rect 1530 -1698 1536 -1692
rect 1530 -1704 1536 -1698
rect 1530 -1710 1536 -1704
rect 1530 -1716 1536 -1710
rect 1530 -1722 1536 -1716
rect 1530 -1728 1536 -1722
rect 1530 -1734 1536 -1728
rect 1530 -1740 1536 -1734
rect 1530 -1746 1536 -1740
rect 1530 -1752 1536 -1746
rect 1530 -1758 1536 -1752
rect 1530 -1764 1536 -1758
rect 1530 -1770 1536 -1764
rect 1530 -1776 1536 -1770
rect 1530 -1782 1536 -1776
rect 1530 -1788 1536 -1782
rect 1530 -1794 1536 -1788
rect 1530 -1800 1536 -1794
rect 1530 -1806 1536 -1800
rect 1530 -1812 1536 -1806
rect 1530 -1818 1536 -1812
rect 1530 -1824 1536 -1818
rect 1530 -1830 1536 -1824
rect 1530 -1836 1536 -1830
rect 1530 -1842 1536 -1836
rect 1530 -1848 1536 -1842
rect 1530 -1854 1536 -1848
rect 1530 -1860 1536 -1854
rect 1530 -1866 1536 -1860
rect 1530 -1872 1536 -1866
rect 1530 -1878 1536 -1872
rect 1530 -1884 1536 -1878
rect 1530 -1890 1536 -1884
rect 1530 -1896 1536 -1890
rect 1530 -1902 1536 -1896
rect 1530 -1908 1536 -1902
rect 1530 -1914 1536 -1908
rect 1530 -1920 1536 -1914
rect 1530 -1926 1536 -1920
rect 1530 -1932 1536 -1926
rect 1530 -1938 1536 -1932
rect 1530 -1944 1536 -1938
rect 1530 -1950 1536 -1944
rect 1530 -1956 1536 -1950
rect 1530 -1962 1536 -1956
rect 1530 -1968 1536 -1962
rect 1530 -1974 1536 -1968
rect 1530 -1980 1536 -1974
rect 1530 -1986 1536 -1980
rect 1530 -1992 1536 -1986
rect 1530 -1998 1536 -1992
rect 1530 -2004 1536 -1998
rect 1530 -2010 1536 -2004
rect 1530 -2016 1536 -2010
rect 1530 -2022 1536 -2016
rect 1530 -2028 1536 -2022
rect 1530 -2034 1536 -2028
rect 1530 -2040 1536 -2034
rect 1530 -2046 1536 -2040
rect 1530 -2052 1536 -2046
rect 1530 -2058 1536 -2052
rect 1530 -2064 1536 -2058
rect 1530 -2070 1536 -2064
rect 1530 -2076 1536 -2070
rect 1530 -2082 1536 -2076
rect 1530 -2088 1536 -2082
rect 1530 -2094 1536 -2088
rect 1530 -2100 1536 -2094
rect 1530 -2106 1536 -2100
rect 1530 -2112 1536 -2106
rect 1530 -2118 1536 -2112
rect 1530 -2124 1536 -2118
rect 1530 -2130 1536 -2124
rect 1530 -2136 1536 -2130
rect 1530 -2142 1536 -2136
rect 1530 -2148 1536 -2142
rect 1530 -2154 1536 -2148
rect 1530 -2226 1536 -2220
rect 1530 -2232 1536 -2226
rect 1530 -2238 1536 -2232
rect 1530 -2244 1536 -2238
rect 1530 -2250 1536 -2244
rect 1530 -2256 1536 -2250
rect 1530 -2262 1536 -2256
rect 1530 -2268 1536 -2262
rect 1530 -2274 1536 -2268
rect 1530 -2280 1536 -2274
rect 1530 -2286 1536 -2280
rect 1530 -2292 1536 -2286
rect 1530 -2298 1536 -2292
rect 1530 -2304 1536 -2298
rect 1530 -2310 1536 -2304
rect 1530 -2316 1536 -2310
rect 1530 -2322 1536 -2316
rect 1530 -2328 1536 -2322
rect 1530 -2334 1536 -2328
rect 1530 -2340 1536 -2334
rect 1530 -2346 1536 -2340
rect 1530 -2352 1536 -2346
rect 1530 -2358 1536 -2352
rect 1530 -2364 1536 -2358
rect 1530 -2370 1536 -2364
rect 1530 -2376 1536 -2370
rect 1530 -2382 1536 -2376
rect 1530 -2388 1536 -2382
rect 1530 -2394 1536 -2388
rect 1530 -2400 1536 -2394
rect 1530 -2406 1536 -2400
rect 1530 -2412 1536 -2406
rect 1530 -2418 1536 -2412
rect 1530 -2424 1536 -2418
rect 1530 -2430 1536 -2424
rect 1530 -2436 1536 -2430
rect 1530 -2442 1536 -2436
rect 1530 -2448 1536 -2442
rect 1530 -2454 1536 -2448
rect 1530 -2460 1536 -2454
rect 1530 -2466 1536 -2460
rect 1530 -2472 1536 -2466
rect 1530 -2478 1536 -2472
rect 1530 -2484 1536 -2478
rect 1530 -2490 1536 -2484
rect 1530 -2496 1536 -2490
rect 1530 -2502 1536 -2496
rect 1530 -2508 1536 -2502
rect 1530 -2514 1536 -2508
rect 1530 -2520 1536 -2514
rect 1530 -2526 1536 -2520
rect 1530 -2532 1536 -2526
rect 1530 -2538 1536 -2532
rect 1530 -2544 1536 -2538
rect 1530 -2550 1536 -2544
rect 1530 -2556 1536 -2550
rect 1530 -2562 1536 -2556
rect 1530 -2568 1536 -2562
rect 1530 -2574 1536 -2568
rect 1530 -2580 1536 -2574
rect 1530 -2586 1536 -2580
rect 1530 -2592 1536 -2586
rect 1530 -2598 1536 -2592
rect 1530 -2604 1536 -2598
rect 1530 -2610 1536 -2604
rect 1530 -2616 1536 -2610
rect 1530 -2622 1536 -2616
rect 1530 -2628 1536 -2622
rect 1530 -2634 1536 -2628
rect 1530 -2640 1536 -2634
rect 1530 -2646 1536 -2640
rect 1530 -2652 1536 -2646
rect 1530 -2658 1536 -2652
rect 1530 -2664 1536 -2658
rect 1530 -2670 1536 -2664
rect 1530 -2676 1536 -2670
rect 1530 -2682 1536 -2676
rect 1530 -2688 1536 -2682
rect 1530 -2694 1536 -2688
rect 1530 -2700 1536 -2694
rect 1530 -2706 1536 -2700
rect 1530 -2712 1536 -2706
rect 1530 -2718 1536 -2712
rect 1530 -2724 1536 -2718
rect 1530 -2730 1536 -2724
rect 1530 -2736 1536 -2730
rect 1530 -2742 1536 -2736
rect 1530 -2748 1536 -2742
rect 1530 -2754 1536 -2748
rect 1530 -2760 1536 -2754
rect 1530 -2766 1536 -2760
rect 1530 -2772 1536 -2766
rect 1530 -2778 1536 -2772
rect 1530 -2784 1536 -2778
rect 1530 -2790 1536 -2784
rect 1530 -2874 1536 -2868
rect 1530 -2880 1536 -2874
rect 1530 -2886 1536 -2880
rect 1530 -2892 1536 -2886
rect 1530 -2898 1536 -2892
rect 1530 -2904 1536 -2898
rect 1530 -2910 1536 -2904
rect 1530 -2916 1536 -2910
rect 1530 -2922 1536 -2916
rect 1530 -2928 1536 -2922
rect 1530 -2934 1536 -2928
rect 1530 -2940 1536 -2934
rect 1530 -2946 1536 -2940
rect 1530 -2952 1536 -2946
rect 1530 -2958 1536 -2952
rect 1530 -2964 1536 -2958
rect 1530 -2970 1536 -2964
rect 1530 -2976 1536 -2970
rect 1530 -2982 1536 -2976
rect 1530 -2988 1536 -2982
rect 1530 -2994 1536 -2988
rect 1530 -3000 1536 -2994
rect 1530 -3006 1536 -3000
rect 1530 -3012 1536 -3006
rect 1530 -3018 1536 -3012
rect 1530 -3024 1536 -3018
rect 1530 -3030 1536 -3024
rect 1530 -3036 1536 -3030
rect 1530 -3042 1536 -3036
rect 1530 -3048 1536 -3042
rect 1530 -3054 1536 -3048
rect 1530 -3060 1536 -3054
rect 1530 -3066 1536 -3060
rect 1530 -3072 1536 -3066
rect 1530 -3078 1536 -3072
rect 1530 -3084 1536 -3078
rect 1530 -3090 1536 -3084
rect 1530 -3096 1536 -3090
rect 1530 -3102 1536 -3096
rect 1530 -3108 1536 -3102
rect 1530 -3114 1536 -3108
rect 1530 -3120 1536 -3114
rect 1530 -3126 1536 -3120
rect 1530 -3132 1536 -3126
rect 1530 -3138 1536 -3132
rect 1530 -3144 1536 -3138
rect 1530 -3150 1536 -3144
rect 1530 -3156 1536 -3150
rect 1530 -3162 1536 -3156
rect 1530 -3168 1536 -3162
rect 1530 -3174 1536 -3168
rect 1530 -3180 1536 -3174
rect 1530 -3186 1536 -3180
rect 1530 -3192 1536 -3186
rect 1530 -3198 1536 -3192
rect 1530 -3204 1536 -3198
rect 1530 -3210 1536 -3204
rect 1530 -3216 1536 -3210
rect 1530 -3222 1536 -3216
rect 1530 -3228 1536 -3222
rect 1530 -3234 1536 -3228
rect 1530 -3276 1536 -3270
rect 1530 -3282 1536 -3276
rect 1530 -3288 1536 -3282
rect 1530 -3294 1536 -3288
rect 1530 -3300 1536 -3294
rect 1530 -3306 1536 -3300
rect 1530 -3312 1536 -3306
rect 1530 -3318 1536 -3312
rect 1530 -3324 1536 -3318
rect 1530 -3330 1536 -3324
rect 1530 -3336 1536 -3330
rect 1530 -3342 1536 -3336
rect 1530 -3348 1536 -3342
rect 1530 -3354 1536 -3348
rect 1530 -3360 1536 -3354
rect 1530 -3366 1536 -3360
rect 1530 -3372 1536 -3366
rect 1530 -3378 1536 -3372
rect 1530 -3384 1536 -3378
rect 1530 -3390 1536 -3384
rect 1530 -3396 1536 -3390
rect 1530 -3402 1536 -3396
rect 1530 -3408 1536 -3402
rect 1530 -3414 1536 -3408
rect 1530 -3420 1536 -3414
rect 1530 -3426 1536 -3420
rect 1530 -3432 1536 -3426
rect 1530 -3438 1536 -3432
rect 1530 -3444 1536 -3438
rect 1530 -3450 1536 -3444
rect 1530 -3456 1536 -3450
rect 1530 -3462 1536 -3456
rect 1530 -3468 1536 -3462
rect 1530 -3474 1536 -3468
rect 1530 -3480 1536 -3474
rect 1536 -1122 1542 -1116
rect 1536 -1128 1542 -1122
rect 1536 -1134 1542 -1128
rect 1536 -1140 1542 -1134
rect 1536 -1146 1542 -1140
rect 1536 -1152 1542 -1146
rect 1536 -1158 1542 -1152
rect 1536 -1164 1542 -1158
rect 1536 -1170 1542 -1164
rect 1536 -1176 1542 -1170
rect 1536 -1182 1542 -1176
rect 1536 -1188 1542 -1182
rect 1536 -1194 1542 -1188
rect 1536 -1200 1542 -1194
rect 1536 -1206 1542 -1200
rect 1536 -1212 1542 -1206
rect 1536 -1218 1542 -1212
rect 1536 -1224 1542 -1218
rect 1536 -1230 1542 -1224
rect 1536 -1236 1542 -1230
rect 1536 -1242 1542 -1236
rect 1536 -1248 1542 -1242
rect 1536 -1254 1542 -1248
rect 1536 -1260 1542 -1254
rect 1536 -1266 1542 -1260
rect 1536 -1272 1542 -1266
rect 1536 -1278 1542 -1272
rect 1536 -1284 1542 -1278
rect 1536 -1290 1542 -1284
rect 1536 -1296 1542 -1290
rect 1536 -1302 1542 -1296
rect 1536 -1308 1542 -1302
rect 1536 -1314 1542 -1308
rect 1536 -1320 1542 -1314
rect 1536 -1326 1542 -1320
rect 1536 -1332 1542 -1326
rect 1536 -1338 1542 -1332
rect 1536 -1344 1542 -1338
rect 1536 -1350 1542 -1344
rect 1536 -1356 1542 -1350
rect 1536 -1362 1542 -1356
rect 1536 -1368 1542 -1362
rect 1536 -1374 1542 -1368
rect 1536 -1380 1542 -1374
rect 1536 -1386 1542 -1380
rect 1536 -1392 1542 -1386
rect 1536 -1398 1542 -1392
rect 1536 -1404 1542 -1398
rect 1536 -1410 1542 -1404
rect 1536 -1416 1542 -1410
rect 1536 -1422 1542 -1416
rect 1536 -1428 1542 -1422
rect 1536 -1434 1542 -1428
rect 1536 -1440 1542 -1434
rect 1536 -1446 1542 -1440
rect 1536 -1452 1542 -1446
rect 1536 -1458 1542 -1452
rect 1536 -1464 1542 -1458
rect 1536 -1470 1542 -1464
rect 1536 -1476 1542 -1470
rect 1536 -1482 1542 -1476
rect 1536 -1488 1542 -1482
rect 1536 -1494 1542 -1488
rect 1536 -1500 1542 -1494
rect 1536 -1506 1542 -1500
rect 1536 -1512 1542 -1506
rect 1536 -1518 1542 -1512
rect 1536 -1524 1542 -1518
rect 1536 -1530 1542 -1524
rect 1536 -1536 1542 -1530
rect 1536 -1542 1542 -1536
rect 1536 -1548 1542 -1542
rect 1536 -1554 1542 -1548
rect 1536 -1560 1542 -1554
rect 1536 -1566 1542 -1560
rect 1536 -1572 1542 -1566
rect 1536 -1578 1542 -1572
rect 1536 -1584 1542 -1578
rect 1536 -1590 1542 -1584
rect 1536 -1596 1542 -1590
rect 1536 -1602 1542 -1596
rect 1536 -1608 1542 -1602
rect 1536 -1614 1542 -1608
rect 1536 -1620 1542 -1614
rect 1536 -1626 1542 -1620
rect 1536 -1632 1542 -1626
rect 1536 -1638 1542 -1632
rect 1536 -1644 1542 -1638
rect 1536 -1650 1542 -1644
rect 1536 -1656 1542 -1650
rect 1536 -1662 1542 -1656
rect 1536 -1668 1542 -1662
rect 1536 -1674 1542 -1668
rect 1536 -1680 1542 -1674
rect 1536 -1686 1542 -1680
rect 1536 -1692 1542 -1686
rect 1536 -1698 1542 -1692
rect 1536 -1704 1542 -1698
rect 1536 -1710 1542 -1704
rect 1536 -1716 1542 -1710
rect 1536 -1722 1542 -1716
rect 1536 -1728 1542 -1722
rect 1536 -1734 1542 -1728
rect 1536 -1740 1542 -1734
rect 1536 -1746 1542 -1740
rect 1536 -1752 1542 -1746
rect 1536 -1758 1542 -1752
rect 1536 -1764 1542 -1758
rect 1536 -1770 1542 -1764
rect 1536 -1776 1542 -1770
rect 1536 -1782 1542 -1776
rect 1536 -1788 1542 -1782
rect 1536 -1794 1542 -1788
rect 1536 -1800 1542 -1794
rect 1536 -1806 1542 -1800
rect 1536 -1812 1542 -1806
rect 1536 -1818 1542 -1812
rect 1536 -1824 1542 -1818
rect 1536 -1830 1542 -1824
rect 1536 -1836 1542 -1830
rect 1536 -1842 1542 -1836
rect 1536 -1848 1542 -1842
rect 1536 -1854 1542 -1848
rect 1536 -1860 1542 -1854
rect 1536 -1866 1542 -1860
rect 1536 -1872 1542 -1866
rect 1536 -1878 1542 -1872
rect 1536 -1884 1542 -1878
rect 1536 -1890 1542 -1884
rect 1536 -1896 1542 -1890
rect 1536 -1902 1542 -1896
rect 1536 -1908 1542 -1902
rect 1536 -1914 1542 -1908
rect 1536 -1920 1542 -1914
rect 1536 -1926 1542 -1920
rect 1536 -1932 1542 -1926
rect 1536 -1938 1542 -1932
rect 1536 -1944 1542 -1938
rect 1536 -1950 1542 -1944
rect 1536 -1956 1542 -1950
rect 1536 -1962 1542 -1956
rect 1536 -1968 1542 -1962
rect 1536 -1974 1542 -1968
rect 1536 -1980 1542 -1974
rect 1536 -1986 1542 -1980
rect 1536 -1992 1542 -1986
rect 1536 -1998 1542 -1992
rect 1536 -2004 1542 -1998
rect 1536 -2010 1542 -2004
rect 1536 -2016 1542 -2010
rect 1536 -2022 1542 -2016
rect 1536 -2028 1542 -2022
rect 1536 -2034 1542 -2028
rect 1536 -2040 1542 -2034
rect 1536 -2046 1542 -2040
rect 1536 -2052 1542 -2046
rect 1536 -2058 1542 -2052
rect 1536 -2064 1542 -2058
rect 1536 -2070 1542 -2064
rect 1536 -2076 1542 -2070
rect 1536 -2082 1542 -2076
rect 1536 -2088 1542 -2082
rect 1536 -2094 1542 -2088
rect 1536 -2100 1542 -2094
rect 1536 -2106 1542 -2100
rect 1536 -2112 1542 -2106
rect 1536 -2118 1542 -2112
rect 1536 -2124 1542 -2118
rect 1536 -2130 1542 -2124
rect 1536 -2136 1542 -2130
rect 1536 -2142 1542 -2136
rect 1536 -2220 1542 -2214
rect 1536 -2226 1542 -2220
rect 1536 -2232 1542 -2226
rect 1536 -2238 1542 -2232
rect 1536 -2244 1542 -2238
rect 1536 -2250 1542 -2244
rect 1536 -2256 1542 -2250
rect 1536 -2262 1542 -2256
rect 1536 -2268 1542 -2262
rect 1536 -2274 1542 -2268
rect 1536 -2280 1542 -2274
rect 1536 -2286 1542 -2280
rect 1536 -2292 1542 -2286
rect 1536 -2298 1542 -2292
rect 1536 -2304 1542 -2298
rect 1536 -2310 1542 -2304
rect 1536 -2316 1542 -2310
rect 1536 -2322 1542 -2316
rect 1536 -2328 1542 -2322
rect 1536 -2334 1542 -2328
rect 1536 -2340 1542 -2334
rect 1536 -2346 1542 -2340
rect 1536 -2352 1542 -2346
rect 1536 -2358 1542 -2352
rect 1536 -2364 1542 -2358
rect 1536 -2370 1542 -2364
rect 1536 -2376 1542 -2370
rect 1536 -2382 1542 -2376
rect 1536 -2388 1542 -2382
rect 1536 -2394 1542 -2388
rect 1536 -2400 1542 -2394
rect 1536 -2406 1542 -2400
rect 1536 -2412 1542 -2406
rect 1536 -2418 1542 -2412
rect 1536 -2424 1542 -2418
rect 1536 -2430 1542 -2424
rect 1536 -2436 1542 -2430
rect 1536 -2442 1542 -2436
rect 1536 -2448 1542 -2442
rect 1536 -2454 1542 -2448
rect 1536 -2460 1542 -2454
rect 1536 -2466 1542 -2460
rect 1536 -2472 1542 -2466
rect 1536 -2478 1542 -2472
rect 1536 -2484 1542 -2478
rect 1536 -2490 1542 -2484
rect 1536 -2496 1542 -2490
rect 1536 -2502 1542 -2496
rect 1536 -2508 1542 -2502
rect 1536 -2514 1542 -2508
rect 1536 -2520 1542 -2514
rect 1536 -2526 1542 -2520
rect 1536 -2532 1542 -2526
rect 1536 -2538 1542 -2532
rect 1536 -2544 1542 -2538
rect 1536 -2550 1542 -2544
rect 1536 -2556 1542 -2550
rect 1536 -2562 1542 -2556
rect 1536 -2568 1542 -2562
rect 1536 -2574 1542 -2568
rect 1536 -2580 1542 -2574
rect 1536 -2586 1542 -2580
rect 1536 -2592 1542 -2586
rect 1536 -2598 1542 -2592
rect 1536 -2604 1542 -2598
rect 1536 -2610 1542 -2604
rect 1536 -2616 1542 -2610
rect 1536 -2622 1542 -2616
rect 1536 -2628 1542 -2622
rect 1536 -2634 1542 -2628
rect 1536 -2640 1542 -2634
rect 1536 -2646 1542 -2640
rect 1536 -2652 1542 -2646
rect 1536 -2658 1542 -2652
rect 1536 -2664 1542 -2658
rect 1536 -2670 1542 -2664
rect 1536 -2676 1542 -2670
rect 1536 -2682 1542 -2676
rect 1536 -2688 1542 -2682
rect 1536 -2694 1542 -2688
rect 1536 -2700 1542 -2694
rect 1536 -2706 1542 -2700
rect 1536 -2712 1542 -2706
rect 1536 -2718 1542 -2712
rect 1536 -2724 1542 -2718
rect 1536 -2730 1542 -2724
rect 1536 -2736 1542 -2730
rect 1536 -2742 1542 -2736
rect 1536 -2748 1542 -2742
rect 1536 -2754 1542 -2748
rect 1536 -2760 1542 -2754
rect 1536 -2766 1542 -2760
rect 1536 -2772 1542 -2766
rect 1536 -2778 1542 -2772
rect 1536 -2784 1542 -2778
rect 1536 -2868 1542 -2862
rect 1536 -2874 1542 -2868
rect 1536 -2880 1542 -2874
rect 1536 -2886 1542 -2880
rect 1536 -2892 1542 -2886
rect 1536 -2898 1542 -2892
rect 1536 -2904 1542 -2898
rect 1536 -2910 1542 -2904
rect 1536 -2916 1542 -2910
rect 1536 -2922 1542 -2916
rect 1536 -2928 1542 -2922
rect 1536 -2934 1542 -2928
rect 1536 -2940 1542 -2934
rect 1536 -2946 1542 -2940
rect 1536 -2952 1542 -2946
rect 1536 -2958 1542 -2952
rect 1536 -2964 1542 -2958
rect 1536 -2970 1542 -2964
rect 1536 -2976 1542 -2970
rect 1536 -2982 1542 -2976
rect 1536 -2988 1542 -2982
rect 1536 -2994 1542 -2988
rect 1536 -3000 1542 -2994
rect 1536 -3006 1542 -3000
rect 1536 -3012 1542 -3006
rect 1536 -3018 1542 -3012
rect 1536 -3024 1542 -3018
rect 1536 -3030 1542 -3024
rect 1536 -3036 1542 -3030
rect 1536 -3042 1542 -3036
rect 1536 -3048 1542 -3042
rect 1536 -3054 1542 -3048
rect 1536 -3060 1542 -3054
rect 1536 -3066 1542 -3060
rect 1536 -3072 1542 -3066
rect 1536 -3078 1542 -3072
rect 1536 -3084 1542 -3078
rect 1536 -3090 1542 -3084
rect 1536 -3096 1542 -3090
rect 1536 -3102 1542 -3096
rect 1536 -3108 1542 -3102
rect 1536 -3114 1542 -3108
rect 1536 -3120 1542 -3114
rect 1536 -3126 1542 -3120
rect 1536 -3132 1542 -3126
rect 1536 -3138 1542 -3132
rect 1536 -3144 1542 -3138
rect 1536 -3150 1542 -3144
rect 1536 -3156 1542 -3150
rect 1536 -3162 1542 -3156
rect 1536 -3168 1542 -3162
rect 1536 -3174 1542 -3168
rect 1536 -3180 1542 -3174
rect 1536 -3186 1542 -3180
rect 1536 -3192 1542 -3186
rect 1536 -3198 1542 -3192
rect 1536 -3204 1542 -3198
rect 1536 -3210 1542 -3204
rect 1536 -3216 1542 -3210
rect 1536 -3222 1542 -3216
rect 1536 -3228 1542 -3222
rect 1536 -3234 1542 -3228
rect 1536 -3276 1542 -3270
rect 1536 -3282 1542 -3276
rect 1536 -3288 1542 -3282
rect 1536 -3294 1542 -3288
rect 1536 -3300 1542 -3294
rect 1536 -3306 1542 -3300
rect 1536 -3312 1542 -3306
rect 1536 -3318 1542 -3312
rect 1536 -3324 1542 -3318
rect 1536 -3330 1542 -3324
rect 1536 -3336 1542 -3330
rect 1536 -3342 1542 -3336
rect 1536 -3348 1542 -3342
rect 1536 -3354 1542 -3348
rect 1536 -3360 1542 -3354
rect 1536 -3366 1542 -3360
rect 1536 -3372 1542 -3366
rect 1536 -3378 1542 -3372
rect 1536 -3384 1542 -3378
rect 1536 -3390 1542 -3384
rect 1536 -3396 1542 -3390
rect 1536 -3402 1542 -3396
rect 1536 -3408 1542 -3402
rect 1536 -3414 1542 -3408
rect 1536 -3420 1542 -3414
rect 1536 -3426 1542 -3420
rect 1536 -3432 1542 -3426
rect 1536 -3438 1542 -3432
rect 1536 -3444 1542 -3438
rect 1536 -3450 1542 -3444
rect 1536 -3456 1542 -3450
rect 1536 -3462 1542 -3456
rect 1536 -3468 1542 -3462
rect 1536 -3474 1542 -3468
rect 1536 -3480 1542 -3474
rect 1542 -1110 1548 -1104
rect 1542 -1116 1548 -1110
rect 1542 -1122 1548 -1116
rect 1542 -1128 1548 -1122
rect 1542 -1134 1548 -1128
rect 1542 -1140 1548 -1134
rect 1542 -1146 1548 -1140
rect 1542 -1152 1548 -1146
rect 1542 -1158 1548 -1152
rect 1542 -1164 1548 -1158
rect 1542 -1170 1548 -1164
rect 1542 -1176 1548 -1170
rect 1542 -1182 1548 -1176
rect 1542 -1188 1548 -1182
rect 1542 -1194 1548 -1188
rect 1542 -1200 1548 -1194
rect 1542 -1206 1548 -1200
rect 1542 -1212 1548 -1206
rect 1542 -1218 1548 -1212
rect 1542 -1224 1548 -1218
rect 1542 -1230 1548 -1224
rect 1542 -1236 1548 -1230
rect 1542 -1242 1548 -1236
rect 1542 -1248 1548 -1242
rect 1542 -1254 1548 -1248
rect 1542 -1260 1548 -1254
rect 1542 -1266 1548 -1260
rect 1542 -1272 1548 -1266
rect 1542 -1278 1548 -1272
rect 1542 -1284 1548 -1278
rect 1542 -1290 1548 -1284
rect 1542 -1296 1548 -1290
rect 1542 -1302 1548 -1296
rect 1542 -1308 1548 -1302
rect 1542 -1314 1548 -1308
rect 1542 -1320 1548 -1314
rect 1542 -1326 1548 -1320
rect 1542 -1332 1548 -1326
rect 1542 -1338 1548 -1332
rect 1542 -1344 1548 -1338
rect 1542 -1350 1548 -1344
rect 1542 -1356 1548 -1350
rect 1542 -1362 1548 -1356
rect 1542 -1368 1548 -1362
rect 1542 -1374 1548 -1368
rect 1542 -1380 1548 -1374
rect 1542 -1386 1548 -1380
rect 1542 -1392 1548 -1386
rect 1542 -1398 1548 -1392
rect 1542 -1404 1548 -1398
rect 1542 -1410 1548 -1404
rect 1542 -1416 1548 -1410
rect 1542 -1422 1548 -1416
rect 1542 -1428 1548 -1422
rect 1542 -1434 1548 -1428
rect 1542 -1440 1548 -1434
rect 1542 -1446 1548 -1440
rect 1542 -1452 1548 -1446
rect 1542 -1458 1548 -1452
rect 1542 -1464 1548 -1458
rect 1542 -1470 1548 -1464
rect 1542 -1476 1548 -1470
rect 1542 -1482 1548 -1476
rect 1542 -1488 1548 -1482
rect 1542 -1494 1548 -1488
rect 1542 -1500 1548 -1494
rect 1542 -1506 1548 -1500
rect 1542 -1512 1548 -1506
rect 1542 -1518 1548 -1512
rect 1542 -1524 1548 -1518
rect 1542 -1530 1548 -1524
rect 1542 -1536 1548 -1530
rect 1542 -1542 1548 -1536
rect 1542 -1548 1548 -1542
rect 1542 -1554 1548 -1548
rect 1542 -1560 1548 -1554
rect 1542 -1566 1548 -1560
rect 1542 -1572 1548 -1566
rect 1542 -1578 1548 -1572
rect 1542 -1584 1548 -1578
rect 1542 -1590 1548 -1584
rect 1542 -1596 1548 -1590
rect 1542 -1602 1548 -1596
rect 1542 -1608 1548 -1602
rect 1542 -1614 1548 -1608
rect 1542 -1620 1548 -1614
rect 1542 -1626 1548 -1620
rect 1542 -1632 1548 -1626
rect 1542 -1638 1548 -1632
rect 1542 -1644 1548 -1638
rect 1542 -1650 1548 -1644
rect 1542 -1656 1548 -1650
rect 1542 -1662 1548 -1656
rect 1542 -1668 1548 -1662
rect 1542 -1674 1548 -1668
rect 1542 -1680 1548 -1674
rect 1542 -1686 1548 -1680
rect 1542 -1692 1548 -1686
rect 1542 -1698 1548 -1692
rect 1542 -1704 1548 -1698
rect 1542 -1710 1548 -1704
rect 1542 -1716 1548 -1710
rect 1542 -1722 1548 -1716
rect 1542 -1728 1548 -1722
rect 1542 -1734 1548 -1728
rect 1542 -1740 1548 -1734
rect 1542 -1746 1548 -1740
rect 1542 -1752 1548 -1746
rect 1542 -1758 1548 -1752
rect 1542 -1764 1548 -1758
rect 1542 -1770 1548 -1764
rect 1542 -1776 1548 -1770
rect 1542 -1782 1548 -1776
rect 1542 -1788 1548 -1782
rect 1542 -1794 1548 -1788
rect 1542 -1800 1548 -1794
rect 1542 -1806 1548 -1800
rect 1542 -1812 1548 -1806
rect 1542 -1818 1548 -1812
rect 1542 -1824 1548 -1818
rect 1542 -1830 1548 -1824
rect 1542 -1836 1548 -1830
rect 1542 -1842 1548 -1836
rect 1542 -1848 1548 -1842
rect 1542 -1854 1548 -1848
rect 1542 -1860 1548 -1854
rect 1542 -1866 1548 -1860
rect 1542 -1872 1548 -1866
rect 1542 -1878 1548 -1872
rect 1542 -1884 1548 -1878
rect 1542 -1890 1548 -1884
rect 1542 -1896 1548 -1890
rect 1542 -1902 1548 -1896
rect 1542 -1908 1548 -1902
rect 1542 -1914 1548 -1908
rect 1542 -1920 1548 -1914
rect 1542 -1926 1548 -1920
rect 1542 -1932 1548 -1926
rect 1542 -1938 1548 -1932
rect 1542 -1944 1548 -1938
rect 1542 -1950 1548 -1944
rect 1542 -1956 1548 -1950
rect 1542 -1962 1548 -1956
rect 1542 -1968 1548 -1962
rect 1542 -1974 1548 -1968
rect 1542 -1980 1548 -1974
rect 1542 -1986 1548 -1980
rect 1542 -1992 1548 -1986
rect 1542 -1998 1548 -1992
rect 1542 -2004 1548 -1998
rect 1542 -2010 1548 -2004
rect 1542 -2016 1548 -2010
rect 1542 -2022 1548 -2016
rect 1542 -2028 1548 -2022
rect 1542 -2034 1548 -2028
rect 1542 -2040 1548 -2034
rect 1542 -2046 1548 -2040
rect 1542 -2052 1548 -2046
rect 1542 -2058 1548 -2052
rect 1542 -2064 1548 -2058
rect 1542 -2070 1548 -2064
rect 1542 -2076 1548 -2070
rect 1542 -2082 1548 -2076
rect 1542 -2088 1548 -2082
rect 1542 -2094 1548 -2088
rect 1542 -2100 1548 -2094
rect 1542 -2106 1548 -2100
rect 1542 -2112 1548 -2106
rect 1542 -2118 1548 -2112
rect 1542 -2124 1548 -2118
rect 1542 -2130 1548 -2124
rect 1542 -2136 1548 -2130
rect 1542 -2208 1548 -2202
rect 1542 -2214 1548 -2208
rect 1542 -2220 1548 -2214
rect 1542 -2226 1548 -2220
rect 1542 -2232 1548 -2226
rect 1542 -2238 1548 -2232
rect 1542 -2244 1548 -2238
rect 1542 -2250 1548 -2244
rect 1542 -2256 1548 -2250
rect 1542 -2262 1548 -2256
rect 1542 -2268 1548 -2262
rect 1542 -2274 1548 -2268
rect 1542 -2280 1548 -2274
rect 1542 -2286 1548 -2280
rect 1542 -2292 1548 -2286
rect 1542 -2298 1548 -2292
rect 1542 -2304 1548 -2298
rect 1542 -2310 1548 -2304
rect 1542 -2316 1548 -2310
rect 1542 -2322 1548 -2316
rect 1542 -2328 1548 -2322
rect 1542 -2334 1548 -2328
rect 1542 -2340 1548 -2334
rect 1542 -2346 1548 -2340
rect 1542 -2352 1548 -2346
rect 1542 -2358 1548 -2352
rect 1542 -2364 1548 -2358
rect 1542 -2370 1548 -2364
rect 1542 -2376 1548 -2370
rect 1542 -2382 1548 -2376
rect 1542 -2388 1548 -2382
rect 1542 -2394 1548 -2388
rect 1542 -2400 1548 -2394
rect 1542 -2406 1548 -2400
rect 1542 -2412 1548 -2406
rect 1542 -2418 1548 -2412
rect 1542 -2424 1548 -2418
rect 1542 -2430 1548 -2424
rect 1542 -2436 1548 -2430
rect 1542 -2442 1548 -2436
rect 1542 -2448 1548 -2442
rect 1542 -2454 1548 -2448
rect 1542 -2460 1548 -2454
rect 1542 -2466 1548 -2460
rect 1542 -2472 1548 -2466
rect 1542 -2478 1548 -2472
rect 1542 -2484 1548 -2478
rect 1542 -2490 1548 -2484
rect 1542 -2496 1548 -2490
rect 1542 -2502 1548 -2496
rect 1542 -2508 1548 -2502
rect 1542 -2514 1548 -2508
rect 1542 -2520 1548 -2514
rect 1542 -2526 1548 -2520
rect 1542 -2532 1548 -2526
rect 1542 -2538 1548 -2532
rect 1542 -2544 1548 -2538
rect 1542 -2550 1548 -2544
rect 1542 -2556 1548 -2550
rect 1542 -2562 1548 -2556
rect 1542 -2568 1548 -2562
rect 1542 -2574 1548 -2568
rect 1542 -2580 1548 -2574
rect 1542 -2586 1548 -2580
rect 1542 -2592 1548 -2586
rect 1542 -2598 1548 -2592
rect 1542 -2604 1548 -2598
rect 1542 -2610 1548 -2604
rect 1542 -2616 1548 -2610
rect 1542 -2622 1548 -2616
rect 1542 -2628 1548 -2622
rect 1542 -2634 1548 -2628
rect 1542 -2640 1548 -2634
rect 1542 -2646 1548 -2640
rect 1542 -2652 1548 -2646
rect 1542 -2658 1548 -2652
rect 1542 -2664 1548 -2658
rect 1542 -2670 1548 -2664
rect 1542 -2676 1548 -2670
rect 1542 -2682 1548 -2676
rect 1542 -2688 1548 -2682
rect 1542 -2694 1548 -2688
rect 1542 -2700 1548 -2694
rect 1542 -2706 1548 -2700
rect 1542 -2712 1548 -2706
rect 1542 -2718 1548 -2712
rect 1542 -2724 1548 -2718
rect 1542 -2730 1548 -2724
rect 1542 -2736 1548 -2730
rect 1542 -2742 1548 -2736
rect 1542 -2748 1548 -2742
rect 1542 -2754 1548 -2748
rect 1542 -2760 1548 -2754
rect 1542 -2766 1548 -2760
rect 1542 -2772 1548 -2766
rect 1542 -2778 1548 -2772
rect 1542 -2784 1548 -2778
rect 1542 -2868 1548 -2862
rect 1542 -2874 1548 -2868
rect 1542 -2880 1548 -2874
rect 1542 -2886 1548 -2880
rect 1542 -2892 1548 -2886
rect 1542 -2898 1548 -2892
rect 1542 -2904 1548 -2898
rect 1542 -2910 1548 -2904
rect 1542 -2916 1548 -2910
rect 1542 -2922 1548 -2916
rect 1542 -2928 1548 -2922
rect 1542 -2934 1548 -2928
rect 1542 -2940 1548 -2934
rect 1542 -2946 1548 -2940
rect 1542 -2952 1548 -2946
rect 1542 -2958 1548 -2952
rect 1542 -2964 1548 -2958
rect 1542 -2970 1548 -2964
rect 1542 -2976 1548 -2970
rect 1542 -2982 1548 -2976
rect 1542 -2988 1548 -2982
rect 1542 -2994 1548 -2988
rect 1542 -3000 1548 -2994
rect 1542 -3006 1548 -3000
rect 1542 -3012 1548 -3006
rect 1542 -3018 1548 -3012
rect 1542 -3024 1548 -3018
rect 1542 -3030 1548 -3024
rect 1542 -3036 1548 -3030
rect 1542 -3042 1548 -3036
rect 1542 -3048 1548 -3042
rect 1542 -3054 1548 -3048
rect 1542 -3060 1548 -3054
rect 1542 -3066 1548 -3060
rect 1542 -3072 1548 -3066
rect 1542 -3078 1548 -3072
rect 1542 -3084 1548 -3078
rect 1542 -3090 1548 -3084
rect 1542 -3096 1548 -3090
rect 1542 -3102 1548 -3096
rect 1542 -3108 1548 -3102
rect 1542 -3114 1548 -3108
rect 1542 -3120 1548 -3114
rect 1542 -3126 1548 -3120
rect 1542 -3132 1548 -3126
rect 1542 -3138 1548 -3132
rect 1542 -3144 1548 -3138
rect 1542 -3150 1548 -3144
rect 1542 -3156 1548 -3150
rect 1542 -3162 1548 -3156
rect 1542 -3168 1548 -3162
rect 1542 -3174 1548 -3168
rect 1542 -3180 1548 -3174
rect 1542 -3186 1548 -3180
rect 1542 -3192 1548 -3186
rect 1542 -3198 1548 -3192
rect 1542 -3204 1548 -3198
rect 1542 -3210 1548 -3204
rect 1542 -3216 1548 -3210
rect 1542 -3222 1548 -3216
rect 1542 -3228 1548 -3222
rect 1542 -3234 1548 -3228
rect 1542 -3276 1548 -3270
rect 1542 -3282 1548 -3276
rect 1542 -3288 1548 -3282
rect 1542 -3294 1548 -3288
rect 1542 -3300 1548 -3294
rect 1542 -3306 1548 -3300
rect 1542 -3312 1548 -3306
rect 1542 -3318 1548 -3312
rect 1542 -3324 1548 -3318
rect 1542 -3330 1548 -3324
rect 1542 -3336 1548 -3330
rect 1542 -3342 1548 -3336
rect 1542 -3348 1548 -3342
rect 1542 -3354 1548 -3348
rect 1542 -3360 1548 -3354
rect 1542 -3366 1548 -3360
rect 1542 -3372 1548 -3366
rect 1542 -3378 1548 -3372
rect 1542 -3384 1548 -3378
rect 1542 -3390 1548 -3384
rect 1542 -3396 1548 -3390
rect 1542 -3402 1548 -3396
rect 1542 -3408 1548 -3402
rect 1542 -3414 1548 -3408
rect 1542 -3420 1548 -3414
rect 1542 -3426 1548 -3420
rect 1542 -3432 1548 -3426
rect 1542 -3438 1548 -3432
rect 1542 -3444 1548 -3438
rect 1542 -3450 1548 -3444
rect 1542 -3456 1548 -3450
rect 1542 -3462 1548 -3456
rect 1542 -3468 1548 -3462
rect 1542 -3474 1548 -3468
rect 1548 -1098 1554 -1092
rect 1548 -1104 1554 -1098
rect 1548 -1110 1554 -1104
rect 1548 -1116 1554 -1110
rect 1548 -1122 1554 -1116
rect 1548 -1128 1554 -1122
rect 1548 -1134 1554 -1128
rect 1548 -1140 1554 -1134
rect 1548 -1146 1554 -1140
rect 1548 -1152 1554 -1146
rect 1548 -1158 1554 -1152
rect 1548 -1164 1554 -1158
rect 1548 -1170 1554 -1164
rect 1548 -1176 1554 -1170
rect 1548 -1182 1554 -1176
rect 1548 -1188 1554 -1182
rect 1548 -1194 1554 -1188
rect 1548 -1200 1554 -1194
rect 1548 -1206 1554 -1200
rect 1548 -1212 1554 -1206
rect 1548 -1218 1554 -1212
rect 1548 -1224 1554 -1218
rect 1548 -1230 1554 -1224
rect 1548 -1236 1554 -1230
rect 1548 -1242 1554 -1236
rect 1548 -1248 1554 -1242
rect 1548 -1254 1554 -1248
rect 1548 -1260 1554 -1254
rect 1548 -1266 1554 -1260
rect 1548 -1272 1554 -1266
rect 1548 -1278 1554 -1272
rect 1548 -1284 1554 -1278
rect 1548 -1290 1554 -1284
rect 1548 -1296 1554 -1290
rect 1548 -1302 1554 -1296
rect 1548 -1308 1554 -1302
rect 1548 -1314 1554 -1308
rect 1548 -1320 1554 -1314
rect 1548 -1326 1554 -1320
rect 1548 -1332 1554 -1326
rect 1548 -1338 1554 -1332
rect 1548 -1344 1554 -1338
rect 1548 -1350 1554 -1344
rect 1548 -1356 1554 -1350
rect 1548 -1362 1554 -1356
rect 1548 -1368 1554 -1362
rect 1548 -1374 1554 -1368
rect 1548 -1380 1554 -1374
rect 1548 -1386 1554 -1380
rect 1548 -1392 1554 -1386
rect 1548 -1398 1554 -1392
rect 1548 -1404 1554 -1398
rect 1548 -1410 1554 -1404
rect 1548 -1416 1554 -1410
rect 1548 -1422 1554 -1416
rect 1548 -1428 1554 -1422
rect 1548 -1434 1554 -1428
rect 1548 -1440 1554 -1434
rect 1548 -1446 1554 -1440
rect 1548 -1452 1554 -1446
rect 1548 -1458 1554 -1452
rect 1548 -1464 1554 -1458
rect 1548 -1470 1554 -1464
rect 1548 -1476 1554 -1470
rect 1548 -1482 1554 -1476
rect 1548 -1488 1554 -1482
rect 1548 -1494 1554 -1488
rect 1548 -1500 1554 -1494
rect 1548 -1506 1554 -1500
rect 1548 -1512 1554 -1506
rect 1548 -1518 1554 -1512
rect 1548 -1524 1554 -1518
rect 1548 -1530 1554 -1524
rect 1548 -1536 1554 -1530
rect 1548 -1542 1554 -1536
rect 1548 -1548 1554 -1542
rect 1548 -1554 1554 -1548
rect 1548 -1560 1554 -1554
rect 1548 -1566 1554 -1560
rect 1548 -1572 1554 -1566
rect 1548 -1578 1554 -1572
rect 1548 -1584 1554 -1578
rect 1548 -1590 1554 -1584
rect 1548 -1596 1554 -1590
rect 1548 -1602 1554 -1596
rect 1548 -1608 1554 -1602
rect 1548 -1614 1554 -1608
rect 1548 -1620 1554 -1614
rect 1548 -1626 1554 -1620
rect 1548 -1632 1554 -1626
rect 1548 -1638 1554 -1632
rect 1548 -1644 1554 -1638
rect 1548 -1650 1554 -1644
rect 1548 -1656 1554 -1650
rect 1548 -1662 1554 -1656
rect 1548 -1668 1554 -1662
rect 1548 -1674 1554 -1668
rect 1548 -1680 1554 -1674
rect 1548 -1686 1554 -1680
rect 1548 -1692 1554 -1686
rect 1548 -1698 1554 -1692
rect 1548 -1704 1554 -1698
rect 1548 -1710 1554 -1704
rect 1548 -1716 1554 -1710
rect 1548 -1722 1554 -1716
rect 1548 -1728 1554 -1722
rect 1548 -1734 1554 -1728
rect 1548 -1740 1554 -1734
rect 1548 -1746 1554 -1740
rect 1548 -1752 1554 -1746
rect 1548 -1758 1554 -1752
rect 1548 -1764 1554 -1758
rect 1548 -1770 1554 -1764
rect 1548 -1776 1554 -1770
rect 1548 -1782 1554 -1776
rect 1548 -1788 1554 -1782
rect 1548 -1794 1554 -1788
rect 1548 -1800 1554 -1794
rect 1548 -1806 1554 -1800
rect 1548 -1812 1554 -1806
rect 1548 -1818 1554 -1812
rect 1548 -1824 1554 -1818
rect 1548 -1830 1554 -1824
rect 1548 -1836 1554 -1830
rect 1548 -1842 1554 -1836
rect 1548 -1848 1554 -1842
rect 1548 -1854 1554 -1848
rect 1548 -1860 1554 -1854
rect 1548 -1866 1554 -1860
rect 1548 -1872 1554 -1866
rect 1548 -1878 1554 -1872
rect 1548 -1884 1554 -1878
rect 1548 -1890 1554 -1884
rect 1548 -1896 1554 -1890
rect 1548 -1902 1554 -1896
rect 1548 -1908 1554 -1902
rect 1548 -1914 1554 -1908
rect 1548 -1920 1554 -1914
rect 1548 -1926 1554 -1920
rect 1548 -1932 1554 -1926
rect 1548 -1938 1554 -1932
rect 1548 -1944 1554 -1938
rect 1548 -1950 1554 -1944
rect 1548 -1956 1554 -1950
rect 1548 -1962 1554 -1956
rect 1548 -1968 1554 -1962
rect 1548 -1974 1554 -1968
rect 1548 -1980 1554 -1974
rect 1548 -1986 1554 -1980
rect 1548 -1992 1554 -1986
rect 1548 -1998 1554 -1992
rect 1548 -2004 1554 -1998
rect 1548 -2010 1554 -2004
rect 1548 -2016 1554 -2010
rect 1548 -2022 1554 -2016
rect 1548 -2028 1554 -2022
rect 1548 -2034 1554 -2028
rect 1548 -2040 1554 -2034
rect 1548 -2046 1554 -2040
rect 1548 -2052 1554 -2046
rect 1548 -2058 1554 -2052
rect 1548 -2064 1554 -2058
rect 1548 -2070 1554 -2064
rect 1548 -2076 1554 -2070
rect 1548 -2082 1554 -2076
rect 1548 -2088 1554 -2082
rect 1548 -2094 1554 -2088
rect 1548 -2100 1554 -2094
rect 1548 -2106 1554 -2100
rect 1548 -2112 1554 -2106
rect 1548 -2118 1554 -2112
rect 1548 -2124 1554 -2118
rect 1548 -2130 1554 -2124
rect 1548 -2202 1554 -2196
rect 1548 -2208 1554 -2202
rect 1548 -2214 1554 -2208
rect 1548 -2220 1554 -2214
rect 1548 -2226 1554 -2220
rect 1548 -2232 1554 -2226
rect 1548 -2238 1554 -2232
rect 1548 -2244 1554 -2238
rect 1548 -2250 1554 -2244
rect 1548 -2256 1554 -2250
rect 1548 -2262 1554 -2256
rect 1548 -2268 1554 -2262
rect 1548 -2274 1554 -2268
rect 1548 -2280 1554 -2274
rect 1548 -2286 1554 -2280
rect 1548 -2292 1554 -2286
rect 1548 -2298 1554 -2292
rect 1548 -2304 1554 -2298
rect 1548 -2310 1554 -2304
rect 1548 -2316 1554 -2310
rect 1548 -2322 1554 -2316
rect 1548 -2328 1554 -2322
rect 1548 -2334 1554 -2328
rect 1548 -2340 1554 -2334
rect 1548 -2346 1554 -2340
rect 1548 -2352 1554 -2346
rect 1548 -2358 1554 -2352
rect 1548 -2364 1554 -2358
rect 1548 -2370 1554 -2364
rect 1548 -2376 1554 -2370
rect 1548 -2382 1554 -2376
rect 1548 -2388 1554 -2382
rect 1548 -2394 1554 -2388
rect 1548 -2400 1554 -2394
rect 1548 -2406 1554 -2400
rect 1548 -2412 1554 -2406
rect 1548 -2418 1554 -2412
rect 1548 -2424 1554 -2418
rect 1548 -2430 1554 -2424
rect 1548 -2436 1554 -2430
rect 1548 -2442 1554 -2436
rect 1548 -2448 1554 -2442
rect 1548 -2454 1554 -2448
rect 1548 -2460 1554 -2454
rect 1548 -2466 1554 -2460
rect 1548 -2472 1554 -2466
rect 1548 -2478 1554 -2472
rect 1548 -2484 1554 -2478
rect 1548 -2490 1554 -2484
rect 1548 -2496 1554 -2490
rect 1548 -2502 1554 -2496
rect 1548 -2508 1554 -2502
rect 1548 -2514 1554 -2508
rect 1548 -2520 1554 -2514
rect 1548 -2526 1554 -2520
rect 1548 -2532 1554 -2526
rect 1548 -2538 1554 -2532
rect 1548 -2544 1554 -2538
rect 1548 -2550 1554 -2544
rect 1548 -2556 1554 -2550
rect 1548 -2562 1554 -2556
rect 1548 -2568 1554 -2562
rect 1548 -2574 1554 -2568
rect 1548 -2580 1554 -2574
rect 1548 -2586 1554 -2580
rect 1548 -2592 1554 -2586
rect 1548 -2598 1554 -2592
rect 1548 -2604 1554 -2598
rect 1548 -2610 1554 -2604
rect 1548 -2616 1554 -2610
rect 1548 -2622 1554 -2616
rect 1548 -2628 1554 -2622
rect 1548 -2634 1554 -2628
rect 1548 -2640 1554 -2634
rect 1548 -2646 1554 -2640
rect 1548 -2652 1554 -2646
rect 1548 -2658 1554 -2652
rect 1548 -2664 1554 -2658
rect 1548 -2670 1554 -2664
rect 1548 -2676 1554 -2670
rect 1548 -2682 1554 -2676
rect 1548 -2688 1554 -2682
rect 1548 -2694 1554 -2688
rect 1548 -2700 1554 -2694
rect 1548 -2706 1554 -2700
rect 1548 -2712 1554 -2706
rect 1548 -2718 1554 -2712
rect 1548 -2724 1554 -2718
rect 1548 -2730 1554 -2724
rect 1548 -2736 1554 -2730
rect 1548 -2742 1554 -2736
rect 1548 -2748 1554 -2742
rect 1548 -2754 1554 -2748
rect 1548 -2760 1554 -2754
rect 1548 -2766 1554 -2760
rect 1548 -2772 1554 -2766
rect 1548 -2778 1554 -2772
rect 1548 -2862 1554 -2856
rect 1548 -2868 1554 -2862
rect 1548 -2874 1554 -2868
rect 1548 -2880 1554 -2874
rect 1548 -2886 1554 -2880
rect 1548 -2892 1554 -2886
rect 1548 -2898 1554 -2892
rect 1548 -2904 1554 -2898
rect 1548 -2910 1554 -2904
rect 1548 -2916 1554 -2910
rect 1548 -2922 1554 -2916
rect 1548 -2928 1554 -2922
rect 1548 -2934 1554 -2928
rect 1548 -2940 1554 -2934
rect 1548 -2946 1554 -2940
rect 1548 -2952 1554 -2946
rect 1548 -2958 1554 -2952
rect 1548 -2964 1554 -2958
rect 1548 -2970 1554 -2964
rect 1548 -2976 1554 -2970
rect 1548 -2982 1554 -2976
rect 1548 -2988 1554 -2982
rect 1548 -2994 1554 -2988
rect 1548 -3000 1554 -2994
rect 1548 -3006 1554 -3000
rect 1548 -3012 1554 -3006
rect 1548 -3018 1554 -3012
rect 1548 -3024 1554 -3018
rect 1548 -3030 1554 -3024
rect 1548 -3036 1554 -3030
rect 1548 -3042 1554 -3036
rect 1548 -3048 1554 -3042
rect 1548 -3054 1554 -3048
rect 1548 -3060 1554 -3054
rect 1548 -3066 1554 -3060
rect 1548 -3072 1554 -3066
rect 1548 -3078 1554 -3072
rect 1548 -3084 1554 -3078
rect 1548 -3090 1554 -3084
rect 1548 -3096 1554 -3090
rect 1548 -3102 1554 -3096
rect 1548 -3108 1554 -3102
rect 1548 -3114 1554 -3108
rect 1548 -3120 1554 -3114
rect 1548 -3126 1554 -3120
rect 1548 -3132 1554 -3126
rect 1548 -3138 1554 -3132
rect 1548 -3144 1554 -3138
rect 1548 -3150 1554 -3144
rect 1548 -3156 1554 -3150
rect 1548 -3162 1554 -3156
rect 1548 -3168 1554 -3162
rect 1548 -3174 1554 -3168
rect 1548 -3180 1554 -3174
rect 1548 -3186 1554 -3180
rect 1548 -3192 1554 -3186
rect 1548 -3198 1554 -3192
rect 1548 -3204 1554 -3198
rect 1548 -3210 1554 -3204
rect 1548 -3216 1554 -3210
rect 1548 -3222 1554 -3216
rect 1548 -3228 1554 -3222
rect 1548 -3234 1554 -3228
rect 1548 -3276 1554 -3270
rect 1548 -3282 1554 -3276
rect 1548 -3288 1554 -3282
rect 1548 -3294 1554 -3288
rect 1548 -3300 1554 -3294
rect 1548 -3306 1554 -3300
rect 1548 -3312 1554 -3306
rect 1548 -3318 1554 -3312
rect 1548 -3324 1554 -3318
rect 1548 -3330 1554 -3324
rect 1548 -3336 1554 -3330
rect 1548 -3342 1554 -3336
rect 1548 -3348 1554 -3342
rect 1548 -3354 1554 -3348
rect 1548 -3360 1554 -3354
rect 1548 -3366 1554 -3360
rect 1548 -3372 1554 -3366
rect 1548 -3378 1554 -3372
rect 1548 -3384 1554 -3378
rect 1548 -3390 1554 -3384
rect 1548 -3396 1554 -3390
rect 1548 -3402 1554 -3396
rect 1548 -3408 1554 -3402
rect 1548 -3414 1554 -3408
rect 1548 -3420 1554 -3414
rect 1548 -3426 1554 -3420
rect 1548 -3432 1554 -3426
rect 1548 -3438 1554 -3432
rect 1548 -3444 1554 -3438
rect 1548 -3450 1554 -3444
rect 1548 -3456 1554 -3450
rect 1548 -3462 1554 -3456
rect 1548 -3468 1554 -3462
rect 1548 -3474 1554 -3468
rect 1554 -1092 1560 -1086
rect 1554 -1098 1560 -1092
rect 1554 -1104 1560 -1098
rect 1554 -1110 1560 -1104
rect 1554 -1116 1560 -1110
rect 1554 -1122 1560 -1116
rect 1554 -1128 1560 -1122
rect 1554 -1134 1560 -1128
rect 1554 -1140 1560 -1134
rect 1554 -1146 1560 -1140
rect 1554 -1152 1560 -1146
rect 1554 -1158 1560 -1152
rect 1554 -1164 1560 -1158
rect 1554 -1170 1560 -1164
rect 1554 -1176 1560 -1170
rect 1554 -1182 1560 -1176
rect 1554 -1188 1560 -1182
rect 1554 -1194 1560 -1188
rect 1554 -1200 1560 -1194
rect 1554 -1206 1560 -1200
rect 1554 -1212 1560 -1206
rect 1554 -1218 1560 -1212
rect 1554 -1224 1560 -1218
rect 1554 -1230 1560 -1224
rect 1554 -1236 1560 -1230
rect 1554 -1242 1560 -1236
rect 1554 -1248 1560 -1242
rect 1554 -1254 1560 -1248
rect 1554 -1260 1560 -1254
rect 1554 -1266 1560 -1260
rect 1554 -1272 1560 -1266
rect 1554 -1278 1560 -1272
rect 1554 -1284 1560 -1278
rect 1554 -1290 1560 -1284
rect 1554 -1296 1560 -1290
rect 1554 -1302 1560 -1296
rect 1554 -1308 1560 -1302
rect 1554 -1314 1560 -1308
rect 1554 -1320 1560 -1314
rect 1554 -1326 1560 -1320
rect 1554 -1332 1560 -1326
rect 1554 -1338 1560 -1332
rect 1554 -1344 1560 -1338
rect 1554 -1350 1560 -1344
rect 1554 -1356 1560 -1350
rect 1554 -1362 1560 -1356
rect 1554 -1368 1560 -1362
rect 1554 -1374 1560 -1368
rect 1554 -1380 1560 -1374
rect 1554 -1386 1560 -1380
rect 1554 -1392 1560 -1386
rect 1554 -1398 1560 -1392
rect 1554 -1404 1560 -1398
rect 1554 -1410 1560 -1404
rect 1554 -1416 1560 -1410
rect 1554 -1422 1560 -1416
rect 1554 -1428 1560 -1422
rect 1554 -1434 1560 -1428
rect 1554 -1440 1560 -1434
rect 1554 -1446 1560 -1440
rect 1554 -1452 1560 -1446
rect 1554 -1458 1560 -1452
rect 1554 -1464 1560 -1458
rect 1554 -1470 1560 -1464
rect 1554 -1476 1560 -1470
rect 1554 -1482 1560 -1476
rect 1554 -1488 1560 -1482
rect 1554 -1494 1560 -1488
rect 1554 -1500 1560 -1494
rect 1554 -1506 1560 -1500
rect 1554 -1512 1560 -1506
rect 1554 -1518 1560 -1512
rect 1554 -1524 1560 -1518
rect 1554 -1530 1560 -1524
rect 1554 -1536 1560 -1530
rect 1554 -1542 1560 -1536
rect 1554 -1548 1560 -1542
rect 1554 -1554 1560 -1548
rect 1554 -1560 1560 -1554
rect 1554 -1566 1560 -1560
rect 1554 -1572 1560 -1566
rect 1554 -1578 1560 -1572
rect 1554 -1584 1560 -1578
rect 1554 -1590 1560 -1584
rect 1554 -1596 1560 -1590
rect 1554 -1602 1560 -1596
rect 1554 -1608 1560 -1602
rect 1554 -1614 1560 -1608
rect 1554 -1620 1560 -1614
rect 1554 -1626 1560 -1620
rect 1554 -1632 1560 -1626
rect 1554 -1638 1560 -1632
rect 1554 -1644 1560 -1638
rect 1554 -1650 1560 -1644
rect 1554 -1656 1560 -1650
rect 1554 -1662 1560 -1656
rect 1554 -1668 1560 -1662
rect 1554 -1674 1560 -1668
rect 1554 -1680 1560 -1674
rect 1554 -1686 1560 -1680
rect 1554 -1692 1560 -1686
rect 1554 -1698 1560 -1692
rect 1554 -1704 1560 -1698
rect 1554 -1710 1560 -1704
rect 1554 -1716 1560 -1710
rect 1554 -1722 1560 -1716
rect 1554 -1728 1560 -1722
rect 1554 -1734 1560 -1728
rect 1554 -1740 1560 -1734
rect 1554 -1746 1560 -1740
rect 1554 -1752 1560 -1746
rect 1554 -1758 1560 -1752
rect 1554 -1764 1560 -1758
rect 1554 -1770 1560 -1764
rect 1554 -1776 1560 -1770
rect 1554 -1782 1560 -1776
rect 1554 -1788 1560 -1782
rect 1554 -1794 1560 -1788
rect 1554 -1800 1560 -1794
rect 1554 -1806 1560 -1800
rect 1554 -1812 1560 -1806
rect 1554 -1818 1560 -1812
rect 1554 -1824 1560 -1818
rect 1554 -1830 1560 -1824
rect 1554 -1836 1560 -1830
rect 1554 -1842 1560 -1836
rect 1554 -1848 1560 -1842
rect 1554 -1854 1560 -1848
rect 1554 -1860 1560 -1854
rect 1554 -1866 1560 -1860
rect 1554 -1872 1560 -1866
rect 1554 -1878 1560 -1872
rect 1554 -1884 1560 -1878
rect 1554 -1890 1560 -1884
rect 1554 -1896 1560 -1890
rect 1554 -1902 1560 -1896
rect 1554 -1908 1560 -1902
rect 1554 -1914 1560 -1908
rect 1554 -1920 1560 -1914
rect 1554 -1926 1560 -1920
rect 1554 -1932 1560 -1926
rect 1554 -1938 1560 -1932
rect 1554 -1944 1560 -1938
rect 1554 -1950 1560 -1944
rect 1554 -1956 1560 -1950
rect 1554 -1962 1560 -1956
rect 1554 -1968 1560 -1962
rect 1554 -1974 1560 -1968
rect 1554 -1980 1560 -1974
rect 1554 -1986 1560 -1980
rect 1554 -1992 1560 -1986
rect 1554 -1998 1560 -1992
rect 1554 -2004 1560 -1998
rect 1554 -2010 1560 -2004
rect 1554 -2016 1560 -2010
rect 1554 -2022 1560 -2016
rect 1554 -2028 1560 -2022
rect 1554 -2034 1560 -2028
rect 1554 -2040 1560 -2034
rect 1554 -2046 1560 -2040
rect 1554 -2052 1560 -2046
rect 1554 -2058 1560 -2052
rect 1554 -2064 1560 -2058
rect 1554 -2070 1560 -2064
rect 1554 -2076 1560 -2070
rect 1554 -2082 1560 -2076
rect 1554 -2088 1560 -2082
rect 1554 -2094 1560 -2088
rect 1554 -2100 1560 -2094
rect 1554 -2106 1560 -2100
rect 1554 -2112 1560 -2106
rect 1554 -2118 1560 -2112
rect 1554 -2124 1560 -2118
rect 1554 -2196 1560 -2190
rect 1554 -2202 1560 -2196
rect 1554 -2208 1560 -2202
rect 1554 -2214 1560 -2208
rect 1554 -2220 1560 -2214
rect 1554 -2226 1560 -2220
rect 1554 -2232 1560 -2226
rect 1554 -2238 1560 -2232
rect 1554 -2244 1560 -2238
rect 1554 -2250 1560 -2244
rect 1554 -2256 1560 -2250
rect 1554 -2262 1560 -2256
rect 1554 -2268 1560 -2262
rect 1554 -2274 1560 -2268
rect 1554 -2280 1560 -2274
rect 1554 -2286 1560 -2280
rect 1554 -2292 1560 -2286
rect 1554 -2298 1560 -2292
rect 1554 -2304 1560 -2298
rect 1554 -2310 1560 -2304
rect 1554 -2316 1560 -2310
rect 1554 -2322 1560 -2316
rect 1554 -2328 1560 -2322
rect 1554 -2334 1560 -2328
rect 1554 -2340 1560 -2334
rect 1554 -2346 1560 -2340
rect 1554 -2352 1560 -2346
rect 1554 -2358 1560 -2352
rect 1554 -2364 1560 -2358
rect 1554 -2370 1560 -2364
rect 1554 -2376 1560 -2370
rect 1554 -2382 1560 -2376
rect 1554 -2388 1560 -2382
rect 1554 -2394 1560 -2388
rect 1554 -2400 1560 -2394
rect 1554 -2406 1560 -2400
rect 1554 -2412 1560 -2406
rect 1554 -2418 1560 -2412
rect 1554 -2424 1560 -2418
rect 1554 -2430 1560 -2424
rect 1554 -2436 1560 -2430
rect 1554 -2442 1560 -2436
rect 1554 -2448 1560 -2442
rect 1554 -2454 1560 -2448
rect 1554 -2460 1560 -2454
rect 1554 -2466 1560 -2460
rect 1554 -2472 1560 -2466
rect 1554 -2478 1560 -2472
rect 1554 -2484 1560 -2478
rect 1554 -2490 1560 -2484
rect 1554 -2496 1560 -2490
rect 1554 -2502 1560 -2496
rect 1554 -2508 1560 -2502
rect 1554 -2514 1560 -2508
rect 1554 -2520 1560 -2514
rect 1554 -2526 1560 -2520
rect 1554 -2532 1560 -2526
rect 1554 -2538 1560 -2532
rect 1554 -2544 1560 -2538
rect 1554 -2550 1560 -2544
rect 1554 -2556 1560 -2550
rect 1554 -2562 1560 -2556
rect 1554 -2568 1560 -2562
rect 1554 -2574 1560 -2568
rect 1554 -2580 1560 -2574
rect 1554 -2586 1560 -2580
rect 1554 -2592 1560 -2586
rect 1554 -2598 1560 -2592
rect 1554 -2604 1560 -2598
rect 1554 -2610 1560 -2604
rect 1554 -2616 1560 -2610
rect 1554 -2622 1560 -2616
rect 1554 -2628 1560 -2622
rect 1554 -2634 1560 -2628
rect 1554 -2640 1560 -2634
rect 1554 -2646 1560 -2640
rect 1554 -2652 1560 -2646
rect 1554 -2658 1560 -2652
rect 1554 -2664 1560 -2658
rect 1554 -2670 1560 -2664
rect 1554 -2676 1560 -2670
rect 1554 -2682 1560 -2676
rect 1554 -2688 1560 -2682
rect 1554 -2694 1560 -2688
rect 1554 -2700 1560 -2694
rect 1554 -2706 1560 -2700
rect 1554 -2712 1560 -2706
rect 1554 -2718 1560 -2712
rect 1554 -2724 1560 -2718
rect 1554 -2730 1560 -2724
rect 1554 -2736 1560 -2730
rect 1554 -2742 1560 -2736
rect 1554 -2748 1560 -2742
rect 1554 -2754 1560 -2748
rect 1554 -2760 1560 -2754
rect 1554 -2766 1560 -2760
rect 1554 -2772 1560 -2766
rect 1554 -2778 1560 -2772
rect 1554 -2856 1560 -2850
rect 1554 -2862 1560 -2856
rect 1554 -2868 1560 -2862
rect 1554 -2874 1560 -2868
rect 1554 -2880 1560 -2874
rect 1554 -2886 1560 -2880
rect 1554 -2892 1560 -2886
rect 1554 -2898 1560 -2892
rect 1554 -2904 1560 -2898
rect 1554 -2910 1560 -2904
rect 1554 -2916 1560 -2910
rect 1554 -2922 1560 -2916
rect 1554 -2928 1560 -2922
rect 1554 -2934 1560 -2928
rect 1554 -2940 1560 -2934
rect 1554 -2946 1560 -2940
rect 1554 -2952 1560 -2946
rect 1554 -2958 1560 -2952
rect 1554 -2964 1560 -2958
rect 1554 -2970 1560 -2964
rect 1554 -2976 1560 -2970
rect 1554 -2982 1560 -2976
rect 1554 -2988 1560 -2982
rect 1554 -2994 1560 -2988
rect 1554 -3000 1560 -2994
rect 1554 -3006 1560 -3000
rect 1554 -3012 1560 -3006
rect 1554 -3018 1560 -3012
rect 1554 -3024 1560 -3018
rect 1554 -3030 1560 -3024
rect 1554 -3036 1560 -3030
rect 1554 -3042 1560 -3036
rect 1554 -3048 1560 -3042
rect 1554 -3054 1560 -3048
rect 1554 -3060 1560 -3054
rect 1554 -3066 1560 -3060
rect 1554 -3072 1560 -3066
rect 1554 -3078 1560 -3072
rect 1554 -3084 1560 -3078
rect 1554 -3090 1560 -3084
rect 1554 -3096 1560 -3090
rect 1554 -3102 1560 -3096
rect 1554 -3108 1560 -3102
rect 1554 -3114 1560 -3108
rect 1554 -3120 1560 -3114
rect 1554 -3126 1560 -3120
rect 1554 -3132 1560 -3126
rect 1554 -3138 1560 -3132
rect 1554 -3144 1560 -3138
rect 1554 -3150 1560 -3144
rect 1554 -3156 1560 -3150
rect 1554 -3162 1560 -3156
rect 1554 -3168 1560 -3162
rect 1554 -3174 1560 -3168
rect 1554 -3180 1560 -3174
rect 1554 -3186 1560 -3180
rect 1554 -3192 1560 -3186
rect 1554 -3198 1560 -3192
rect 1554 -3204 1560 -3198
rect 1554 -3210 1560 -3204
rect 1554 -3216 1560 -3210
rect 1554 -3222 1560 -3216
rect 1554 -3228 1560 -3222
rect 1554 -3234 1560 -3228
rect 1554 -3276 1560 -3270
rect 1554 -3282 1560 -3276
rect 1554 -3288 1560 -3282
rect 1554 -3294 1560 -3288
rect 1554 -3300 1560 -3294
rect 1554 -3306 1560 -3300
rect 1554 -3312 1560 -3306
rect 1554 -3318 1560 -3312
rect 1554 -3324 1560 -3318
rect 1554 -3330 1560 -3324
rect 1554 -3336 1560 -3330
rect 1554 -3342 1560 -3336
rect 1554 -3348 1560 -3342
rect 1554 -3354 1560 -3348
rect 1554 -3360 1560 -3354
rect 1554 -3366 1560 -3360
rect 1554 -3372 1560 -3366
rect 1554 -3378 1560 -3372
rect 1554 -3384 1560 -3378
rect 1554 -3390 1560 -3384
rect 1554 -3396 1560 -3390
rect 1554 -3402 1560 -3396
rect 1554 -3408 1560 -3402
rect 1554 -3414 1560 -3408
rect 1554 -3420 1560 -3414
rect 1554 -3426 1560 -3420
rect 1554 -3432 1560 -3426
rect 1554 -3438 1560 -3432
rect 1554 -3444 1560 -3438
rect 1554 -3450 1560 -3444
rect 1554 -3456 1560 -3450
rect 1554 -3462 1560 -3456
rect 1554 -3468 1560 -3462
rect 1554 -3474 1560 -3468
rect 1560 -1080 1566 -1074
rect 1560 -1086 1566 -1080
rect 1560 -1092 1566 -1086
rect 1560 -1098 1566 -1092
rect 1560 -1104 1566 -1098
rect 1560 -1110 1566 -1104
rect 1560 -1116 1566 -1110
rect 1560 -1122 1566 -1116
rect 1560 -1128 1566 -1122
rect 1560 -1134 1566 -1128
rect 1560 -1140 1566 -1134
rect 1560 -1146 1566 -1140
rect 1560 -1152 1566 -1146
rect 1560 -1158 1566 -1152
rect 1560 -1164 1566 -1158
rect 1560 -1170 1566 -1164
rect 1560 -1176 1566 -1170
rect 1560 -1182 1566 -1176
rect 1560 -1188 1566 -1182
rect 1560 -1194 1566 -1188
rect 1560 -1200 1566 -1194
rect 1560 -1206 1566 -1200
rect 1560 -1212 1566 -1206
rect 1560 -1218 1566 -1212
rect 1560 -1224 1566 -1218
rect 1560 -1230 1566 -1224
rect 1560 -1236 1566 -1230
rect 1560 -1242 1566 -1236
rect 1560 -1248 1566 -1242
rect 1560 -1254 1566 -1248
rect 1560 -1260 1566 -1254
rect 1560 -1266 1566 -1260
rect 1560 -1272 1566 -1266
rect 1560 -1278 1566 -1272
rect 1560 -1284 1566 -1278
rect 1560 -1290 1566 -1284
rect 1560 -1296 1566 -1290
rect 1560 -1302 1566 -1296
rect 1560 -1308 1566 -1302
rect 1560 -1314 1566 -1308
rect 1560 -1320 1566 -1314
rect 1560 -1326 1566 -1320
rect 1560 -1332 1566 -1326
rect 1560 -1338 1566 -1332
rect 1560 -1344 1566 -1338
rect 1560 -1350 1566 -1344
rect 1560 -1356 1566 -1350
rect 1560 -1362 1566 -1356
rect 1560 -1368 1566 -1362
rect 1560 -1374 1566 -1368
rect 1560 -1380 1566 -1374
rect 1560 -1386 1566 -1380
rect 1560 -1392 1566 -1386
rect 1560 -1398 1566 -1392
rect 1560 -1404 1566 -1398
rect 1560 -1410 1566 -1404
rect 1560 -1416 1566 -1410
rect 1560 -1422 1566 -1416
rect 1560 -1428 1566 -1422
rect 1560 -1434 1566 -1428
rect 1560 -1440 1566 -1434
rect 1560 -1446 1566 -1440
rect 1560 -1452 1566 -1446
rect 1560 -1458 1566 -1452
rect 1560 -1464 1566 -1458
rect 1560 -1470 1566 -1464
rect 1560 -1476 1566 -1470
rect 1560 -1482 1566 -1476
rect 1560 -1488 1566 -1482
rect 1560 -1494 1566 -1488
rect 1560 -1500 1566 -1494
rect 1560 -1506 1566 -1500
rect 1560 -1512 1566 -1506
rect 1560 -1518 1566 -1512
rect 1560 -1524 1566 -1518
rect 1560 -1530 1566 -1524
rect 1560 -1536 1566 -1530
rect 1560 -1542 1566 -1536
rect 1560 -1548 1566 -1542
rect 1560 -1554 1566 -1548
rect 1560 -1560 1566 -1554
rect 1560 -1566 1566 -1560
rect 1560 -1572 1566 -1566
rect 1560 -1578 1566 -1572
rect 1560 -1584 1566 -1578
rect 1560 -1590 1566 -1584
rect 1560 -1596 1566 -1590
rect 1560 -1602 1566 -1596
rect 1560 -1608 1566 -1602
rect 1560 -1614 1566 -1608
rect 1560 -1620 1566 -1614
rect 1560 -1626 1566 -1620
rect 1560 -1632 1566 -1626
rect 1560 -1638 1566 -1632
rect 1560 -1644 1566 -1638
rect 1560 -1650 1566 -1644
rect 1560 -1656 1566 -1650
rect 1560 -1662 1566 -1656
rect 1560 -1668 1566 -1662
rect 1560 -1674 1566 -1668
rect 1560 -1680 1566 -1674
rect 1560 -1686 1566 -1680
rect 1560 -1692 1566 -1686
rect 1560 -1698 1566 -1692
rect 1560 -1704 1566 -1698
rect 1560 -1710 1566 -1704
rect 1560 -1716 1566 -1710
rect 1560 -1722 1566 -1716
rect 1560 -1728 1566 -1722
rect 1560 -1734 1566 -1728
rect 1560 -1740 1566 -1734
rect 1560 -1746 1566 -1740
rect 1560 -1752 1566 -1746
rect 1560 -1758 1566 -1752
rect 1560 -1764 1566 -1758
rect 1560 -1770 1566 -1764
rect 1560 -1776 1566 -1770
rect 1560 -1782 1566 -1776
rect 1560 -1788 1566 -1782
rect 1560 -1794 1566 -1788
rect 1560 -1800 1566 -1794
rect 1560 -1806 1566 -1800
rect 1560 -1812 1566 -1806
rect 1560 -1818 1566 -1812
rect 1560 -1824 1566 -1818
rect 1560 -1830 1566 -1824
rect 1560 -1836 1566 -1830
rect 1560 -1842 1566 -1836
rect 1560 -1848 1566 -1842
rect 1560 -1854 1566 -1848
rect 1560 -1860 1566 -1854
rect 1560 -1866 1566 -1860
rect 1560 -1872 1566 -1866
rect 1560 -1878 1566 -1872
rect 1560 -1884 1566 -1878
rect 1560 -1890 1566 -1884
rect 1560 -1896 1566 -1890
rect 1560 -1902 1566 -1896
rect 1560 -1908 1566 -1902
rect 1560 -1914 1566 -1908
rect 1560 -1920 1566 -1914
rect 1560 -1926 1566 -1920
rect 1560 -1932 1566 -1926
rect 1560 -1938 1566 -1932
rect 1560 -1944 1566 -1938
rect 1560 -1950 1566 -1944
rect 1560 -1956 1566 -1950
rect 1560 -1962 1566 -1956
rect 1560 -1968 1566 -1962
rect 1560 -1974 1566 -1968
rect 1560 -1980 1566 -1974
rect 1560 -1986 1566 -1980
rect 1560 -1992 1566 -1986
rect 1560 -1998 1566 -1992
rect 1560 -2004 1566 -1998
rect 1560 -2010 1566 -2004
rect 1560 -2016 1566 -2010
rect 1560 -2022 1566 -2016
rect 1560 -2028 1566 -2022
rect 1560 -2034 1566 -2028
rect 1560 -2040 1566 -2034
rect 1560 -2046 1566 -2040
rect 1560 -2052 1566 -2046
rect 1560 -2058 1566 -2052
rect 1560 -2064 1566 -2058
rect 1560 -2070 1566 -2064
rect 1560 -2076 1566 -2070
rect 1560 -2082 1566 -2076
rect 1560 -2088 1566 -2082
rect 1560 -2094 1566 -2088
rect 1560 -2100 1566 -2094
rect 1560 -2106 1566 -2100
rect 1560 -2112 1566 -2106
rect 1560 -2118 1566 -2112
rect 1560 -2190 1566 -2184
rect 1560 -2196 1566 -2190
rect 1560 -2202 1566 -2196
rect 1560 -2208 1566 -2202
rect 1560 -2214 1566 -2208
rect 1560 -2220 1566 -2214
rect 1560 -2226 1566 -2220
rect 1560 -2232 1566 -2226
rect 1560 -2238 1566 -2232
rect 1560 -2244 1566 -2238
rect 1560 -2250 1566 -2244
rect 1560 -2256 1566 -2250
rect 1560 -2262 1566 -2256
rect 1560 -2268 1566 -2262
rect 1560 -2274 1566 -2268
rect 1560 -2280 1566 -2274
rect 1560 -2286 1566 -2280
rect 1560 -2292 1566 -2286
rect 1560 -2298 1566 -2292
rect 1560 -2304 1566 -2298
rect 1560 -2310 1566 -2304
rect 1560 -2316 1566 -2310
rect 1560 -2322 1566 -2316
rect 1560 -2328 1566 -2322
rect 1560 -2334 1566 -2328
rect 1560 -2340 1566 -2334
rect 1560 -2346 1566 -2340
rect 1560 -2352 1566 -2346
rect 1560 -2358 1566 -2352
rect 1560 -2364 1566 -2358
rect 1560 -2370 1566 -2364
rect 1560 -2376 1566 -2370
rect 1560 -2382 1566 -2376
rect 1560 -2388 1566 -2382
rect 1560 -2394 1566 -2388
rect 1560 -2400 1566 -2394
rect 1560 -2406 1566 -2400
rect 1560 -2412 1566 -2406
rect 1560 -2418 1566 -2412
rect 1560 -2424 1566 -2418
rect 1560 -2430 1566 -2424
rect 1560 -2436 1566 -2430
rect 1560 -2442 1566 -2436
rect 1560 -2448 1566 -2442
rect 1560 -2454 1566 -2448
rect 1560 -2460 1566 -2454
rect 1560 -2466 1566 -2460
rect 1560 -2472 1566 -2466
rect 1560 -2478 1566 -2472
rect 1560 -2484 1566 -2478
rect 1560 -2490 1566 -2484
rect 1560 -2496 1566 -2490
rect 1560 -2502 1566 -2496
rect 1560 -2508 1566 -2502
rect 1560 -2514 1566 -2508
rect 1560 -2520 1566 -2514
rect 1560 -2526 1566 -2520
rect 1560 -2532 1566 -2526
rect 1560 -2538 1566 -2532
rect 1560 -2544 1566 -2538
rect 1560 -2550 1566 -2544
rect 1560 -2556 1566 -2550
rect 1560 -2562 1566 -2556
rect 1560 -2568 1566 -2562
rect 1560 -2574 1566 -2568
rect 1560 -2580 1566 -2574
rect 1560 -2586 1566 -2580
rect 1560 -2592 1566 -2586
rect 1560 -2598 1566 -2592
rect 1560 -2604 1566 -2598
rect 1560 -2610 1566 -2604
rect 1560 -2616 1566 -2610
rect 1560 -2622 1566 -2616
rect 1560 -2628 1566 -2622
rect 1560 -2634 1566 -2628
rect 1560 -2640 1566 -2634
rect 1560 -2646 1566 -2640
rect 1560 -2652 1566 -2646
rect 1560 -2658 1566 -2652
rect 1560 -2664 1566 -2658
rect 1560 -2670 1566 -2664
rect 1560 -2676 1566 -2670
rect 1560 -2682 1566 -2676
rect 1560 -2688 1566 -2682
rect 1560 -2694 1566 -2688
rect 1560 -2700 1566 -2694
rect 1560 -2706 1566 -2700
rect 1560 -2712 1566 -2706
rect 1560 -2718 1566 -2712
rect 1560 -2724 1566 -2718
rect 1560 -2730 1566 -2724
rect 1560 -2736 1566 -2730
rect 1560 -2742 1566 -2736
rect 1560 -2748 1566 -2742
rect 1560 -2754 1566 -2748
rect 1560 -2760 1566 -2754
rect 1560 -2766 1566 -2760
rect 1560 -2772 1566 -2766
rect 1560 -2856 1566 -2850
rect 1560 -2862 1566 -2856
rect 1560 -2868 1566 -2862
rect 1560 -2874 1566 -2868
rect 1560 -2880 1566 -2874
rect 1560 -2886 1566 -2880
rect 1560 -2892 1566 -2886
rect 1560 -2898 1566 -2892
rect 1560 -2904 1566 -2898
rect 1560 -2910 1566 -2904
rect 1560 -2916 1566 -2910
rect 1560 -2922 1566 -2916
rect 1560 -2928 1566 -2922
rect 1560 -2934 1566 -2928
rect 1560 -2940 1566 -2934
rect 1560 -2946 1566 -2940
rect 1560 -2952 1566 -2946
rect 1560 -2958 1566 -2952
rect 1560 -2964 1566 -2958
rect 1560 -2970 1566 -2964
rect 1560 -2976 1566 -2970
rect 1560 -2982 1566 -2976
rect 1560 -2988 1566 -2982
rect 1560 -2994 1566 -2988
rect 1560 -3000 1566 -2994
rect 1560 -3006 1566 -3000
rect 1560 -3012 1566 -3006
rect 1560 -3018 1566 -3012
rect 1560 -3024 1566 -3018
rect 1560 -3030 1566 -3024
rect 1560 -3036 1566 -3030
rect 1560 -3042 1566 -3036
rect 1560 -3048 1566 -3042
rect 1560 -3054 1566 -3048
rect 1560 -3060 1566 -3054
rect 1560 -3066 1566 -3060
rect 1560 -3072 1566 -3066
rect 1560 -3078 1566 -3072
rect 1560 -3084 1566 -3078
rect 1560 -3090 1566 -3084
rect 1560 -3096 1566 -3090
rect 1560 -3102 1566 -3096
rect 1560 -3108 1566 -3102
rect 1560 -3114 1566 -3108
rect 1560 -3120 1566 -3114
rect 1560 -3126 1566 -3120
rect 1560 -3132 1566 -3126
rect 1560 -3138 1566 -3132
rect 1560 -3144 1566 -3138
rect 1560 -3150 1566 -3144
rect 1560 -3156 1566 -3150
rect 1560 -3162 1566 -3156
rect 1560 -3168 1566 -3162
rect 1560 -3174 1566 -3168
rect 1560 -3180 1566 -3174
rect 1560 -3186 1566 -3180
rect 1560 -3192 1566 -3186
rect 1560 -3198 1566 -3192
rect 1560 -3204 1566 -3198
rect 1560 -3210 1566 -3204
rect 1560 -3216 1566 -3210
rect 1560 -3222 1566 -3216
rect 1560 -3228 1566 -3222
rect 1560 -3234 1566 -3228
rect 1560 -3276 1566 -3270
rect 1560 -3282 1566 -3276
rect 1560 -3288 1566 -3282
rect 1560 -3294 1566 -3288
rect 1560 -3300 1566 -3294
rect 1560 -3306 1566 -3300
rect 1560 -3312 1566 -3306
rect 1560 -3318 1566 -3312
rect 1560 -3324 1566 -3318
rect 1560 -3330 1566 -3324
rect 1560 -3336 1566 -3330
rect 1560 -3342 1566 -3336
rect 1560 -3348 1566 -3342
rect 1560 -3354 1566 -3348
rect 1560 -3360 1566 -3354
rect 1560 -3366 1566 -3360
rect 1560 -3372 1566 -3366
rect 1560 -3378 1566 -3372
rect 1560 -3384 1566 -3378
rect 1560 -3390 1566 -3384
rect 1560 -3396 1566 -3390
rect 1560 -3402 1566 -3396
rect 1560 -3408 1566 -3402
rect 1560 -3414 1566 -3408
rect 1560 -3420 1566 -3414
rect 1560 -3426 1566 -3420
rect 1560 -3432 1566 -3426
rect 1560 -3438 1566 -3432
rect 1560 -3444 1566 -3438
rect 1560 -3450 1566 -3444
rect 1560 -3456 1566 -3450
rect 1560 -3462 1566 -3456
rect 1560 -3468 1566 -3462
rect 1560 -3474 1566 -3468
rect 1566 -1068 1572 -1062
rect 1566 -1074 1572 -1068
rect 1566 -1080 1572 -1074
rect 1566 -1086 1572 -1080
rect 1566 -1092 1572 -1086
rect 1566 -1098 1572 -1092
rect 1566 -1104 1572 -1098
rect 1566 -1110 1572 -1104
rect 1566 -1116 1572 -1110
rect 1566 -1122 1572 -1116
rect 1566 -1128 1572 -1122
rect 1566 -1134 1572 -1128
rect 1566 -1140 1572 -1134
rect 1566 -1146 1572 -1140
rect 1566 -1152 1572 -1146
rect 1566 -1158 1572 -1152
rect 1566 -1164 1572 -1158
rect 1566 -1170 1572 -1164
rect 1566 -1176 1572 -1170
rect 1566 -1182 1572 -1176
rect 1566 -1188 1572 -1182
rect 1566 -1194 1572 -1188
rect 1566 -1200 1572 -1194
rect 1566 -1206 1572 -1200
rect 1566 -1212 1572 -1206
rect 1566 -1218 1572 -1212
rect 1566 -1224 1572 -1218
rect 1566 -1230 1572 -1224
rect 1566 -1236 1572 -1230
rect 1566 -1242 1572 -1236
rect 1566 -1248 1572 -1242
rect 1566 -1254 1572 -1248
rect 1566 -1260 1572 -1254
rect 1566 -1266 1572 -1260
rect 1566 -1272 1572 -1266
rect 1566 -1278 1572 -1272
rect 1566 -1284 1572 -1278
rect 1566 -1290 1572 -1284
rect 1566 -1296 1572 -1290
rect 1566 -1302 1572 -1296
rect 1566 -1308 1572 -1302
rect 1566 -1314 1572 -1308
rect 1566 -1320 1572 -1314
rect 1566 -1326 1572 -1320
rect 1566 -1332 1572 -1326
rect 1566 -1338 1572 -1332
rect 1566 -1344 1572 -1338
rect 1566 -1350 1572 -1344
rect 1566 -1356 1572 -1350
rect 1566 -1362 1572 -1356
rect 1566 -1368 1572 -1362
rect 1566 -1374 1572 -1368
rect 1566 -1380 1572 -1374
rect 1566 -1386 1572 -1380
rect 1566 -1392 1572 -1386
rect 1566 -1398 1572 -1392
rect 1566 -1404 1572 -1398
rect 1566 -1410 1572 -1404
rect 1566 -1416 1572 -1410
rect 1566 -1422 1572 -1416
rect 1566 -1428 1572 -1422
rect 1566 -1434 1572 -1428
rect 1566 -1440 1572 -1434
rect 1566 -1446 1572 -1440
rect 1566 -1452 1572 -1446
rect 1566 -1458 1572 -1452
rect 1566 -1464 1572 -1458
rect 1566 -1470 1572 -1464
rect 1566 -1476 1572 -1470
rect 1566 -1482 1572 -1476
rect 1566 -1488 1572 -1482
rect 1566 -1494 1572 -1488
rect 1566 -1500 1572 -1494
rect 1566 -1506 1572 -1500
rect 1566 -1512 1572 -1506
rect 1566 -1518 1572 -1512
rect 1566 -1524 1572 -1518
rect 1566 -1530 1572 -1524
rect 1566 -1536 1572 -1530
rect 1566 -1542 1572 -1536
rect 1566 -1548 1572 -1542
rect 1566 -1554 1572 -1548
rect 1566 -1560 1572 -1554
rect 1566 -1566 1572 -1560
rect 1566 -1572 1572 -1566
rect 1566 -1578 1572 -1572
rect 1566 -1584 1572 -1578
rect 1566 -1590 1572 -1584
rect 1566 -1596 1572 -1590
rect 1566 -1602 1572 -1596
rect 1566 -1608 1572 -1602
rect 1566 -1614 1572 -1608
rect 1566 -1620 1572 -1614
rect 1566 -1626 1572 -1620
rect 1566 -1632 1572 -1626
rect 1566 -1638 1572 -1632
rect 1566 -1644 1572 -1638
rect 1566 -1650 1572 -1644
rect 1566 -1656 1572 -1650
rect 1566 -1662 1572 -1656
rect 1566 -1668 1572 -1662
rect 1566 -1674 1572 -1668
rect 1566 -1680 1572 -1674
rect 1566 -1686 1572 -1680
rect 1566 -1692 1572 -1686
rect 1566 -1698 1572 -1692
rect 1566 -1704 1572 -1698
rect 1566 -1710 1572 -1704
rect 1566 -1716 1572 -1710
rect 1566 -1722 1572 -1716
rect 1566 -1728 1572 -1722
rect 1566 -1734 1572 -1728
rect 1566 -1740 1572 -1734
rect 1566 -1746 1572 -1740
rect 1566 -1752 1572 -1746
rect 1566 -1758 1572 -1752
rect 1566 -1764 1572 -1758
rect 1566 -1770 1572 -1764
rect 1566 -1776 1572 -1770
rect 1566 -1782 1572 -1776
rect 1566 -1788 1572 -1782
rect 1566 -1794 1572 -1788
rect 1566 -1800 1572 -1794
rect 1566 -1806 1572 -1800
rect 1566 -1812 1572 -1806
rect 1566 -1818 1572 -1812
rect 1566 -1824 1572 -1818
rect 1566 -1830 1572 -1824
rect 1566 -1836 1572 -1830
rect 1566 -1842 1572 -1836
rect 1566 -1848 1572 -1842
rect 1566 -1854 1572 -1848
rect 1566 -1860 1572 -1854
rect 1566 -1866 1572 -1860
rect 1566 -1872 1572 -1866
rect 1566 -1878 1572 -1872
rect 1566 -1884 1572 -1878
rect 1566 -1890 1572 -1884
rect 1566 -1896 1572 -1890
rect 1566 -1902 1572 -1896
rect 1566 -1908 1572 -1902
rect 1566 -1914 1572 -1908
rect 1566 -1920 1572 -1914
rect 1566 -1926 1572 -1920
rect 1566 -1932 1572 -1926
rect 1566 -1938 1572 -1932
rect 1566 -1944 1572 -1938
rect 1566 -1950 1572 -1944
rect 1566 -1956 1572 -1950
rect 1566 -1962 1572 -1956
rect 1566 -1968 1572 -1962
rect 1566 -1974 1572 -1968
rect 1566 -1980 1572 -1974
rect 1566 -1986 1572 -1980
rect 1566 -1992 1572 -1986
rect 1566 -1998 1572 -1992
rect 1566 -2004 1572 -1998
rect 1566 -2010 1572 -2004
rect 1566 -2016 1572 -2010
rect 1566 -2022 1572 -2016
rect 1566 -2028 1572 -2022
rect 1566 -2034 1572 -2028
rect 1566 -2040 1572 -2034
rect 1566 -2046 1572 -2040
rect 1566 -2052 1572 -2046
rect 1566 -2058 1572 -2052
rect 1566 -2064 1572 -2058
rect 1566 -2070 1572 -2064
rect 1566 -2076 1572 -2070
rect 1566 -2082 1572 -2076
rect 1566 -2088 1572 -2082
rect 1566 -2094 1572 -2088
rect 1566 -2100 1572 -2094
rect 1566 -2106 1572 -2100
rect 1566 -2184 1572 -2178
rect 1566 -2190 1572 -2184
rect 1566 -2196 1572 -2190
rect 1566 -2202 1572 -2196
rect 1566 -2208 1572 -2202
rect 1566 -2214 1572 -2208
rect 1566 -2220 1572 -2214
rect 1566 -2226 1572 -2220
rect 1566 -2232 1572 -2226
rect 1566 -2238 1572 -2232
rect 1566 -2244 1572 -2238
rect 1566 -2250 1572 -2244
rect 1566 -2256 1572 -2250
rect 1566 -2262 1572 -2256
rect 1566 -2268 1572 -2262
rect 1566 -2274 1572 -2268
rect 1566 -2280 1572 -2274
rect 1566 -2286 1572 -2280
rect 1566 -2292 1572 -2286
rect 1566 -2298 1572 -2292
rect 1566 -2304 1572 -2298
rect 1566 -2310 1572 -2304
rect 1566 -2316 1572 -2310
rect 1566 -2322 1572 -2316
rect 1566 -2328 1572 -2322
rect 1566 -2334 1572 -2328
rect 1566 -2340 1572 -2334
rect 1566 -2346 1572 -2340
rect 1566 -2352 1572 -2346
rect 1566 -2358 1572 -2352
rect 1566 -2364 1572 -2358
rect 1566 -2370 1572 -2364
rect 1566 -2376 1572 -2370
rect 1566 -2382 1572 -2376
rect 1566 -2388 1572 -2382
rect 1566 -2394 1572 -2388
rect 1566 -2400 1572 -2394
rect 1566 -2406 1572 -2400
rect 1566 -2412 1572 -2406
rect 1566 -2418 1572 -2412
rect 1566 -2424 1572 -2418
rect 1566 -2430 1572 -2424
rect 1566 -2436 1572 -2430
rect 1566 -2442 1572 -2436
rect 1566 -2448 1572 -2442
rect 1566 -2454 1572 -2448
rect 1566 -2460 1572 -2454
rect 1566 -2466 1572 -2460
rect 1566 -2472 1572 -2466
rect 1566 -2478 1572 -2472
rect 1566 -2484 1572 -2478
rect 1566 -2490 1572 -2484
rect 1566 -2496 1572 -2490
rect 1566 -2502 1572 -2496
rect 1566 -2508 1572 -2502
rect 1566 -2514 1572 -2508
rect 1566 -2520 1572 -2514
rect 1566 -2526 1572 -2520
rect 1566 -2532 1572 -2526
rect 1566 -2538 1572 -2532
rect 1566 -2544 1572 -2538
rect 1566 -2550 1572 -2544
rect 1566 -2556 1572 -2550
rect 1566 -2562 1572 -2556
rect 1566 -2568 1572 -2562
rect 1566 -2574 1572 -2568
rect 1566 -2580 1572 -2574
rect 1566 -2586 1572 -2580
rect 1566 -2592 1572 -2586
rect 1566 -2598 1572 -2592
rect 1566 -2604 1572 -2598
rect 1566 -2610 1572 -2604
rect 1566 -2616 1572 -2610
rect 1566 -2622 1572 -2616
rect 1566 -2628 1572 -2622
rect 1566 -2634 1572 -2628
rect 1566 -2640 1572 -2634
rect 1566 -2646 1572 -2640
rect 1566 -2652 1572 -2646
rect 1566 -2658 1572 -2652
rect 1566 -2664 1572 -2658
rect 1566 -2670 1572 -2664
rect 1566 -2676 1572 -2670
rect 1566 -2682 1572 -2676
rect 1566 -2688 1572 -2682
rect 1566 -2694 1572 -2688
rect 1566 -2700 1572 -2694
rect 1566 -2706 1572 -2700
rect 1566 -2712 1572 -2706
rect 1566 -2718 1572 -2712
rect 1566 -2724 1572 -2718
rect 1566 -2730 1572 -2724
rect 1566 -2736 1572 -2730
rect 1566 -2742 1572 -2736
rect 1566 -2748 1572 -2742
rect 1566 -2754 1572 -2748
rect 1566 -2760 1572 -2754
rect 1566 -2766 1572 -2760
rect 1566 -2850 1572 -2844
rect 1566 -2856 1572 -2850
rect 1566 -2862 1572 -2856
rect 1566 -2868 1572 -2862
rect 1566 -2874 1572 -2868
rect 1566 -2880 1572 -2874
rect 1566 -2886 1572 -2880
rect 1566 -2892 1572 -2886
rect 1566 -2898 1572 -2892
rect 1566 -2904 1572 -2898
rect 1566 -2910 1572 -2904
rect 1566 -2916 1572 -2910
rect 1566 -2922 1572 -2916
rect 1566 -2928 1572 -2922
rect 1566 -2934 1572 -2928
rect 1566 -2940 1572 -2934
rect 1566 -2946 1572 -2940
rect 1566 -2952 1572 -2946
rect 1566 -2958 1572 -2952
rect 1566 -2964 1572 -2958
rect 1566 -2970 1572 -2964
rect 1566 -2976 1572 -2970
rect 1566 -2982 1572 -2976
rect 1566 -2988 1572 -2982
rect 1566 -2994 1572 -2988
rect 1566 -3000 1572 -2994
rect 1566 -3006 1572 -3000
rect 1566 -3012 1572 -3006
rect 1566 -3018 1572 -3012
rect 1566 -3024 1572 -3018
rect 1566 -3030 1572 -3024
rect 1566 -3036 1572 -3030
rect 1566 -3042 1572 -3036
rect 1566 -3048 1572 -3042
rect 1566 -3054 1572 -3048
rect 1566 -3060 1572 -3054
rect 1566 -3066 1572 -3060
rect 1566 -3072 1572 -3066
rect 1566 -3078 1572 -3072
rect 1566 -3084 1572 -3078
rect 1566 -3090 1572 -3084
rect 1566 -3096 1572 -3090
rect 1566 -3102 1572 -3096
rect 1566 -3108 1572 -3102
rect 1566 -3114 1572 -3108
rect 1566 -3120 1572 -3114
rect 1566 -3126 1572 -3120
rect 1566 -3132 1572 -3126
rect 1566 -3138 1572 -3132
rect 1566 -3144 1572 -3138
rect 1566 -3150 1572 -3144
rect 1566 -3156 1572 -3150
rect 1566 -3162 1572 -3156
rect 1566 -3168 1572 -3162
rect 1566 -3174 1572 -3168
rect 1566 -3180 1572 -3174
rect 1566 -3186 1572 -3180
rect 1566 -3192 1572 -3186
rect 1566 -3198 1572 -3192
rect 1566 -3204 1572 -3198
rect 1566 -3210 1572 -3204
rect 1566 -3216 1572 -3210
rect 1566 -3222 1572 -3216
rect 1566 -3228 1572 -3222
rect 1566 -3234 1572 -3228
rect 1566 -3276 1572 -3270
rect 1566 -3282 1572 -3276
rect 1566 -3288 1572 -3282
rect 1566 -3294 1572 -3288
rect 1566 -3300 1572 -3294
rect 1566 -3306 1572 -3300
rect 1566 -3312 1572 -3306
rect 1566 -3318 1572 -3312
rect 1566 -3324 1572 -3318
rect 1566 -3330 1572 -3324
rect 1566 -3336 1572 -3330
rect 1566 -3342 1572 -3336
rect 1566 -3348 1572 -3342
rect 1566 -3354 1572 -3348
rect 1566 -3360 1572 -3354
rect 1566 -3366 1572 -3360
rect 1566 -3372 1572 -3366
rect 1566 -3378 1572 -3372
rect 1566 -3384 1572 -3378
rect 1566 -3390 1572 -3384
rect 1566 -3396 1572 -3390
rect 1566 -3402 1572 -3396
rect 1566 -3408 1572 -3402
rect 1566 -3414 1572 -3408
rect 1566 -3420 1572 -3414
rect 1566 -3426 1572 -3420
rect 1566 -3432 1572 -3426
rect 1566 -3438 1572 -3432
rect 1566 -3444 1572 -3438
rect 1566 -3450 1572 -3444
rect 1566 -3456 1572 -3450
rect 1566 -3462 1572 -3456
rect 1566 -3468 1572 -3462
rect 1572 -1062 1578 -1056
rect 1572 -1068 1578 -1062
rect 1572 -1074 1578 -1068
rect 1572 -1080 1578 -1074
rect 1572 -1086 1578 -1080
rect 1572 -1092 1578 -1086
rect 1572 -1098 1578 -1092
rect 1572 -1104 1578 -1098
rect 1572 -1110 1578 -1104
rect 1572 -1116 1578 -1110
rect 1572 -1122 1578 -1116
rect 1572 -1128 1578 -1122
rect 1572 -1134 1578 -1128
rect 1572 -1140 1578 -1134
rect 1572 -1146 1578 -1140
rect 1572 -1152 1578 -1146
rect 1572 -1158 1578 -1152
rect 1572 -1164 1578 -1158
rect 1572 -1170 1578 -1164
rect 1572 -1176 1578 -1170
rect 1572 -1182 1578 -1176
rect 1572 -1188 1578 -1182
rect 1572 -1194 1578 -1188
rect 1572 -1200 1578 -1194
rect 1572 -1206 1578 -1200
rect 1572 -1212 1578 -1206
rect 1572 -1218 1578 -1212
rect 1572 -1224 1578 -1218
rect 1572 -1230 1578 -1224
rect 1572 -1236 1578 -1230
rect 1572 -1242 1578 -1236
rect 1572 -1248 1578 -1242
rect 1572 -1254 1578 -1248
rect 1572 -1260 1578 -1254
rect 1572 -1266 1578 -1260
rect 1572 -1272 1578 -1266
rect 1572 -1278 1578 -1272
rect 1572 -1284 1578 -1278
rect 1572 -1290 1578 -1284
rect 1572 -1296 1578 -1290
rect 1572 -1302 1578 -1296
rect 1572 -1308 1578 -1302
rect 1572 -1314 1578 -1308
rect 1572 -1320 1578 -1314
rect 1572 -1326 1578 -1320
rect 1572 -1332 1578 -1326
rect 1572 -1338 1578 -1332
rect 1572 -1344 1578 -1338
rect 1572 -1350 1578 -1344
rect 1572 -1356 1578 -1350
rect 1572 -1362 1578 -1356
rect 1572 -1368 1578 -1362
rect 1572 -1374 1578 -1368
rect 1572 -1380 1578 -1374
rect 1572 -1386 1578 -1380
rect 1572 -1392 1578 -1386
rect 1572 -1398 1578 -1392
rect 1572 -1404 1578 -1398
rect 1572 -1410 1578 -1404
rect 1572 -1416 1578 -1410
rect 1572 -1422 1578 -1416
rect 1572 -1428 1578 -1422
rect 1572 -1434 1578 -1428
rect 1572 -1440 1578 -1434
rect 1572 -1446 1578 -1440
rect 1572 -1452 1578 -1446
rect 1572 -1458 1578 -1452
rect 1572 -1464 1578 -1458
rect 1572 -1470 1578 -1464
rect 1572 -1476 1578 -1470
rect 1572 -1482 1578 -1476
rect 1572 -1488 1578 -1482
rect 1572 -1494 1578 -1488
rect 1572 -1500 1578 -1494
rect 1572 -1506 1578 -1500
rect 1572 -1512 1578 -1506
rect 1572 -1518 1578 -1512
rect 1572 -1524 1578 -1518
rect 1572 -1530 1578 -1524
rect 1572 -1536 1578 -1530
rect 1572 -1542 1578 -1536
rect 1572 -1548 1578 -1542
rect 1572 -1554 1578 -1548
rect 1572 -1560 1578 -1554
rect 1572 -1566 1578 -1560
rect 1572 -1572 1578 -1566
rect 1572 -1578 1578 -1572
rect 1572 -1584 1578 -1578
rect 1572 -1590 1578 -1584
rect 1572 -1596 1578 -1590
rect 1572 -1602 1578 -1596
rect 1572 -1608 1578 -1602
rect 1572 -1614 1578 -1608
rect 1572 -1620 1578 -1614
rect 1572 -1626 1578 -1620
rect 1572 -1632 1578 -1626
rect 1572 -1638 1578 -1632
rect 1572 -1644 1578 -1638
rect 1572 -1650 1578 -1644
rect 1572 -1656 1578 -1650
rect 1572 -1662 1578 -1656
rect 1572 -1668 1578 -1662
rect 1572 -1674 1578 -1668
rect 1572 -1680 1578 -1674
rect 1572 -1686 1578 -1680
rect 1572 -1692 1578 -1686
rect 1572 -1698 1578 -1692
rect 1572 -1704 1578 -1698
rect 1572 -1710 1578 -1704
rect 1572 -1716 1578 -1710
rect 1572 -1722 1578 -1716
rect 1572 -1728 1578 -1722
rect 1572 -1734 1578 -1728
rect 1572 -1740 1578 -1734
rect 1572 -1746 1578 -1740
rect 1572 -1752 1578 -1746
rect 1572 -1758 1578 -1752
rect 1572 -1764 1578 -1758
rect 1572 -1770 1578 -1764
rect 1572 -1776 1578 -1770
rect 1572 -1782 1578 -1776
rect 1572 -1788 1578 -1782
rect 1572 -1794 1578 -1788
rect 1572 -1800 1578 -1794
rect 1572 -1806 1578 -1800
rect 1572 -1812 1578 -1806
rect 1572 -1818 1578 -1812
rect 1572 -1824 1578 -1818
rect 1572 -1830 1578 -1824
rect 1572 -1836 1578 -1830
rect 1572 -1842 1578 -1836
rect 1572 -1848 1578 -1842
rect 1572 -1854 1578 -1848
rect 1572 -1860 1578 -1854
rect 1572 -1866 1578 -1860
rect 1572 -1872 1578 -1866
rect 1572 -1878 1578 -1872
rect 1572 -1884 1578 -1878
rect 1572 -1890 1578 -1884
rect 1572 -1896 1578 -1890
rect 1572 -1902 1578 -1896
rect 1572 -1908 1578 -1902
rect 1572 -1914 1578 -1908
rect 1572 -1920 1578 -1914
rect 1572 -1926 1578 -1920
rect 1572 -1932 1578 -1926
rect 1572 -1938 1578 -1932
rect 1572 -1944 1578 -1938
rect 1572 -1950 1578 -1944
rect 1572 -1956 1578 -1950
rect 1572 -1962 1578 -1956
rect 1572 -1968 1578 -1962
rect 1572 -1974 1578 -1968
rect 1572 -1980 1578 -1974
rect 1572 -1986 1578 -1980
rect 1572 -1992 1578 -1986
rect 1572 -1998 1578 -1992
rect 1572 -2004 1578 -1998
rect 1572 -2010 1578 -2004
rect 1572 -2016 1578 -2010
rect 1572 -2022 1578 -2016
rect 1572 -2028 1578 -2022
rect 1572 -2034 1578 -2028
rect 1572 -2040 1578 -2034
rect 1572 -2046 1578 -2040
rect 1572 -2052 1578 -2046
rect 1572 -2058 1578 -2052
rect 1572 -2064 1578 -2058
rect 1572 -2070 1578 -2064
rect 1572 -2076 1578 -2070
rect 1572 -2082 1578 -2076
rect 1572 -2088 1578 -2082
rect 1572 -2094 1578 -2088
rect 1572 -2100 1578 -2094
rect 1572 -2172 1578 -2166
rect 1572 -2178 1578 -2172
rect 1572 -2184 1578 -2178
rect 1572 -2190 1578 -2184
rect 1572 -2196 1578 -2190
rect 1572 -2202 1578 -2196
rect 1572 -2208 1578 -2202
rect 1572 -2214 1578 -2208
rect 1572 -2220 1578 -2214
rect 1572 -2226 1578 -2220
rect 1572 -2232 1578 -2226
rect 1572 -2238 1578 -2232
rect 1572 -2244 1578 -2238
rect 1572 -2250 1578 -2244
rect 1572 -2256 1578 -2250
rect 1572 -2262 1578 -2256
rect 1572 -2268 1578 -2262
rect 1572 -2274 1578 -2268
rect 1572 -2280 1578 -2274
rect 1572 -2286 1578 -2280
rect 1572 -2292 1578 -2286
rect 1572 -2298 1578 -2292
rect 1572 -2304 1578 -2298
rect 1572 -2310 1578 -2304
rect 1572 -2316 1578 -2310
rect 1572 -2322 1578 -2316
rect 1572 -2328 1578 -2322
rect 1572 -2334 1578 -2328
rect 1572 -2340 1578 -2334
rect 1572 -2346 1578 -2340
rect 1572 -2352 1578 -2346
rect 1572 -2358 1578 -2352
rect 1572 -2364 1578 -2358
rect 1572 -2370 1578 -2364
rect 1572 -2376 1578 -2370
rect 1572 -2382 1578 -2376
rect 1572 -2388 1578 -2382
rect 1572 -2394 1578 -2388
rect 1572 -2400 1578 -2394
rect 1572 -2406 1578 -2400
rect 1572 -2412 1578 -2406
rect 1572 -2418 1578 -2412
rect 1572 -2424 1578 -2418
rect 1572 -2430 1578 -2424
rect 1572 -2436 1578 -2430
rect 1572 -2442 1578 -2436
rect 1572 -2448 1578 -2442
rect 1572 -2454 1578 -2448
rect 1572 -2460 1578 -2454
rect 1572 -2466 1578 -2460
rect 1572 -2472 1578 -2466
rect 1572 -2478 1578 -2472
rect 1572 -2484 1578 -2478
rect 1572 -2490 1578 -2484
rect 1572 -2496 1578 -2490
rect 1572 -2502 1578 -2496
rect 1572 -2508 1578 -2502
rect 1572 -2514 1578 -2508
rect 1572 -2520 1578 -2514
rect 1572 -2526 1578 -2520
rect 1572 -2532 1578 -2526
rect 1572 -2538 1578 -2532
rect 1572 -2544 1578 -2538
rect 1572 -2550 1578 -2544
rect 1572 -2556 1578 -2550
rect 1572 -2562 1578 -2556
rect 1572 -2568 1578 -2562
rect 1572 -2574 1578 -2568
rect 1572 -2580 1578 -2574
rect 1572 -2586 1578 -2580
rect 1572 -2592 1578 -2586
rect 1572 -2598 1578 -2592
rect 1572 -2604 1578 -2598
rect 1572 -2610 1578 -2604
rect 1572 -2616 1578 -2610
rect 1572 -2622 1578 -2616
rect 1572 -2628 1578 -2622
rect 1572 -2634 1578 -2628
rect 1572 -2640 1578 -2634
rect 1572 -2646 1578 -2640
rect 1572 -2652 1578 -2646
rect 1572 -2658 1578 -2652
rect 1572 -2664 1578 -2658
rect 1572 -2670 1578 -2664
rect 1572 -2676 1578 -2670
rect 1572 -2682 1578 -2676
rect 1572 -2688 1578 -2682
rect 1572 -2694 1578 -2688
rect 1572 -2700 1578 -2694
rect 1572 -2706 1578 -2700
rect 1572 -2712 1578 -2706
rect 1572 -2718 1578 -2712
rect 1572 -2724 1578 -2718
rect 1572 -2730 1578 -2724
rect 1572 -2736 1578 -2730
rect 1572 -2742 1578 -2736
rect 1572 -2748 1578 -2742
rect 1572 -2754 1578 -2748
rect 1572 -2760 1578 -2754
rect 1572 -2766 1578 -2760
rect 1572 -2844 1578 -2838
rect 1572 -2850 1578 -2844
rect 1572 -2856 1578 -2850
rect 1572 -2862 1578 -2856
rect 1572 -2868 1578 -2862
rect 1572 -2874 1578 -2868
rect 1572 -2880 1578 -2874
rect 1572 -2886 1578 -2880
rect 1572 -2892 1578 -2886
rect 1572 -2898 1578 -2892
rect 1572 -2904 1578 -2898
rect 1572 -2910 1578 -2904
rect 1572 -2916 1578 -2910
rect 1572 -2922 1578 -2916
rect 1572 -2928 1578 -2922
rect 1572 -2934 1578 -2928
rect 1572 -2940 1578 -2934
rect 1572 -2946 1578 -2940
rect 1572 -2952 1578 -2946
rect 1572 -2958 1578 -2952
rect 1572 -2964 1578 -2958
rect 1572 -2970 1578 -2964
rect 1572 -2976 1578 -2970
rect 1572 -2982 1578 -2976
rect 1572 -2988 1578 -2982
rect 1572 -2994 1578 -2988
rect 1572 -3000 1578 -2994
rect 1572 -3006 1578 -3000
rect 1572 -3012 1578 -3006
rect 1572 -3018 1578 -3012
rect 1572 -3024 1578 -3018
rect 1572 -3030 1578 -3024
rect 1572 -3036 1578 -3030
rect 1572 -3042 1578 -3036
rect 1572 -3048 1578 -3042
rect 1572 -3054 1578 -3048
rect 1572 -3060 1578 -3054
rect 1572 -3066 1578 -3060
rect 1572 -3072 1578 -3066
rect 1572 -3078 1578 -3072
rect 1572 -3084 1578 -3078
rect 1572 -3090 1578 -3084
rect 1572 -3096 1578 -3090
rect 1572 -3102 1578 -3096
rect 1572 -3108 1578 -3102
rect 1572 -3114 1578 -3108
rect 1572 -3120 1578 -3114
rect 1572 -3126 1578 -3120
rect 1572 -3132 1578 -3126
rect 1572 -3138 1578 -3132
rect 1572 -3144 1578 -3138
rect 1572 -3150 1578 -3144
rect 1572 -3156 1578 -3150
rect 1572 -3162 1578 -3156
rect 1572 -3168 1578 -3162
rect 1572 -3174 1578 -3168
rect 1572 -3180 1578 -3174
rect 1572 -3186 1578 -3180
rect 1572 -3192 1578 -3186
rect 1572 -3198 1578 -3192
rect 1572 -3204 1578 -3198
rect 1572 -3210 1578 -3204
rect 1572 -3216 1578 -3210
rect 1572 -3222 1578 -3216
rect 1572 -3228 1578 -3222
rect 1572 -3234 1578 -3228
rect 1572 -3276 1578 -3270
rect 1572 -3282 1578 -3276
rect 1572 -3288 1578 -3282
rect 1572 -3294 1578 -3288
rect 1572 -3300 1578 -3294
rect 1572 -3306 1578 -3300
rect 1572 -3312 1578 -3306
rect 1572 -3318 1578 -3312
rect 1572 -3324 1578 -3318
rect 1572 -3330 1578 -3324
rect 1572 -3336 1578 -3330
rect 1572 -3342 1578 -3336
rect 1572 -3348 1578 -3342
rect 1572 -3354 1578 -3348
rect 1572 -3360 1578 -3354
rect 1572 -3366 1578 -3360
rect 1572 -3372 1578 -3366
rect 1572 -3378 1578 -3372
rect 1572 -3384 1578 -3378
rect 1572 -3390 1578 -3384
rect 1572 -3396 1578 -3390
rect 1572 -3402 1578 -3396
rect 1572 -3408 1578 -3402
rect 1572 -3414 1578 -3408
rect 1572 -3420 1578 -3414
rect 1572 -3426 1578 -3420
rect 1572 -3432 1578 -3426
rect 1572 -3438 1578 -3432
rect 1572 -3444 1578 -3438
rect 1572 -3450 1578 -3444
rect 1572 -3456 1578 -3450
rect 1572 -3462 1578 -3456
rect 1572 -3468 1578 -3462
rect 1578 -1050 1584 -1044
rect 1578 -1056 1584 -1050
rect 1578 -1062 1584 -1056
rect 1578 -1068 1584 -1062
rect 1578 -1074 1584 -1068
rect 1578 -1080 1584 -1074
rect 1578 -1086 1584 -1080
rect 1578 -1092 1584 -1086
rect 1578 -1098 1584 -1092
rect 1578 -1104 1584 -1098
rect 1578 -1110 1584 -1104
rect 1578 -1116 1584 -1110
rect 1578 -1122 1584 -1116
rect 1578 -1128 1584 -1122
rect 1578 -1134 1584 -1128
rect 1578 -1140 1584 -1134
rect 1578 -1146 1584 -1140
rect 1578 -1152 1584 -1146
rect 1578 -1158 1584 -1152
rect 1578 -1164 1584 -1158
rect 1578 -1170 1584 -1164
rect 1578 -1176 1584 -1170
rect 1578 -1182 1584 -1176
rect 1578 -1188 1584 -1182
rect 1578 -1194 1584 -1188
rect 1578 -1200 1584 -1194
rect 1578 -1206 1584 -1200
rect 1578 -1212 1584 -1206
rect 1578 -1218 1584 -1212
rect 1578 -1224 1584 -1218
rect 1578 -1230 1584 -1224
rect 1578 -1236 1584 -1230
rect 1578 -1242 1584 -1236
rect 1578 -1248 1584 -1242
rect 1578 -1254 1584 -1248
rect 1578 -1260 1584 -1254
rect 1578 -1266 1584 -1260
rect 1578 -1272 1584 -1266
rect 1578 -1278 1584 -1272
rect 1578 -1284 1584 -1278
rect 1578 -1290 1584 -1284
rect 1578 -1296 1584 -1290
rect 1578 -1302 1584 -1296
rect 1578 -1308 1584 -1302
rect 1578 -1314 1584 -1308
rect 1578 -1320 1584 -1314
rect 1578 -1326 1584 -1320
rect 1578 -1332 1584 -1326
rect 1578 -1338 1584 -1332
rect 1578 -1344 1584 -1338
rect 1578 -1350 1584 -1344
rect 1578 -1356 1584 -1350
rect 1578 -1362 1584 -1356
rect 1578 -1368 1584 -1362
rect 1578 -1374 1584 -1368
rect 1578 -1380 1584 -1374
rect 1578 -1386 1584 -1380
rect 1578 -1392 1584 -1386
rect 1578 -1398 1584 -1392
rect 1578 -1404 1584 -1398
rect 1578 -1410 1584 -1404
rect 1578 -1416 1584 -1410
rect 1578 -1422 1584 -1416
rect 1578 -1428 1584 -1422
rect 1578 -1434 1584 -1428
rect 1578 -1440 1584 -1434
rect 1578 -1446 1584 -1440
rect 1578 -1452 1584 -1446
rect 1578 -1458 1584 -1452
rect 1578 -1464 1584 -1458
rect 1578 -1470 1584 -1464
rect 1578 -1476 1584 -1470
rect 1578 -1482 1584 -1476
rect 1578 -1488 1584 -1482
rect 1578 -1494 1584 -1488
rect 1578 -1500 1584 -1494
rect 1578 -1506 1584 -1500
rect 1578 -1512 1584 -1506
rect 1578 -1518 1584 -1512
rect 1578 -1524 1584 -1518
rect 1578 -1530 1584 -1524
rect 1578 -1536 1584 -1530
rect 1578 -1542 1584 -1536
rect 1578 -1548 1584 -1542
rect 1578 -1554 1584 -1548
rect 1578 -1560 1584 -1554
rect 1578 -1566 1584 -1560
rect 1578 -1572 1584 -1566
rect 1578 -1578 1584 -1572
rect 1578 -1584 1584 -1578
rect 1578 -1590 1584 -1584
rect 1578 -1596 1584 -1590
rect 1578 -1602 1584 -1596
rect 1578 -1608 1584 -1602
rect 1578 -1614 1584 -1608
rect 1578 -1620 1584 -1614
rect 1578 -1626 1584 -1620
rect 1578 -1632 1584 -1626
rect 1578 -1638 1584 -1632
rect 1578 -1644 1584 -1638
rect 1578 -1650 1584 -1644
rect 1578 -1656 1584 -1650
rect 1578 -1662 1584 -1656
rect 1578 -1668 1584 -1662
rect 1578 -1674 1584 -1668
rect 1578 -1680 1584 -1674
rect 1578 -1686 1584 -1680
rect 1578 -1692 1584 -1686
rect 1578 -1698 1584 -1692
rect 1578 -1704 1584 -1698
rect 1578 -1710 1584 -1704
rect 1578 -1716 1584 -1710
rect 1578 -1722 1584 -1716
rect 1578 -1728 1584 -1722
rect 1578 -1734 1584 -1728
rect 1578 -1740 1584 -1734
rect 1578 -1746 1584 -1740
rect 1578 -1752 1584 -1746
rect 1578 -1758 1584 -1752
rect 1578 -1764 1584 -1758
rect 1578 -1770 1584 -1764
rect 1578 -1776 1584 -1770
rect 1578 -1782 1584 -1776
rect 1578 -1788 1584 -1782
rect 1578 -1794 1584 -1788
rect 1578 -1800 1584 -1794
rect 1578 -1806 1584 -1800
rect 1578 -1812 1584 -1806
rect 1578 -1818 1584 -1812
rect 1578 -1824 1584 -1818
rect 1578 -1830 1584 -1824
rect 1578 -1836 1584 -1830
rect 1578 -1842 1584 -1836
rect 1578 -1848 1584 -1842
rect 1578 -1854 1584 -1848
rect 1578 -1860 1584 -1854
rect 1578 -1866 1584 -1860
rect 1578 -1872 1584 -1866
rect 1578 -1878 1584 -1872
rect 1578 -1884 1584 -1878
rect 1578 -1890 1584 -1884
rect 1578 -1896 1584 -1890
rect 1578 -1902 1584 -1896
rect 1578 -1908 1584 -1902
rect 1578 -1914 1584 -1908
rect 1578 -1920 1584 -1914
rect 1578 -1926 1584 -1920
rect 1578 -1932 1584 -1926
rect 1578 -1938 1584 -1932
rect 1578 -1944 1584 -1938
rect 1578 -1950 1584 -1944
rect 1578 -1956 1584 -1950
rect 1578 -1962 1584 -1956
rect 1578 -1968 1584 -1962
rect 1578 -1974 1584 -1968
rect 1578 -1980 1584 -1974
rect 1578 -1986 1584 -1980
rect 1578 -1992 1584 -1986
rect 1578 -1998 1584 -1992
rect 1578 -2004 1584 -1998
rect 1578 -2010 1584 -2004
rect 1578 -2016 1584 -2010
rect 1578 -2022 1584 -2016
rect 1578 -2028 1584 -2022
rect 1578 -2034 1584 -2028
rect 1578 -2040 1584 -2034
rect 1578 -2046 1584 -2040
rect 1578 -2052 1584 -2046
rect 1578 -2058 1584 -2052
rect 1578 -2064 1584 -2058
rect 1578 -2070 1584 -2064
rect 1578 -2076 1584 -2070
rect 1578 -2082 1584 -2076
rect 1578 -2088 1584 -2082
rect 1578 -2094 1584 -2088
rect 1578 -2166 1584 -2160
rect 1578 -2172 1584 -2166
rect 1578 -2178 1584 -2172
rect 1578 -2184 1584 -2178
rect 1578 -2190 1584 -2184
rect 1578 -2196 1584 -2190
rect 1578 -2202 1584 -2196
rect 1578 -2208 1584 -2202
rect 1578 -2214 1584 -2208
rect 1578 -2220 1584 -2214
rect 1578 -2226 1584 -2220
rect 1578 -2232 1584 -2226
rect 1578 -2238 1584 -2232
rect 1578 -2244 1584 -2238
rect 1578 -2250 1584 -2244
rect 1578 -2256 1584 -2250
rect 1578 -2262 1584 -2256
rect 1578 -2268 1584 -2262
rect 1578 -2274 1584 -2268
rect 1578 -2280 1584 -2274
rect 1578 -2286 1584 -2280
rect 1578 -2292 1584 -2286
rect 1578 -2298 1584 -2292
rect 1578 -2304 1584 -2298
rect 1578 -2310 1584 -2304
rect 1578 -2316 1584 -2310
rect 1578 -2322 1584 -2316
rect 1578 -2328 1584 -2322
rect 1578 -2334 1584 -2328
rect 1578 -2340 1584 -2334
rect 1578 -2346 1584 -2340
rect 1578 -2352 1584 -2346
rect 1578 -2358 1584 -2352
rect 1578 -2364 1584 -2358
rect 1578 -2370 1584 -2364
rect 1578 -2376 1584 -2370
rect 1578 -2382 1584 -2376
rect 1578 -2388 1584 -2382
rect 1578 -2394 1584 -2388
rect 1578 -2400 1584 -2394
rect 1578 -2406 1584 -2400
rect 1578 -2412 1584 -2406
rect 1578 -2418 1584 -2412
rect 1578 -2424 1584 -2418
rect 1578 -2430 1584 -2424
rect 1578 -2436 1584 -2430
rect 1578 -2442 1584 -2436
rect 1578 -2448 1584 -2442
rect 1578 -2454 1584 -2448
rect 1578 -2460 1584 -2454
rect 1578 -2466 1584 -2460
rect 1578 -2472 1584 -2466
rect 1578 -2478 1584 -2472
rect 1578 -2484 1584 -2478
rect 1578 -2490 1584 -2484
rect 1578 -2496 1584 -2490
rect 1578 -2502 1584 -2496
rect 1578 -2508 1584 -2502
rect 1578 -2514 1584 -2508
rect 1578 -2520 1584 -2514
rect 1578 -2526 1584 -2520
rect 1578 -2532 1584 -2526
rect 1578 -2538 1584 -2532
rect 1578 -2544 1584 -2538
rect 1578 -2550 1584 -2544
rect 1578 -2556 1584 -2550
rect 1578 -2562 1584 -2556
rect 1578 -2568 1584 -2562
rect 1578 -2574 1584 -2568
rect 1578 -2580 1584 -2574
rect 1578 -2586 1584 -2580
rect 1578 -2592 1584 -2586
rect 1578 -2598 1584 -2592
rect 1578 -2604 1584 -2598
rect 1578 -2610 1584 -2604
rect 1578 -2616 1584 -2610
rect 1578 -2622 1584 -2616
rect 1578 -2628 1584 -2622
rect 1578 -2634 1584 -2628
rect 1578 -2640 1584 -2634
rect 1578 -2646 1584 -2640
rect 1578 -2652 1584 -2646
rect 1578 -2658 1584 -2652
rect 1578 -2664 1584 -2658
rect 1578 -2670 1584 -2664
rect 1578 -2676 1584 -2670
rect 1578 -2682 1584 -2676
rect 1578 -2688 1584 -2682
rect 1578 -2694 1584 -2688
rect 1578 -2700 1584 -2694
rect 1578 -2706 1584 -2700
rect 1578 -2712 1584 -2706
rect 1578 -2718 1584 -2712
rect 1578 -2724 1584 -2718
rect 1578 -2730 1584 -2724
rect 1578 -2736 1584 -2730
rect 1578 -2742 1584 -2736
rect 1578 -2748 1584 -2742
rect 1578 -2754 1584 -2748
rect 1578 -2760 1584 -2754
rect 1578 -2844 1584 -2838
rect 1578 -2850 1584 -2844
rect 1578 -2856 1584 -2850
rect 1578 -2862 1584 -2856
rect 1578 -2868 1584 -2862
rect 1578 -2874 1584 -2868
rect 1578 -2880 1584 -2874
rect 1578 -2886 1584 -2880
rect 1578 -2892 1584 -2886
rect 1578 -2898 1584 -2892
rect 1578 -2904 1584 -2898
rect 1578 -2910 1584 -2904
rect 1578 -2916 1584 -2910
rect 1578 -2922 1584 -2916
rect 1578 -2928 1584 -2922
rect 1578 -2934 1584 -2928
rect 1578 -2940 1584 -2934
rect 1578 -2946 1584 -2940
rect 1578 -2952 1584 -2946
rect 1578 -2958 1584 -2952
rect 1578 -2964 1584 -2958
rect 1578 -2970 1584 -2964
rect 1578 -2976 1584 -2970
rect 1578 -2982 1584 -2976
rect 1578 -2988 1584 -2982
rect 1578 -2994 1584 -2988
rect 1578 -3000 1584 -2994
rect 1578 -3006 1584 -3000
rect 1578 -3012 1584 -3006
rect 1578 -3018 1584 -3012
rect 1578 -3024 1584 -3018
rect 1578 -3030 1584 -3024
rect 1578 -3036 1584 -3030
rect 1578 -3042 1584 -3036
rect 1578 -3048 1584 -3042
rect 1578 -3054 1584 -3048
rect 1578 -3060 1584 -3054
rect 1578 -3066 1584 -3060
rect 1578 -3072 1584 -3066
rect 1578 -3078 1584 -3072
rect 1578 -3084 1584 -3078
rect 1578 -3090 1584 -3084
rect 1578 -3096 1584 -3090
rect 1578 -3102 1584 -3096
rect 1578 -3108 1584 -3102
rect 1578 -3114 1584 -3108
rect 1578 -3120 1584 -3114
rect 1578 -3126 1584 -3120
rect 1578 -3132 1584 -3126
rect 1578 -3138 1584 -3132
rect 1578 -3144 1584 -3138
rect 1578 -3150 1584 -3144
rect 1578 -3156 1584 -3150
rect 1578 -3162 1584 -3156
rect 1578 -3168 1584 -3162
rect 1578 -3174 1584 -3168
rect 1578 -3180 1584 -3174
rect 1578 -3186 1584 -3180
rect 1578 -3192 1584 -3186
rect 1578 -3198 1584 -3192
rect 1578 -3204 1584 -3198
rect 1578 -3210 1584 -3204
rect 1578 -3216 1584 -3210
rect 1578 -3222 1584 -3216
rect 1578 -3228 1584 -3222
rect 1578 -3234 1584 -3228
rect 1578 -3276 1584 -3270
rect 1578 -3282 1584 -3276
rect 1578 -3288 1584 -3282
rect 1578 -3294 1584 -3288
rect 1578 -3300 1584 -3294
rect 1578 -3306 1584 -3300
rect 1578 -3312 1584 -3306
rect 1578 -3318 1584 -3312
rect 1578 -3324 1584 -3318
rect 1578 -3330 1584 -3324
rect 1578 -3336 1584 -3330
rect 1578 -3342 1584 -3336
rect 1578 -3348 1584 -3342
rect 1578 -3354 1584 -3348
rect 1578 -3360 1584 -3354
rect 1578 -3366 1584 -3360
rect 1578 -3372 1584 -3366
rect 1578 -3378 1584 -3372
rect 1578 -3384 1584 -3378
rect 1578 -3390 1584 -3384
rect 1578 -3396 1584 -3390
rect 1578 -3402 1584 -3396
rect 1578 -3408 1584 -3402
rect 1578 -3414 1584 -3408
rect 1578 -3420 1584 -3414
rect 1578 -3426 1584 -3420
rect 1578 -3432 1584 -3426
rect 1578 -3438 1584 -3432
rect 1578 -3444 1584 -3438
rect 1578 -3450 1584 -3444
rect 1578 -3456 1584 -3450
rect 1578 -3462 1584 -3456
rect 1578 -3468 1584 -3462
rect 1584 -1044 1590 -1038
rect 1584 -1050 1590 -1044
rect 1584 -1056 1590 -1050
rect 1584 -1062 1590 -1056
rect 1584 -1068 1590 -1062
rect 1584 -1074 1590 -1068
rect 1584 -1080 1590 -1074
rect 1584 -1086 1590 -1080
rect 1584 -1092 1590 -1086
rect 1584 -1098 1590 -1092
rect 1584 -1104 1590 -1098
rect 1584 -1110 1590 -1104
rect 1584 -1116 1590 -1110
rect 1584 -1122 1590 -1116
rect 1584 -1128 1590 -1122
rect 1584 -1134 1590 -1128
rect 1584 -1140 1590 -1134
rect 1584 -1146 1590 -1140
rect 1584 -1152 1590 -1146
rect 1584 -1158 1590 -1152
rect 1584 -1164 1590 -1158
rect 1584 -1170 1590 -1164
rect 1584 -1176 1590 -1170
rect 1584 -1182 1590 -1176
rect 1584 -1188 1590 -1182
rect 1584 -1194 1590 -1188
rect 1584 -1200 1590 -1194
rect 1584 -1206 1590 -1200
rect 1584 -1212 1590 -1206
rect 1584 -1218 1590 -1212
rect 1584 -1224 1590 -1218
rect 1584 -1230 1590 -1224
rect 1584 -1236 1590 -1230
rect 1584 -1242 1590 -1236
rect 1584 -1248 1590 -1242
rect 1584 -1254 1590 -1248
rect 1584 -1260 1590 -1254
rect 1584 -1266 1590 -1260
rect 1584 -1272 1590 -1266
rect 1584 -1278 1590 -1272
rect 1584 -1284 1590 -1278
rect 1584 -1290 1590 -1284
rect 1584 -1296 1590 -1290
rect 1584 -1302 1590 -1296
rect 1584 -1308 1590 -1302
rect 1584 -1314 1590 -1308
rect 1584 -1320 1590 -1314
rect 1584 -1326 1590 -1320
rect 1584 -1332 1590 -1326
rect 1584 -1338 1590 -1332
rect 1584 -1344 1590 -1338
rect 1584 -1350 1590 -1344
rect 1584 -1356 1590 -1350
rect 1584 -1362 1590 -1356
rect 1584 -1368 1590 -1362
rect 1584 -1374 1590 -1368
rect 1584 -1380 1590 -1374
rect 1584 -1386 1590 -1380
rect 1584 -1392 1590 -1386
rect 1584 -1398 1590 -1392
rect 1584 -1404 1590 -1398
rect 1584 -1410 1590 -1404
rect 1584 -1416 1590 -1410
rect 1584 -1422 1590 -1416
rect 1584 -1428 1590 -1422
rect 1584 -1434 1590 -1428
rect 1584 -1440 1590 -1434
rect 1584 -1446 1590 -1440
rect 1584 -1452 1590 -1446
rect 1584 -1458 1590 -1452
rect 1584 -1464 1590 -1458
rect 1584 -1470 1590 -1464
rect 1584 -1476 1590 -1470
rect 1584 -1482 1590 -1476
rect 1584 -1488 1590 -1482
rect 1584 -1494 1590 -1488
rect 1584 -1500 1590 -1494
rect 1584 -1506 1590 -1500
rect 1584 -1512 1590 -1506
rect 1584 -1518 1590 -1512
rect 1584 -1524 1590 -1518
rect 1584 -1530 1590 -1524
rect 1584 -1536 1590 -1530
rect 1584 -1542 1590 -1536
rect 1584 -1548 1590 -1542
rect 1584 -1554 1590 -1548
rect 1584 -1560 1590 -1554
rect 1584 -1566 1590 -1560
rect 1584 -1572 1590 -1566
rect 1584 -1578 1590 -1572
rect 1584 -1584 1590 -1578
rect 1584 -1590 1590 -1584
rect 1584 -1596 1590 -1590
rect 1584 -1602 1590 -1596
rect 1584 -1608 1590 -1602
rect 1584 -1614 1590 -1608
rect 1584 -1620 1590 -1614
rect 1584 -1626 1590 -1620
rect 1584 -1632 1590 -1626
rect 1584 -1638 1590 -1632
rect 1584 -1644 1590 -1638
rect 1584 -1650 1590 -1644
rect 1584 -1656 1590 -1650
rect 1584 -1662 1590 -1656
rect 1584 -1668 1590 -1662
rect 1584 -1674 1590 -1668
rect 1584 -1680 1590 -1674
rect 1584 -1686 1590 -1680
rect 1584 -1692 1590 -1686
rect 1584 -1698 1590 -1692
rect 1584 -1704 1590 -1698
rect 1584 -1710 1590 -1704
rect 1584 -1716 1590 -1710
rect 1584 -1722 1590 -1716
rect 1584 -1728 1590 -1722
rect 1584 -1734 1590 -1728
rect 1584 -1740 1590 -1734
rect 1584 -1746 1590 -1740
rect 1584 -1752 1590 -1746
rect 1584 -1758 1590 -1752
rect 1584 -1764 1590 -1758
rect 1584 -1770 1590 -1764
rect 1584 -1776 1590 -1770
rect 1584 -1782 1590 -1776
rect 1584 -1788 1590 -1782
rect 1584 -1794 1590 -1788
rect 1584 -1800 1590 -1794
rect 1584 -1806 1590 -1800
rect 1584 -1812 1590 -1806
rect 1584 -1818 1590 -1812
rect 1584 -1824 1590 -1818
rect 1584 -1830 1590 -1824
rect 1584 -1836 1590 -1830
rect 1584 -1842 1590 -1836
rect 1584 -1848 1590 -1842
rect 1584 -1854 1590 -1848
rect 1584 -1860 1590 -1854
rect 1584 -1866 1590 -1860
rect 1584 -1872 1590 -1866
rect 1584 -1878 1590 -1872
rect 1584 -1884 1590 -1878
rect 1584 -1890 1590 -1884
rect 1584 -1896 1590 -1890
rect 1584 -1902 1590 -1896
rect 1584 -1908 1590 -1902
rect 1584 -1914 1590 -1908
rect 1584 -1920 1590 -1914
rect 1584 -1926 1590 -1920
rect 1584 -1932 1590 -1926
rect 1584 -1938 1590 -1932
rect 1584 -1944 1590 -1938
rect 1584 -1950 1590 -1944
rect 1584 -1956 1590 -1950
rect 1584 -1962 1590 -1956
rect 1584 -1968 1590 -1962
rect 1584 -1974 1590 -1968
rect 1584 -1980 1590 -1974
rect 1584 -1986 1590 -1980
rect 1584 -1992 1590 -1986
rect 1584 -1998 1590 -1992
rect 1584 -2004 1590 -1998
rect 1584 -2010 1590 -2004
rect 1584 -2016 1590 -2010
rect 1584 -2022 1590 -2016
rect 1584 -2028 1590 -2022
rect 1584 -2034 1590 -2028
rect 1584 -2040 1590 -2034
rect 1584 -2046 1590 -2040
rect 1584 -2052 1590 -2046
rect 1584 -2058 1590 -2052
rect 1584 -2064 1590 -2058
rect 1584 -2070 1590 -2064
rect 1584 -2076 1590 -2070
rect 1584 -2082 1590 -2076
rect 1584 -2088 1590 -2082
rect 1584 -2160 1590 -2154
rect 1584 -2166 1590 -2160
rect 1584 -2172 1590 -2166
rect 1584 -2178 1590 -2172
rect 1584 -2184 1590 -2178
rect 1584 -2190 1590 -2184
rect 1584 -2196 1590 -2190
rect 1584 -2202 1590 -2196
rect 1584 -2208 1590 -2202
rect 1584 -2214 1590 -2208
rect 1584 -2220 1590 -2214
rect 1584 -2226 1590 -2220
rect 1584 -2232 1590 -2226
rect 1584 -2238 1590 -2232
rect 1584 -2244 1590 -2238
rect 1584 -2250 1590 -2244
rect 1584 -2256 1590 -2250
rect 1584 -2262 1590 -2256
rect 1584 -2268 1590 -2262
rect 1584 -2274 1590 -2268
rect 1584 -2280 1590 -2274
rect 1584 -2286 1590 -2280
rect 1584 -2292 1590 -2286
rect 1584 -2298 1590 -2292
rect 1584 -2304 1590 -2298
rect 1584 -2310 1590 -2304
rect 1584 -2316 1590 -2310
rect 1584 -2322 1590 -2316
rect 1584 -2328 1590 -2322
rect 1584 -2334 1590 -2328
rect 1584 -2340 1590 -2334
rect 1584 -2346 1590 -2340
rect 1584 -2352 1590 -2346
rect 1584 -2358 1590 -2352
rect 1584 -2364 1590 -2358
rect 1584 -2370 1590 -2364
rect 1584 -2376 1590 -2370
rect 1584 -2382 1590 -2376
rect 1584 -2388 1590 -2382
rect 1584 -2394 1590 -2388
rect 1584 -2400 1590 -2394
rect 1584 -2406 1590 -2400
rect 1584 -2412 1590 -2406
rect 1584 -2418 1590 -2412
rect 1584 -2424 1590 -2418
rect 1584 -2430 1590 -2424
rect 1584 -2436 1590 -2430
rect 1584 -2442 1590 -2436
rect 1584 -2448 1590 -2442
rect 1584 -2454 1590 -2448
rect 1584 -2460 1590 -2454
rect 1584 -2466 1590 -2460
rect 1584 -2472 1590 -2466
rect 1584 -2478 1590 -2472
rect 1584 -2484 1590 -2478
rect 1584 -2490 1590 -2484
rect 1584 -2496 1590 -2490
rect 1584 -2502 1590 -2496
rect 1584 -2508 1590 -2502
rect 1584 -2514 1590 -2508
rect 1584 -2520 1590 -2514
rect 1584 -2526 1590 -2520
rect 1584 -2532 1590 -2526
rect 1584 -2538 1590 -2532
rect 1584 -2544 1590 -2538
rect 1584 -2550 1590 -2544
rect 1584 -2556 1590 -2550
rect 1584 -2562 1590 -2556
rect 1584 -2568 1590 -2562
rect 1584 -2574 1590 -2568
rect 1584 -2580 1590 -2574
rect 1584 -2586 1590 -2580
rect 1584 -2592 1590 -2586
rect 1584 -2598 1590 -2592
rect 1584 -2604 1590 -2598
rect 1584 -2610 1590 -2604
rect 1584 -2616 1590 -2610
rect 1584 -2622 1590 -2616
rect 1584 -2628 1590 -2622
rect 1584 -2634 1590 -2628
rect 1584 -2640 1590 -2634
rect 1584 -2646 1590 -2640
rect 1584 -2652 1590 -2646
rect 1584 -2658 1590 -2652
rect 1584 -2664 1590 -2658
rect 1584 -2670 1590 -2664
rect 1584 -2676 1590 -2670
rect 1584 -2682 1590 -2676
rect 1584 -2688 1590 -2682
rect 1584 -2694 1590 -2688
rect 1584 -2700 1590 -2694
rect 1584 -2706 1590 -2700
rect 1584 -2712 1590 -2706
rect 1584 -2718 1590 -2712
rect 1584 -2724 1590 -2718
rect 1584 -2730 1590 -2724
rect 1584 -2736 1590 -2730
rect 1584 -2742 1590 -2736
rect 1584 -2748 1590 -2742
rect 1584 -2754 1590 -2748
rect 1584 -2838 1590 -2832
rect 1584 -2844 1590 -2838
rect 1584 -2850 1590 -2844
rect 1584 -2856 1590 -2850
rect 1584 -2862 1590 -2856
rect 1584 -2868 1590 -2862
rect 1584 -2874 1590 -2868
rect 1584 -2880 1590 -2874
rect 1584 -2886 1590 -2880
rect 1584 -2892 1590 -2886
rect 1584 -2898 1590 -2892
rect 1584 -2904 1590 -2898
rect 1584 -2910 1590 -2904
rect 1584 -2916 1590 -2910
rect 1584 -2922 1590 -2916
rect 1584 -2928 1590 -2922
rect 1584 -2934 1590 -2928
rect 1584 -2940 1590 -2934
rect 1584 -2946 1590 -2940
rect 1584 -2952 1590 -2946
rect 1584 -2958 1590 -2952
rect 1584 -2964 1590 -2958
rect 1584 -2970 1590 -2964
rect 1584 -2976 1590 -2970
rect 1584 -2982 1590 -2976
rect 1584 -2988 1590 -2982
rect 1584 -2994 1590 -2988
rect 1584 -3000 1590 -2994
rect 1584 -3006 1590 -3000
rect 1584 -3012 1590 -3006
rect 1584 -3018 1590 -3012
rect 1584 -3024 1590 -3018
rect 1584 -3030 1590 -3024
rect 1584 -3036 1590 -3030
rect 1584 -3042 1590 -3036
rect 1584 -3048 1590 -3042
rect 1584 -3054 1590 -3048
rect 1584 -3060 1590 -3054
rect 1584 -3066 1590 -3060
rect 1584 -3072 1590 -3066
rect 1584 -3078 1590 -3072
rect 1584 -3084 1590 -3078
rect 1584 -3090 1590 -3084
rect 1584 -3096 1590 -3090
rect 1584 -3102 1590 -3096
rect 1584 -3108 1590 -3102
rect 1584 -3114 1590 -3108
rect 1584 -3120 1590 -3114
rect 1584 -3126 1590 -3120
rect 1584 -3132 1590 -3126
rect 1584 -3138 1590 -3132
rect 1584 -3144 1590 -3138
rect 1584 -3150 1590 -3144
rect 1584 -3156 1590 -3150
rect 1584 -3162 1590 -3156
rect 1584 -3168 1590 -3162
rect 1584 -3174 1590 -3168
rect 1584 -3180 1590 -3174
rect 1584 -3186 1590 -3180
rect 1584 -3192 1590 -3186
rect 1584 -3198 1590 -3192
rect 1584 -3204 1590 -3198
rect 1584 -3210 1590 -3204
rect 1584 -3216 1590 -3210
rect 1584 -3222 1590 -3216
rect 1584 -3228 1590 -3222
rect 1584 -3234 1590 -3228
rect 1584 -3276 1590 -3270
rect 1584 -3282 1590 -3276
rect 1584 -3288 1590 -3282
rect 1584 -3294 1590 -3288
rect 1584 -3300 1590 -3294
rect 1584 -3306 1590 -3300
rect 1584 -3312 1590 -3306
rect 1584 -3318 1590 -3312
rect 1584 -3324 1590 -3318
rect 1584 -3330 1590 -3324
rect 1584 -3336 1590 -3330
rect 1584 -3342 1590 -3336
rect 1584 -3348 1590 -3342
rect 1584 -3354 1590 -3348
rect 1584 -3360 1590 -3354
rect 1584 -3366 1590 -3360
rect 1584 -3372 1590 -3366
rect 1584 -3378 1590 -3372
rect 1584 -3384 1590 -3378
rect 1584 -3390 1590 -3384
rect 1584 -3396 1590 -3390
rect 1584 -3402 1590 -3396
rect 1584 -3408 1590 -3402
rect 1584 -3414 1590 -3408
rect 1584 -3420 1590 -3414
rect 1584 -3426 1590 -3420
rect 1584 -3432 1590 -3426
rect 1584 -3438 1590 -3432
rect 1584 -3444 1590 -3438
rect 1584 -3450 1590 -3444
rect 1584 -3456 1590 -3450
rect 1584 -3462 1590 -3456
rect 1590 -1032 1596 -1026
rect 1590 -1038 1596 -1032
rect 1590 -1044 1596 -1038
rect 1590 -1050 1596 -1044
rect 1590 -1056 1596 -1050
rect 1590 -1062 1596 -1056
rect 1590 -1068 1596 -1062
rect 1590 -1074 1596 -1068
rect 1590 -1080 1596 -1074
rect 1590 -1086 1596 -1080
rect 1590 -1092 1596 -1086
rect 1590 -1098 1596 -1092
rect 1590 -1104 1596 -1098
rect 1590 -1110 1596 -1104
rect 1590 -1116 1596 -1110
rect 1590 -1122 1596 -1116
rect 1590 -1128 1596 -1122
rect 1590 -1134 1596 -1128
rect 1590 -1140 1596 -1134
rect 1590 -1146 1596 -1140
rect 1590 -1152 1596 -1146
rect 1590 -1158 1596 -1152
rect 1590 -1164 1596 -1158
rect 1590 -1170 1596 -1164
rect 1590 -1176 1596 -1170
rect 1590 -1182 1596 -1176
rect 1590 -1188 1596 -1182
rect 1590 -1194 1596 -1188
rect 1590 -1200 1596 -1194
rect 1590 -1206 1596 -1200
rect 1590 -1212 1596 -1206
rect 1590 -1218 1596 -1212
rect 1590 -1224 1596 -1218
rect 1590 -1230 1596 -1224
rect 1590 -1236 1596 -1230
rect 1590 -1242 1596 -1236
rect 1590 -1248 1596 -1242
rect 1590 -1254 1596 -1248
rect 1590 -1260 1596 -1254
rect 1590 -1266 1596 -1260
rect 1590 -1272 1596 -1266
rect 1590 -1278 1596 -1272
rect 1590 -1284 1596 -1278
rect 1590 -1290 1596 -1284
rect 1590 -1296 1596 -1290
rect 1590 -1302 1596 -1296
rect 1590 -1308 1596 -1302
rect 1590 -1314 1596 -1308
rect 1590 -1320 1596 -1314
rect 1590 -1326 1596 -1320
rect 1590 -1332 1596 -1326
rect 1590 -1338 1596 -1332
rect 1590 -1344 1596 -1338
rect 1590 -1350 1596 -1344
rect 1590 -1356 1596 -1350
rect 1590 -1362 1596 -1356
rect 1590 -1368 1596 -1362
rect 1590 -1374 1596 -1368
rect 1590 -1380 1596 -1374
rect 1590 -1386 1596 -1380
rect 1590 -1392 1596 -1386
rect 1590 -1398 1596 -1392
rect 1590 -1404 1596 -1398
rect 1590 -1410 1596 -1404
rect 1590 -1416 1596 -1410
rect 1590 -1422 1596 -1416
rect 1590 -1428 1596 -1422
rect 1590 -1434 1596 -1428
rect 1590 -1440 1596 -1434
rect 1590 -1446 1596 -1440
rect 1590 -1452 1596 -1446
rect 1590 -1458 1596 -1452
rect 1590 -1464 1596 -1458
rect 1590 -1470 1596 -1464
rect 1590 -1476 1596 -1470
rect 1590 -1482 1596 -1476
rect 1590 -1488 1596 -1482
rect 1590 -1494 1596 -1488
rect 1590 -1500 1596 -1494
rect 1590 -1506 1596 -1500
rect 1590 -1512 1596 -1506
rect 1590 -1518 1596 -1512
rect 1590 -1524 1596 -1518
rect 1590 -1530 1596 -1524
rect 1590 -1536 1596 -1530
rect 1590 -1542 1596 -1536
rect 1590 -1548 1596 -1542
rect 1590 -1554 1596 -1548
rect 1590 -1560 1596 -1554
rect 1590 -1566 1596 -1560
rect 1590 -1572 1596 -1566
rect 1590 -1578 1596 -1572
rect 1590 -1584 1596 -1578
rect 1590 -1590 1596 -1584
rect 1590 -1596 1596 -1590
rect 1590 -1602 1596 -1596
rect 1590 -1608 1596 -1602
rect 1590 -1614 1596 -1608
rect 1590 -1620 1596 -1614
rect 1590 -1626 1596 -1620
rect 1590 -1632 1596 -1626
rect 1590 -1638 1596 -1632
rect 1590 -1644 1596 -1638
rect 1590 -1650 1596 -1644
rect 1590 -1656 1596 -1650
rect 1590 -1662 1596 -1656
rect 1590 -1668 1596 -1662
rect 1590 -1674 1596 -1668
rect 1590 -1680 1596 -1674
rect 1590 -1686 1596 -1680
rect 1590 -1692 1596 -1686
rect 1590 -1698 1596 -1692
rect 1590 -1704 1596 -1698
rect 1590 -1710 1596 -1704
rect 1590 -1716 1596 -1710
rect 1590 -1722 1596 -1716
rect 1590 -1728 1596 -1722
rect 1590 -1734 1596 -1728
rect 1590 -1740 1596 -1734
rect 1590 -1746 1596 -1740
rect 1590 -1752 1596 -1746
rect 1590 -1758 1596 -1752
rect 1590 -1764 1596 -1758
rect 1590 -1770 1596 -1764
rect 1590 -1776 1596 -1770
rect 1590 -1782 1596 -1776
rect 1590 -1788 1596 -1782
rect 1590 -1794 1596 -1788
rect 1590 -1800 1596 -1794
rect 1590 -1806 1596 -1800
rect 1590 -1812 1596 -1806
rect 1590 -1818 1596 -1812
rect 1590 -1824 1596 -1818
rect 1590 -1830 1596 -1824
rect 1590 -1836 1596 -1830
rect 1590 -1842 1596 -1836
rect 1590 -1848 1596 -1842
rect 1590 -1854 1596 -1848
rect 1590 -1860 1596 -1854
rect 1590 -1866 1596 -1860
rect 1590 -1872 1596 -1866
rect 1590 -1878 1596 -1872
rect 1590 -1884 1596 -1878
rect 1590 -1890 1596 -1884
rect 1590 -1896 1596 -1890
rect 1590 -1902 1596 -1896
rect 1590 -1908 1596 -1902
rect 1590 -1914 1596 -1908
rect 1590 -1920 1596 -1914
rect 1590 -1926 1596 -1920
rect 1590 -1932 1596 -1926
rect 1590 -1938 1596 -1932
rect 1590 -1944 1596 -1938
rect 1590 -1950 1596 -1944
rect 1590 -1956 1596 -1950
rect 1590 -1962 1596 -1956
rect 1590 -1968 1596 -1962
rect 1590 -1974 1596 -1968
rect 1590 -1980 1596 -1974
rect 1590 -1986 1596 -1980
rect 1590 -1992 1596 -1986
rect 1590 -1998 1596 -1992
rect 1590 -2004 1596 -1998
rect 1590 -2010 1596 -2004
rect 1590 -2016 1596 -2010
rect 1590 -2022 1596 -2016
rect 1590 -2028 1596 -2022
rect 1590 -2034 1596 -2028
rect 1590 -2040 1596 -2034
rect 1590 -2046 1596 -2040
rect 1590 -2052 1596 -2046
rect 1590 -2058 1596 -2052
rect 1590 -2064 1596 -2058
rect 1590 -2070 1596 -2064
rect 1590 -2076 1596 -2070
rect 1590 -2082 1596 -2076
rect 1590 -2154 1596 -2148
rect 1590 -2160 1596 -2154
rect 1590 -2166 1596 -2160
rect 1590 -2172 1596 -2166
rect 1590 -2178 1596 -2172
rect 1590 -2184 1596 -2178
rect 1590 -2190 1596 -2184
rect 1590 -2196 1596 -2190
rect 1590 -2202 1596 -2196
rect 1590 -2208 1596 -2202
rect 1590 -2214 1596 -2208
rect 1590 -2220 1596 -2214
rect 1590 -2226 1596 -2220
rect 1590 -2232 1596 -2226
rect 1590 -2238 1596 -2232
rect 1590 -2244 1596 -2238
rect 1590 -2250 1596 -2244
rect 1590 -2256 1596 -2250
rect 1590 -2262 1596 -2256
rect 1590 -2268 1596 -2262
rect 1590 -2274 1596 -2268
rect 1590 -2280 1596 -2274
rect 1590 -2286 1596 -2280
rect 1590 -2292 1596 -2286
rect 1590 -2298 1596 -2292
rect 1590 -2304 1596 -2298
rect 1590 -2310 1596 -2304
rect 1590 -2316 1596 -2310
rect 1590 -2322 1596 -2316
rect 1590 -2328 1596 -2322
rect 1590 -2334 1596 -2328
rect 1590 -2340 1596 -2334
rect 1590 -2346 1596 -2340
rect 1590 -2352 1596 -2346
rect 1590 -2358 1596 -2352
rect 1590 -2364 1596 -2358
rect 1590 -2370 1596 -2364
rect 1590 -2376 1596 -2370
rect 1590 -2382 1596 -2376
rect 1590 -2388 1596 -2382
rect 1590 -2394 1596 -2388
rect 1590 -2400 1596 -2394
rect 1590 -2406 1596 -2400
rect 1590 -2412 1596 -2406
rect 1590 -2418 1596 -2412
rect 1590 -2424 1596 -2418
rect 1590 -2430 1596 -2424
rect 1590 -2436 1596 -2430
rect 1590 -2442 1596 -2436
rect 1590 -2448 1596 -2442
rect 1590 -2454 1596 -2448
rect 1590 -2460 1596 -2454
rect 1590 -2466 1596 -2460
rect 1590 -2472 1596 -2466
rect 1590 -2478 1596 -2472
rect 1590 -2484 1596 -2478
rect 1590 -2490 1596 -2484
rect 1590 -2496 1596 -2490
rect 1590 -2502 1596 -2496
rect 1590 -2508 1596 -2502
rect 1590 -2514 1596 -2508
rect 1590 -2520 1596 -2514
rect 1590 -2526 1596 -2520
rect 1590 -2532 1596 -2526
rect 1590 -2538 1596 -2532
rect 1590 -2544 1596 -2538
rect 1590 -2550 1596 -2544
rect 1590 -2556 1596 -2550
rect 1590 -2562 1596 -2556
rect 1590 -2568 1596 -2562
rect 1590 -2574 1596 -2568
rect 1590 -2580 1596 -2574
rect 1590 -2586 1596 -2580
rect 1590 -2592 1596 -2586
rect 1590 -2598 1596 -2592
rect 1590 -2604 1596 -2598
rect 1590 -2610 1596 -2604
rect 1590 -2616 1596 -2610
rect 1590 -2622 1596 -2616
rect 1590 -2628 1596 -2622
rect 1590 -2634 1596 -2628
rect 1590 -2640 1596 -2634
rect 1590 -2646 1596 -2640
rect 1590 -2652 1596 -2646
rect 1590 -2658 1596 -2652
rect 1590 -2664 1596 -2658
rect 1590 -2670 1596 -2664
rect 1590 -2676 1596 -2670
rect 1590 -2682 1596 -2676
rect 1590 -2688 1596 -2682
rect 1590 -2694 1596 -2688
rect 1590 -2700 1596 -2694
rect 1590 -2706 1596 -2700
rect 1590 -2712 1596 -2706
rect 1590 -2718 1596 -2712
rect 1590 -2724 1596 -2718
rect 1590 -2730 1596 -2724
rect 1590 -2736 1596 -2730
rect 1590 -2742 1596 -2736
rect 1590 -2748 1596 -2742
rect 1590 -2754 1596 -2748
rect 1590 -2832 1596 -2826
rect 1590 -2838 1596 -2832
rect 1590 -2844 1596 -2838
rect 1590 -2850 1596 -2844
rect 1590 -2856 1596 -2850
rect 1590 -2862 1596 -2856
rect 1590 -2868 1596 -2862
rect 1590 -2874 1596 -2868
rect 1590 -2880 1596 -2874
rect 1590 -2886 1596 -2880
rect 1590 -2892 1596 -2886
rect 1590 -2898 1596 -2892
rect 1590 -2904 1596 -2898
rect 1590 -2910 1596 -2904
rect 1590 -2916 1596 -2910
rect 1590 -2922 1596 -2916
rect 1590 -2928 1596 -2922
rect 1590 -2934 1596 -2928
rect 1590 -2940 1596 -2934
rect 1590 -2946 1596 -2940
rect 1590 -2952 1596 -2946
rect 1590 -2958 1596 -2952
rect 1590 -2964 1596 -2958
rect 1590 -2970 1596 -2964
rect 1590 -2976 1596 -2970
rect 1590 -2982 1596 -2976
rect 1590 -2988 1596 -2982
rect 1590 -2994 1596 -2988
rect 1590 -3000 1596 -2994
rect 1590 -3006 1596 -3000
rect 1590 -3012 1596 -3006
rect 1590 -3018 1596 -3012
rect 1590 -3024 1596 -3018
rect 1590 -3030 1596 -3024
rect 1590 -3036 1596 -3030
rect 1590 -3042 1596 -3036
rect 1590 -3048 1596 -3042
rect 1590 -3054 1596 -3048
rect 1590 -3060 1596 -3054
rect 1590 -3066 1596 -3060
rect 1590 -3072 1596 -3066
rect 1590 -3078 1596 -3072
rect 1590 -3084 1596 -3078
rect 1590 -3090 1596 -3084
rect 1590 -3096 1596 -3090
rect 1590 -3102 1596 -3096
rect 1590 -3108 1596 -3102
rect 1590 -3114 1596 -3108
rect 1590 -3120 1596 -3114
rect 1590 -3126 1596 -3120
rect 1590 -3132 1596 -3126
rect 1590 -3138 1596 -3132
rect 1590 -3144 1596 -3138
rect 1590 -3150 1596 -3144
rect 1590 -3156 1596 -3150
rect 1590 -3162 1596 -3156
rect 1590 -3168 1596 -3162
rect 1590 -3174 1596 -3168
rect 1590 -3180 1596 -3174
rect 1590 -3186 1596 -3180
rect 1590 -3192 1596 -3186
rect 1590 -3198 1596 -3192
rect 1590 -3204 1596 -3198
rect 1590 -3210 1596 -3204
rect 1590 -3216 1596 -3210
rect 1590 -3222 1596 -3216
rect 1590 -3228 1596 -3222
rect 1590 -3234 1596 -3228
rect 1590 -3276 1596 -3270
rect 1590 -3282 1596 -3276
rect 1590 -3288 1596 -3282
rect 1590 -3294 1596 -3288
rect 1590 -3300 1596 -3294
rect 1590 -3306 1596 -3300
rect 1590 -3312 1596 -3306
rect 1590 -3318 1596 -3312
rect 1590 -3324 1596 -3318
rect 1590 -3330 1596 -3324
rect 1590 -3336 1596 -3330
rect 1590 -3342 1596 -3336
rect 1590 -3348 1596 -3342
rect 1590 -3354 1596 -3348
rect 1590 -3360 1596 -3354
rect 1590 -3366 1596 -3360
rect 1590 -3372 1596 -3366
rect 1590 -3378 1596 -3372
rect 1590 -3384 1596 -3378
rect 1590 -3390 1596 -3384
rect 1590 -3396 1596 -3390
rect 1590 -3402 1596 -3396
rect 1590 -3408 1596 -3402
rect 1590 -3414 1596 -3408
rect 1590 -3420 1596 -3414
rect 1590 -3426 1596 -3420
rect 1590 -3432 1596 -3426
rect 1590 -3438 1596 -3432
rect 1590 -3444 1596 -3438
rect 1590 -3450 1596 -3444
rect 1590 -3456 1596 -3450
rect 1590 -3462 1596 -3456
rect 1596 -1020 1602 -1014
rect 1596 -1026 1602 -1020
rect 1596 -1032 1602 -1026
rect 1596 -1038 1602 -1032
rect 1596 -1044 1602 -1038
rect 1596 -1050 1602 -1044
rect 1596 -1056 1602 -1050
rect 1596 -1062 1602 -1056
rect 1596 -1068 1602 -1062
rect 1596 -1074 1602 -1068
rect 1596 -1080 1602 -1074
rect 1596 -1086 1602 -1080
rect 1596 -1092 1602 -1086
rect 1596 -1098 1602 -1092
rect 1596 -1104 1602 -1098
rect 1596 -1110 1602 -1104
rect 1596 -1116 1602 -1110
rect 1596 -1122 1602 -1116
rect 1596 -1128 1602 -1122
rect 1596 -1134 1602 -1128
rect 1596 -1140 1602 -1134
rect 1596 -1146 1602 -1140
rect 1596 -1152 1602 -1146
rect 1596 -1158 1602 -1152
rect 1596 -1164 1602 -1158
rect 1596 -1170 1602 -1164
rect 1596 -1176 1602 -1170
rect 1596 -1182 1602 -1176
rect 1596 -1188 1602 -1182
rect 1596 -1194 1602 -1188
rect 1596 -1200 1602 -1194
rect 1596 -1206 1602 -1200
rect 1596 -1212 1602 -1206
rect 1596 -1218 1602 -1212
rect 1596 -1224 1602 -1218
rect 1596 -1230 1602 -1224
rect 1596 -1236 1602 -1230
rect 1596 -1242 1602 -1236
rect 1596 -1248 1602 -1242
rect 1596 -1254 1602 -1248
rect 1596 -1260 1602 -1254
rect 1596 -1266 1602 -1260
rect 1596 -1272 1602 -1266
rect 1596 -1278 1602 -1272
rect 1596 -1284 1602 -1278
rect 1596 -1290 1602 -1284
rect 1596 -1296 1602 -1290
rect 1596 -1302 1602 -1296
rect 1596 -1308 1602 -1302
rect 1596 -1314 1602 -1308
rect 1596 -1320 1602 -1314
rect 1596 -1326 1602 -1320
rect 1596 -1332 1602 -1326
rect 1596 -1338 1602 -1332
rect 1596 -1344 1602 -1338
rect 1596 -1350 1602 -1344
rect 1596 -1356 1602 -1350
rect 1596 -1362 1602 -1356
rect 1596 -1368 1602 -1362
rect 1596 -1374 1602 -1368
rect 1596 -1380 1602 -1374
rect 1596 -1386 1602 -1380
rect 1596 -1392 1602 -1386
rect 1596 -1398 1602 -1392
rect 1596 -1404 1602 -1398
rect 1596 -1410 1602 -1404
rect 1596 -1416 1602 -1410
rect 1596 -1422 1602 -1416
rect 1596 -1428 1602 -1422
rect 1596 -1434 1602 -1428
rect 1596 -1440 1602 -1434
rect 1596 -1446 1602 -1440
rect 1596 -1452 1602 -1446
rect 1596 -1458 1602 -1452
rect 1596 -1464 1602 -1458
rect 1596 -1470 1602 -1464
rect 1596 -1476 1602 -1470
rect 1596 -1482 1602 -1476
rect 1596 -1488 1602 -1482
rect 1596 -1494 1602 -1488
rect 1596 -1500 1602 -1494
rect 1596 -1506 1602 -1500
rect 1596 -1512 1602 -1506
rect 1596 -1518 1602 -1512
rect 1596 -1524 1602 -1518
rect 1596 -1530 1602 -1524
rect 1596 -1536 1602 -1530
rect 1596 -1542 1602 -1536
rect 1596 -1548 1602 -1542
rect 1596 -1554 1602 -1548
rect 1596 -1560 1602 -1554
rect 1596 -1566 1602 -1560
rect 1596 -1572 1602 -1566
rect 1596 -1578 1602 -1572
rect 1596 -1584 1602 -1578
rect 1596 -1590 1602 -1584
rect 1596 -1596 1602 -1590
rect 1596 -1602 1602 -1596
rect 1596 -1608 1602 -1602
rect 1596 -1614 1602 -1608
rect 1596 -1620 1602 -1614
rect 1596 -1626 1602 -1620
rect 1596 -1632 1602 -1626
rect 1596 -1638 1602 -1632
rect 1596 -1644 1602 -1638
rect 1596 -1650 1602 -1644
rect 1596 -1656 1602 -1650
rect 1596 -1662 1602 -1656
rect 1596 -1668 1602 -1662
rect 1596 -1674 1602 -1668
rect 1596 -1680 1602 -1674
rect 1596 -1686 1602 -1680
rect 1596 -1692 1602 -1686
rect 1596 -1698 1602 -1692
rect 1596 -1704 1602 -1698
rect 1596 -1710 1602 -1704
rect 1596 -1716 1602 -1710
rect 1596 -1722 1602 -1716
rect 1596 -1728 1602 -1722
rect 1596 -1734 1602 -1728
rect 1596 -1740 1602 -1734
rect 1596 -1746 1602 -1740
rect 1596 -1752 1602 -1746
rect 1596 -1758 1602 -1752
rect 1596 -1764 1602 -1758
rect 1596 -1770 1602 -1764
rect 1596 -1776 1602 -1770
rect 1596 -1782 1602 -1776
rect 1596 -1788 1602 -1782
rect 1596 -1794 1602 -1788
rect 1596 -1800 1602 -1794
rect 1596 -1806 1602 -1800
rect 1596 -1812 1602 -1806
rect 1596 -1818 1602 -1812
rect 1596 -1824 1602 -1818
rect 1596 -1830 1602 -1824
rect 1596 -1836 1602 -1830
rect 1596 -1842 1602 -1836
rect 1596 -1848 1602 -1842
rect 1596 -1854 1602 -1848
rect 1596 -1860 1602 -1854
rect 1596 -1866 1602 -1860
rect 1596 -1872 1602 -1866
rect 1596 -1878 1602 -1872
rect 1596 -1884 1602 -1878
rect 1596 -1890 1602 -1884
rect 1596 -1896 1602 -1890
rect 1596 -1902 1602 -1896
rect 1596 -1908 1602 -1902
rect 1596 -1914 1602 -1908
rect 1596 -1920 1602 -1914
rect 1596 -1926 1602 -1920
rect 1596 -1932 1602 -1926
rect 1596 -1938 1602 -1932
rect 1596 -1944 1602 -1938
rect 1596 -1950 1602 -1944
rect 1596 -1956 1602 -1950
rect 1596 -1962 1602 -1956
rect 1596 -1968 1602 -1962
rect 1596 -1974 1602 -1968
rect 1596 -1980 1602 -1974
rect 1596 -1986 1602 -1980
rect 1596 -1992 1602 -1986
rect 1596 -1998 1602 -1992
rect 1596 -2004 1602 -1998
rect 1596 -2010 1602 -2004
rect 1596 -2016 1602 -2010
rect 1596 -2022 1602 -2016
rect 1596 -2028 1602 -2022
rect 1596 -2034 1602 -2028
rect 1596 -2040 1602 -2034
rect 1596 -2046 1602 -2040
rect 1596 -2052 1602 -2046
rect 1596 -2058 1602 -2052
rect 1596 -2064 1602 -2058
rect 1596 -2070 1602 -2064
rect 1596 -2148 1602 -2142
rect 1596 -2154 1602 -2148
rect 1596 -2160 1602 -2154
rect 1596 -2166 1602 -2160
rect 1596 -2172 1602 -2166
rect 1596 -2178 1602 -2172
rect 1596 -2184 1602 -2178
rect 1596 -2190 1602 -2184
rect 1596 -2196 1602 -2190
rect 1596 -2202 1602 -2196
rect 1596 -2208 1602 -2202
rect 1596 -2214 1602 -2208
rect 1596 -2220 1602 -2214
rect 1596 -2226 1602 -2220
rect 1596 -2232 1602 -2226
rect 1596 -2238 1602 -2232
rect 1596 -2244 1602 -2238
rect 1596 -2250 1602 -2244
rect 1596 -2256 1602 -2250
rect 1596 -2262 1602 -2256
rect 1596 -2268 1602 -2262
rect 1596 -2274 1602 -2268
rect 1596 -2280 1602 -2274
rect 1596 -2286 1602 -2280
rect 1596 -2292 1602 -2286
rect 1596 -2298 1602 -2292
rect 1596 -2304 1602 -2298
rect 1596 -2310 1602 -2304
rect 1596 -2316 1602 -2310
rect 1596 -2322 1602 -2316
rect 1596 -2328 1602 -2322
rect 1596 -2334 1602 -2328
rect 1596 -2340 1602 -2334
rect 1596 -2346 1602 -2340
rect 1596 -2352 1602 -2346
rect 1596 -2358 1602 -2352
rect 1596 -2364 1602 -2358
rect 1596 -2370 1602 -2364
rect 1596 -2376 1602 -2370
rect 1596 -2382 1602 -2376
rect 1596 -2388 1602 -2382
rect 1596 -2394 1602 -2388
rect 1596 -2400 1602 -2394
rect 1596 -2406 1602 -2400
rect 1596 -2412 1602 -2406
rect 1596 -2418 1602 -2412
rect 1596 -2424 1602 -2418
rect 1596 -2430 1602 -2424
rect 1596 -2436 1602 -2430
rect 1596 -2442 1602 -2436
rect 1596 -2448 1602 -2442
rect 1596 -2454 1602 -2448
rect 1596 -2460 1602 -2454
rect 1596 -2466 1602 -2460
rect 1596 -2472 1602 -2466
rect 1596 -2478 1602 -2472
rect 1596 -2484 1602 -2478
rect 1596 -2490 1602 -2484
rect 1596 -2496 1602 -2490
rect 1596 -2502 1602 -2496
rect 1596 -2508 1602 -2502
rect 1596 -2514 1602 -2508
rect 1596 -2520 1602 -2514
rect 1596 -2526 1602 -2520
rect 1596 -2532 1602 -2526
rect 1596 -2538 1602 -2532
rect 1596 -2544 1602 -2538
rect 1596 -2550 1602 -2544
rect 1596 -2556 1602 -2550
rect 1596 -2562 1602 -2556
rect 1596 -2568 1602 -2562
rect 1596 -2574 1602 -2568
rect 1596 -2580 1602 -2574
rect 1596 -2586 1602 -2580
rect 1596 -2592 1602 -2586
rect 1596 -2598 1602 -2592
rect 1596 -2604 1602 -2598
rect 1596 -2610 1602 -2604
rect 1596 -2616 1602 -2610
rect 1596 -2622 1602 -2616
rect 1596 -2628 1602 -2622
rect 1596 -2634 1602 -2628
rect 1596 -2640 1602 -2634
rect 1596 -2646 1602 -2640
rect 1596 -2652 1602 -2646
rect 1596 -2658 1602 -2652
rect 1596 -2664 1602 -2658
rect 1596 -2670 1602 -2664
rect 1596 -2676 1602 -2670
rect 1596 -2682 1602 -2676
rect 1596 -2688 1602 -2682
rect 1596 -2694 1602 -2688
rect 1596 -2700 1602 -2694
rect 1596 -2706 1602 -2700
rect 1596 -2712 1602 -2706
rect 1596 -2718 1602 -2712
rect 1596 -2724 1602 -2718
rect 1596 -2730 1602 -2724
rect 1596 -2736 1602 -2730
rect 1596 -2742 1602 -2736
rect 1596 -2748 1602 -2742
rect 1596 -2832 1602 -2826
rect 1596 -2838 1602 -2832
rect 1596 -2844 1602 -2838
rect 1596 -2850 1602 -2844
rect 1596 -2856 1602 -2850
rect 1596 -2862 1602 -2856
rect 1596 -2868 1602 -2862
rect 1596 -2874 1602 -2868
rect 1596 -2880 1602 -2874
rect 1596 -2886 1602 -2880
rect 1596 -2892 1602 -2886
rect 1596 -2898 1602 -2892
rect 1596 -2904 1602 -2898
rect 1596 -2910 1602 -2904
rect 1596 -2916 1602 -2910
rect 1596 -2922 1602 -2916
rect 1596 -2928 1602 -2922
rect 1596 -2934 1602 -2928
rect 1596 -2940 1602 -2934
rect 1596 -2946 1602 -2940
rect 1596 -2952 1602 -2946
rect 1596 -2958 1602 -2952
rect 1596 -2964 1602 -2958
rect 1596 -2970 1602 -2964
rect 1596 -2976 1602 -2970
rect 1596 -2982 1602 -2976
rect 1596 -2988 1602 -2982
rect 1596 -2994 1602 -2988
rect 1596 -3000 1602 -2994
rect 1596 -3006 1602 -3000
rect 1596 -3012 1602 -3006
rect 1596 -3018 1602 -3012
rect 1596 -3024 1602 -3018
rect 1596 -3030 1602 -3024
rect 1596 -3036 1602 -3030
rect 1596 -3042 1602 -3036
rect 1596 -3048 1602 -3042
rect 1596 -3054 1602 -3048
rect 1596 -3060 1602 -3054
rect 1596 -3066 1602 -3060
rect 1596 -3072 1602 -3066
rect 1596 -3078 1602 -3072
rect 1596 -3084 1602 -3078
rect 1596 -3090 1602 -3084
rect 1596 -3096 1602 -3090
rect 1596 -3102 1602 -3096
rect 1596 -3108 1602 -3102
rect 1596 -3114 1602 -3108
rect 1596 -3120 1602 -3114
rect 1596 -3126 1602 -3120
rect 1596 -3132 1602 -3126
rect 1596 -3138 1602 -3132
rect 1596 -3144 1602 -3138
rect 1596 -3150 1602 -3144
rect 1596 -3156 1602 -3150
rect 1596 -3162 1602 -3156
rect 1596 -3168 1602 -3162
rect 1596 -3174 1602 -3168
rect 1596 -3180 1602 -3174
rect 1596 -3186 1602 -3180
rect 1596 -3192 1602 -3186
rect 1596 -3198 1602 -3192
rect 1596 -3204 1602 -3198
rect 1596 -3210 1602 -3204
rect 1596 -3216 1602 -3210
rect 1596 -3222 1602 -3216
rect 1596 -3228 1602 -3222
rect 1596 -3234 1602 -3228
rect 1596 -3276 1602 -3270
rect 1596 -3282 1602 -3276
rect 1596 -3288 1602 -3282
rect 1596 -3294 1602 -3288
rect 1596 -3300 1602 -3294
rect 1596 -3306 1602 -3300
rect 1596 -3312 1602 -3306
rect 1596 -3318 1602 -3312
rect 1596 -3324 1602 -3318
rect 1596 -3330 1602 -3324
rect 1596 -3336 1602 -3330
rect 1596 -3342 1602 -3336
rect 1596 -3348 1602 -3342
rect 1596 -3354 1602 -3348
rect 1596 -3360 1602 -3354
rect 1596 -3366 1602 -3360
rect 1596 -3372 1602 -3366
rect 1596 -3378 1602 -3372
rect 1596 -3384 1602 -3378
rect 1596 -3390 1602 -3384
rect 1596 -3396 1602 -3390
rect 1596 -3402 1602 -3396
rect 1596 -3408 1602 -3402
rect 1596 -3414 1602 -3408
rect 1596 -3420 1602 -3414
rect 1596 -3426 1602 -3420
rect 1596 -3432 1602 -3426
rect 1596 -3438 1602 -3432
rect 1596 -3444 1602 -3438
rect 1596 -3450 1602 -3444
rect 1596 -3456 1602 -3450
rect 1596 -3462 1602 -3456
rect 1602 -1014 1608 -1008
rect 1602 -1020 1608 -1014
rect 1602 -1026 1608 -1020
rect 1602 -1032 1608 -1026
rect 1602 -1038 1608 -1032
rect 1602 -1044 1608 -1038
rect 1602 -1050 1608 -1044
rect 1602 -1056 1608 -1050
rect 1602 -1062 1608 -1056
rect 1602 -1068 1608 -1062
rect 1602 -1074 1608 -1068
rect 1602 -1080 1608 -1074
rect 1602 -1086 1608 -1080
rect 1602 -1092 1608 -1086
rect 1602 -1098 1608 -1092
rect 1602 -1104 1608 -1098
rect 1602 -1110 1608 -1104
rect 1602 -1116 1608 -1110
rect 1602 -1122 1608 -1116
rect 1602 -1128 1608 -1122
rect 1602 -1134 1608 -1128
rect 1602 -1140 1608 -1134
rect 1602 -1146 1608 -1140
rect 1602 -1152 1608 -1146
rect 1602 -1158 1608 -1152
rect 1602 -1164 1608 -1158
rect 1602 -1170 1608 -1164
rect 1602 -1176 1608 -1170
rect 1602 -1182 1608 -1176
rect 1602 -1188 1608 -1182
rect 1602 -1194 1608 -1188
rect 1602 -1200 1608 -1194
rect 1602 -1206 1608 -1200
rect 1602 -1212 1608 -1206
rect 1602 -1218 1608 -1212
rect 1602 -1224 1608 -1218
rect 1602 -1230 1608 -1224
rect 1602 -1236 1608 -1230
rect 1602 -1242 1608 -1236
rect 1602 -1248 1608 -1242
rect 1602 -1254 1608 -1248
rect 1602 -1260 1608 -1254
rect 1602 -1266 1608 -1260
rect 1602 -1272 1608 -1266
rect 1602 -1278 1608 -1272
rect 1602 -1284 1608 -1278
rect 1602 -1290 1608 -1284
rect 1602 -1296 1608 -1290
rect 1602 -1302 1608 -1296
rect 1602 -1308 1608 -1302
rect 1602 -1314 1608 -1308
rect 1602 -1320 1608 -1314
rect 1602 -1326 1608 -1320
rect 1602 -1332 1608 -1326
rect 1602 -1338 1608 -1332
rect 1602 -1344 1608 -1338
rect 1602 -1350 1608 -1344
rect 1602 -1356 1608 -1350
rect 1602 -1362 1608 -1356
rect 1602 -1368 1608 -1362
rect 1602 -1374 1608 -1368
rect 1602 -1380 1608 -1374
rect 1602 -1386 1608 -1380
rect 1602 -1392 1608 -1386
rect 1602 -1398 1608 -1392
rect 1602 -1404 1608 -1398
rect 1602 -1410 1608 -1404
rect 1602 -1416 1608 -1410
rect 1602 -1422 1608 -1416
rect 1602 -1428 1608 -1422
rect 1602 -1434 1608 -1428
rect 1602 -1440 1608 -1434
rect 1602 -1446 1608 -1440
rect 1602 -1452 1608 -1446
rect 1602 -1458 1608 -1452
rect 1602 -1464 1608 -1458
rect 1602 -1470 1608 -1464
rect 1602 -1476 1608 -1470
rect 1602 -1482 1608 -1476
rect 1602 -1488 1608 -1482
rect 1602 -1494 1608 -1488
rect 1602 -1500 1608 -1494
rect 1602 -1506 1608 -1500
rect 1602 -1512 1608 -1506
rect 1602 -1518 1608 -1512
rect 1602 -1524 1608 -1518
rect 1602 -1530 1608 -1524
rect 1602 -1536 1608 -1530
rect 1602 -1542 1608 -1536
rect 1602 -1548 1608 -1542
rect 1602 -1554 1608 -1548
rect 1602 -1560 1608 -1554
rect 1602 -1566 1608 -1560
rect 1602 -1572 1608 -1566
rect 1602 -1578 1608 -1572
rect 1602 -1584 1608 -1578
rect 1602 -1590 1608 -1584
rect 1602 -1596 1608 -1590
rect 1602 -1602 1608 -1596
rect 1602 -1608 1608 -1602
rect 1602 -1614 1608 -1608
rect 1602 -1620 1608 -1614
rect 1602 -1626 1608 -1620
rect 1602 -1632 1608 -1626
rect 1602 -1638 1608 -1632
rect 1602 -1644 1608 -1638
rect 1602 -1650 1608 -1644
rect 1602 -1656 1608 -1650
rect 1602 -1662 1608 -1656
rect 1602 -1668 1608 -1662
rect 1602 -1674 1608 -1668
rect 1602 -1680 1608 -1674
rect 1602 -1686 1608 -1680
rect 1602 -1692 1608 -1686
rect 1602 -1698 1608 -1692
rect 1602 -1704 1608 -1698
rect 1602 -1710 1608 -1704
rect 1602 -1716 1608 -1710
rect 1602 -1722 1608 -1716
rect 1602 -1728 1608 -1722
rect 1602 -1734 1608 -1728
rect 1602 -1740 1608 -1734
rect 1602 -1746 1608 -1740
rect 1602 -1752 1608 -1746
rect 1602 -1758 1608 -1752
rect 1602 -1764 1608 -1758
rect 1602 -1770 1608 -1764
rect 1602 -1776 1608 -1770
rect 1602 -1782 1608 -1776
rect 1602 -1788 1608 -1782
rect 1602 -1794 1608 -1788
rect 1602 -1800 1608 -1794
rect 1602 -1806 1608 -1800
rect 1602 -1812 1608 -1806
rect 1602 -1818 1608 -1812
rect 1602 -1824 1608 -1818
rect 1602 -1830 1608 -1824
rect 1602 -1836 1608 -1830
rect 1602 -1842 1608 -1836
rect 1602 -1848 1608 -1842
rect 1602 -1854 1608 -1848
rect 1602 -1860 1608 -1854
rect 1602 -1866 1608 -1860
rect 1602 -1872 1608 -1866
rect 1602 -1878 1608 -1872
rect 1602 -1884 1608 -1878
rect 1602 -1890 1608 -1884
rect 1602 -1896 1608 -1890
rect 1602 -1902 1608 -1896
rect 1602 -1908 1608 -1902
rect 1602 -1914 1608 -1908
rect 1602 -1920 1608 -1914
rect 1602 -1926 1608 -1920
rect 1602 -1932 1608 -1926
rect 1602 -1938 1608 -1932
rect 1602 -1944 1608 -1938
rect 1602 -1950 1608 -1944
rect 1602 -1956 1608 -1950
rect 1602 -1962 1608 -1956
rect 1602 -1968 1608 -1962
rect 1602 -1974 1608 -1968
rect 1602 -1980 1608 -1974
rect 1602 -1986 1608 -1980
rect 1602 -1992 1608 -1986
rect 1602 -1998 1608 -1992
rect 1602 -2004 1608 -1998
rect 1602 -2010 1608 -2004
rect 1602 -2016 1608 -2010
rect 1602 -2022 1608 -2016
rect 1602 -2028 1608 -2022
rect 1602 -2034 1608 -2028
rect 1602 -2040 1608 -2034
rect 1602 -2046 1608 -2040
rect 1602 -2052 1608 -2046
rect 1602 -2058 1608 -2052
rect 1602 -2064 1608 -2058
rect 1602 -2136 1608 -2130
rect 1602 -2142 1608 -2136
rect 1602 -2148 1608 -2142
rect 1602 -2154 1608 -2148
rect 1602 -2160 1608 -2154
rect 1602 -2166 1608 -2160
rect 1602 -2172 1608 -2166
rect 1602 -2178 1608 -2172
rect 1602 -2184 1608 -2178
rect 1602 -2190 1608 -2184
rect 1602 -2196 1608 -2190
rect 1602 -2202 1608 -2196
rect 1602 -2208 1608 -2202
rect 1602 -2214 1608 -2208
rect 1602 -2220 1608 -2214
rect 1602 -2226 1608 -2220
rect 1602 -2232 1608 -2226
rect 1602 -2238 1608 -2232
rect 1602 -2244 1608 -2238
rect 1602 -2250 1608 -2244
rect 1602 -2256 1608 -2250
rect 1602 -2262 1608 -2256
rect 1602 -2268 1608 -2262
rect 1602 -2274 1608 -2268
rect 1602 -2280 1608 -2274
rect 1602 -2286 1608 -2280
rect 1602 -2292 1608 -2286
rect 1602 -2298 1608 -2292
rect 1602 -2304 1608 -2298
rect 1602 -2310 1608 -2304
rect 1602 -2316 1608 -2310
rect 1602 -2322 1608 -2316
rect 1602 -2328 1608 -2322
rect 1602 -2334 1608 -2328
rect 1602 -2340 1608 -2334
rect 1602 -2346 1608 -2340
rect 1602 -2352 1608 -2346
rect 1602 -2358 1608 -2352
rect 1602 -2364 1608 -2358
rect 1602 -2370 1608 -2364
rect 1602 -2376 1608 -2370
rect 1602 -2382 1608 -2376
rect 1602 -2388 1608 -2382
rect 1602 -2394 1608 -2388
rect 1602 -2400 1608 -2394
rect 1602 -2406 1608 -2400
rect 1602 -2412 1608 -2406
rect 1602 -2418 1608 -2412
rect 1602 -2424 1608 -2418
rect 1602 -2430 1608 -2424
rect 1602 -2436 1608 -2430
rect 1602 -2442 1608 -2436
rect 1602 -2448 1608 -2442
rect 1602 -2454 1608 -2448
rect 1602 -2460 1608 -2454
rect 1602 -2466 1608 -2460
rect 1602 -2472 1608 -2466
rect 1602 -2478 1608 -2472
rect 1602 -2484 1608 -2478
rect 1602 -2490 1608 -2484
rect 1602 -2496 1608 -2490
rect 1602 -2502 1608 -2496
rect 1602 -2508 1608 -2502
rect 1602 -2514 1608 -2508
rect 1602 -2520 1608 -2514
rect 1602 -2526 1608 -2520
rect 1602 -2532 1608 -2526
rect 1602 -2538 1608 -2532
rect 1602 -2544 1608 -2538
rect 1602 -2550 1608 -2544
rect 1602 -2556 1608 -2550
rect 1602 -2562 1608 -2556
rect 1602 -2568 1608 -2562
rect 1602 -2574 1608 -2568
rect 1602 -2580 1608 -2574
rect 1602 -2586 1608 -2580
rect 1602 -2592 1608 -2586
rect 1602 -2598 1608 -2592
rect 1602 -2604 1608 -2598
rect 1602 -2610 1608 -2604
rect 1602 -2616 1608 -2610
rect 1602 -2622 1608 -2616
rect 1602 -2628 1608 -2622
rect 1602 -2634 1608 -2628
rect 1602 -2640 1608 -2634
rect 1602 -2646 1608 -2640
rect 1602 -2652 1608 -2646
rect 1602 -2658 1608 -2652
rect 1602 -2664 1608 -2658
rect 1602 -2670 1608 -2664
rect 1602 -2676 1608 -2670
rect 1602 -2682 1608 -2676
rect 1602 -2688 1608 -2682
rect 1602 -2694 1608 -2688
rect 1602 -2700 1608 -2694
rect 1602 -2706 1608 -2700
rect 1602 -2712 1608 -2706
rect 1602 -2718 1608 -2712
rect 1602 -2724 1608 -2718
rect 1602 -2730 1608 -2724
rect 1602 -2736 1608 -2730
rect 1602 -2742 1608 -2736
rect 1602 -2748 1608 -2742
rect 1602 -2826 1608 -2820
rect 1602 -2832 1608 -2826
rect 1602 -2838 1608 -2832
rect 1602 -2844 1608 -2838
rect 1602 -2850 1608 -2844
rect 1602 -2856 1608 -2850
rect 1602 -2862 1608 -2856
rect 1602 -2868 1608 -2862
rect 1602 -2874 1608 -2868
rect 1602 -2880 1608 -2874
rect 1602 -2886 1608 -2880
rect 1602 -2892 1608 -2886
rect 1602 -2898 1608 -2892
rect 1602 -2904 1608 -2898
rect 1602 -2910 1608 -2904
rect 1602 -2916 1608 -2910
rect 1602 -2922 1608 -2916
rect 1602 -2928 1608 -2922
rect 1602 -2934 1608 -2928
rect 1602 -2940 1608 -2934
rect 1602 -2946 1608 -2940
rect 1602 -2952 1608 -2946
rect 1602 -2958 1608 -2952
rect 1602 -2964 1608 -2958
rect 1602 -2970 1608 -2964
rect 1602 -2976 1608 -2970
rect 1602 -2982 1608 -2976
rect 1602 -2988 1608 -2982
rect 1602 -2994 1608 -2988
rect 1602 -3000 1608 -2994
rect 1602 -3006 1608 -3000
rect 1602 -3012 1608 -3006
rect 1602 -3018 1608 -3012
rect 1602 -3024 1608 -3018
rect 1602 -3030 1608 -3024
rect 1602 -3036 1608 -3030
rect 1602 -3042 1608 -3036
rect 1602 -3048 1608 -3042
rect 1602 -3054 1608 -3048
rect 1602 -3060 1608 -3054
rect 1602 -3066 1608 -3060
rect 1602 -3072 1608 -3066
rect 1602 -3078 1608 -3072
rect 1602 -3084 1608 -3078
rect 1602 -3090 1608 -3084
rect 1602 -3096 1608 -3090
rect 1602 -3102 1608 -3096
rect 1602 -3108 1608 -3102
rect 1602 -3114 1608 -3108
rect 1602 -3120 1608 -3114
rect 1602 -3126 1608 -3120
rect 1602 -3132 1608 -3126
rect 1602 -3138 1608 -3132
rect 1602 -3144 1608 -3138
rect 1602 -3150 1608 -3144
rect 1602 -3156 1608 -3150
rect 1602 -3162 1608 -3156
rect 1602 -3168 1608 -3162
rect 1602 -3174 1608 -3168
rect 1602 -3180 1608 -3174
rect 1602 -3186 1608 -3180
rect 1602 -3192 1608 -3186
rect 1602 -3198 1608 -3192
rect 1602 -3204 1608 -3198
rect 1602 -3210 1608 -3204
rect 1602 -3216 1608 -3210
rect 1602 -3222 1608 -3216
rect 1602 -3228 1608 -3222
rect 1602 -3234 1608 -3228
rect 1602 -3276 1608 -3270
rect 1602 -3282 1608 -3276
rect 1602 -3288 1608 -3282
rect 1602 -3294 1608 -3288
rect 1602 -3300 1608 -3294
rect 1602 -3306 1608 -3300
rect 1602 -3312 1608 -3306
rect 1602 -3318 1608 -3312
rect 1602 -3324 1608 -3318
rect 1602 -3330 1608 -3324
rect 1602 -3336 1608 -3330
rect 1602 -3342 1608 -3336
rect 1602 -3348 1608 -3342
rect 1602 -3354 1608 -3348
rect 1602 -3360 1608 -3354
rect 1602 -3366 1608 -3360
rect 1602 -3372 1608 -3366
rect 1602 -3378 1608 -3372
rect 1602 -3384 1608 -3378
rect 1602 -3390 1608 -3384
rect 1602 -3396 1608 -3390
rect 1602 -3402 1608 -3396
rect 1602 -3408 1608 -3402
rect 1602 -3414 1608 -3408
rect 1602 -3420 1608 -3414
rect 1602 -3426 1608 -3420
rect 1602 -3432 1608 -3426
rect 1602 -3438 1608 -3432
rect 1602 -3444 1608 -3438
rect 1602 -3450 1608 -3444
rect 1602 -3456 1608 -3450
rect 1608 -1002 1614 -996
rect 1608 -1008 1614 -1002
rect 1608 -1014 1614 -1008
rect 1608 -1020 1614 -1014
rect 1608 -1026 1614 -1020
rect 1608 -1032 1614 -1026
rect 1608 -1038 1614 -1032
rect 1608 -1044 1614 -1038
rect 1608 -1050 1614 -1044
rect 1608 -1056 1614 -1050
rect 1608 -1062 1614 -1056
rect 1608 -1068 1614 -1062
rect 1608 -1074 1614 -1068
rect 1608 -1080 1614 -1074
rect 1608 -1086 1614 -1080
rect 1608 -1092 1614 -1086
rect 1608 -1098 1614 -1092
rect 1608 -1104 1614 -1098
rect 1608 -1110 1614 -1104
rect 1608 -1116 1614 -1110
rect 1608 -1122 1614 -1116
rect 1608 -1128 1614 -1122
rect 1608 -1134 1614 -1128
rect 1608 -1140 1614 -1134
rect 1608 -1146 1614 -1140
rect 1608 -1152 1614 -1146
rect 1608 -1158 1614 -1152
rect 1608 -1164 1614 -1158
rect 1608 -1170 1614 -1164
rect 1608 -1176 1614 -1170
rect 1608 -1182 1614 -1176
rect 1608 -1188 1614 -1182
rect 1608 -1194 1614 -1188
rect 1608 -1200 1614 -1194
rect 1608 -1206 1614 -1200
rect 1608 -1212 1614 -1206
rect 1608 -1218 1614 -1212
rect 1608 -1224 1614 -1218
rect 1608 -1230 1614 -1224
rect 1608 -1236 1614 -1230
rect 1608 -1242 1614 -1236
rect 1608 -1248 1614 -1242
rect 1608 -1254 1614 -1248
rect 1608 -1260 1614 -1254
rect 1608 -1266 1614 -1260
rect 1608 -1272 1614 -1266
rect 1608 -1278 1614 -1272
rect 1608 -1284 1614 -1278
rect 1608 -1290 1614 -1284
rect 1608 -1296 1614 -1290
rect 1608 -1302 1614 -1296
rect 1608 -1308 1614 -1302
rect 1608 -1314 1614 -1308
rect 1608 -1320 1614 -1314
rect 1608 -1326 1614 -1320
rect 1608 -1332 1614 -1326
rect 1608 -1338 1614 -1332
rect 1608 -1344 1614 -1338
rect 1608 -1350 1614 -1344
rect 1608 -1356 1614 -1350
rect 1608 -1362 1614 -1356
rect 1608 -1368 1614 -1362
rect 1608 -1374 1614 -1368
rect 1608 -1380 1614 -1374
rect 1608 -1386 1614 -1380
rect 1608 -1392 1614 -1386
rect 1608 -1398 1614 -1392
rect 1608 -1404 1614 -1398
rect 1608 -1410 1614 -1404
rect 1608 -1416 1614 -1410
rect 1608 -1422 1614 -1416
rect 1608 -1428 1614 -1422
rect 1608 -1434 1614 -1428
rect 1608 -1440 1614 -1434
rect 1608 -1446 1614 -1440
rect 1608 -1452 1614 -1446
rect 1608 -1458 1614 -1452
rect 1608 -1464 1614 -1458
rect 1608 -1470 1614 -1464
rect 1608 -1476 1614 -1470
rect 1608 -1482 1614 -1476
rect 1608 -1488 1614 -1482
rect 1608 -1494 1614 -1488
rect 1608 -1500 1614 -1494
rect 1608 -1506 1614 -1500
rect 1608 -1512 1614 -1506
rect 1608 -1518 1614 -1512
rect 1608 -1524 1614 -1518
rect 1608 -1530 1614 -1524
rect 1608 -1536 1614 -1530
rect 1608 -1542 1614 -1536
rect 1608 -1548 1614 -1542
rect 1608 -1554 1614 -1548
rect 1608 -1560 1614 -1554
rect 1608 -1566 1614 -1560
rect 1608 -1572 1614 -1566
rect 1608 -1578 1614 -1572
rect 1608 -1584 1614 -1578
rect 1608 -1590 1614 -1584
rect 1608 -1596 1614 -1590
rect 1608 -1602 1614 -1596
rect 1608 -1608 1614 -1602
rect 1608 -1614 1614 -1608
rect 1608 -1620 1614 -1614
rect 1608 -1626 1614 -1620
rect 1608 -1632 1614 -1626
rect 1608 -1638 1614 -1632
rect 1608 -1644 1614 -1638
rect 1608 -1650 1614 -1644
rect 1608 -1656 1614 -1650
rect 1608 -1662 1614 -1656
rect 1608 -1668 1614 -1662
rect 1608 -1674 1614 -1668
rect 1608 -1680 1614 -1674
rect 1608 -1686 1614 -1680
rect 1608 -1692 1614 -1686
rect 1608 -1698 1614 -1692
rect 1608 -1704 1614 -1698
rect 1608 -1710 1614 -1704
rect 1608 -1716 1614 -1710
rect 1608 -1722 1614 -1716
rect 1608 -1728 1614 -1722
rect 1608 -1734 1614 -1728
rect 1608 -1740 1614 -1734
rect 1608 -1746 1614 -1740
rect 1608 -1752 1614 -1746
rect 1608 -1758 1614 -1752
rect 1608 -1764 1614 -1758
rect 1608 -1770 1614 -1764
rect 1608 -1776 1614 -1770
rect 1608 -1782 1614 -1776
rect 1608 -1788 1614 -1782
rect 1608 -1794 1614 -1788
rect 1608 -1800 1614 -1794
rect 1608 -1806 1614 -1800
rect 1608 -1812 1614 -1806
rect 1608 -1818 1614 -1812
rect 1608 -1824 1614 -1818
rect 1608 -1830 1614 -1824
rect 1608 -1836 1614 -1830
rect 1608 -1842 1614 -1836
rect 1608 -1848 1614 -1842
rect 1608 -1854 1614 -1848
rect 1608 -1860 1614 -1854
rect 1608 -1866 1614 -1860
rect 1608 -1872 1614 -1866
rect 1608 -1878 1614 -1872
rect 1608 -1884 1614 -1878
rect 1608 -1890 1614 -1884
rect 1608 -1896 1614 -1890
rect 1608 -1902 1614 -1896
rect 1608 -1908 1614 -1902
rect 1608 -1914 1614 -1908
rect 1608 -1920 1614 -1914
rect 1608 -1926 1614 -1920
rect 1608 -1932 1614 -1926
rect 1608 -1938 1614 -1932
rect 1608 -1944 1614 -1938
rect 1608 -1950 1614 -1944
rect 1608 -1956 1614 -1950
rect 1608 -1962 1614 -1956
rect 1608 -1968 1614 -1962
rect 1608 -1974 1614 -1968
rect 1608 -1980 1614 -1974
rect 1608 -1986 1614 -1980
rect 1608 -1992 1614 -1986
rect 1608 -1998 1614 -1992
rect 1608 -2004 1614 -1998
rect 1608 -2010 1614 -2004
rect 1608 -2016 1614 -2010
rect 1608 -2022 1614 -2016
rect 1608 -2028 1614 -2022
rect 1608 -2034 1614 -2028
rect 1608 -2040 1614 -2034
rect 1608 -2046 1614 -2040
rect 1608 -2052 1614 -2046
rect 1608 -2058 1614 -2052
rect 1608 -2130 1614 -2124
rect 1608 -2136 1614 -2130
rect 1608 -2142 1614 -2136
rect 1608 -2148 1614 -2142
rect 1608 -2154 1614 -2148
rect 1608 -2160 1614 -2154
rect 1608 -2166 1614 -2160
rect 1608 -2172 1614 -2166
rect 1608 -2178 1614 -2172
rect 1608 -2184 1614 -2178
rect 1608 -2190 1614 -2184
rect 1608 -2196 1614 -2190
rect 1608 -2202 1614 -2196
rect 1608 -2208 1614 -2202
rect 1608 -2214 1614 -2208
rect 1608 -2220 1614 -2214
rect 1608 -2226 1614 -2220
rect 1608 -2232 1614 -2226
rect 1608 -2238 1614 -2232
rect 1608 -2244 1614 -2238
rect 1608 -2250 1614 -2244
rect 1608 -2256 1614 -2250
rect 1608 -2262 1614 -2256
rect 1608 -2268 1614 -2262
rect 1608 -2274 1614 -2268
rect 1608 -2280 1614 -2274
rect 1608 -2286 1614 -2280
rect 1608 -2292 1614 -2286
rect 1608 -2298 1614 -2292
rect 1608 -2304 1614 -2298
rect 1608 -2310 1614 -2304
rect 1608 -2316 1614 -2310
rect 1608 -2322 1614 -2316
rect 1608 -2328 1614 -2322
rect 1608 -2334 1614 -2328
rect 1608 -2340 1614 -2334
rect 1608 -2346 1614 -2340
rect 1608 -2352 1614 -2346
rect 1608 -2358 1614 -2352
rect 1608 -2364 1614 -2358
rect 1608 -2370 1614 -2364
rect 1608 -2376 1614 -2370
rect 1608 -2382 1614 -2376
rect 1608 -2388 1614 -2382
rect 1608 -2394 1614 -2388
rect 1608 -2400 1614 -2394
rect 1608 -2406 1614 -2400
rect 1608 -2412 1614 -2406
rect 1608 -2418 1614 -2412
rect 1608 -2424 1614 -2418
rect 1608 -2430 1614 -2424
rect 1608 -2436 1614 -2430
rect 1608 -2442 1614 -2436
rect 1608 -2448 1614 -2442
rect 1608 -2454 1614 -2448
rect 1608 -2460 1614 -2454
rect 1608 -2466 1614 -2460
rect 1608 -2472 1614 -2466
rect 1608 -2478 1614 -2472
rect 1608 -2484 1614 -2478
rect 1608 -2490 1614 -2484
rect 1608 -2496 1614 -2490
rect 1608 -2502 1614 -2496
rect 1608 -2508 1614 -2502
rect 1608 -2514 1614 -2508
rect 1608 -2520 1614 -2514
rect 1608 -2526 1614 -2520
rect 1608 -2532 1614 -2526
rect 1608 -2538 1614 -2532
rect 1608 -2544 1614 -2538
rect 1608 -2550 1614 -2544
rect 1608 -2556 1614 -2550
rect 1608 -2562 1614 -2556
rect 1608 -2568 1614 -2562
rect 1608 -2574 1614 -2568
rect 1608 -2580 1614 -2574
rect 1608 -2586 1614 -2580
rect 1608 -2592 1614 -2586
rect 1608 -2598 1614 -2592
rect 1608 -2604 1614 -2598
rect 1608 -2610 1614 -2604
rect 1608 -2616 1614 -2610
rect 1608 -2622 1614 -2616
rect 1608 -2628 1614 -2622
rect 1608 -2634 1614 -2628
rect 1608 -2640 1614 -2634
rect 1608 -2646 1614 -2640
rect 1608 -2652 1614 -2646
rect 1608 -2658 1614 -2652
rect 1608 -2664 1614 -2658
rect 1608 -2670 1614 -2664
rect 1608 -2676 1614 -2670
rect 1608 -2682 1614 -2676
rect 1608 -2688 1614 -2682
rect 1608 -2694 1614 -2688
rect 1608 -2700 1614 -2694
rect 1608 -2706 1614 -2700
rect 1608 -2712 1614 -2706
rect 1608 -2718 1614 -2712
rect 1608 -2724 1614 -2718
rect 1608 -2730 1614 -2724
rect 1608 -2736 1614 -2730
rect 1608 -2742 1614 -2736
rect 1608 -2820 1614 -2814
rect 1608 -2826 1614 -2820
rect 1608 -2832 1614 -2826
rect 1608 -2838 1614 -2832
rect 1608 -2844 1614 -2838
rect 1608 -2850 1614 -2844
rect 1608 -2856 1614 -2850
rect 1608 -2862 1614 -2856
rect 1608 -2868 1614 -2862
rect 1608 -2874 1614 -2868
rect 1608 -2880 1614 -2874
rect 1608 -2886 1614 -2880
rect 1608 -2892 1614 -2886
rect 1608 -2898 1614 -2892
rect 1608 -2904 1614 -2898
rect 1608 -2910 1614 -2904
rect 1608 -2916 1614 -2910
rect 1608 -2922 1614 -2916
rect 1608 -2928 1614 -2922
rect 1608 -2934 1614 -2928
rect 1608 -2940 1614 -2934
rect 1608 -2946 1614 -2940
rect 1608 -2952 1614 -2946
rect 1608 -2958 1614 -2952
rect 1608 -2964 1614 -2958
rect 1608 -2970 1614 -2964
rect 1608 -2976 1614 -2970
rect 1608 -2982 1614 -2976
rect 1608 -2988 1614 -2982
rect 1608 -2994 1614 -2988
rect 1608 -3000 1614 -2994
rect 1608 -3006 1614 -3000
rect 1608 -3012 1614 -3006
rect 1608 -3018 1614 -3012
rect 1608 -3024 1614 -3018
rect 1608 -3030 1614 -3024
rect 1608 -3036 1614 -3030
rect 1608 -3042 1614 -3036
rect 1608 -3048 1614 -3042
rect 1608 -3054 1614 -3048
rect 1608 -3060 1614 -3054
rect 1608 -3066 1614 -3060
rect 1608 -3072 1614 -3066
rect 1608 -3078 1614 -3072
rect 1608 -3084 1614 -3078
rect 1608 -3090 1614 -3084
rect 1608 -3096 1614 -3090
rect 1608 -3102 1614 -3096
rect 1608 -3108 1614 -3102
rect 1608 -3114 1614 -3108
rect 1608 -3120 1614 -3114
rect 1608 -3126 1614 -3120
rect 1608 -3132 1614 -3126
rect 1608 -3138 1614 -3132
rect 1608 -3144 1614 -3138
rect 1608 -3150 1614 -3144
rect 1608 -3156 1614 -3150
rect 1608 -3162 1614 -3156
rect 1608 -3168 1614 -3162
rect 1608 -3174 1614 -3168
rect 1608 -3180 1614 -3174
rect 1608 -3186 1614 -3180
rect 1608 -3192 1614 -3186
rect 1608 -3198 1614 -3192
rect 1608 -3204 1614 -3198
rect 1608 -3210 1614 -3204
rect 1608 -3216 1614 -3210
rect 1608 -3222 1614 -3216
rect 1608 -3228 1614 -3222
rect 1608 -3234 1614 -3228
rect 1608 -3276 1614 -3270
rect 1608 -3282 1614 -3276
rect 1608 -3288 1614 -3282
rect 1608 -3294 1614 -3288
rect 1608 -3300 1614 -3294
rect 1608 -3306 1614 -3300
rect 1608 -3312 1614 -3306
rect 1608 -3318 1614 -3312
rect 1608 -3324 1614 -3318
rect 1608 -3330 1614 -3324
rect 1608 -3336 1614 -3330
rect 1608 -3342 1614 -3336
rect 1608 -3348 1614 -3342
rect 1608 -3354 1614 -3348
rect 1608 -3360 1614 -3354
rect 1608 -3366 1614 -3360
rect 1608 -3372 1614 -3366
rect 1608 -3378 1614 -3372
rect 1608 -3384 1614 -3378
rect 1608 -3390 1614 -3384
rect 1608 -3396 1614 -3390
rect 1608 -3402 1614 -3396
rect 1608 -3408 1614 -3402
rect 1608 -3414 1614 -3408
rect 1608 -3420 1614 -3414
rect 1608 -3426 1614 -3420
rect 1608 -3432 1614 -3426
rect 1608 -3438 1614 -3432
rect 1608 -3444 1614 -3438
rect 1608 -3450 1614 -3444
rect 1608 -3456 1614 -3450
rect 1614 -996 1620 -990
rect 1614 -1002 1620 -996
rect 1614 -1008 1620 -1002
rect 1614 -1014 1620 -1008
rect 1614 -1020 1620 -1014
rect 1614 -1026 1620 -1020
rect 1614 -1032 1620 -1026
rect 1614 -1038 1620 -1032
rect 1614 -1044 1620 -1038
rect 1614 -1050 1620 -1044
rect 1614 -1056 1620 -1050
rect 1614 -1062 1620 -1056
rect 1614 -1068 1620 -1062
rect 1614 -1074 1620 -1068
rect 1614 -1080 1620 -1074
rect 1614 -1086 1620 -1080
rect 1614 -1092 1620 -1086
rect 1614 -1098 1620 -1092
rect 1614 -1104 1620 -1098
rect 1614 -1110 1620 -1104
rect 1614 -1116 1620 -1110
rect 1614 -1122 1620 -1116
rect 1614 -1128 1620 -1122
rect 1614 -1134 1620 -1128
rect 1614 -1140 1620 -1134
rect 1614 -1146 1620 -1140
rect 1614 -1152 1620 -1146
rect 1614 -1158 1620 -1152
rect 1614 -1164 1620 -1158
rect 1614 -1170 1620 -1164
rect 1614 -1176 1620 -1170
rect 1614 -1182 1620 -1176
rect 1614 -1188 1620 -1182
rect 1614 -1194 1620 -1188
rect 1614 -1200 1620 -1194
rect 1614 -1206 1620 -1200
rect 1614 -1212 1620 -1206
rect 1614 -1218 1620 -1212
rect 1614 -1224 1620 -1218
rect 1614 -1230 1620 -1224
rect 1614 -1236 1620 -1230
rect 1614 -1242 1620 -1236
rect 1614 -1248 1620 -1242
rect 1614 -1254 1620 -1248
rect 1614 -1260 1620 -1254
rect 1614 -1266 1620 -1260
rect 1614 -1272 1620 -1266
rect 1614 -1278 1620 -1272
rect 1614 -1284 1620 -1278
rect 1614 -1290 1620 -1284
rect 1614 -1296 1620 -1290
rect 1614 -1302 1620 -1296
rect 1614 -1308 1620 -1302
rect 1614 -1314 1620 -1308
rect 1614 -1320 1620 -1314
rect 1614 -1326 1620 -1320
rect 1614 -1332 1620 -1326
rect 1614 -1338 1620 -1332
rect 1614 -1344 1620 -1338
rect 1614 -1350 1620 -1344
rect 1614 -1356 1620 -1350
rect 1614 -1362 1620 -1356
rect 1614 -1368 1620 -1362
rect 1614 -1374 1620 -1368
rect 1614 -1380 1620 -1374
rect 1614 -1386 1620 -1380
rect 1614 -1392 1620 -1386
rect 1614 -1398 1620 -1392
rect 1614 -1404 1620 -1398
rect 1614 -1410 1620 -1404
rect 1614 -1416 1620 -1410
rect 1614 -1422 1620 -1416
rect 1614 -1428 1620 -1422
rect 1614 -1434 1620 -1428
rect 1614 -1440 1620 -1434
rect 1614 -1446 1620 -1440
rect 1614 -1452 1620 -1446
rect 1614 -1458 1620 -1452
rect 1614 -1464 1620 -1458
rect 1614 -1470 1620 -1464
rect 1614 -1476 1620 -1470
rect 1614 -1482 1620 -1476
rect 1614 -1488 1620 -1482
rect 1614 -1494 1620 -1488
rect 1614 -1500 1620 -1494
rect 1614 -1506 1620 -1500
rect 1614 -1512 1620 -1506
rect 1614 -1518 1620 -1512
rect 1614 -1524 1620 -1518
rect 1614 -1530 1620 -1524
rect 1614 -1536 1620 -1530
rect 1614 -1542 1620 -1536
rect 1614 -1548 1620 -1542
rect 1614 -1554 1620 -1548
rect 1614 -1560 1620 -1554
rect 1614 -1566 1620 -1560
rect 1614 -1572 1620 -1566
rect 1614 -1578 1620 -1572
rect 1614 -1584 1620 -1578
rect 1614 -1590 1620 -1584
rect 1614 -1596 1620 -1590
rect 1614 -1602 1620 -1596
rect 1614 -1608 1620 -1602
rect 1614 -1614 1620 -1608
rect 1614 -1620 1620 -1614
rect 1614 -1626 1620 -1620
rect 1614 -1632 1620 -1626
rect 1614 -1638 1620 -1632
rect 1614 -1644 1620 -1638
rect 1614 -1650 1620 -1644
rect 1614 -1656 1620 -1650
rect 1614 -1662 1620 -1656
rect 1614 -1668 1620 -1662
rect 1614 -1674 1620 -1668
rect 1614 -1680 1620 -1674
rect 1614 -1686 1620 -1680
rect 1614 -1692 1620 -1686
rect 1614 -1698 1620 -1692
rect 1614 -1704 1620 -1698
rect 1614 -1710 1620 -1704
rect 1614 -1716 1620 -1710
rect 1614 -1722 1620 -1716
rect 1614 -1728 1620 -1722
rect 1614 -1734 1620 -1728
rect 1614 -1740 1620 -1734
rect 1614 -1746 1620 -1740
rect 1614 -1752 1620 -1746
rect 1614 -1758 1620 -1752
rect 1614 -1764 1620 -1758
rect 1614 -1770 1620 -1764
rect 1614 -1776 1620 -1770
rect 1614 -1782 1620 -1776
rect 1614 -1788 1620 -1782
rect 1614 -1794 1620 -1788
rect 1614 -1800 1620 -1794
rect 1614 -1806 1620 -1800
rect 1614 -1812 1620 -1806
rect 1614 -1818 1620 -1812
rect 1614 -1824 1620 -1818
rect 1614 -1830 1620 -1824
rect 1614 -1836 1620 -1830
rect 1614 -1842 1620 -1836
rect 1614 -1848 1620 -1842
rect 1614 -1854 1620 -1848
rect 1614 -1860 1620 -1854
rect 1614 -1866 1620 -1860
rect 1614 -1872 1620 -1866
rect 1614 -1878 1620 -1872
rect 1614 -1884 1620 -1878
rect 1614 -1890 1620 -1884
rect 1614 -1896 1620 -1890
rect 1614 -1902 1620 -1896
rect 1614 -1908 1620 -1902
rect 1614 -1914 1620 -1908
rect 1614 -1920 1620 -1914
rect 1614 -1926 1620 -1920
rect 1614 -1932 1620 -1926
rect 1614 -1938 1620 -1932
rect 1614 -1944 1620 -1938
rect 1614 -1950 1620 -1944
rect 1614 -1956 1620 -1950
rect 1614 -1962 1620 -1956
rect 1614 -1968 1620 -1962
rect 1614 -1974 1620 -1968
rect 1614 -1980 1620 -1974
rect 1614 -1986 1620 -1980
rect 1614 -1992 1620 -1986
rect 1614 -1998 1620 -1992
rect 1614 -2004 1620 -1998
rect 1614 -2010 1620 -2004
rect 1614 -2016 1620 -2010
rect 1614 -2022 1620 -2016
rect 1614 -2028 1620 -2022
rect 1614 -2034 1620 -2028
rect 1614 -2040 1620 -2034
rect 1614 -2046 1620 -2040
rect 1614 -2052 1620 -2046
rect 1614 -2124 1620 -2118
rect 1614 -2130 1620 -2124
rect 1614 -2136 1620 -2130
rect 1614 -2142 1620 -2136
rect 1614 -2148 1620 -2142
rect 1614 -2154 1620 -2148
rect 1614 -2160 1620 -2154
rect 1614 -2166 1620 -2160
rect 1614 -2172 1620 -2166
rect 1614 -2178 1620 -2172
rect 1614 -2184 1620 -2178
rect 1614 -2190 1620 -2184
rect 1614 -2196 1620 -2190
rect 1614 -2202 1620 -2196
rect 1614 -2208 1620 -2202
rect 1614 -2214 1620 -2208
rect 1614 -2220 1620 -2214
rect 1614 -2226 1620 -2220
rect 1614 -2232 1620 -2226
rect 1614 -2238 1620 -2232
rect 1614 -2244 1620 -2238
rect 1614 -2250 1620 -2244
rect 1614 -2256 1620 -2250
rect 1614 -2262 1620 -2256
rect 1614 -2268 1620 -2262
rect 1614 -2274 1620 -2268
rect 1614 -2280 1620 -2274
rect 1614 -2286 1620 -2280
rect 1614 -2292 1620 -2286
rect 1614 -2298 1620 -2292
rect 1614 -2304 1620 -2298
rect 1614 -2310 1620 -2304
rect 1614 -2316 1620 -2310
rect 1614 -2322 1620 -2316
rect 1614 -2328 1620 -2322
rect 1614 -2334 1620 -2328
rect 1614 -2340 1620 -2334
rect 1614 -2346 1620 -2340
rect 1614 -2352 1620 -2346
rect 1614 -2358 1620 -2352
rect 1614 -2364 1620 -2358
rect 1614 -2370 1620 -2364
rect 1614 -2376 1620 -2370
rect 1614 -2382 1620 -2376
rect 1614 -2388 1620 -2382
rect 1614 -2394 1620 -2388
rect 1614 -2400 1620 -2394
rect 1614 -2406 1620 -2400
rect 1614 -2412 1620 -2406
rect 1614 -2418 1620 -2412
rect 1614 -2424 1620 -2418
rect 1614 -2430 1620 -2424
rect 1614 -2436 1620 -2430
rect 1614 -2442 1620 -2436
rect 1614 -2448 1620 -2442
rect 1614 -2454 1620 -2448
rect 1614 -2460 1620 -2454
rect 1614 -2466 1620 -2460
rect 1614 -2472 1620 -2466
rect 1614 -2478 1620 -2472
rect 1614 -2484 1620 -2478
rect 1614 -2490 1620 -2484
rect 1614 -2496 1620 -2490
rect 1614 -2502 1620 -2496
rect 1614 -2508 1620 -2502
rect 1614 -2514 1620 -2508
rect 1614 -2520 1620 -2514
rect 1614 -2526 1620 -2520
rect 1614 -2532 1620 -2526
rect 1614 -2538 1620 -2532
rect 1614 -2544 1620 -2538
rect 1614 -2550 1620 -2544
rect 1614 -2556 1620 -2550
rect 1614 -2562 1620 -2556
rect 1614 -2568 1620 -2562
rect 1614 -2574 1620 -2568
rect 1614 -2580 1620 -2574
rect 1614 -2586 1620 -2580
rect 1614 -2592 1620 -2586
rect 1614 -2598 1620 -2592
rect 1614 -2604 1620 -2598
rect 1614 -2610 1620 -2604
rect 1614 -2616 1620 -2610
rect 1614 -2622 1620 -2616
rect 1614 -2628 1620 -2622
rect 1614 -2634 1620 -2628
rect 1614 -2640 1620 -2634
rect 1614 -2646 1620 -2640
rect 1614 -2652 1620 -2646
rect 1614 -2658 1620 -2652
rect 1614 -2664 1620 -2658
rect 1614 -2670 1620 -2664
rect 1614 -2676 1620 -2670
rect 1614 -2682 1620 -2676
rect 1614 -2688 1620 -2682
rect 1614 -2694 1620 -2688
rect 1614 -2700 1620 -2694
rect 1614 -2706 1620 -2700
rect 1614 -2712 1620 -2706
rect 1614 -2718 1620 -2712
rect 1614 -2724 1620 -2718
rect 1614 -2730 1620 -2724
rect 1614 -2736 1620 -2730
rect 1614 -2820 1620 -2814
rect 1614 -2826 1620 -2820
rect 1614 -2832 1620 -2826
rect 1614 -2838 1620 -2832
rect 1614 -2844 1620 -2838
rect 1614 -2850 1620 -2844
rect 1614 -2856 1620 -2850
rect 1614 -2862 1620 -2856
rect 1614 -2868 1620 -2862
rect 1614 -2874 1620 -2868
rect 1614 -2880 1620 -2874
rect 1614 -2886 1620 -2880
rect 1614 -2892 1620 -2886
rect 1614 -2898 1620 -2892
rect 1614 -2904 1620 -2898
rect 1614 -2910 1620 -2904
rect 1614 -2916 1620 -2910
rect 1614 -2922 1620 -2916
rect 1614 -2928 1620 -2922
rect 1614 -2934 1620 -2928
rect 1614 -2940 1620 -2934
rect 1614 -2946 1620 -2940
rect 1614 -2952 1620 -2946
rect 1614 -2958 1620 -2952
rect 1614 -2964 1620 -2958
rect 1614 -2970 1620 -2964
rect 1614 -2976 1620 -2970
rect 1614 -2982 1620 -2976
rect 1614 -2988 1620 -2982
rect 1614 -2994 1620 -2988
rect 1614 -3000 1620 -2994
rect 1614 -3006 1620 -3000
rect 1614 -3012 1620 -3006
rect 1614 -3018 1620 -3012
rect 1614 -3024 1620 -3018
rect 1614 -3030 1620 -3024
rect 1614 -3036 1620 -3030
rect 1614 -3042 1620 -3036
rect 1614 -3048 1620 -3042
rect 1614 -3054 1620 -3048
rect 1614 -3060 1620 -3054
rect 1614 -3066 1620 -3060
rect 1614 -3072 1620 -3066
rect 1614 -3078 1620 -3072
rect 1614 -3084 1620 -3078
rect 1614 -3090 1620 -3084
rect 1614 -3096 1620 -3090
rect 1614 -3102 1620 -3096
rect 1614 -3108 1620 -3102
rect 1614 -3114 1620 -3108
rect 1614 -3120 1620 -3114
rect 1614 -3126 1620 -3120
rect 1614 -3132 1620 -3126
rect 1614 -3138 1620 -3132
rect 1614 -3144 1620 -3138
rect 1614 -3150 1620 -3144
rect 1614 -3156 1620 -3150
rect 1614 -3162 1620 -3156
rect 1614 -3168 1620 -3162
rect 1614 -3174 1620 -3168
rect 1614 -3180 1620 -3174
rect 1614 -3186 1620 -3180
rect 1614 -3192 1620 -3186
rect 1614 -3198 1620 -3192
rect 1614 -3204 1620 -3198
rect 1614 -3210 1620 -3204
rect 1614 -3216 1620 -3210
rect 1614 -3222 1620 -3216
rect 1614 -3228 1620 -3222
rect 1614 -3234 1620 -3228
rect 1614 -3276 1620 -3270
rect 1614 -3282 1620 -3276
rect 1614 -3288 1620 -3282
rect 1614 -3294 1620 -3288
rect 1614 -3300 1620 -3294
rect 1614 -3306 1620 -3300
rect 1614 -3312 1620 -3306
rect 1614 -3318 1620 -3312
rect 1614 -3324 1620 -3318
rect 1614 -3330 1620 -3324
rect 1614 -3336 1620 -3330
rect 1614 -3342 1620 -3336
rect 1614 -3348 1620 -3342
rect 1614 -3354 1620 -3348
rect 1614 -3360 1620 -3354
rect 1614 -3366 1620 -3360
rect 1614 -3372 1620 -3366
rect 1614 -3378 1620 -3372
rect 1614 -3384 1620 -3378
rect 1614 -3390 1620 -3384
rect 1614 -3396 1620 -3390
rect 1614 -3402 1620 -3396
rect 1614 -3408 1620 -3402
rect 1614 -3414 1620 -3408
rect 1614 -3420 1620 -3414
rect 1614 -3426 1620 -3420
rect 1614 -3432 1620 -3426
rect 1614 -3438 1620 -3432
rect 1614 -3444 1620 -3438
rect 1614 -3450 1620 -3444
rect 1614 -3456 1620 -3450
rect 1620 -984 1626 -978
rect 1620 -990 1626 -984
rect 1620 -996 1626 -990
rect 1620 -1002 1626 -996
rect 1620 -1008 1626 -1002
rect 1620 -1014 1626 -1008
rect 1620 -1020 1626 -1014
rect 1620 -1026 1626 -1020
rect 1620 -1032 1626 -1026
rect 1620 -1038 1626 -1032
rect 1620 -1044 1626 -1038
rect 1620 -1050 1626 -1044
rect 1620 -1056 1626 -1050
rect 1620 -1062 1626 -1056
rect 1620 -1068 1626 -1062
rect 1620 -1074 1626 -1068
rect 1620 -1080 1626 -1074
rect 1620 -1086 1626 -1080
rect 1620 -1092 1626 -1086
rect 1620 -1098 1626 -1092
rect 1620 -1104 1626 -1098
rect 1620 -1110 1626 -1104
rect 1620 -1116 1626 -1110
rect 1620 -1122 1626 -1116
rect 1620 -1128 1626 -1122
rect 1620 -1134 1626 -1128
rect 1620 -1140 1626 -1134
rect 1620 -1146 1626 -1140
rect 1620 -1152 1626 -1146
rect 1620 -1158 1626 -1152
rect 1620 -1164 1626 -1158
rect 1620 -1170 1626 -1164
rect 1620 -1176 1626 -1170
rect 1620 -1182 1626 -1176
rect 1620 -1188 1626 -1182
rect 1620 -1194 1626 -1188
rect 1620 -1200 1626 -1194
rect 1620 -1206 1626 -1200
rect 1620 -1212 1626 -1206
rect 1620 -1218 1626 -1212
rect 1620 -1224 1626 -1218
rect 1620 -1230 1626 -1224
rect 1620 -1236 1626 -1230
rect 1620 -1242 1626 -1236
rect 1620 -1248 1626 -1242
rect 1620 -1254 1626 -1248
rect 1620 -1260 1626 -1254
rect 1620 -1266 1626 -1260
rect 1620 -1272 1626 -1266
rect 1620 -1278 1626 -1272
rect 1620 -1284 1626 -1278
rect 1620 -1290 1626 -1284
rect 1620 -1296 1626 -1290
rect 1620 -1302 1626 -1296
rect 1620 -1308 1626 -1302
rect 1620 -1314 1626 -1308
rect 1620 -1320 1626 -1314
rect 1620 -1326 1626 -1320
rect 1620 -1332 1626 -1326
rect 1620 -1338 1626 -1332
rect 1620 -1344 1626 -1338
rect 1620 -1350 1626 -1344
rect 1620 -1356 1626 -1350
rect 1620 -1362 1626 -1356
rect 1620 -1368 1626 -1362
rect 1620 -1374 1626 -1368
rect 1620 -1380 1626 -1374
rect 1620 -1386 1626 -1380
rect 1620 -1392 1626 -1386
rect 1620 -1398 1626 -1392
rect 1620 -1404 1626 -1398
rect 1620 -1410 1626 -1404
rect 1620 -1416 1626 -1410
rect 1620 -1422 1626 -1416
rect 1620 -1428 1626 -1422
rect 1620 -1434 1626 -1428
rect 1620 -1440 1626 -1434
rect 1620 -1446 1626 -1440
rect 1620 -1452 1626 -1446
rect 1620 -1458 1626 -1452
rect 1620 -1464 1626 -1458
rect 1620 -1470 1626 -1464
rect 1620 -1476 1626 -1470
rect 1620 -1482 1626 -1476
rect 1620 -1488 1626 -1482
rect 1620 -1494 1626 -1488
rect 1620 -1500 1626 -1494
rect 1620 -1506 1626 -1500
rect 1620 -1512 1626 -1506
rect 1620 -1518 1626 -1512
rect 1620 -1524 1626 -1518
rect 1620 -1530 1626 -1524
rect 1620 -1536 1626 -1530
rect 1620 -1542 1626 -1536
rect 1620 -1548 1626 -1542
rect 1620 -1554 1626 -1548
rect 1620 -1560 1626 -1554
rect 1620 -1566 1626 -1560
rect 1620 -1572 1626 -1566
rect 1620 -1578 1626 -1572
rect 1620 -1584 1626 -1578
rect 1620 -1590 1626 -1584
rect 1620 -1596 1626 -1590
rect 1620 -1602 1626 -1596
rect 1620 -1608 1626 -1602
rect 1620 -1614 1626 -1608
rect 1620 -1620 1626 -1614
rect 1620 -1626 1626 -1620
rect 1620 -1632 1626 -1626
rect 1620 -1638 1626 -1632
rect 1620 -1644 1626 -1638
rect 1620 -1650 1626 -1644
rect 1620 -1656 1626 -1650
rect 1620 -1662 1626 -1656
rect 1620 -1668 1626 -1662
rect 1620 -1674 1626 -1668
rect 1620 -1680 1626 -1674
rect 1620 -1686 1626 -1680
rect 1620 -1692 1626 -1686
rect 1620 -1698 1626 -1692
rect 1620 -1704 1626 -1698
rect 1620 -1710 1626 -1704
rect 1620 -1716 1626 -1710
rect 1620 -1722 1626 -1716
rect 1620 -1728 1626 -1722
rect 1620 -1734 1626 -1728
rect 1620 -1740 1626 -1734
rect 1620 -1746 1626 -1740
rect 1620 -1752 1626 -1746
rect 1620 -1758 1626 -1752
rect 1620 -1764 1626 -1758
rect 1620 -1770 1626 -1764
rect 1620 -1776 1626 -1770
rect 1620 -1782 1626 -1776
rect 1620 -1788 1626 -1782
rect 1620 -1794 1626 -1788
rect 1620 -1800 1626 -1794
rect 1620 -1806 1626 -1800
rect 1620 -1812 1626 -1806
rect 1620 -1818 1626 -1812
rect 1620 -1824 1626 -1818
rect 1620 -1830 1626 -1824
rect 1620 -1836 1626 -1830
rect 1620 -1842 1626 -1836
rect 1620 -1848 1626 -1842
rect 1620 -1854 1626 -1848
rect 1620 -1860 1626 -1854
rect 1620 -1866 1626 -1860
rect 1620 -1872 1626 -1866
rect 1620 -1878 1626 -1872
rect 1620 -1884 1626 -1878
rect 1620 -1890 1626 -1884
rect 1620 -1896 1626 -1890
rect 1620 -1902 1626 -1896
rect 1620 -1908 1626 -1902
rect 1620 -1914 1626 -1908
rect 1620 -1920 1626 -1914
rect 1620 -1926 1626 -1920
rect 1620 -1932 1626 -1926
rect 1620 -1938 1626 -1932
rect 1620 -1944 1626 -1938
rect 1620 -1950 1626 -1944
rect 1620 -1956 1626 -1950
rect 1620 -1962 1626 -1956
rect 1620 -1968 1626 -1962
rect 1620 -1974 1626 -1968
rect 1620 -1980 1626 -1974
rect 1620 -1986 1626 -1980
rect 1620 -1992 1626 -1986
rect 1620 -1998 1626 -1992
rect 1620 -2004 1626 -1998
rect 1620 -2010 1626 -2004
rect 1620 -2016 1626 -2010
rect 1620 -2022 1626 -2016
rect 1620 -2028 1626 -2022
rect 1620 -2034 1626 -2028
rect 1620 -2040 1626 -2034
rect 1620 -2046 1626 -2040
rect 1620 -2118 1626 -2112
rect 1620 -2124 1626 -2118
rect 1620 -2130 1626 -2124
rect 1620 -2136 1626 -2130
rect 1620 -2142 1626 -2136
rect 1620 -2148 1626 -2142
rect 1620 -2154 1626 -2148
rect 1620 -2160 1626 -2154
rect 1620 -2166 1626 -2160
rect 1620 -2172 1626 -2166
rect 1620 -2178 1626 -2172
rect 1620 -2184 1626 -2178
rect 1620 -2190 1626 -2184
rect 1620 -2196 1626 -2190
rect 1620 -2202 1626 -2196
rect 1620 -2208 1626 -2202
rect 1620 -2214 1626 -2208
rect 1620 -2220 1626 -2214
rect 1620 -2226 1626 -2220
rect 1620 -2232 1626 -2226
rect 1620 -2238 1626 -2232
rect 1620 -2244 1626 -2238
rect 1620 -2250 1626 -2244
rect 1620 -2256 1626 -2250
rect 1620 -2262 1626 -2256
rect 1620 -2268 1626 -2262
rect 1620 -2274 1626 -2268
rect 1620 -2280 1626 -2274
rect 1620 -2286 1626 -2280
rect 1620 -2292 1626 -2286
rect 1620 -2298 1626 -2292
rect 1620 -2304 1626 -2298
rect 1620 -2310 1626 -2304
rect 1620 -2316 1626 -2310
rect 1620 -2322 1626 -2316
rect 1620 -2328 1626 -2322
rect 1620 -2334 1626 -2328
rect 1620 -2340 1626 -2334
rect 1620 -2346 1626 -2340
rect 1620 -2352 1626 -2346
rect 1620 -2358 1626 -2352
rect 1620 -2364 1626 -2358
rect 1620 -2370 1626 -2364
rect 1620 -2376 1626 -2370
rect 1620 -2382 1626 -2376
rect 1620 -2388 1626 -2382
rect 1620 -2394 1626 -2388
rect 1620 -2400 1626 -2394
rect 1620 -2406 1626 -2400
rect 1620 -2412 1626 -2406
rect 1620 -2418 1626 -2412
rect 1620 -2424 1626 -2418
rect 1620 -2430 1626 -2424
rect 1620 -2436 1626 -2430
rect 1620 -2442 1626 -2436
rect 1620 -2448 1626 -2442
rect 1620 -2454 1626 -2448
rect 1620 -2460 1626 -2454
rect 1620 -2466 1626 -2460
rect 1620 -2472 1626 -2466
rect 1620 -2478 1626 -2472
rect 1620 -2484 1626 -2478
rect 1620 -2490 1626 -2484
rect 1620 -2496 1626 -2490
rect 1620 -2502 1626 -2496
rect 1620 -2508 1626 -2502
rect 1620 -2514 1626 -2508
rect 1620 -2520 1626 -2514
rect 1620 -2526 1626 -2520
rect 1620 -2532 1626 -2526
rect 1620 -2538 1626 -2532
rect 1620 -2544 1626 -2538
rect 1620 -2550 1626 -2544
rect 1620 -2556 1626 -2550
rect 1620 -2562 1626 -2556
rect 1620 -2568 1626 -2562
rect 1620 -2574 1626 -2568
rect 1620 -2580 1626 -2574
rect 1620 -2586 1626 -2580
rect 1620 -2592 1626 -2586
rect 1620 -2598 1626 -2592
rect 1620 -2604 1626 -2598
rect 1620 -2610 1626 -2604
rect 1620 -2616 1626 -2610
rect 1620 -2622 1626 -2616
rect 1620 -2628 1626 -2622
rect 1620 -2634 1626 -2628
rect 1620 -2640 1626 -2634
rect 1620 -2646 1626 -2640
rect 1620 -2652 1626 -2646
rect 1620 -2658 1626 -2652
rect 1620 -2664 1626 -2658
rect 1620 -2670 1626 -2664
rect 1620 -2676 1626 -2670
rect 1620 -2682 1626 -2676
rect 1620 -2688 1626 -2682
rect 1620 -2694 1626 -2688
rect 1620 -2700 1626 -2694
rect 1620 -2706 1626 -2700
rect 1620 -2712 1626 -2706
rect 1620 -2718 1626 -2712
rect 1620 -2724 1626 -2718
rect 1620 -2730 1626 -2724
rect 1620 -2736 1626 -2730
rect 1620 -2814 1626 -2808
rect 1620 -2820 1626 -2814
rect 1620 -2826 1626 -2820
rect 1620 -2832 1626 -2826
rect 1620 -2838 1626 -2832
rect 1620 -2844 1626 -2838
rect 1620 -2850 1626 -2844
rect 1620 -2856 1626 -2850
rect 1620 -2862 1626 -2856
rect 1620 -2868 1626 -2862
rect 1620 -2874 1626 -2868
rect 1620 -2880 1626 -2874
rect 1620 -2886 1626 -2880
rect 1620 -2892 1626 -2886
rect 1620 -2898 1626 -2892
rect 1620 -2904 1626 -2898
rect 1620 -2910 1626 -2904
rect 1620 -2916 1626 -2910
rect 1620 -2922 1626 -2916
rect 1620 -2928 1626 -2922
rect 1620 -2934 1626 -2928
rect 1620 -2940 1626 -2934
rect 1620 -2946 1626 -2940
rect 1620 -2952 1626 -2946
rect 1620 -2958 1626 -2952
rect 1620 -2964 1626 -2958
rect 1620 -2970 1626 -2964
rect 1620 -2976 1626 -2970
rect 1620 -2982 1626 -2976
rect 1620 -2988 1626 -2982
rect 1620 -2994 1626 -2988
rect 1620 -3000 1626 -2994
rect 1620 -3006 1626 -3000
rect 1620 -3012 1626 -3006
rect 1620 -3018 1626 -3012
rect 1620 -3024 1626 -3018
rect 1620 -3030 1626 -3024
rect 1620 -3036 1626 -3030
rect 1620 -3042 1626 -3036
rect 1620 -3048 1626 -3042
rect 1620 -3054 1626 -3048
rect 1620 -3060 1626 -3054
rect 1620 -3066 1626 -3060
rect 1620 -3072 1626 -3066
rect 1620 -3078 1626 -3072
rect 1620 -3084 1626 -3078
rect 1620 -3090 1626 -3084
rect 1620 -3096 1626 -3090
rect 1620 -3102 1626 -3096
rect 1620 -3108 1626 -3102
rect 1620 -3114 1626 -3108
rect 1620 -3120 1626 -3114
rect 1620 -3126 1626 -3120
rect 1620 -3132 1626 -3126
rect 1620 -3138 1626 -3132
rect 1620 -3144 1626 -3138
rect 1620 -3150 1626 -3144
rect 1620 -3156 1626 -3150
rect 1620 -3162 1626 -3156
rect 1620 -3168 1626 -3162
rect 1620 -3174 1626 -3168
rect 1620 -3180 1626 -3174
rect 1620 -3186 1626 -3180
rect 1620 -3192 1626 -3186
rect 1620 -3198 1626 -3192
rect 1620 -3204 1626 -3198
rect 1620 -3210 1626 -3204
rect 1620 -3216 1626 -3210
rect 1620 -3222 1626 -3216
rect 1620 -3228 1626 -3222
rect 1620 -3234 1626 -3228
rect 1620 -3276 1626 -3270
rect 1620 -3282 1626 -3276
rect 1620 -3288 1626 -3282
rect 1620 -3294 1626 -3288
rect 1620 -3300 1626 -3294
rect 1620 -3306 1626 -3300
rect 1620 -3312 1626 -3306
rect 1620 -3318 1626 -3312
rect 1620 -3324 1626 -3318
rect 1620 -3330 1626 -3324
rect 1620 -3336 1626 -3330
rect 1620 -3342 1626 -3336
rect 1620 -3348 1626 -3342
rect 1620 -3354 1626 -3348
rect 1620 -3360 1626 -3354
rect 1620 -3366 1626 -3360
rect 1620 -3372 1626 -3366
rect 1620 -3378 1626 -3372
rect 1620 -3384 1626 -3378
rect 1620 -3390 1626 -3384
rect 1620 -3396 1626 -3390
rect 1620 -3402 1626 -3396
rect 1620 -3408 1626 -3402
rect 1620 -3414 1626 -3408
rect 1620 -3420 1626 -3414
rect 1620 -3426 1626 -3420
rect 1620 -3432 1626 -3426
rect 1620 -3438 1626 -3432
rect 1620 -3444 1626 -3438
rect 1620 -3450 1626 -3444
rect 1626 -978 1632 -972
rect 1626 -984 1632 -978
rect 1626 -990 1632 -984
rect 1626 -996 1632 -990
rect 1626 -1002 1632 -996
rect 1626 -1008 1632 -1002
rect 1626 -1014 1632 -1008
rect 1626 -1020 1632 -1014
rect 1626 -1026 1632 -1020
rect 1626 -1032 1632 -1026
rect 1626 -1038 1632 -1032
rect 1626 -1044 1632 -1038
rect 1626 -1050 1632 -1044
rect 1626 -1056 1632 -1050
rect 1626 -1062 1632 -1056
rect 1626 -1068 1632 -1062
rect 1626 -1074 1632 -1068
rect 1626 -1080 1632 -1074
rect 1626 -1086 1632 -1080
rect 1626 -1092 1632 -1086
rect 1626 -1098 1632 -1092
rect 1626 -1104 1632 -1098
rect 1626 -1110 1632 -1104
rect 1626 -1116 1632 -1110
rect 1626 -1122 1632 -1116
rect 1626 -1128 1632 -1122
rect 1626 -1134 1632 -1128
rect 1626 -1140 1632 -1134
rect 1626 -1146 1632 -1140
rect 1626 -1152 1632 -1146
rect 1626 -1158 1632 -1152
rect 1626 -1164 1632 -1158
rect 1626 -1170 1632 -1164
rect 1626 -1176 1632 -1170
rect 1626 -1182 1632 -1176
rect 1626 -1188 1632 -1182
rect 1626 -1194 1632 -1188
rect 1626 -1200 1632 -1194
rect 1626 -1206 1632 -1200
rect 1626 -1212 1632 -1206
rect 1626 -1218 1632 -1212
rect 1626 -1224 1632 -1218
rect 1626 -1230 1632 -1224
rect 1626 -1236 1632 -1230
rect 1626 -1242 1632 -1236
rect 1626 -1248 1632 -1242
rect 1626 -1254 1632 -1248
rect 1626 -1260 1632 -1254
rect 1626 -1266 1632 -1260
rect 1626 -1272 1632 -1266
rect 1626 -1278 1632 -1272
rect 1626 -1284 1632 -1278
rect 1626 -1290 1632 -1284
rect 1626 -1296 1632 -1290
rect 1626 -1302 1632 -1296
rect 1626 -1308 1632 -1302
rect 1626 -1314 1632 -1308
rect 1626 -1320 1632 -1314
rect 1626 -1326 1632 -1320
rect 1626 -1332 1632 -1326
rect 1626 -1338 1632 -1332
rect 1626 -1344 1632 -1338
rect 1626 -1350 1632 -1344
rect 1626 -1356 1632 -1350
rect 1626 -1362 1632 -1356
rect 1626 -1368 1632 -1362
rect 1626 -1374 1632 -1368
rect 1626 -1380 1632 -1374
rect 1626 -1386 1632 -1380
rect 1626 -1392 1632 -1386
rect 1626 -1398 1632 -1392
rect 1626 -1404 1632 -1398
rect 1626 -1410 1632 -1404
rect 1626 -1416 1632 -1410
rect 1626 -1422 1632 -1416
rect 1626 -1428 1632 -1422
rect 1626 -1434 1632 -1428
rect 1626 -1440 1632 -1434
rect 1626 -1446 1632 -1440
rect 1626 -1452 1632 -1446
rect 1626 -1458 1632 -1452
rect 1626 -1464 1632 -1458
rect 1626 -1470 1632 -1464
rect 1626 -1476 1632 -1470
rect 1626 -1482 1632 -1476
rect 1626 -1488 1632 -1482
rect 1626 -1494 1632 -1488
rect 1626 -1500 1632 -1494
rect 1626 -1506 1632 -1500
rect 1626 -1512 1632 -1506
rect 1626 -1518 1632 -1512
rect 1626 -1524 1632 -1518
rect 1626 -1530 1632 -1524
rect 1626 -1536 1632 -1530
rect 1626 -1542 1632 -1536
rect 1626 -1548 1632 -1542
rect 1626 -1554 1632 -1548
rect 1626 -1560 1632 -1554
rect 1626 -1566 1632 -1560
rect 1626 -1572 1632 -1566
rect 1626 -1578 1632 -1572
rect 1626 -1584 1632 -1578
rect 1626 -1590 1632 -1584
rect 1626 -1596 1632 -1590
rect 1626 -1602 1632 -1596
rect 1626 -1608 1632 -1602
rect 1626 -1614 1632 -1608
rect 1626 -1620 1632 -1614
rect 1626 -1626 1632 -1620
rect 1626 -1632 1632 -1626
rect 1626 -1638 1632 -1632
rect 1626 -1644 1632 -1638
rect 1626 -1650 1632 -1644
rect 1626 -1656 1632 -1650
rect 1626 -1662 1632 -1656
rect 1626 -1668 1632 -1662
rect 1626 -1674 1632 -1668
rect 1626 -1680 1632 -1674
rect 1626 -1686 1632 -1680
rect 1626 -1692 1632 -1686
rect 1626 -1698 1632 -1692
rect 1626 -1704 1632 -1698
rect 1626 -1710 1632 -1704
rect 1626 -1716 1632 -1710
rect 1626 -1722 1632 -1716
rect 1626 -1728 1632 -1722
rect 1626 -1734 1632 -1728
rect 1626 -1740 1632 -1734
rect 1626 -1746 1632 -1740
rect 1626 -1752 1632 -1746
rect 1626 -1758 1632 -1752
rect 1626 -1764 1632 -1758
rect 1626 -1770 1632 -1764
rect 1626 -1776 1632 -1770
rect 1626 -1782 1632 -1776
rect 1626 -1788 1632 -1782
rect 1626 -1794 1632 -1788
rect 1626 -1800 1632 -1794
rect 1626 -1806 1632 -1800
rect 1626 -1812 1632 -1806
rect 1626 -1818 1632 -1812
rect 1626 -1824 1632 -1818
rect 1626 -1830 1632 -1824
rect 1626 -1836 1632 -1830
rect 1626 -1842 1632 -1836
rect 1626 -1848 1632 -1842
rect 1626 -1854 1632 -1848
rect 1626 -1860 1632 -1854
rect 1626 -1866 1632 -1860
rect 1626 -1872 1632 -1866
rect 1626 -1878 1632 -1872
rect 1626 -1884 1632 -1878
rect 1626 -1890 1632 -1884
rect 1626 -1896 1632 -1890
rect 1626 -1902 1632 -1896
rect 1626 -1908 1632 -1902
rect 1626 -1914 1632 -1908
rect 1626 -1920 1632 -1914
rect 1626 -1926 1632 -1920
rect 1626 -1932 1632 -1926
rect 1626 -1938 1632 -1932
rect 1626 -1944 1632 -1938
rect 1626 -1950 1632 -1944
rect 1626 -1956 1632 -1950
rect 1626 -1962 1632 -1956
rect 1626 -1968 1632 -1962
rect 1626 -1974 1632 -1968
rect 1626 -1980 1632 -1974
rect 1626 -1986 1632 -1980
rect 1626 -1992 1632 -1986
rect 1626 -1998 1632 -1992
rect 1626 -2004 1632 -1998
rect 1626 -2010 1632 -2004
rect 1626 -2016 1632 -2010
rect 1626 -2022 1632 -2016
rect 1626 -2028 1632 -2022
rect 1626 -2034 1632 -2028
rect 1626 -2040 1632 -2034
rect 1626 -2112 1632 -2106
rect 1626 -2118 1632 -2112
rect 1626 -2124 1632 -2118
rect 1626 -2130 1632 -2124
rect 1626 -2136 1632 -2130
rect 1626 -2142 1632 -2136
rect 1626 -2148 1632 -2142
rect 1626 -2154 1632 -2148
rect 1626 -2160 1632 -2154
rect 1626 -2166 1632 -2160
rect 1626 -2172 1632 -2166
rect 1626 -2178 1632 -2172
rect 1626 -2184 1632 -2178
rect 1626 -2190 1632 -2184
rect 1626 -2196 1632 -2190
rect 1626 -2202 1632 -2196
rect 1626 -2208 1632 -2202
rect 1626 -2214 1632 -2208
rect 1626 -2220 1632 -2214
rect 1626 -2226 1632 -2220
rect 1626 -2232 1632 -2226
rect 1626 -2238 1632 -2232
rect 1626 -2244 1632 -2238
rect 1626 -2250 1632 -2244
rect 1626 -2256 1632 -2250
rect 1626 -2262 1632 -2256
rect 1626 -2268 1632 -2262
rect 1626 -2274 1632 -2268
rect 1626 -2280 1632 -2274
rect 1626 -2286 1632 -2280
rect 1626 -2292 1632 -2286
rect 1626 -2298 1632 -2292
rect 1626 -2304 1632 -2298
rect 1626 -2310 1632 -2304
rect 1626 -2316 1632 -2310
rect 1626 -2322 1632 -2316
rect 1626 -2328 1632 -2322
rect 1626 -2334 1632 -2328
rect 1626 -2340 1632 -2334
rect 1626 -2346 1632 -2340
rect 1626 -2352 1632 -2346
rect 1626 -2358 1632 -2352
rect 1626 -2364 1632 -2358
rect 1626 -2370 1632 -2364
rect 1626 -2376 1632 -2370
rect 1626 -2382 1632 -2376
rect 1626 -2388 1632 -2382
rect 1626 -2394 1632 -2388
rect 1626 -2400 1632 -2394
rect 1626 -2406 1632 -2400
rect 1626 -2412 1632 -2406
rect 1626 -2418 1632 -2412
rect 1626 -2424 1632 -2418
rect 1626 -2430 1632 -2424
rect 1626 -2436 1632 -2430
rect 1626 -2442 1632 -2436
rect 1626 -2448 1632 -2442
rect 1626 -2454 1632 -2448
rect 1626 -2460 1632 -2454
rect 1626 -2466 1632 -2460
rect 1626 -2472 1632 -2466
rect 1626 -2478 1632 -2472
rect 1626 -2484 1632 -2478
rect 1626 -2490 1632 -2484
rect 1626 -2496 1632 -2490
rect 1626 -2502 1632 -2496
rect 1626 -2508 1632 -2502
rect 1626 -2514 1632 -2508
rect 1626 -2520 1632 -2514
rect 1626 -2526 1632 -2520
rect 1626 -2532 1632 -2526
rect 1626 -2538 1632 -2532
rect 1626 -2544 1632 -2538
rect 1626 -2550 1632 -2544
rect 1626 -2556 1632 -2550
rect 1626 -2562 1632 -2556
rect 1626 -2568 1632 -2562
rect 1626 -2574 1632 -2568
rect 1626 -2580 1632 -2574
rect 1626 -2586 1632 -2580
rect 1626 -2592 1632 -2586
rect 1626 -2598 1632 -2592
rect 1626 -2604 1632 -2598
rect 1626 -2610 1632 -2604
rect 1626 -2616 1632 -2610
rect 1626 -2622 1632 -2616
rect 1626 -2628 1632 -2622
rect 1626 -2634 1632 -2628
rect 1626 -2640 1632 -2634
rect 1626 -2646 1632 -2640
rect 1626 -2652 1632 -2646
rect 1626 -2658 1632 -2652
rect 1626 -2664 1632 -2658
rect 1626 -2670 1632 -2664
rect 1626 -2676 1632 -2670
rect 1626 -2682 1632 -2676
rect 1626 -2688 1632 -2682
rect 1626 -2694 1632 -2688
rect 1626 -2700 1632 -2694
rect 1626 -2706 1632 -2700
rect 1626 -2712 1632 -2706
rect 1626 -2718 1632 -2712
rect 1626 -2724 1632 -2718
rect 1626 -2730 1632 -2724
rect 1626 -2808 1632 -2802
rect 1626 -2814 1632 -2808
rect 1626 -2820 1632 -2814
rect 1626 -2826 1632 -2820
rect 1626 -2832 1632 -2826
rect 1626 -2838 1632 -2832
rect 1626 -2844 1632 -2838
rect 1626 -2850 1632 -2844
rect 1626 -2856 1632 -2850
rect 1626 -2862 1632 -2856
rect 1626 -2868 1632 -2862
rect 1626 -2874 1632 -2868
rect 1626 -2880 1632 -2874
rect 1626 -2886 1632 -2880
rect 1626 -2892 1632 -2886
rect 1626 -2898 1632 -2892
rect 1626 -2904 1632 -2898
rect 1626 -2910 1632 -2904
rect 1626 -2916 1632 -2910
rect 1626 -2922 1632 -2916
rect 1626 -2928 1632 -2922
rect 1626 -2934 1632 -2928
rect 1626 -2940 1632 -2934
rect 1626 -2946 1632 -2940
rect 1626 -2952 1632 -2946
rect 1626 -2958 1632 -2952
rect 1626 -2964 1632 -2958
rect 1626 -2970 1632 -2964
rect 1626 -2976 1632 -2970
rect 1626 -2982 1632 -2976
rect 1626 -2988 1632 -2982
rect 1626 -2994 1632 -2988
rect 1626 -3000 1632 -2994
rect 1626 -3006 1632 -3000
rect 1626 -3012 1632 -3006
rect 1626 -3018 1632 -3012
rect 1626 -3024 1632 -3018
rect 1626 -3030 1632 -3024
rect 1626 -3036 1632 -3030
rect 1626 -3042 1632 -3036
rect 1626 -3048 1632 -3042
rect 1626 -3054 1632 -3048
rect 1626 -3060 1632 -3054
rect 1626 -3066 1632 -3060
rect 1626 -3072 1632 -3066
rect 1626 -3078 1632 -3072
rect 1626 -3084 1632 -3078
rect 1626 -3090 1632 -3084
rect 1626 -3096 1632 -3090
rect 1626 -3102 1632 -3096
rect 1626 -3108 1632 -3102
rect 1626 -3114 1632 -3108
rect 1626 -3120 1632 -3114
rect 1626 -3126 1632 -3120
rect 1626 -3132 1632 -3126
rect 1626 -3138 1632 -3132
rect 1626 -3144 1632 -3138
rect 1626 -3150 1632 -3144
rect 1626 -3156 1632 -3150
rect 1626 -3162 1632 -3156
rect 1626 -3168 1632 -3162
rect 1626 -3174 1632 -3168
rect 1626 -3180 1632 -3174
rect 1626 -3186 1632 -3180
rect 1626 -3192 1632 -3186
rect 1626 -3198 1632 -3192
rect 1626 -3204 1632 -3198
rect 1626 -3210 1632 -3204
rect 1626 -3216 1632 -3210
rect 1626 -3222 1632 -3216
rect 1626 -3228 1632 -3222
rect 1626 -3234 1632 -3228
rect 1626 -3276 1632 -3270
rect 1626 -3282 1632 -3276
rect 1626 -3288 1632 -3282
rect 1626 -3294 1632 -3288
rect 1626 -3300 1632 -3294
rect 1626 -3306 1632 -3300
rect 1626 -3312 1632 -3306
rect 1626 -3318 1632 -3312
rect 1626 -3324 1632 -3318
rect 1626 -3330 1632 -3324
rect 1626 -3336 1632 -3330
rect 1626 -3342 1632 -3336
rect 1626 -3348 1632 -3342
rect 1626 -3354 1632 -3348
rect 1626 -3360 1632 -3354
rect 1626 -3366 1632 -3360
rect 1626 -3372 1632 -3366
rect 1626 -3378 1632 -3372
rect 1626 -3384 1632 -3378
rect 1626 -3390 1632 -3384
rect 1626 -3396 1632 -3390
rect 1626 -3402 1632 -3396
rect 1626 -3408 1632 -3402
rect 1626 -3414 1632 -3408
rect 1626 -3420 1632 -3414
rect 1626 -3426 1632 -3420
rect 1626 -3432 1632 -3426
rect 1626 -3438 1632 -3432
rect 1626 -3444 1632 -3438
rect 1626 -3450 1632 -3444
rect 1632 -966 1638 -960
rect 1632 -972 1638 -966
rect 1632 -978 1638 -972
rect 1632 -984 1638 -978
rect 1632 -990 1638 -984
rect 1632 -996 1638 -990
rect 1632 -1002 1638 -996
rect 1632 -1008 1638 -1002
rect 1632 -1014 1638 -1008
rect 1632 -1020 1638 -1014
rect 1632 -1026 1638 -1020
rect 1632 -1032 1638 -1026
rect 1632 -1038 1638 -1032
rect 1632 -1044 1638 -1038
rect 1632 -1050 1638 -1044
rect 1632 -1056 1638 -1050
rect 1632 -1062 1638 -1056
rect 1632 -1068 1638 -1062
rect 1632 -1074 1638 -1068
rect 1632 -1080 1638 -1074
rect 1632 -1086 1638 -1080
rect 1632 -1092 1638 -1086
rect 1632 -1098 1638 -1092
rect 1632 -1104 1638 -1098
rect 1632 -1110 1638 -1104
rect 1632 -1116 1638 -1110
rect 1632 -1122 1638 -1116
rect 1632 -1128 1638 -1122
rect 1632 -1134 1638 -1128
rect 1632 -1140 1638 -1134
rect 1632 -1146 1638 -1140
rect 1632 -1152 1638 -1146
rect 1632 -1158 1638 -1152
rect 1632 -1164 1638 -1158
rect 1632 -1170 1638 -1164
rect 1632 -1176 1638 -1170
rect 1632 -1182 1638 -1176
rect 1632 -1188 1638 -1182
rect 1632 -1194 1638 -1188
rect 1632 -1200 1638 -1194
rect 1632 -1206 1638 -1200
rect 1632 -1212 1638 -1206
rect 1632 -1218 1638 -1212
rect 1632 -1224 1638 -1218
rect 1632 -1230 1638 -1224
rect 1632 -1236 1638 -1230
rect 1632 -1242 1638 -1236
rect 1632 -1248 1638 -1242
rect 1632 -1254 1638 -1248
rect 1632 -1260 1638 -1254
rect 1632 -1266 1638 -1260
rect 1632 -1272 1638 -1266
rect 1632 -1278 1638 -1272
rect 1632 -1284 1638 -1278
rect 1632 -1290 1638 -1284
rect 1632 -1296 1638 -1290
rect 1632 -1302 1638 -1296
rect 1632 -1308 1638 -1302
rect 1632 -1314 1638 -1308
rect 1632 -1320 1638 -1314
rect 1632 -1326 1638 -1320
rect 1632 -1332 1638 -1326
rect 1632 -1338 1638 -1332
rect 1632 -1344 1638 -1338
rect 1632 -1350 1638 -1344
rect 1632 -1356 1638 -1350
rect 1632 -1362 1638 -1356
rect 1632 -1368 1638 -1362
rect 1632 -1374 1638 -1368
rect 1632 -1380 1638 -1374
rect 1632 -1386 1638 -1380
rect 1632 -1392 1638 -1386
rect 1632 -1398 1638 -1392
rect 1632 -1404 1638 -1398
rect 1632 -1410 1638 -1404
rect 1632 -1416 1638 -1410
rect 1632 -1422 1638 -1416
rect 1632 -1428 1638 -1422
rect 1632 -1434 1638 -1428
rect 1632 -1440 1638 -1434
rect 1632 -1446 1638 -1440
rect 1632 -1452 1638 -1446
rect 1632 -1458 1638 -1452
rect 1632 -1464 1638 -1458
rect 1632 -1470 1638 -1464
rect 1632 -1476 1638 -1470
rect 1632 -1482 1638 -1476
rect 1632 -1488 1638 -1482
rect 1632 -1494 1638 -1488
rect 1632 -1500 1638 -1494
rect 1632 -1506 1638 -1500
rect 1632 -1512 1638 -1506
rect 1632 -1518 1638 -1512
rect 1632 -1524 1638 -1518
rect 1632 -1530 1638 -1524
rect 1632 -1536 1638 -1530
rect 1632 -1542 1638 -1536
rect 1632 -1548 1638 -1542
rect 1632 -1554 1638 -1548
rect 1632 -1560 1638 -1554
rect 1632 -1566 1638 -1560
rect 1632 -1572 1638 -1566
rect 1632 -1578 1638 -1572
rect 1632 -1584 1638 -1578
rect 1632 -1590 1638 -1584
rect 1632 -1596 1638 -1590
rect 1632 -1602 1638 -1596
rect 1632 -1608 1638 -1602
rect 1632 -1614 1638 -1608
rect 1632 -1620 1638 -1614
rect 1632 -1626 1638 -1620
rect 1632 -1632 1638 -1626
rect 1632 -1638 1638 -1632
rect 1632 -1644 1638 -1638
rect 1632 -1650 1638 -1644
rect 1632 -1656 1638 -1650
rect 1632 -1662 1638 -1656
rect 1632 -1668 1638 -1662
rect 1632 -1674 1638 -1668
rect 1632 -1680 1638 -1674
rect 1632 -1686 1638 -1680
rect 1632 -1692 1638 -1686
rect 1632 -1698 1638 -1692
rect 1632 -1704 1638 -1698
rect 1632 -1710 1638 -1704
rect 1632 -1716 1638 -1710
rect 1632 -1722 1638 -1716
rect 1632 -1728 1638 -1722
rect 1632 -1734 1638 -1728
rect 1632 -1740 1638 -1734
rect 1632 -1746 1638 -1740
rect 1632 -1752 1638 -1746
rect 1632 -1758 1638 -1752
rect 1632 -1764 1638 -1758
rect 1632 -1770 1638 -1764
rect 1632 -1776 1638 -1770
rect 1632 -1782 1638 -1776
rect 1632 -1788 1638 -1782
rect 1632 -1794 1638 -1788
rect 1632 -1800 1638 -1794
rect 1632 -1806 1638 -1800
rect 1632 -1812 1638 -1806
rect 1632 -1818 1638 -1812
rect 1632 -1824 1638 -1818
rect 1632 -1830 1638 -1824
rect 1632 -1836 1638 -1830
rect 1632 -1842 1638 -1836
rect 1632 -1848 1638 -1842
rect 1632 -1854 1638 -1848
rect 1632 -1860 1638 -1854
rect 1632 -1866 1638 -1860
rect 1632 -1872 1638 -1866
rect 1632 -1878 1638 -1872
rect 1632 -1884 1638 -1878
rect 1632 -1890 1638 -1884
rect 1632 -1896 1638 -1890
rect 1632 -1902 1638 -1896
rect 1632 -1908 1638 -1902
rect 1632 -1914 1638 -1908
rect 1632 -1920 1638 -1914
rect 1632 -1926 1638 -1920
rect 1632 -1932 1638 -1926
rect 1632 -1938 1638 -1932
rect 1632 -1944 1638 -1938
rect 1632 -1950 1638 -1944
rect 1632 -1956 1638 -1950
rect 1632 -1962 1638 -1956
rect 1632 -1968 1638 -1962
rect 1632 -1974 1638 -1968
rect 1632 -1980 1638 -1974
rect 1632 -1986 1638 -1980
rect 1632 -1992 1638 -1986
rect 1632 -1998 1638 -1992
rect 1632 -2004 1638 -1998
rect 1632 -2010 1638 -2004
rect 1632 -2016 1638 -2010
rect 1632 -2022 1638 -2016
rect 1632 -2028 1638 -2022
rect 1632 -2106 1638 -2100
rect 1632 -2112 1638 -2106
rect 1632 -2118 1638 -2112
rect 1632 -2124 1638 -2118
rect 1632 -2130 1638 -2124
rect 1632 -2136 1638 -2130
rect 1632 -2142 1638 -2136
rect 1632 -2148 1638 -2142
rect 1632 -2154 1638 -2148
rect 1632 -2160 1638 -2154
rect 1632 -2166 1638 -2160
rect 1632 -2172 1638 -2166
rect 1632 -2178 1638 -2172
rect 1632 -2184 1638 -2178
rect 1632 -2190 1638 -2184
rect 1632 -2196 1638 -2190
rect 1632 -2202 1638 -2196
rect 1632 -2208 1638 -2202
rect 1632 -2214 1638 -2208
rect 1632 -2220 1638 -2214
rect 1632 -2226 1638 -2220
rect 1632 -2232 1638 -2226
rect 1632 -2238 1638 -2232
rect 1632 -2244 1638 -2238
rect 1632 -2250 1638 -2244
rect 1632 -2256 1638 -2250
rect 1632 -2262 1638 -2256
rect 1632 -2268 1638 -2262
rect 1632 -2274 1638 -2268
rect 1632 -2280 1638 -2274
rect 1632 -2286 1638 -2280
rect 1632 -2292 1638 -2286
rect 1632 -2298 1638 -2292
rect 1632 -2304 1638 -2298
rect 1632 -2310 1638 -2304
rect 1632 -2316 1638 -2310
rect 1632 -2322 1638 -2316
rect 1632 -2328 1638 -2322
rect 1632 -2334 1638 -2328
rect 1632 -2340 1638 -2334
rect 1632 -2346 1638 -2340
rect 1632 -2352 1638 -2346
rect 1632 -2358 1638 -2352
rect 1632 -2364 1638 -2358
rect 1632 -2370 1638 -2364
rect 1632 -2376 1638 -2370
rect 1632 -2382 1638 -2376
rect 1632 -2388 1638 -2382
rect 1632 -2394 1638 -2388
rect 1632 -2400 1638 -2394
rect 1632 -2406 1638 -2400
rect 1632 -2412 1638 -2406
rect 1632 -2418 1638 -2412
rect 1632 -2424 1638 -2418
rect 1632 -2430 1638 -2424
rect 1632 -2436 1638 -2430
rect 1632 -2442 1638 -2436
rect 1632 -2448 1638 -2442
rect 1632 -2454 1638 -2448
rect 1632 -2460 1638 -2454
rect 1632 -2466 1638 -2460
rect 1632 -2472 1638 -2466
rect 1632 -2478 1638 -2472
rect 1632 -2484 1638 -2478
rect 1632 -2490 1638 -2484
rect 1632 -2496 1638 -2490
rect 1632 -2502 1638 -2496
rect 1632 -2508 1638 -2502
rect 1632 -2514 1638 -2508
rect 1632 -2520 1638 -2514
rect 1632 -2526 1638 -2520
rect 1632 -2532 1638 -2526
rect 1632 -2538 1638 -2532
rect 1632 -2544 1638 -2538
rect 1632 -2550 1638 -2544
rect 1632 -2556 1638 -2550
rect 1632 -2562 1638 -2556
rect 1632 -2568 1638 -2562
rect 1632 -2574 1638 -2568
rect 1632 -2580 1638 -2574
rect 1632 -2586 1638 -2580
rect 1632 -2592 1638 -2586
rect 1632 -2598 1638 -2592
rect 1632 -2604 1638 -2598
rect 1632 -2610 1638 -2604
rect 1632 -2616 1638 -2610
rect 1632 -2622 1638 -2616
rect 1632 -2628 1638 -2622
rect 1632 -2634 1638 -2628
rect 1632 -2640 1638 -2634
rect 1632 -2646 1638 -2640
rect 1632 -2652 1638 -2646
rect 1632 -2658 1638 -2652
rect 1632 -2664 1638 -2658
rect 1632 -2670 1638 -2664
rect 1632 -2676 1638 -2670
rect 1632 -2682 1638 -2676
rect 1632 -2688 1638 -2682
rect 1632 -2694 1638 -2688
rect 1632 -2700 1638 -2694
rect 1632 -2706 1638 -2700
rect 1632 -2712 1638 -2706
rect 1632 -2718 1638 -2712
rect 1632 -2724 1638 -2718
rect 1632 -2730 1638 -2724
rect 1632 -2808 1638 -2802
rect 1632 -2814 1638 -2808
rect 1632 -2820 1638 -2814
rect 1632 -2826 1638 -2820
rect 1632 -2832 1638 -2826
rect 1632 -2838 1638 -2832
rect 1632 -2844 1638 -2838
rect 1632 -2850 1638 -2844
rect 1632 -2856 1638 -2850
rect 1632 -2862 1638 -2856
rect 1632 -2868 1638 -2862
rect 1632 -2874 1638 -2868
rect 1632 -2880 1638 -2874
rect 1632 -2886 1638 -2880
rect 1632 -2892 1638 -2886
rect 1632 -2898 1638 -2892
rect 1632 -2904 1638 -2898
rect 1632 -2910 1638 -2904
rect 1632 -2916 1638 -2910
rect 1632 -2922 1638 -2916
rect 1632 -2928 1638 -2922
rect 1632 -2934 1638 -2928
rect 1632 -2940 1638 -2934
rect 1632 -2946 1638 -2940
rect 1632 -2952 1638 -2946
rect 1632 -2958 1638 -2952
rect 1632 -2964 1638 -2958
rect 1632 -2970 1638 -2964
rect 1632 -2976 1638 -2970
rect 1632 -2982 1638 -2976
rect 1632 -2988 1638 -2982
rect 1632 -2994 1638 -2988
rect 1632 -3000 1638 -2994
rect 1632 -3006 1638 -3000
rect 1632 -3012 1638 -3006
rect 1632 -3018 1638 -3012
rect 1632 -3024 1638 -3018
rect 1632 -3030 1638 -3024
rect 1632 -3036 1638 -3030
rect 1632 -3042 1638 -3036
rect 1632 -3048 1638 -3042
rect 1632 -3054 1638 -3048
rect 1632 -3060 1638 -3054
rect 1632 -3066 1638 -3060
rect 1632 -3072 1638 -3066
rect 1632 -3078 1638 -3072
rect 1632 -3084 1638 -3078
rect 1632 -3090 1638 -3084
rect 1632 -3096 1638 -3090
rect 1632 -3102 1638 -3096
rect 1632 -3108 1638 -3102
rect 1632 -3114 1638 -3108
rect 1632 -3120 1638 -3114
rect 1632 -3126 1638 -3120
rect 1632 -3132 1638 -3126
rect 1632 -3138 1638 -3132
rect 1632 -3144 1638 -3138
rect 1632 -3150 1638 -3144
rect 1632 -3156 1638 -3150
rect 1632 -3162 1638 -3156
rect 1632 -3168 1638 -3162
rect 1632 -3174 1638 -3168
rect 1632 -3180 1638 -3174
rect 1632 -3186 1638 -3180
rect 1632 -3192 1638 -3186
rect 1632 -3198 1638 -3192
rect 1632 -3204 1638 -3198
rect 1632 -3210 1638 -3204
rect 1632 -3216 1638 -3210
rect 1632 -3222 1638 -3216
rect 1632 -3228 1638 -3222
rect 1632 -3234 1638 -3228
rect 1632 -3276 1638 -3270
rect 1632 -3282 1638 -3276
rect 1632 -3288 1638 -3282
rect 1632 -3294 1638 -3288
rect 1632 -3300 1638 -3294
rect 1632 -3306 1638 -3300
rect 1632 -3312 1638 -3306
rect 1632 -3318 1638 -3312
rect 1632 -3324 1638 -3318
rect 1632 -3330 1638 -3324
rect 1632 -3336 1638 -3330
rect 1632 -3342 1638 -3336
rect 1632 -3348 1638 -3342
rect 1632 -3354 1638 -3348
rect 1632 -3360 1638 -3354
rect 1632 -3366 1638 -3360
rect 1632 -3372 1638 -3366
rect 1632 -3378 1638 -3372
rect 1632 -3384 1638 -3378
rect 1632 -3390 1638 -3384
rect 1632 -3396 1638 -3390
rect 1632 -3402 1638 -3396
rect 1632 -3408 1638 -3402
rect 1632 -3414 1638 -3408
rect 1632 -3420 1638 -3414
rect 1632 -3426 1638 -3420
rect 1632 -3432 1638 -3426
rect 1632 -3438 1638 -3432
rect 1632 -3444 1638 -3438
rect 1632 -3450 1638 -3444
rect 1638 -954 1644 -948
rect 1638 -960 1644 -954
rect 1638 -966 1644 -960
rect 1638 -972 1644 -966
rect 1638 -978 1644 -972
rect 1638 -984 1644 -978
rect 1638 -990 1644 -984
rect 1638 -996 1644 -990
rect 1638 -1002 1644 -996
rect 1638 -1008 1644 -1002
rect 1638 -1014 1644 -1008
rect 1638 -1020 1644 -1014
rect 1638 -1026 1644 -1020
rect 1638 -1032 1644 -1026
rect 1638 -1038 1644 -1032
rect 1638 -1044 1644 -1038
rect 1638 -1050 1644 -1044
rect 1638 -1056 1644 -1050
rect 1638 -1062 1644 -1056
rect 1638 -1068 1644 -1062
rect 1638 -1074 1644 -1068
rect 1638 -1080 1644 -1074
rect 1638 -1086 1644 -1080
rect 1638 -1092 1644 -1086
rect 1638 -1098 1644 -1092
rect 1638 -1104 1644 -1098
rect 1638 -1110 1644 -1104
rect 1638 -1116 1644 -1110
rect 1638 -1122 1644 -1116
rect 1638 -1128 1644 -1122
rect 1638 -1134 1644 -1128
rect 1638 -1140 1644 -1134
rect 1638 -1146 1644 -1140
rect 1638 -1152 1644 -1146
rect 1638 -1158 1644 -1152
rect 1638 -1164 1644 -1158
rect 1638 -1170 1644 -1164
rect 1638 -1176 1644 -1170
rect 1638 -1182 1644 -1176
rect 1638 -1188 1644 -1182
rect 1638 -1194 1644 -1188
rect 1638 -1200 1644 -1194
rect 1638 -1206 1644 -1200
rect 1638 -1212 1644 -1206
rect 1638 -1218 1644 -1212
rect 1638 -1224 1644 -1218
rect 1638 -1230 1644 -1224
rect 1638 -1236 1644 -1230
rect 1638 -1242 1644 -1236
rect 1638 -1248 1644 -1242
rect 1638 -1254 1644 -1248
rect 1638 -1260 1644 -1254
rect 1638 -1266 1644 -1260
rect 1638 -1272 1644 -1266
rect 1638 -1278 1644 -1272
rect 1638 -1284 1644 -1278
rect 1638 -1290 1644 -1284
rect 1638 -1296 1644 -1290
rect 1638 -1302 1644 -1296
rect 1638 -1308 1644 -1302
rect 1638 -1314 1644 -1308
rect 1638 -1320 1644 -1314
rect 1638 -1326 1644 -1320
rect 1638 -1332 1644 -1326
rect 1638 -1338 1644 -1332
rect 1638 -1344 1644 -1338
rect 1638 -1350 1644 -1344
rect 1638 -1356 1644 -1350
rect 1638 -1362 1644 -1356
rect 1638 -1368 1644 -1362
rect 1638 -1374 1644 -1368
rect 1638 -1380 1644 -1374
rect 1638 -1386 1644 -1380
rect 1638 -1392 1644 -1386
rect 1638 -1398 1644 -1392
rect 1638 -1404 1644 -1398
rect 1638 -1410 1644 -1404
rect 1638 -1416 1644 -1410
rect 1638 -1422 1644 -1416
rect 1638 -1428 1644 -1422
rect 1638 -1434 1644 -1428
rect 1638 -1440 1644 -1434
rect 1638 -1446 1644 -1440
rect 1638 -1452 1644 -1446
rect 1638 -1458 1644 -1452
rect 1638 -1464 1644 -1458
rect 1638 -1470 1644 -1464
rect 1638 -1476 1644 -1470
rect 1638 -1482 1644 -1476
rect 1638 -1488 1644 -1482
rect 1638 -1494 1644 -1488
rect 1638 -1500 1644 -1494
rect 1638 -1506 1644 -1500
rect 1638 -1512 1644 -1506
rect 1638 -1518 1644 -1512
rect 1638 -1524 1644 -1518
rect 1638 -1530 1644 -1524
rect 1638 -1536 1644 -1530
rect 1638 -1542 1644 -1536
rect 1638 -1548 1644 -1542
rect 1638 -1554 1644 -1548
rect 1638 -1560 1644 -1554
rect 1638 -1566 1644 -1560
rect 1638 -1572 1644 -1566
rect 1638 -1578 1644 -1572
rect 1638 -1584 1644 -1578
rect 1638 -1590 1644 -1584
rect 1638 -1596 1644 -1590
rect 1638 -1602 1644 -1596
rect 1638 -1608 1644 -1602
rect 1638 -1614 1644 -1608
rect 1638 -1620 1644 -1614
rect 1638 -1626 1644 -1620
rect 1638 -1632 1644 -1626
rect 1638 -1638 1644 -1632
rect 1638 -1644 1644 -1638
rect 1638 -1650 1644 -1644
rect 1638 -1656 1644 -1650
rect 1638 -1662 1644 -1656
rect 1638 -1668 1644 -1662
rect 1638 -1674 1644 -1668
rect 1638 -1680 1644 -1674
rect 1638 -1686 1644 -1680
rect 1638 -1692 1644 -1686
rect 1638 -1698 1644 -1692
rect 1638 -1704 1644 -1698
rect 1638 -1710 1644 -1704
rect 1638 -1716 1644 -1710
rect 1638 -1722 1644 -1716
rect 1638 -1728 1644 -1722
rect 1638 -1734 1644 -1728
rect 1638 -1740 1644 -1734
rect 1638 -1746 1644 -1740
rect 1638 -1752 1644 -1746
rect 1638 -1758 1644 -1752
rect 1638 -1764 1644 -1758
rect 1638 -1770 1644 -1764
rect 1638 -1776 1644 -1770
rect 1638 -1782 1644 -1776
rect 1638 -1788 1644 -1782
rect 1638 -1794 1644 -1788
rect 1638 -1800 1644 -1794
rect 1638 -1806 1644 -1800
rect 1638 -1812 1644 -1806
rect 1638 -1818 1644 -1812
rect 1638 -1824 1644 -1818
rect 1638 -1830 1644 -1824
rect 1638 -1836 1644 -1830
rect 1638 -1842 1644 -1836
rect 1638 -1848 1644 -1842
rect 1638 -1854 1644 -1848
rect 1638 -1860 1644 -1854
rect 1638 -1866 1644 -1860
rect 1638 -1872 1644 -1866
rect 1638 -1878 1644 -1872
rect 1638 -1884 1644 -1878
rect 1638 -1890 1644 -1884
rect 1638 -1896 1644 -1890
rect 1638 -1902 1644 -1896
rect 1638 -1908 1644 -1902
rect 1638 -1914 1644 -1908
rect 1638 -1920 1644 -1914
rect 1638 -1926 1644 -1920
rect 1638 -1932 1644 -1926
rect 1638 -1938 1644 -1932
rect 1638 -1944 1644 -1938
rect 1638 -1950 1644 -1944
rect 1638 -1956 1644 -1950
rect 1638 -1962 1644 -1956
rect 1638 -1968 1644 -1962
rect 1638 -1974 1644 -1968
rect 1638 -1980 1644 -1974
rect 1638 -1986 1644 -1980
rect 1638 -1992 1644 -1986
rect 1638 -1998 1644 -1992
rect 1638 -2004 1644 -1998
rect 1638 -2010 1644 -2004
rect 1638 -2016 1644 -2010
rect 1638 -2022 1644 -2016
rect 1638 -2100 1644 -2094
rect 1638 -2106 1644 -2100
rect 1638 -2112 1644 -2106
rect 1638 -2118 1644 -2112
rect 1638 -2124 1644 -2118
rect 1638 -2130 1644 -2124
rect 1638 -2136 1644 -2130
rect 1638 -2142 1644 -2136
rect 1638 -2148 1644 -2142
rect 1638 -2154 1644 -2148
rect 1638 -2160 1644 -2154
rect 1638 -2166 1644 -2160
rect 1638 -2172 1644 -2166
rect 1638 -2178 1644 -2172
rect 1638 -2184 1644 -2178
rect 1638 -2190 1644 -2184
rect 1638 -2196 1644 -2190
rect 1638 -2202 1644 -2196
rect 1638 -2208 1644 -2202
rect 1638 -2214 1644 -2208
rect 1638 -2220 1644 -2214
rect 1638 -2226 1644 -2220
rect 1638 -2232 1644 -2226
rect 1638 -2238 1644 -2232
rect 1638 -2244 1644 -2238
rect 1638 -2250 1644 -2244
rect 1638 -2256 1644 -2250
rect 1638 -2262 1644 -2256
rect 1638 -2268 1644 -2262
rect 1638 -2274 1644 -2268
rect 1638 -2280 1644 -2274
rect 1638 -2286 1644 -2280
rect 1638 -2292 1644 -2286
rect 1638 -2298 1644 -2292
rect 1638 -2304 1644 -2298
rect 1638 -2310 1644 -2304
rect 1638 -2316 1644 -2310
rect 1638 -2322 1644 -2316
rect 1638 -2328 1644 -2322
rect 1638 -2334 1644 -2328
rect 1638 -2340 1644 -2334
rect 1638 -2346 1644 -2340
rect 1638 -2352 1644 -2346
rect 1638 -2358 1644 -2352
rect 1638 -2364 1644 -2358
rect 1638 -2370 1644 -2364
rect 1638 -2376 1644 -2370
rect 1638 -2382 1644 -2376
rect 1638 -2388 1644 -2382
rect 1638 -2394 1644 -2388
rect 1638 -2400 1644 -2394
rect 1638 -2406 1644 -2400
rect 1638 -2412 1644 -2406
rect 1638 -2418 1644 -2412
rect 1638 -2424 1644 -2418
rect 1638 -2430 1644 -2424
rect 1638 -2436 1644 -2430
rect 1638 -2442 1644 -2436
rect 1638 -2448 1644 -2442
rect 1638 -2454 1644 -2448
rect 1638 -2460 1644 -2454
rect 1638 -2466 1644 -2460
rect 1638 -2472 1644 -2466
rect 1638 -2478 1644 -2472
rect 1638 -2484 1644 -2478
rect 1638 -2490 1644 -2484
rect 1638 -2496 1644 -2490
rect 1638 -2502 1644 -2496
rect 1638 -2508 1644 -2502
rect 1638 -2514 1644 -2508
rect 1638 -2520 1644 -2514
rect 1638 -2526 1644 -2520
rect 1638 -2532 1644 -2526
rect 1638 -2538 1644 -2532
rect 1638 -2544 1644 -2538
rect 1638 -2550 1644 -2544
rect 1638 -2556 1644 -2550
rect 1638 -2562 1644 -2556
rect 1638 -2568 1644 -2562
rect 1638 -2574 1644 -2568
rect 1638 -2580 1644 -2574
rect 1638 -2586 1644 -2580
rect 1638 -2592 1644 -2586
rect 1638 -2598 1644 -2592
rect 1638 -2604 1644 -2598
rect 1638 -2610 1644 -2604
rect 1638 -2616 1644 -2610
rect 1638 -2622 1644 -2616
rect 1638 -2628 1644 -2622
rect 1638 -2634 1644 -2628
rect 1638 -2640 1644 -2634
rect 1638 -2646 1644 -2640
rect 1638 -2652 1644 -2646
rect 1638 -2658 1644 -2652
rect 1638 -2664 1644 -2658
rect 1638 -2670 1644 -2664
rect 1638 -2676 1644 -2670
rect 1638 -2682 1644 -2676
rect 1638 -2688 1644 -2682
rect 1638 -2694 1644 -2688
rect 1638 -2700 1644 -2694
rect 1638 -2706 1644 -2700
rect 1638 -2712 1644 -2706
rect 1638 -2718 1644 -2712
rect 1638 -2724 1644 -2718
rect 1638 -2802 1644 -2796
rect 1638 -2808 1644 -2802
rect 1638 -2814 1644 -2808
rect 1638 -2820 1644 -2814
rect 1638 -2826 1644 -2820
rect 1638 -2832 1644 -2826
rect 1638 -2838 1644 -2832
rect 1638 -2844 1644 -2838
rect 1638 -2850 1644 -2844
rect 1638 -2856 1644 -2850
rect 1638 -2862 1644 -2856
rect 1638 -2868 1644 -2862
rect 1638 -2874 1644 -2868
rect 1638 -2880 1644 -2874
rect 1638 -2886 1644 -2880
rect 1638 -2892 1644 -2886
rect 1638 -2898 1644 -2892
rect 1638 -2904 1644 -2898
rect 1638 -2910 1644 -2904
rect 1638 -2916 1644 -2910
rect 1638 -2922 1644 -2916
rect 1638 -2928 1644 -2922
rect 1638 -2934 1644 -2928
rect 1638 -2940 1644 -2934
rect 1638 -2946 1644 -2940
rect 1638 -2952 1644 -2946
rect 1638 -2958 1644 -2952
rect 1638 -2964 1644 -2958
rect 1638 -2970 1644 -2964
rect 1638 -2976 1644 -2970
rect 1638 -2982 1644 -2976
rect 1638 -2988 1644 -2982
rect 1638 -2994 1644 -2988
rect 1638 -3000 1644 -2994
rect 1638 -3006 1644 -3000
rect 1638 -3012 1644 -3006
rect 1638 -3018 1644 -3012
rect 1638 -3024 1644 -3018
rect 1638 -3030 1644 -3024
rect 1638 -3036 1644 -3030
rect 1638 -3042 1644 -3036
rect 1638 -3048 1644 -3042
rect 1638 -3054 1644 -3048
rect 1638 -3060 1644 -3054
rect 1638 -3066 1644 -3060
rect 1638 -3072 1644 -3066
rect 1638 -3078 1644 -3072
rect 1638 -3084 1644 -3078
rect 1638 -3090 1644 -3084
rect 1638 -3096 1644 -3090
rect 1638 -3102 1644 -3096
rect 1638 -3108 1644 -3102
rect 1638 -3114 1644 -3108
rect 1638 -3120 1644 -3114
rect 1638 -3126 1644 -3120
rect 1638 -3132 1644 -3126
rect 1638 -3138 1644 -3132
rect 1638 -3144 1644 -3138
rect 1638 -3150 1644 -3144
rect 1638 -3156 1644 -3150
rect 1638 -3162 1644 -3156
rect 1638 -3168 1644 -3162
rect 1638 -3174 1644 -3168
rect 1638 -3180 1644 -3174
rect 1638 -3186 1644 -3180
rect 1638 -3192 1644 -3186
rect 1638 -3198 1644 -3192
rect 1638 -3204 1644 -3198
rect 1638 -3210 1644 -3204
rect 1638 -3216 1644 -3210
rect 1638 -3222 1644 -3216
rect 1638 -3228 1644 -3222
rect 1638 -3234 1644 -3228
rect 1638 -3276 1644 -3270
rect 1638 -3282 1644 -3276
rect 1638 -3288 1644 -3282
rect 1638 -3294 1644 -3288
rect 1638 -3300 1644 -3294
rect 1638 -3306 1644 -3300
rect 1638 -3312 1644 -3306
rect 1638 -3318 1644 -3312
rect 1638 -3324 1644 -3318
rect 1638 -3330 1644 -3324
rect 1638 -3336 1644 -3330
rect 1638 -3342 1644 -3336
rect 1638 -3348 1644 -3342
rect 1638 -3354 1644 -3348
rect 1638 -3360 1644 -3354
rect 1638 -3366 1644 -3360
rect 1638 -3372 1644 -3366
rect 1638 -3378 1644 -3372
rect 1638 -3384 1644 -3378
rect 1638 -3390 1644 -3384
rect 1638 -3396 1644 -3390
rect 1638 -3402 1644 -3396
rect 1638 -3408 1644 -3402
rect 1638 -3414 1644 -3408
rect 1638 -3420 1644 -3414
rect 1638 -3426 1644 -3420
rect 1638 -3432 1644 -3426
rect 1638 -3438 1644 -3432
rect 1638 -3444 1644 -3438
rect 1644 -948 1650 -942
rect 1644 -954 1650 -948
rect 1644 -960 1650 -954
rect 1644 -966 1650 -960
rect 1644 -972 1650 -966
rect 1644 -978 1650 -972
rect 1644 -984 1650 -978
rect 1644 -990 1650 -984
rect 1644 -996 1650 -990
rect 1644 -1002 1650 -996
rect 1644 -1008 1650 -1002
rect 1644 -1014 1650 -1008
rect 1644 -1020 1650 -1014
rect 1644 -1026 1650 -1020
rect 1644 -1032 1650 -1026
rect 1644 -1038 1650 -1032
rect 1644 -1044 1650 -1038
rect 1644 -1050 1650 -1044
rect 1644 -1056 1650 -1050
rect 1644 -1062 1650 -1056
rect 1644 -1068 1650 -1062
rect 1644 -1074 1650 -1068
rect 1644 -1080 1650 -1074
rect 1644 -1086 1650 -1080
rect 1644 -1092 1650 -1086
rect 1644 -1098 1650 -1092
rect 1644 -1104 1650 -1098
rect 1644 -1110 1650 -1104
rect 1644 -1116 1650 -1110
rect 1644 -1122 1650 -1116
rect 1644 -1128 1650 -1122
rect 1644 -1134 1650 -1128
rect 1644 -1140 1650 -1134
rect 1644 -1146 1650 -1140
rect 1644 -1152 1650 -1146
rect 1644 -1158 1650 -1152
rect 1644 -1164 1650 -1158
rect 1644 -1170 1650 -1164
rect 1644 -1176 1650 -1170
rect 1644 -1182 1650 -1176
rect 1644 -1188 1650 -1182
rect 1644 -1194 1650 -1188
rect 1644 -1200 1650 -1194
rect 1644 -1206 1650 -1200
rect 1644 -1212 1650 -1206
rect 1644 -1218 1650 -1212
rect 1644 -1224 1650 -1218
rect 1644 -1230 1650 -1224
rect 1644 -1236 1650 -1230
rect 1644 -1242 1650 -1236
rect 1644 -1248 1650 -1242
rect 1644 -1254 1650 -1248
rect 1644 -1260 1650 -1254
rect 1644 -1266 1650 -1260
rect 1644 -1272 1650 -1266
rect 1644 -1278 1650 -1272
rect 1644 -1284 1650 -1278
rect 1644 -1290 1650 -1284
rect 1644 -1296 1650 -1290
rect 1644 -1302 1650 -1296
rect 1644 -1308 1650 -1302
rect 1644 -1314 1650 -1308
rect 1644 -1320 1650 -1314
rect 1644 -1326 1650 -1320
rect 1644 -1332 1650 -1326
rect 1644 -1338 1650 -1332
rect 1644 -1344 1650 -1338
rect 1644 -1350 1650 -1344
rect 1644 -1356 1650 -1350
rect 1644 -1362 1650 -1356
rect 1644 -1368 1650 -1362
rect 1644 -1374 1650 -1368
rect 1644 -1380 1650 -1374
rect 1644 -1386 1650 -1380
rect 1644 -1392 1650 -1386
rect 1644 -1398 1650 -1392
rect 1644 -1404 1650 -1398
rect 1644 -1410 1650 -1404
rect 1644 -1416 1650 -1410
rect 1644 -1422 1650 -1416
rect 1644 -1428 1650 -1422
rect 1644 -1434 1650 -1428
rect 1644 -1440 1650 -1434
rect 1644 -1446 1650 -1440
rect 1644 -1452 1650 -1446
rect 1644 -1458 1650 -1452
rect 1644 -1464 1650 -1458
rect 1644 -1470 1650 -1464
rect 1644 -1476 1650 -1470
rect 1644 -1482 1650 -1476
rect 1644 -1488 1650 -1482
rect 1644 -1494 1650 -1488
rect 1644 -1500 1650 -1494
rect 1644 -1506 1650 -1500
rect 1644 -1512 1650 -1506
rect 1644 -1518 1650 -1512
rect 1644 -1524 1650 -1518
rect 1644 -1530 1650 -1524
rect 1644 -1536 1650 -1530
rect 1644 -1542 1650 -1536
rect 1644 -1548 1650 -1542
rect 1644 -1554 1650 -1548
rect 1644 -1560 1650 -1554
rect 1644 -1566 1650 -1560
rect 1644 -1572 1650 -1566
rect 1644 -1578 1650 -1572
rect 1644 -1584 1650 -1578
rect 1644 -1590 1650 -1584
rect 1644 -1596 1650 -1590
rect 1644 -1602 1650 -1596
rect 1644 -1608 1650 -1602
rect 1644 -1614 1650 -1608
rect 1644 -1620 1650 -1614
rect 1644 -1626 1650 -1620
rect 1644 -1632 1650 -1626
rect 1644 -1638 1650 -1632
rect 1644 -1644 1650 -1638
rect 1644 -1650 1650 -1644
rect 1644 -1656 1650 -1650
rect 1644 -1662 1650 -1656
rect 1644 -1668 1650 -1662
rect 1644 -1674 1650 -1668
rect 1644 -1680 1650 -1674
rect 1644 -1686 1650 -1680
rect 1644 -1692 1650 -1686
rect 1644 -1698 1650 -1692
rect 1644 -1704 1650 -1698
rect 1644 -1710 1650 -1704
rect 1644 -1716 1650 -1710
rect 1644 -1722 1650 -1716
rect 1644 -1728 1650 -1722
rect 1644 -1734 1650 -1728
rect 1644 -1740 1650 -1734
rect 1644 -1746 1650 -1740
rect 1644 -1752 1650 -1746
rect 1644 -1758 1650 -1752
rect 1644 -1764 1650 -1758
rect 1644 -1770 1650 -1764
rect 1644 -1776 1650 -1770
rect 1644 -1782 1650 -1776
rect 1644 -1788 1650 -1782
rect 1644 -1794 1650 -1788
rect 1644 -1800 1650 -1794
rect 1644 -1806 1650 -1800
rect 1644 -1812 1650 -1806
rect 1644 -1818 1650 -1812
rect 1644 -1824 1650 -1818
rect 1644 -1830 1650 -1824
rect 1644 -1836 1650 -1830
rect 1644 -1842 1650 -1836
rect 1644 -1848 1650 -1842
rect 1644 -1854 1650 -1848
rect 1644 -1860 1650 -1854
rect 1644 -1866 1650 -1860
rect 1644 -1872 1650 -1866
rect 1644 -1878 1650 -1872
rect 1644 -1884 1650 -1878
rect 1644 -1890 1650 -1884
rect 1644 -1896 1650 -1890
rect 1644 -1902 1650 -1896
rect 1644 -1908 1650 -1902
rect 1644 -1914 1650 -1908
rect 1644 -1920 1650 -1914
rect 1644 -1926 1650 -1920
rect 1644 -1932 1650 -1926
rect 1644 -1938 1650 -1932
rect 1644 -1944 1650 -1938
rect 1644 -1950 1650 -1944
rect 1644 -1956 1650 -1950
rect 1644 -1962 1650 -1956
rect 1644 -1968 1650 -1962
rect 1644 -1974 1650 -1968
rect 1644 -1980 1650 -1974
rect 1644 -1986 1650 -1980
rect 1644 -1992 1650 -1986
rect 1644 -1998 1650 -1992
rect 1644 -2004 1650 -1998
rect 1644 -2010 1650 -2004
rect 1644 -2016 1650 -2010
rect 1644 -2094 1650 -2088
rect 1644 -2100 1650 -2094
rect 1644 -2106 1650 -2100
rect 1644 -2112 1650 -2106
rect 1644 -2118 1650 -2112
rect 1644 -2124 1650 -2118
rect 1644 -2130 1650 -2124
rect 1644 -2136 1650 -2130
rect 1644 -2142 1650 -2136
rect 1644 -2148 1650 -2142
rect 1644 -2154 1650 -2148
rect 1644 -2160 1650 -2154
rect 1644 -2166 1650 -2160
rect 1644 -2172 1650 -2166
rect 1644 -2178 1650 -2172
rect 1644 -2184 1650 -2178
rect 1644 -2190 1650 -2184
rect 1644 -2196 1650 -2190
rect 1644 -2202 1650 -2196
rect 1644 -2208 1650 -2202
rect 1644 -2214 1650 -2208
rect 1644 -2220 1650 -2214
rect 1644 -2226 1650 -2220
rect 1644 -2232 1650 -2226
rect 1644 -2238 1650 -2232
rect 1644 -2244 1650 -2238
rect 1644 -2250 1650 -2244
rect 1644 -2256 1650 -2250
rect 1644 -2262 1650 -2256
rect 1644 -2268 1650 -2262
rect 1644 -2274 1650 -2268
rect 1644 -2280 1650 -2274
rect 1644 -2286 1650 -2280
rect 1644 -2292 1650 -2286
rect 1644 -2298 1650 -2292
rect 1644 -2304 1650 -2298
rect 1644 -2310 1650 -2304
rect 1644 -2316 1650 -2310
rect 1644 -2322 1650 -2316
rect 1644 -2328 1650 -2322
rect 1644 -2334 1650 -2328
rect 1644 -2340 1650 -2334
rect 1644 -2346 1650 -2340
rect 1644 -2352 1650 -2346
rect 1644 -2358 1650 -2352
rect 1644 -2364 1650 -2358
rect 1644 -2370 1650 -2364
rect 1644 -2376 1650 -2370
rect 1644 -2382 1650 -2376
rect 1644 -2388 1650 -2382
rect 1644 -2394 1650 -2388
rect 1644 -2400 1650 -2394
rect 1644 -2406 1650 -2400
rect 1644 -2412 1650 -2406
rect 1644 -2418 1650 -2412
rect 1644 -2424 1650 -2418
rect 1644 -2430 1650 -2424
rect 1644 -2436 1650 -2430
rect 1644 -2442 1650 -2436
rect 1644 -2448 1650 -2442
rect 1644 -2454 1650 -2448
rect 1644 -2460 1650 -2454
rect 1644 -2466 1650 -2460
rect 1644 -2472 1650 -2466
rect 1644 -2478 1650 -2472
rect 1644 -2484 1650 -2478
rect 1644 -2490 1650 -2484
rect 1644 -2496 1650 -2490
rect 1644 -2502 1650 -2496
rect 1644 -2508 1650 -2502
rect 1644 -2514 1650 -2508
rect 1644 -2520 1650 -2514
rect 1644 -2526 1650 -2520
rect 1644 -2532 1650 -2526
rect 1644 -2538 1650 -2532
rect 1644 -2544 1650 -2538
rect 1644 -2550 1650 -2544
rect 1644 -2556 1650 -2550
rect 1644 -2562 1650 -2556
rect 1644 -2568 1650 -2562
rect 1644 -2574 1650 -2568
rect 1644 -2580 1650 -2574
rect 1644 -2586 1650 -2580
rect 1644 -2592 1650 -2586
rect 1644 -2598 1650 -2592
rect 1644 -2604 1650 -2598
rect 1644 -2610 1650 -2604
rect 1644 -2616 1650 -2610
rect 1644 -2622 1650 -2616
rect 1644 -2628 1650 -2622
rect 1644 -2634 1650 -2628
rect 1644 -2640 1650 -2634
rect 1644 -2646 1650 -2640
rect 1644 -2652 1650 -2646
rect 1644 -2658 1650 -2652
rect 1644 -2664 1650 -2658
rect 1644 -2670 1650 -2664
rect 1644 -2676 1650 -2670
rect 1644 -2682 1650 -2676
rect 1644 -2688 1650 -2682
rect 1644 -2694 1650 -2688
rect 1644 -2700 1650 -2694
rect 1644 -2706 1650 -2700
rect 1644 -2712 1650 -2706
rect 1644 -2718 1650 -2712
rect 1644 -2802 1650 -2796
rect 1644 -2808 1650 -2802
rect 1644 -2814 1650 -2808
rect 1644 -2820 1650 -2814
rect 1644 -2826 1650 -2820
rect 1644 -2832 1650 -2826
rect 1644 -2838 1650 -2832
rect 1644 -2844 1650 -2838
rect 1644 -2850 1650 -2844
rect 1644 -2856 1650 -2850
rect 1644 -2862 1650 -2856
rect 1644 -2868 1650 -2862
rect 1644 -2874 1650 -2868
rect 1644 -2880 1650 -2874
rect 1644 -2886 1650 -2880
rect 1644 -2892 1650 -2886
rect 1644 -2898 1650 -2892
rect 1644 -2904 1650 -2898
rect 1644 -2910 1650 -2904
rect 1644 -2916 1650 -2910
rect 1644 -2922 1650 -2916
rect 1644 -2928 1650 -2922
rect 1644 -2934 1650 -2928
rect 1644 -2940 1650 -2934
rect 1644 -2946 1650 -2940
rect 1644 -2952 1650 -2946
rect 1644 -2958 1650 -2952
rect 1644 -2964 1650 -2958
rect 1644 -2970 1650 -2964
rect 1644 -2976 1650 -2970
rect 1644 -2982 1650 -2976
rect 1644 -2988 1650 -2982
rect 1644 -2994 1650 -2988
rect 1644 -3000 1650 -2994
rect 1644 -3006 1650 -3000
rect 1644 -3012 1650 -3006
rect 1644 -3018 1650 -3012
rect 1644 -3024 1650 -3018
rect 1644 -3030 1650 -3024
rect 1644 -3036 1650 -3030
rect 1644 -3042 1650 -3036
rect 1644 -3048 1650 -3042
rect 1644 -3054 1650 -3048
rect 1644 -3060 1650 -3054
rect 1644 -3066 1650 -3060
rect 1644 -3072 1650 -3066
rect 1644 -3078 1650 -3072
rect 1644 -3084 1650 -3078
rect 1644 -3090 1650 -3084
rect 1644 -3096 1650 -3090
rect 1644 -3102 1650 -3096
rect 1644 -3108 1650 -3102
rect 1644 -3114 1650 -3108
rect 1644 -3120 1650 -3114
rect 1644 -3126 1650 -3120
rect 1644 -3132 1650 -3126
rect 1644 -3138 1650 -3132
rect 1644 -3144 1650 -3138
rect 1644 -3150 1650 -3144
rect 1644 -3156 1650 -3150
rect 1644 -3162 1650 -3156
rect 1644 -3168 1650 -3162
rect 1644 -3174 1650 -3168
rect 1644 -3180 1650 -3174
rect 1644 -3186 1650 -3180
rect 1644 -3192 1650 -3186
rect 1644 -3198 1650 -3192
rect 1644 -3204 1650 -3198
rect 1644 -3210 1650 -3204
rect 1644 -3216 1650 -3210
rect 1644 -3222 1650 -3216
rect 1644 -3228 1650 -3222
rect 1644 -3234 1650 -3228
rect 1644 -3276 1650 -3270
rect 1644 -3282 1650 -3276
rect 1644 -3288 1650 -3282
rect 1644 -3294 1650 -3288
rect 1644 -3300 1650 -3294
rect 1644 -3306 1650 -3300
rect 1644 -3312 1650 -3306
rect 1644 -3318 1650 -3312
rect 1644 -3324 1650 -3318
rect 1644 -3330 1650 -3324
rect 1644 -3336 1650 -3330
rect 1644 -3342 1650 -3336
rect 1644 -3348 1650 -3342
rect 1644 -3354 1650 -3348
rect 1644 -3360 1650 -3354
rect 1644 -3366 1650 -3360
rect 1644 -3372 1650 -3366
rect 1644 -3378 1650 -3372
rect 1644 -3384 1650 -3378
rect 1644 -3390 1650 -3384
rect 1644 -3396 1650 -3390
rect 1644 -3402 1650 -3396
rect 1644 -3408 1650 -3402
rect 1644 -3414 1650 -3408
rect 1644 -3420 1650 -3414
rect 1644 -3426 1650 -3420
rect 1644 -3432 1650 -3426
rect 1644 -3438 1650 -3432
rect 1644 -3444 1650 -3438
rect 1650 -936 1656 -930
rect 1650 -942 1656 -936
rect 1650 -948 1656 -942
rect 1650 -954 1656 -948
rect 1650 -960 1656 -954
rect 1650 -966 1656 -960
rect 1650 -972 1656 -966
rect 1650 -978 1656 -972
rect 1650 -984 1656 -978
rect 1650 -990 1656 -984
rect 1650 -996 1656 -990
rect 1650 -1002 1656 -996
rect 1650 -1008 1656 -1002
rect 1650 -1014 1656 -1008
rect 1650 -1020 1656 -1014
rect 1650 -1026 1656 -1020
rect 1650 -1032 1656 -1026
rect 1650 -1038 1656 -1032
rect 1650 -1044 1656 -1038
rect 1650 -1050 1656 -1044
rect 1650 -1056 1656 -1050
rect 1650 -1062 1656 -1056
rect 1650 -1068 1656 -1062
rect 1650 -1074 1656 -1068
rect 1650 -1080 1656 -1074
rect 1650 -1086 1656 -1080
rect 1650 -1092 1656 -1086
rect 1650 -1098 1656 -1092
rect 1650 -1104 1656 -1098
rect 1650 -1110 1656 -1104
rect 1650 -1116 1656 -1110
rect 1650 -1122 1656 -1116
rect 1650 -1128 1656 -1122
rect 1650 -1134 1656 -1128
rect 1650 -1140 1656 -1134
rect 1650 -1146 1656 -1140
rect 1650 -1152 1656 -1146
rect 1650 -1158 1656 -1152
rect 1650 -1164 1656 -1158
rect 1650 -1170 1656 -1164
rect 1650 -1176 1656 -1170
rect 1650 -1182 1656 -1176
rect 1650 -1188 1656 -1182
rect 1650 -1194 1656 -1188
rect 1650 -1200 1656 -1194
rect 1650 -1206 1656 -1200
rect 1650 -1212 1656 -1206
rect 1650 -1218 1656 -1212
rect 1650 -1224 1656 -1218
rect 1650 -1230 1656 -1224
rect 1650 -1236 1656 -1230
rect 1650 -1242 1656 -1236
rect 1650 -1248 1656 -1242
rect 1650 -1254 1656 -1248
rect 1650 -1260 1656 -1254
rect 1650 -1266 1656 -1260
rect 1650 -1272 1656 -1266
rect 1650 -1278 1656 -1272
rect 1650 -1284 1656 -1278
rect 1650 -1290 1656 -1284
rect 1650 -1296 1656 -1290
rect 1650 -1302 1656 -1296
rect 1650 -1308 1656 -1302
rect 1650 -1314 1656 -1308
rect 1650 -1320 1656 -1314
rect 1650 -1326 1656 -1320
rect 1650 -1332 1656 -1326
rect 1650 -1338 1656 -1332
rect 1650 -1344 1656 -1338
rect 1650 -1350 1656 -1344
rect 1650 -1356 1656 -1350
rect 1650 -1362 1656 -1356
rect 1650 -1368 1656 -1362
rect 1650 -1374 1656 -1368
rect 1650 -1380 1656 -1374
rect 1650 -1386 1656 -1380
rect 1650 -1392 1656 -1386
rect 1650 -1398 1656 -1392
rect 1650 -1404 1656 -1398
rect 1650 -1410 1656 -1404
rect 1650 -1416 1656 -1410
rect 1650 -1422 1656 -1416
rect 1650 -1428 1656 -1422
rect 1650 -1434 1656 -1428
rect 1650 -1440 1656 -1434
rect 1650 -1446 1656 -1440
rect 1650 -1452 1656 -1446
rect 1650 -1458 1656 -1452
rect 1650 -1464 1656 -1458
rect 1650 -1470 1656 -1464
rect 1650 -1476 1656 -1470
rect 1650 -1482 1656 -1476
rect 1650 -1488 1656 -1482
rect 1650 -1494 1656 -1488
rect 1650 -1500 1656 -1494
rect 1650 -1506 1656 -1500
rect 1650 -1512 1656 -1506
rect 1650 -1518 1656 -1512
rect 1650 -1524 1656 -1518
rect 1650 -1530 1656 -1524
rect 1650 -1536 1656 -1530
rect 1650 -1542 1656 -1536
rect 1650 -1548 1656 -1542
rect 1650 -1554 1656 -1548
rect 1650 -1560 1656 -1554
rect 1650 -1566 1656 -1560
rect 1650 -1572 1656 -1566
rect 1650 -1578 1656 -1572
rect 1650 -1584 1656 -1578
rect 1650 -1590 1656 -1584
rect 1650 -1596 1656 -1590
rect 1650 -1602 1656 -1596
rect 1650 -1608 1656 -1602
rect 1650 -1614 1656 -1608
rect 1650 -1620 1656 -1614
rect 1650 -1626 1656 -1620
rect 1650 -1632 1656 -1626
rect 1650 -1638 1656 -1632
rect 1650 -1644 1656 -1638
rect 1650 -1650 1656 -1644
rect 1650 -1656 1656 -1650
rect 1650 -1662 1656 -1656
rect 1650 -1668 1656 -1662
rect 1650 -1674 1656 -1668
rect 1650 -1680 1656 -1674
rect 1650 -1686 1656 -1680
rect 1650 -1692 1656 -1686
rect 1650 -1698 1656 -1692
rect 1650 -1704 1656 -1698
rect 1650 -1710 1656 -1704
rect 1650 -1716 1656 -1710
rect 1650 -1722 1656 -1716
rect 1650 -1728 1656 -1722
rect 1650 -1734 1656 -1728
rect 1650 -1740 1656 -1734
rect 1650 -1746 1656 -1740
rect 1650 -1752 1656 -1746
rect 1650 -1758 1656 -1752
rect 1650 -1764 1656 -1758
rect 1650 -1770 1656 -1764
rect 1650 -1776 1656 -1770
rect 1650 -1782 1656 -1776
rect 1650 -1788 1656 -1782
rect 1650 -1794 1656 -1788
rect 1650 -1800 1656 -1794
rect 1650 -1806 1656 -1800
rect 1650 -1812 1656 -1806
rect 1650 -1818 1656 -1812
rect 1650 -1824 1656 -1818
rect 1650 -1830 1656 -1824
rect 1650 -1836 1656 -1830
rect 1650 -1842 1656 -1836
rect 1650 -1848 1656 -1842
rect 1650 -1854 1656 -1848
rect 1650 -1860 1656 -1854
rect 1650 -1866 1656 -1860
rect 1650 -1872 1656 -1866
rect 1650 -1878 1656 -1872
rect 1650 -1884 1656 -1878
rect 1650 -1890 1656 -1884
rect 1650 -1896 1656 -1890
rect 1650 -1902 1656 -1896
rect 1650 -1908 1656 -1902
rect 1650 -1914 1656 -1908
rect 1650 -1920 1656 -1914
rect 1650 -1926 1656 -1920
rect 1650 -1932 1656 -1926
rect 1650 -1938 1656 -1932
rect 1650 -1944 1656 -1938
rect 1650 -1950 1656 -1944
rect 1650 -1956 1656 -1950
rect 1650 -1962 1656 -1956
rect 1650 -1968 1656 -1962
rect 1650 -1974 1656 -1968
rect 1650 -1980 1656 -1974
rect 1650 -1986 1656 -1980
rect 1650 -1992 1656 -1986
rect 1650 -1998 1656 -1992
rect 1650 -2004 1656 -1998
rect 1650 -2010 1656 -2004
rect 1650 -2082 1656 -2076
rect 1650 -2088 1656 -2082
rect 1650 -2094 1656 -2088
rect 1650 -2100 1656 -2094
rect 1650 -2106 1656 -2100
rect 1650 -2112 1656 -2106
rect 1650 -2118 1656 -2112
rect 1650 -2124 1656 -2118
rect 1650 -2130 1656 -2124
rect 1650 -2136 1656 -2130
rect 1650 -2142 1656 -2136
rect 1650 -2148 1656 -2142
rect 1650 -2154 1656 -2148
rect 1650 -2160 1656 -2154
rect 1650 -2166 1656 -2160
rect 1650 -2172 1656 -2166
rect 1650 -2178 1656 -2172
rect 1650 -2184 1656 -2178
rect 1650 -2190 1656 -2184
rect 1650 -2196 1656 -2190
rect 1650 -2202 1656 -2196
rect 1650 -2208 1656 -2202
rect 1650 -2214 1656 -2208
rect 1650 -2220 1656 -2214
rect 1650 -2226 1656 -2220
rect 1650 -2232 1656 -2226
rect 1650 -2238 1656 -2232
rect 1650 -2244 1656 -2238
rect 1650 -2250 1656 -2244
rect 1650 -2256 1656 -2250
rect 1650 -2262 1656 -2256
rect 1650 -2268 1656 -2262
rect 1650 -2274 1656 -2268
rect 1650 -2280 1656 -2274
rect 1650 -2286 1656 -2280
rect 1650 -2292 1656 -2286
rect 1650 -2298 1656 -2292
rect 1650 -2304 1656 -2298
rect 1650 -2310 1656 -2304
rect 1650 -2316 1656 -2310
rect 1650 -2322 1656 -2316
rect 1650 -2328 1656 -2322
rect 1650 -2334 1656 -2328
rect 1650 -2340 1656 -2334
rect 1650 -2346 1656 -2340
rect 1650 -2352 1656 -2346
rect 1650 -2358 1656 -2352
rect 1650 -2364 1656 -2358
rect 1650 -2370 1656 -2364
rect 1650 -2376 1656 -2370
rect 1650 -2382 1656 -2376
rect 1650 -2388 1656 -2382
rect 1650 -2394 1656 -2388
rect 1650 -2400 1656 -2394
rect 1650 -2406 1656 -2400
rect 1650 -2412 1656 -2406
rect 1650 -2418 1656 -2412
rect 1650 -2424 1656 -2418
rect 1650 -2430 1656 -2424
rect 1650 -2436 1656 -2430
rect 1650 -2442 1656 -2436
rect 1650 -2448 1656 -2442
rect 1650 -2454 1656 -2448
rect 1650 -2460 1656 -2454
rect 1650 -2466 1656 -2460
rect 1650 -2472 1656 -2466
rect 1650 -2478 1656 -2472
rect 1650 -2484 1656 -2478
rect 1650 -2490 1656 -2484
rect 1650 -2496 1656 -2490
rect 1650 -2502 1656 -2496
rect 1650 -2508 1656 -2502
rect 1650 -2514 1656 -2508
rect 1650 -2520 1656 -2514
rect 1650 -2526 1656 -2520
rect 1650 -2532 1656 -2526
rect 1650 -2538 1656 -2532
rect 1650 -2544 1656 -2538
rect 1650 -2550 1656 -2544
rect 1650 -2556 1656 -2550
rect 1650 -2562 1656 -2556
rect 1650 -2568 1656 -2562
rect 1650 -2574 1656 -2568
rect 1650 -2580 1656 -2574
rect 1650 -2586 1656 -2580
rect 1650 -2592 1656 -2586
rect 1650 -2598 1656 -2592
rect 1650 -2604 1656 -2598
rect 1650 -2610 1656 -2604
rect 1650 -2616 1656 -2610
rect 1650 -2622 1656 -2616
rect 1650 -2628 1656 -2622
rect 1650 -2634 1656 -2628
rect 1650 -2640 1656 -2634
rect 1650 -2646 1656 -2640
rect 1650 -2652 1656 -2646
rect 1650 -2658 1656 -2652
rect 1650 -2664 1656 -2658
rect 1650 -2670 1656 -2664
rect 1650 -2676 1656 -2670
rect 1650 -2682 1656 -2676
rect 1650 -2688 1656 -2682
rect 1650 -2694 1656 -2688
rect 1650 -2700 1656 -2694
rect 1650 -2706 1656 -2700
rect 1650 -2712 1656 -2706
rect 1650 -2718 1656 -2712
rect 1650 -2796 1656 -2790
rect 1650 -2802 1656 -2796
rect 1650 -2808 1656 -2802
rect 1650 -2814 1656 -2808
rect 1650 -2820 1656 -2814
rect 1650 -2826 1656 -2820
rect 1650 -2832 1656 -2826
rect 1650 -2838 1656 -2832
rect 1650 -2844 1656 -2838
rect 1650 -2850 1656 -2844
rect 1650 -2856 1656 -2850
rect 1650 -2862 1656 -2856
rect 1650 -2868 1656 -2862
rect 1650 -2874 1656 -2868
rect 1650 -2880 1656 -2874
rect 1650 -2886 1656 -2880
rect 1650 -2892 1656 -2886
rect 1650 -2898 1656 -2892
rect 1650 -2904 1656 -2898
rect 1650 -2910 1656 -2904
rect 1650 -2916 1656 -2910
rect 1650 -2922 1656 -2916
rect 1650 -2928 1656 -2922
rect 1650 -2934 1656 -2928
rect 1650 -2940 1656 -2934
rect 1650 -2946 1656 -2940
rect 1650 -2952 1656 -2946
rect 1650 -2958 1656 -2952
rect 1650 -2964 1656 -2958
rect 1650 -2970 1656 -2964
rect 1650 -2976 1656 -2970
rect 1650 -2982 1656 -2976
rect 1650 -2988 1656 -2982
rect 1650 -2994 1656 -2988
rect 1650 -3000 1656 -2994
rect 1650 -3006 1656 -3000
rect 1650 -3012 1656 -3006
rect 1650 -3018 1656 -3012
rect 1650 -3024 1656 -3018
rect 1650 -3030 1656 -3024
rect 1650 -3036 1656 -3030
rect 1650 -3042 1656 -3036
rect 1650 -3048 1656 -3042
rect 1650 -3054 1656 -3048
rect 1650 -3060 1656 -3054
rect 1650 -3066 1656 -3060
rect 1650 -3072 1656 -3066
rect 1650 -3078 1656 -3072
rect 1650 -3084 1656 -3078
rect 1650 -3090 1656 -3084
rect 1650 -3096 1656 -3090
rect 1650 -3102 1656 -3096
rect 1650 -3108 1656 -3102
rect 1650 -3114 1656 -3108
rect 1650 -3120 1656 -3114
rect 1650 -3126 1656 -3120
rect 1650 -3132 1656 -3126
rect 1650 -3138 1656 -3132
rect 1650 -3144 1656 -3138
rect 1650 -3150 1656 -3144
rect 1650 -3156 1656 -3150
rect 1650 -3162 1656 -3156
rect 1650 -3168 1656 -3162
rect 1650 -3174 1656 -3168
rect 1650 -3180 1656 -3174
rect 1650 -3186 1656 -3180
rect 1650 -3192 1656 -3186
rect 1650 -3198 1656 -3192
rect 1650 -3204 1656 -3198
rect 1650 -3210 1656 -3204
rect 1650 -3216 1656 -3210
rect 1650 -3222 1656 -3216
rect 1650 -3228 1656 -3222
rect 1650 -3234 1656 -3228
rect 1650 -3276 1656 -3270
rect 1650 -3282 1656 -3276
rect 1650 -3288 1656 -3282
rect 1650 -3294 1656 -3288
rect 1650 -3300 1656 -3294
rect 1650 -3306 1656 -3300
rect 1650 -3312 1656 -3306
rect 1650 -3318 1656 -3312
rect 1650 -3324 1656 -3318
rect 1650 -3330 1656 -3324
rect 1650 -3336 1656 -3330
rect 1650 -3342 1656 -3336
rect 1650 -3348 1656 -3342
rect 1650 -3354 1656 -3348
rect 1650 -3360 1656 -3354
rect 1650 -3366 1656 -3360
rect 1650 -3372 1656 -3366
rect 1650 -3378 1656 -3372
rect 1650 -3384 1656 -3378
rect 1650 -3390 1656 -3384
rect 1650 -3396 1656 -3390
rect 1650 -3402 1656 -3396
rect 1650 -3408 1656 -3402
rect 1650 -3414 1656 -3408
rect 1650 -3420 1656 -3414
rect 1650 -3426 1656 -3420
rect 1650 -3432 1656 -3426
rect 1650 -3438 1656 -3432
rect 1656 -930 1662 -924
rect 1656 -936 1662 -930
rect 1656 -942 1662 -936
rect 1656 -948 1662 -942
rect 1656 -954 1662 -948
rect 1656 -960 1662 -954
rect 1656 -966 1662 -960
rect 1656 -972 1662 -966
rect 1656 -978 1662 -972
rect 1656 -984 1662 -978
rect 1656 -990 1662 -984
rect 1656 -996 1662 -990
rect 1656 -1002 1662 -996
rect 1656 -1008 1662 -1002
rect 1656 -1014 1662 -1008
rect 1656 -1020 1662 -1014
rect 1656 -1026 1662 -1020
rect 1656 -1032 1662 -1026
rect 1656 -1038 1662 -1032
rect 1656 -1044 1662 -1038
rect 1656 -1050 1662 -1044
rect 1656 -1056 1662 -1050
rect 1656 -1062 1662 -1056
rect 1656 -1068 1662 -1062
rect 1656 -1074 1662 -1068
rect 1656 -1080 1662 -1074
rect 1656 -1086 1662 -1080
rect 1656 -1092 1662 -1086
rect 1656 -1098 1662 -1092
rect 1656 -1104 1662 -1098
rect 1656 -1110 1662 -1104
rect 1656 -1116 1662 -1110
rect 1656 -1122 1662 -1116
rect 1656 -1128 1662 -1122
rect 1656 -1134 1662 -1128
rect 1656 -1140 1662 -1134
rect 1656 -1146 1662 -1140
rect 1656 -1152 1662 -1146
rect 1656 -1158 1662 -1152
rect 1656 -1164 1662 -1158
rect 1656 -1170 1662 -1164
rect 1656 -1176 1662 -1170
rect 1656 -1182 1662 -1176
rect 1656 -1188 1662 -1182
rect 1656 -1194 1662 -1188
rect 1656 -1200 1662 -1194
rect 1656 -1206 1662 -1200
rect 1656 -1212 1662 -1206
rect 1656 -1218 1662 -1212
rect 1656 -1224 1662 -1218
rect 1656 -1230 1662 -1224
rect 1656 -1236 1662 -1230
rect 1656 -1242 1662 -1236
rect 1656 -1248 1662 -1242
rect 1656 -1254 1662 -1248
rect 1656 -1260 1662 -1254
rect 1656 -1266 1662 -1260
rect 1656 -1272 1662 -1266
rect 1656 -1278 1662 -1272
rect 1656 -1284 1662 -1278
rect 1656 -1290 1662 -1284
rect 1656 -1296 1662 -1290
rect 1656 -1302 1662 -1296
rect 1656 -1308 1662 -1302
rect 1656 -1314 1662 -1308
rect 1656 -1320 1662 -1314
rect 1656 -1326 1662 -1320
rect 1656 -1332 1662 -1326
rect 1656 -1338 1662 -1332
rect 1656 -1344 1662 -1338
rect 1656 -1350 1662 -1344
rect 1656 -1356 1662 -1350
rect 1656 -1362 1662 -1356
rect 1656 -1368 1662 -1362
rect 1656 -1374 1662 -1368
rect 1656 -1380 1662 -1374
rect 1656 -1386 1662 -1380
rect 1656 -1392 1662 -1386
rect 1656 -1398 1662 -1392
rect 1656 -1404 1662 -1398
rect 1656 -1410 1662 -1404
rect 1656 -1416 1662 -1410
rect 1656 -1422 1662 -1416
rect 1656 -1428 1662 -1422
rect 1656 -1434 1662 -1428
rect 1656 -1440 1662 -1434
rect 1656 -1446 1662 -1440
rect 1656 -1452 1662 -1446
rect 1656 -1458 1662 -1452
rect 1656 -1464 1662 -1458
rect 1656 -1470 1662 -1464
rect 1656 -1476 1662 -1470
rect 1656 -1482 1662 -1476
rect 1656 -1488 1662 -1482
rect 1656 -1494 1662 -1488
rect 1656 -1500 1662 -1494
rect 1656 -1506 1662 -1500
rect 1656 -1512 1662 -1506
rect 1656 -1518 1662 -1512
rect 1656 -1524 1662 -1518
rect 1656 -1530 1662 -1524
rect 1656 -1536 1662 -1530
rect 1656 -1542 1662 -1536
rect 1656 -1548 1662 -1542
rect 1656 -1554 1662 -1548
rect 1656 -1560 1662 -1554
rect 1656 -1566 1662 -1560
rect 1656 -1572 1662 -1566
rect 1656 -1578 1662 -1572
rect 1656 -1584 1662 -1578
rect 1656 -1590 1662 -1584
rect 1656 -1596 1662 -1590
rect 1656 -1602 1662 -1596
rect 1656 -1608 1662 -1602
rect 1656 -1614 1662 -1608
rect 1656 -1620 1662 -1614
rect 1656 -1626 1662 -1620
rect 1656 -1632 1662 -1626
rect 1656 -1638 1662 -1632
rect 1656 -1644 1662 -1638
rect 1656 -1650 1662 -1644
rect 1656 -1656 1662 -1650
rect 1656 -1662 1662 -1656
rect 1656 -1668 1662 -1662
rect 1656 -1674 1662 -1668
rect 1656 -1680 1662 -1674
rect 1656 -1686 1662 -1680
rect 1656 -1692 1662 -1686
rect 1656 -1698 1662 -1692
rect 1656 -1704 1662 -1698
rect 1656 -1710 1662 -1704
rect 1656 -1716 1662 -1710
rect 1656 -1722 1662 -1716
rect 1656 -1728 1662 -1722
rect 1656 -1734 1662 -1728
rect 1656 -1740 1662 -1734
rect 1656 -1746 1662 -1740
rect 1656 -1752 1662 -1746
rect 1656 -1758 1662 -1752
rect 1656 -1764 1662 -1758
rect 1656 -1770 1662 -1764
rect 1656 -1776 1662 -1770
rect 1656 -1782 1662 -1776
rect 1656 -1788 1662 -1782
rect 1656 -1794 1662 -1788
rect 1656 -1800 1662 -1794
rect 1656 -1806 1662 -1800
rect 1656 -1812 1662 -1806
rect 1656 -1818 1662 -1812
rect 1656 -1824 1662 -1818
rect 1656 -1830 1662 -1824
rect 1656 -1836 1662 -1830
rect 1656 -1842 1662 -1836
rect 1656 -1848 1662 -1842
rect 1656 -1854 1662 -1848
rect 1656 -1860 1662 -1854
rect 1656 -1866 1662 -1860
rect 1656 -1872 1662 -1866
rect 1656 -1878 1662 -1872
rect 1656 -1884 1662 -1878
rect 1656 -1890 1662 -1884
rect 1656 -1896 1662 -1890
rect 1656 -1902 1662 -1896
rect 1656 -1908 1662 -1902
rect 1656 -1914 1662 -1908
rect 1656 -1920 1662 -1914
rect 1656 -1926 1662 -1920
rect 1656 -1932 1662 -1926
rect 1656 -1938 1662 -1932
rect 1656 -1944 1662 -1938
rect 1656 -1950 1662 -1944
rect 1656 -1956 1662 -1950
rect 1656 -1962 1662 -1956
rect 1656 -1968 1662 -1962
rect 1656 -1974 1662 -1968
rect 1656 -1980 1662 -1974
rect 1656 -1986 1662 -1980
rect 1656 -1992 1662 -1986
rect 1656 -1998 1662 -1992
rect 1656 -2004 1662 -1998
rect 1656 -2076 1662 -2070
rect 1656 -2082 1662 -2076
rect 1656 -2088 1662 -2082
rect 1656 -2094 1662 -2088
rect 1656 -2100 1662 -2094
rect 1656 -2106 1662 -2100
rect 1656 -2112 1662 -2106
rect 1656 -2118 1662 -2112
rect 1656 -2124 1662 -2118
rect 1656 -2130 1662 -2124
rect 1656 -2136 1662 -2130
rect 1656 -2142 1662 -2136
rect 1656 -2148 1662 -2142
rect 1656 -2154 1662 -2148
rect 1656 -2160 1662 -2154
rect 1656 -2166 1662 -2160
rect 1656 -2172 1662 -2166
rect 1656 -2178 1662 -2172
rect 1656 -2184 1662 -2178
rect 1656 -2190 1662 -2184
rect 1656 -2196 1662 -2190
rect 1656 -2202 1662 -2196
rect 1656 -2208 1662 -2202
rect 1656 -2214 1662 -2208
rect 1656 -2220 1662 -2214
rect 1656 -2226 1662 -2220
rect 1656 -2232 1662 -2226
rect 1656 -2238 1662 -2232
rect 1656 -2244 1662 -2238
rect 1656 -2250 1662 -2244
rect 1656 -2256 1662 -2250
rect 1656 -2262 1662 -2256
rect 1656 -2268 1662 -2262
rect 1656 -2274 1662 -2268
rect 1656 -2280 1662 -2274
rect 1656 -2286 1662 -2280
rect 1656 -2292 1662 -2286
rect 1656 -2298 1662 -2292
rect 1656 -2304 1662 -2298
rect 1656 -2310 1662 -2304
rect 1656 -2316 1662 -2310
rect 1656 -2322 1662 -2316
rect 1656 -2328 1662 -2322
rect 1656 -2334 1662 -2328
rect 1656 -2340 1662 -2334
rect 1656 -2346 1662 -2340
rect 1656 -2352 1662 -2346
rect 1656 -2358 1662 -2352
rect 1656 -2364 1662 -2358
rect 1656 -2370 1662 -2364
rect 1656 -2376 1662 -2370
rect 1656 -2382 1662 -2376
rect 1656 -2388 1662 -2382
rect 1656 -2394 1662 -2388
rect 1656 -2400 1662 -2394
rect 1656 -2406 1662 -2400
rect 1656 -2412 1662 -2406
rect 1656 -2418 1662 -2412
rect 1656 -2424 1662 -2418
rect 1656 -2430 1662 -2424
rect 1656 -2436 1662 -2430
rect 1656 -2442 1662 -2436
rect 1656 -2448 1662 -2442
rect 1656 -2454 1662 -2448
rect 1656 -2460 1662 -2454
rect 1656 -2466 1662 -2460
rect 1656 -2472 1662 -2466
rect 1656 -2478 1662 -2472
rect 1656 -2484 1662 -2478
rect 1656 -2490 1662 -2484
rect 1656 -2496 1662 -2490
rect 1656 -2502 1662 -2496
rect 1656 -2508 1662 -2502
rect 1656 -2514 1662 -2508
rect 1656 -2520 1662 -2514
rect 1656 -2526 1662 -2520
rect 1656 -2532 1662 -2526
rect 1656 -2538 1662 -2532
rect 1656 -2544 1662 -2538
rect 1656 -2550 1662 -2544
rect 1656 -2556 1662 -2550
rect 1656 -2562 1662 -2556
rect 1656 -2568 1662 -2562
rect 1656 -2574 1662 -2568
rect 1656 -2580 1662 -2574
rect 1656 -2586 1662 -2580
rect 1656 -2592 1662 -2586
rect 1656 -2598 1662 -2592
rect 1656 -2604 1662 -2598
rect 1656 -2610 1662 -2604
rect 1656 -2616 1662 -2610
rect 1656 -2622 1662 -2616
rect 1656 -2628 1662 -2622
rect 1656 -2634 1662 -2628
rect 1656 -2640 1662 -2634
rect 1656 -2646 1662 -2640
rect 1656 -2652 1662 -2646
rect 1656 -2658 1662 -2652
rect 1656 -2664 1662 -2658
rect 1656 -2670 1662 -2664
rect 1656 -2676 1662 -2670
rect 1656 -2682 1662 -2676
rect 1656 -2688 1662 -2682
rect 1656 -2694 1662 -2688
rect 1656 -2700 1662 -2694
rect 1656 -2706 1662 -2700
rect 1656 -2712 1662 -2706
rect 1656 -2790 1662 -2784
rect 1656 -2796 1662 -2790
rect 1656 -2802 1662 -2796
rect 1656 -2808 1662 -2802
rect 1656 -2814 1662 -2808
rect 1656 -2820 1662 -2814
rect 1656 -2826 1662 -2820
rect 1656 -2832 1662 -2826
rect 1656 -2838 1662 -2832
rect 1656 -2844 1662 -2838
rect 1656 -2850 1662 -2844
rect 1656 -2856 1662 -2850
rect 1656 -2862 1662 -2856
rect 1656 -2868 1662 -2862
rect 1656 -2874 1662 -2868
rect 1656 -2880 1662 -2874
rect 1656 -2886 1662 -2880
rect 1656 -2892 1662 -2886
rect 1656 -2898 1662 -2892
rect 1656 -2904 1662 -2898
rect 1656 -2910 1662 -2904
rect 1656 -2916 1662 -2910
rect 1656 -2922 1662 -2916
rect 1656 -2928 1662 -2922
rect 1656 -2934 1662 -2928
rect 1656 -2940 1662 -2934
rect 1656 -2946 1662 -2940
rect 1656 -2952 1662 -2946
rect 1656 -2958 1662 -2952
rect 1656 -2964 1662 -2958
rect 1656 -2970 1662 -2964
rect 1656 -2976 1662 -2970
rect 1656 -2982 1662 -2976
rect 1656 -2988 1662 -2982
rect 1656 -2994 1662 -2988
rect 1656 -3000 1662 -2994
rect 1656 -3006 1662 -3000
rect 1656 -3012 1662 -3006
rect 1656 -3018 1662 -3012
rect 1656 -3024 1662 -3018
rect 1656 -3030 1662 -3024
rect 1656 -3036 1662 -3030
rect 1656 -3042 1662 -3036
rect 1656 -3048 1662 -3042
rect 1656 -3054 1662 -3048
rect 1656 -3060 1662 -3054
rect 1656 -3066 1662 -3060
rect 1656 -3072 1662 -3066
rect 1656 -3078 1662 -3072
rect 1656 -3084 1662 -3078
rect 1656 -3090 1662 -3084
rect 1656 -3096 1662 -3090
rect 1656 -3102 1662 -3096
rect 1656 -3108 1662 -3102
rect 1656 -3114 1662 -3108
rect 1656 -3120 1662 -3114
rect 1656 -3126 1662 -3120
rect 1656 -3132 1662 -3126
rect 1656 -3138 1662 -3132
rect 1656 -3144 1662 -3138
rect 1656 -3150 1662 -3144
rect 1656 -3156 1662 -3150
rect 1656 -3162 1662 -3156
rect 1656 -3168 1662 -3162
rect 1656 -3174 1662 -3168
rect 1656 -3180 1662 -3174
rect 1656 -3186 1662 -3180
rect 1656 -3192 1662 -3186
rect 1656 -3198 1662 -3192
rect 1656 -3204 1662 -3198
rect 1656 -3210 1662 -3204
rect 1656 -3216 1662 -3210
rect 1656 -3222 1662 -3216
rect 1656 -3228 1662 -3222
rect 1656 -3234 1662 -3228
rect 1656 -3276 1662 -3270
rect 1656 -3282 1662 -3276
rect 1656 -3288 1662 -3282
rect 1656 -3294 1662 -3288
rect 1656 -3300 1662 -3294
rect 1656 -3306 1662 -3300
rect 1656 -3312 1662 -3306
rect 1656 -3318 1662 -3312
rect 1656 -3324 1662 -3318
rect 1656 -3330 1662 -3324
rect 1656 -3336 1662 -3330
rect 1656 -3342 1662 -3336
rect 1656 -3348 1662 -3342
rect 1656 -3354 1662 -3348
rect 1656 -3360 1662 -3354
rect 1656 -3366 1662 -3360
rect 1656 -3372 1662 -3366
rect 1656 -3378 1662 -3372
rect 1656 -3384 1662 -3378
rect 1656 -3390 1662 -3384
rect 1656 -3396 1662 -3390
rect 1656 -3402 1662 -3396
rect 1656 -3408 1662 -3402
rect 1656 -3414 1662 -3408
rect 1656 -3420 1662 -3414
rect 1656 -3426 1662 -3420
rect 1656 -3432 1662 -3426
rect 1656 -3438 1662 -3432
rect 1662 -918 1668 -912
rect 1662 -924 1668 -918
rect 1662 -930 1668 -924
rect 1662 -936 1668 -930
rect 1662 -942 1668 -936
rect 1662 -948 1668 -942
rect 1662 -954 1668 -948
rect 1662 -960 1668 -954
rect 1662 -966 1668 -960
rect 1662 -972 1668 -966
rect 1662 -978 1668 -972
rect 1662 -984 1668 -978
rect 1662 -990 1668 -984
rect 1662 -996 1668 -990
rect 1662 -1002 1668 -996
rect 1662 -1008 1668 -1002
rect 1662 -1014 1668 -1008
rect 1662 -1020 1668 -1014
rect 1662 -1026 1668 -1020
rect 1662 -1032 1668 -1026
rect 1662 -1038 1668 -1032
rect 1662 -1044 1668 -1038
rect 1662 -1050 1668 -1044
rect 1662 -1056 1668 -1050
rect 1662 -1062 1668 -1056
rect 1662 -1068 1668 -1062
rect 1662 -1074 1668 -1068
rect 1662 -1080 1668 -1074
rect 1662 -1086 1668 -1080
rect 1662 -1092 1668 -1086
rect 1662 -1098 1668 -1092
rect 1662 -1104 1668 -1098
rect 1662 -1110 1668 -1104
rect 1662 -1116 1668 -1110
rect 1662 -1122 1668 -1116
rect 1662 -1128 1668 -1122
rect 1662 -1134 1668 -1128
rect 1662 -1140 1668 -1134
rect 1662 -1146 1668 -1140
rect 1662 -1152 1668 -1146
rect 1662 -1158 1668 -1152
rect 1662 -1164 1668 -1158
rect 1662 -1170 1668 -1164
rect 1662 -1176 1668 -1170
rect 1662 -1182 1668 -1176
rect 1662 -1188 1668 -1182
rect 1662 -1194 1668 -1188
rect 1662 -1200 1668 -1194
rect 1662 -1206 1668 -1200
rect 1662 -1212 1668 -1206
rect 1662 -1218 1668 -1212
rect 1662 -1224 1668 -1218
rect 1662 -1230 1668 -1224
rect 1662 -1236 1668 -1230
rect 1662 -1242 1668 -1236
rect 1662 -1248 1668 -1242
rect 1662 -1254 1668 -1248
rect 1662 -1260 1668 -1254
rect 1662 -1266 1668 -1260
rect 1662 -1272 1668 -1266
rect 1662 -1278 1668 -1272
rect 1662 -1284 1668 -1278
rect 1662 -1290 1668 -1284
rect 1662 -1296 1668 -1290
rect 1662 -1302 1668 -1296
rect 1662 -1308 1668 -1302
rect 1662 -1314 1668 -1308
rect 1662 -1320 1668 -1314
rect 1662 -1326 1668 -1320
rect 1662 -1332 1668 -1326
rect 1662 -1338 1668 -1332
rect 1662 -1344 1668 -1338
rect 1662 -1350 1668 -1344
rect 1662 -1356 1668 -1350
rect 1662 -1362 1668 -1356
rect 1662 -1368 1668 -1362
rect 1662 -1374 1668 -1368
rect 1662 -1380 1668 -1374
rect 1662 -1386 1668 -1380
rect 1662 -1392 1668 -1386
rect 1662 -1398 1668 -1392
rect 1662 -1404 1668 -1398
rect 1662 -1410 1668 -1404
rect 1662 -1416 1668 -1410
rect 1662 -1422 1668 -1416
rect 1662 -1428 1668 -1422
rect 1662 -1434 1668 -1428
rect 1662 -1440 1668 -1434
rect 1662 -1446 1668 -1440
rect 1662 -1452 1668 -1446
rect 1662 -1458 1668 -1452
rect 1662 -1464 1668 -1458
rect 1662 -1470 1668 -1464
rect 1662 -1476 1668 -1470
rect 1662 -1482 1668 -1476
rect 1662 -1488 1668 -1482
rect 1662 -1494 1668 -1488
rect 1662 -1500 1668 -1494
rect 1662 -1506 1668 -1500
rect 1662 -1512 1668 -1506
rect 1662 -1518 1668 -1512
rect 1662 -1524 1668 -1518
rect 1662 -1530 1668 -1524
rect 1662 -1536 1668 -1530
rect 1662 -1542 1668 -1536
rect 1662 -1548 1668 -1542
rect 1662 -1554 1668 -1548
rect 1662 -1560 1668 -1554
rect 1662 -1566 1668 -1560
rect 1662 -1572 1668 -1566
rect 1662 -1578 1668 -1572
rect 1662 -1584 1668 -1578
rect 1662 -1590 1668 -1584
rect 1662 -1596 1668 -1590
rect 1662 -1602 1668 -1596
rect 1662 -1608 1668 -1602
rect 1662 -1614 1668 -1608
rect 1662 -1620 1668 -1614
rect 1662 -1626 1668 -1620
rect 1662 -1632 1668 -1626
rect 1662 -1638 1668 -1632
rect 1662 -1644 1668 -1638
rect 1662 -1650 1668 -1644
rect 1662 -1656 1668 -1650
rect 1662 -1662 1668 -1656
rect 1662 -1668 1668 -1662
rect 1662 -1674 1668 -1668
rect 1662 -1680 1668 -1674
rect 1662 -1686 1668 -1680
rect 1662 -1692 1668 -1686
rect 1662 -1698 1668 -1692
rect 1662 -1704 1668 -1698
rect 1662 -1710 1668 -1704
rect 1662 -1716 1668 -1710
rect 1662 -1722 1668 -1716
rect 1662 -1728 1668 -1722
rect 1662 -1734 1668 -1728
rect 1662 -1740 1668 -1734
rect 1662 -1746 1668 -1740
rect 1662 -1752 1668 -1746
rect 1662 -1758 1668 -1752
rect 1662 -1764 1668 -1758
rect 1662 -1770 1668 -1764
rect 1662 -1776 1668 -1770
rect 1662 -1782 1668 -1776
rect 1662 -1788 1668 -1782
rect 1662 -1794 1668 -1788
rect 1662 -1800 1668 -1794
rect 1662 -1806 1668 -1800
rect 1662 -1812 1668 -1806
rect 1662 -1818 1668 -1812
rect 1662 -1824 1668 -1818
rect 1662 -1830 1668 -1824
rect 1662 -1836 1668 -1830
rect 1662 -1842 1668 -1836
rect 1662 -1848 1668 -1842
rect 1662 -1854 1668 -1848
rect 1662 -1860 1668 -1854
rect 1662 -1866 1668 -1860
rect 1662 -1872 1668 -1866
rect 1662 -1878 1668 -1872
rect 1662 -1884 1668 -1878
rect 1662 -1890 1668 -1884
rect 1662 -1896 1668 -1890
rect 1662 -1902 1668 -1896
rect 1662 -1908 1668 -1902
rect 1662 -1914 1668 -1908
rect 1662 -1920 1668 -1914
rect 1662 -1926 1668 -1920
rect 1662 -1932 1668 -1926
rect 1662 -1938 1668 -1932
rect 1662 -1944 1668 -1938
rect 1662 -1950 1668 -1944
rect 1662 -1956 1668 -1950
rect 1662 -1962 1668 -1956
rect 1662 -1968 1668 -1962
rect 1662 -1974 1668 -1968
rect 1662 -1980 1668 -1974
rect 1662 -1986 1668 -1980
rect 1662 -1992 1668 -1986
rect 1662 -1998 1668 -1992
rect 1662 -2070 1668 -2064
rect 1662 -2076 1668 -2070
rect 1662 -2082 1668 -2076
rect 1662 -2088 1668 -2082
rect 1662 -2094 1668 -2088
rect 1662 -2100 1668 -2094
rect 1662 -2106 1668 -2100
rect 1662 -2112 1668 -2106
rect 1662 -2118 1668 -2112
rect 1662 -2124 1668 -2118
rect 1662 -2130 1668 -2124
rect 1662 -2136 1668 -2130
rect 1662 -2142 1668 -2136
rect 1662 -2148 1668 -2142
rect 1662 -2154 1668 -2148
rect 1662 -2160 1668 -2154
rect 1662 -2166 1668 -2160
rect 1662 -2172 1668 -2166
rect 1662 -2178 1668 -2172
rect 1662 -2184 1668 -2178
rect 1662 -2190 1668 -2184
rect 1662 -2196 1668 -2190
rect 1662 -2202 1668 -2196
rect 1662 -2208 1668 -2202
rect 1662 -2214 1668 -2208
rect 1662 -2220 1668 -2214
rect 1662 -2226 1668 -2220
rect 1662 -2232 1668 -2226
rect 1662 -2238 1668 -2232
rect 1662 -2244 1668 -2238
rect 1662 -2250 1668 -2244
rect 1662 -2256 1668 -2250
rect 1662 -2262 1668 -2256
rect 1662 -2268 1668 -2262
rect 1662 -2274 1668 -2268
rect 1662 -2280 1668 -2274
rect 1662 -2286 1668 -2280
rect 1662 -2292 1668 -2286
rect 1662 -2298 1668 -2292
rect 1662 -2304 1668 -2298
rect 1662 -2310 1668 -2304
rect 1662 -2316 1668 -2310
rect 1662 -2322 1668 -2316
rect 1662 -2328 1668 -2322
rect 1662 -2334 1668 -2328
rect 1662 -2340 1668 -2334
rect 1662 -2346 1668 -2340
rect 1662 -2352 1668 -2346
rect 1662 -2358 1668 -2352
rect 1662 -2364 1668 -2358
rect 1662 -2370 1668 -2364
rect 1662 -2376 1668 -2370
rect 1662 -2382 1668 -2376
rect 1662 -2388 1668 -2382
rect 1662 -2394 1668 -2388
rect 1662 -2400 1668 -2394
rect 1662 -2406 1668 -2400
rect 1662 -2412 1668 -2406
rect 1662 -2418 1668 -2412
rect 1662 -2424 1668 -2418
rect 1662 -2430 1668 -2424
rect 1662 -2436 1668 -2430
rect 1662 -2442 1668 -2436
rect 1662 -2448 1668 -2442
rect 1662 -2454 1668 -2448
rect 1662 -2460 1668 -2454
rect 1662 -2466 1668 -2460
rect 1662 -2472 1668 -2466
rect 1662 -2478 1668 -2472
rect 1662 -2484 1668 -2478
rect 1662 -2490 1668 -2484
rect 1662 -2496 1668 -2490
rect 1662 -2502 1668 -2496
rect 1662 -2508 1668 -2502
rect 1662 -2514 1668 -2508
rect 1662 -2520 1668 -2514
rect 1662 -2526 1668 -2520
rect 1662 -2532 1668 -2526
rect 1662 -2538 1668 -2532
rect 1662 -2544 1668 -2538
rect 1662 -2550 1668 -2544
rect 1662 -2556 1668 -2550
rect 1662 -2562 1668 -2556
rect 1662 -2568 1668 -2562
rect 1662 -2574 1668 -2568
rect 1662 -2580 1668 -2574
rect 1662 -2586 1668 -2580
rect 1662 -2592 1668 -2586
rect 1662 -2598 1668 -2592
rect 1662 -2604 1668 -2598
rect 1662 -2610 1668 -2604
rect 1662 -2616 1668 -2610
rect 1662 -2622 1668 -2616
rect 1662 -2628 1668 -2622
rect 1662 -2634 1668 -2628
rect 1662 -2640 1668 -2634
rect 1662 -2646 1668 -2640
rect 1662 -2652 1668 -2646
rect 1662 -2658 1668 -2652
rect 1662 -2664 1668 -2658
rect 1662 -2670 1668 -2664
rect 1662 -2676 1668 -2670
rect 1662 -2682 1668 -2676
rect 1662 -2688 1668 -2682
rect 1662 -2694 1668 -2688
rect 1662 -2700 1668 -2694
rect 1662 -2706 1668 -2700
rect 1662 -2712 1668 -2706
rect 1662 -2790 1668 -2784
rect 1662 -2796 1668 -2790
rect 1662 -2802 1668 -2796
rect 1662 -2808 1668 -2802
rect 1662 -2814 1668 -2808
rect 1662 -2820 1668 -2814
rect 1662 -2826 1668 -2820
rect 1662 -2832 1668 -2826
rect 1662 -2838 1668 -2832
rect 1662 -2844 1668 -2838
rect 1662 -2850 1668 -2844
rect 1662 -2856 1668 -2850
rect 1662 -2862 1668 -2856
rect 1662 -2868 1668 -2862
rect 1662 -2874 1668 -2868
rect 1662 -2880 1668 -2874
rect 1662 -2886 1668 -2880
rect 1662 -2892 1668 -2886
rect 1662 -2898 1668 -2892
rect 1662 -2904 1668 -2898
rect 1662 -2910 1668 -2904
rect 1662 -2916 1668 -2910
rect 1662 -2922 1668 -2916
rect 1662 -2928 1668 -2922
rect 1662 -2934 1668 -2928
rect 1662 -2940 1668 -2934
rect 1662 -2946 1668 -2940
rect 1662 -2952 1668 -2946
rect 1662 -2958 1668 -2952
rect 1662 -2964 1668 -2958
rect 1662 -2970 1668 -2964
rect 1662 -2976 1668 -2970
rect 1662 -2982 1668 -2976
rect 1662 -2988 1668 -2982
rect 1662 -2994 1668 -2988
rect 1662 -3000 1668 -2994
rect 1662 -3006 1668 -3000
rect 1662 -3012 1668 -3006
rect 1662 -3018 1668 -3012
rect 1662 -3024 1668 -3018
rect 1662 -3030 1668 -3024
rect 1662 -3036 1668 -3030
rect 1662 -3042 1668 -3036
rect 1662 -3048 1668 -3042
rect 1662 -3054 1668 -3048
rect 1662 -3060 1668 -3054
rect 1662 -3066 1668 -3060
rect 1662 -3072 1668 -3066
rect 1662 -3078 1668 -3072
rect 1662 -3084 1668 -3078
rect 1662 -3090 1668 -3084
rect 1662 -3096 1668 -3090
rect 1662 -3102 1668 -3096
rect 1662 -3108 1668 -3102
rect 1662 -3114 1668 -3108
rect 1662 -3120 1668 -3114
rect 1662 -3126 1668 -3120
rect 1662 -3132 1668 -3126
rect 1662 -3138 1668 -3132
rect 1662 -3144 1668 -3138
rect 1662 -3150 1668 -3144
rect 1662 -3156 1668 -3150
rect 1662 -3162 1668 -3156
rect 1662 -3168 1668 -3162
rect 1662 -3174 1668 -3168
rect 1662 -3180 1668 -3174
rect 1662 -3186 1668 -3180
rect 1662 -3192 1668 -3186
rect 1662 -3198 1668 -3192
rect 1662 -3204 1668 -3198
rect 1662 -3210 1668 -3204
rect 1662 -3216 1668 -3210
rect 1662 -3222 1668 -3216
rect 1662 -3228 1668 -3222
rect 1662 -3234 1668 -3228
rect 1662 -3276 1668 -3270
rect 1662 -3282 1668 -3276
rect 1662 -3288 1668 -3282
rect 1662 -3294 1668 -3288
rect 1662 -3300 1668 -3294
rect 1662 -3306 1668 -3300
rect 1662 -3312 1668 -3306
rect 1662 -3318 1668 -3312
rect 1662 -3324 1668 -3318
rect 1662 -3330 1668 -3324
rect 1662 -3336 1668 -3330
rect 1662 -3342 1668 -3336
rect 1662 -3348 1668 -3342
rect 1662 -3354 1668 -3348
rect 1662 -3360 1668 -3354
rect 1662 -3366 1668 -3360
rect 1662 -3372 1668 -3366
rect 1662 -3378 1668 -3372
rect 1662 -3384 1668 -3378
rect 1662 -3390 1668 -3384
rect 1662 -3396 1668 -3390
rect 1662 -3402 1668 -3396
rect 1662 -3408 1668 -3402
rect 1662 -3414 1668 -3408
rect 1662 -3420 1668 -3414
rect 1662 -3426 1668 -3420
rect 1662 -3432 1668 -3426
rect 1662 -3438 1668 -3432
rect 1668 -912 1674 -906
rect 1668 -918 1674 -912
rect 1668 -924 1674 -918
rect 1668 -930 1674 -924
rect 1668 -936 1674 -930
rect 1668 -942 1674 -936
rect 1668 -948 1674 -942
rect 1668 -954 1674 -948
rect 1668 -960 1674 -954
rect 1668 -966 1674 -960
rect 1668 -972 1674 -966
rect 1668 -978 1674 -972
rect 1668 -984 1674 -978
rect 1668 -990 1674 -984
rect 1668 -996 1674 -990
rect 1668 -1002 1674 -996
rect 1668 -1008 1674 -1002
rect 1668 -1014 1674 -1008
rect 1668 -1020 1674 -1014
rect 1668 -1026 1674 -1020
rect 1668 -1032 1674 -1026
rect 1668 -1038 1674 -1032
rect 1668 -1044 1674 -1038
rect 1668 -1050 1674 -1044
rect 1668 -1056 1674 -1050
rect 1668 -1062 1674 -1056
rect 1668 -1068 1674 -1062
rect 1668 -1074 1674 -1068
rect 1668 -1080 1674 -1074
rect 1668 -1086 1674 -1080
rect 1668 -1092 1674 -1086
rect 1668 -1098 1674 -1092
rect 1668 -1104 1674 -1098
rect 1668 -1110 1674 -1104
rect 1668 -1116 1674 -1110
rect 1668 -1122 1674 -1116
rect 1668 -1128 1674 -1122
rect 1668 -1134 1674 -1128
rect 1668 -1140 1674 -1134
rect 1668 -1146 1674 -1140
rect 1668 -1152 1674 -1146
rect 1668 -1158 1674 -1152
rect 1668 -1164 1674 -1158
rect 1668 -1170 1674 -1164
rect 1668 -1176 1674 -1170
rect 1668 -1182 1674 -1176
rect 1668 -1188 1674 -1182
rect 1668 -1194 1674 -1188
rect 1668 -1200 1674 -1194
rect 1668 -1206 1674 -1200
rect 1668 -1212 1674 -1206
rect 1668 -1218 1674 -1212
rect 1668 -1224 1674 -1218
rect 1668 -1230 1674 -1224
rect 1668 -1236 1674 -1230
rect 1668 -1242 1674 -1236
rect 1668 -1248 1674 -1242
rect 1668 -1254 1674 -1248
rect 1668 -1260 1674 -1254
rect 1668 -1266 1674 -1260
rect 1668 -1272 1674 -1266
rect 1668 -1278 1674 -1272
rect 1668 -1284 1674 -1278
rect 1668 -1290 1674 -1284
rect 1668 -1296 1674 -1290
rect 1668 -1302 1674 -1296
rect 1668 -1308 1674 -1302
rect 1668 -1314 1674 -1308
rect 1668 -1320 1674 -1314
rect 1668 -1326 1674 -1320
rect 1668 -1332 1674 -1326
rect 1668 -1338 1674 -1332
rect 1668 -1344 1674 -1338
rect 1668 -1350 1674 -1344
rect 1668 -1356 1674 -1350
rect 1668 -1362 1674 -1356
rect 1668 -1368 1674 -1362
rect 1668 -1374 1674 -1368
rect 1668 -1380 1674 -1374
rect 1668 -1386 1674 -1380
rect 1668 -1392 1674 -1386
rect 1668 -1398 1674 -1392
rect 1668 -1404 1674 -1398
rect 1668 -1410 1674 -1404
rect 1668 -1416 1674 -1410
rect 1668 -1422 1674 -1416
rect 1668 -1428 1674 -1422
rect 1668 -1434 1674 -1428
rect 1668 -1440 1674 -1434
rect 1668 -1446 1674 -1440
rect 1668 -1452 1674 -1446
rect 1668 -1458 1674 -1452
rect 1668 -1464 1674 -1458
rect 1668 -1470 1674 -1464
rect 1668 -1476 1674 -1470
rect 1668 -1482 1674 -1476
rect 1668 -1488 1674 -1482
rect 1668 -1494 1674 -1488
rect 1668 -1500 1674 -1494
rect 1668 -1506 1674 -1500
rect 1668 -1512 1674 -1506
rect 1668 -1518 1674 -1512
rect 1668 -1524 1674 -1518
rect 1668 -1530 1674 -1524
rect 1668 -1536 1674 -1530
rect 1668 -1542 1674 -1536
rect 1668 -1548 1674 -1542
rect 1668 -1554 1674 -1548
rect 1668 -1560 1674 -1554
rect 1668 -1566 1674 -1560
rect 1668 -1572 1674 -1566
rect 1668 -1578 1674 -1572
rect 1668 -1584 1674 -1578
rect 1668 -1590 1674 -1584
rect 1668 -1596 1674 -1590
rect 1668 -1602 1674 -1596
rect 1668 -1608 1674 -1602
rect 1668 -1614 1674 -1608
rect 1668 -1620 1674 -1614
rect 1668 -1626 1674 -1620
rect 1668 -1632 1674 -1626
rect 1668 -1638 1674 -1632
rect 1668 -1644 1674 -1638
rect 1668 -1650 1674 -1644
rect 1668 -1656 1674 -1650
rect 1668 -1662 1674 -1656
rect 1668 -1668 1674 -1662
rect 1668 -1674 1674 -1668
rect 1668 -1680 1674 -1674
rect 1668 -1686 1674 -1680
rect 1668 -1692 1674 -1686
rect 1668 -1698 1674 -1692
rect 1668 -1704 1674 -1698
rect 1668 -1710 1674 -1704
rect 1668 -1716 1674 -1710
rect 1668 -1722 1674 -1716
rect 1668 -1728 1674 -1722
rect 1668 -1734 1674 -1728
rect 1668 -1740 1674 -1734
rect 1668 -1746 1674 -1740
rect 1668 -1752 1674 -1746
rect 1668 -1758 1674 -1752
rect 1668 -1764 1674 -1758
rect 1668 -1770 1674 -1764
rect 1668 -1776 1674 -1770
rect 1668 -1782 1674 -1776
rect 1668 -1788 1674 -1782
rect 1668 -1794 1674 -1788
rect 1668 -1800 1674 -1794
rect 1668 -1806 1674 -1800
rect 1668 -1812 1674 -1806
rect 1668 -1818 1674 -1812
rect 1668 -1824 1674 -1818
rect 1668 -1830 1674 -1824
rect 1668 -1836 1674 -1830
rect 1668 -1842 1674 -1836
rect 1668 -1848 1674 -1842
rect 1668 -1854 1674 -1848
rect 1668 -1860 1674 -1854
rect 1668 -1866 1674 -1860
rect 1668 -1872 1674 -1866
rect 1668 -1878 1674 -1872
rect 1668 -1884 1674 -1878
rect 1668 -1890 1674 -1884
rect 1668 -1896 1674 -1890
rect 1668 -1902 1674 -1896
rect 1668 -1908 1674 -1902
rect 1668 -1914 1674 -1908
rect 1668 -1920 1674 -1914
rect 1668 -1926 1674 -1920
rect 1668 -1932 1674 -1926
rect 1668 -1938 1674 -1932
rect 1668 -1944 1674 -1938
rect 1668 -1950 1674 -1944
rect 1668 -1956 1674 -1950
rect 1668 -1962 1674 -1956
rect 1668 -1968 1674 -1962
rect 1668 -1974 1674 -1968
rect 1668 -1980 1674 -1974
rect 1668 -1986 1674 -1980
rect 1668 -1992 1674 -1986
rect 1668 -2064 1674 -2058
rect 1668 -2070 1674 -2064
rect 1668 -2076 1674 -2070
rect 1668 -2082 1674 -2076
rect 1668 -2088 1674 -2082
rect 1668 -2094 1674 -2088
rect 1668 -2100 1674 -2094
rect 1668 -2106 1674 -2100
rect 1668 -2112 1674 -2106
rect 1668 -2118 1674 -2112
rect 1668 -2124 1674 -2118
rect 1668 -2130 1674 -2124
rect 1668 -2136 1674 -2130
rect 1668 -2142 1674 -2136
rect 1668 -2148 1674 -2142
rect 1668 -2154 1674 -2148
rect 1668 -2160 1674 -2154
rect 1668 -2166 1674 -2160
rect 1668 -2172 1674 -2166
rect 1668 -2178 1674 -2172
rect 1668 -2184 1674 -2178
rect 1668 -2190 1674 -2184
rect 1668 -2196 1674 -2190
rect 1668 -2202 1674 -2196
rect 1668 -2208 1674 -2202
rect 1668 -2214 1674 -2208
rect 1668 -2220 1674 -2214
rect 1668 -2226 1674 -2220
rect 1668 -2232 1674 -2226
rect 1668 -2238 1674 -2232
rect 1668 -2244 1674 -2238
rect 1668 -2250 1674 -2244
rect 1668 -2256 1674 -2250
rect 1668 -2262 1674 -2256
rect 1668 -2268 1674 -2262
rect 1668 -2274 1674 -2268
rect 1668 -2280 1674 -2274
rect 1668 -2286 1674 -2280
rect 1668 -2292 1674 -2286
rect 1668 -2298 1674 -2292
rect 1668 -2304 1674 -2298
rect 1668 -2310 1674 -2304
rect 1668 -2316 1674 -2310
rect 1668 -2322 1674 -2316
rect 1668 -2328 1674 -2322
rect 1668 -2334 1674 -2328
rect 1668 -2340 1674 -2334
rect 1668 -2346 1674 -2340
rect 1668 -2352 1674 -2346
rect 1668 -2358 1674 -2352
rect 1668 -2364 1674 -2358
rect 1668 -2370 1674 -2364
rect 1668 -2376 1674 -2370
rect 1668 -2382 1674 -2376
rect 1668 -2388 1674 -2382
rect 1668 -2394 1674 -2388
rect 1668 -2400 1674 -2394
rect 1668 -2406 1674 -2400
rect 1668 -2412 1674 -2406
rect 1668 -2418 1674 -2412
rect 1668 -2424 1674 -2418
rect 1668 -2430 1674 -2424
rect 1668 -2436 1674 -2430
rect 1668 -2442 1674 -2436
rect 1668 -2448 1674 -2442
rect 1668 -2454 1674 -2448
rect 1668 -2460 1674 -2454
rect 1668 -2466 1674 -2460
rect 1668 -2472 1674 -2466
rect 1668 -2478 1674 -2472
rect 1668 -2484 1674 -2478
rect 1668 -2490 1674 -2484
rect 1668 -2496 1674 -2490
rect 1668 -2502 1674 -2496
rect 1668 -2508 1674 -2502
rect 1668 -2514 1674 -2508
rect 1668 -2520 1674 -2514
rect 1668 -2526 1674 -2520
rect 1668 -2532 1674 -2526
rect 1668 -2538 1674 -2532
rect 1668 -2544 1674 -2538
rect 1668 -2550 1674 -2544
rect 1668 -2556 1674 -2550
rect 1668 -2562 1674 -2556
rect 1668 -2568 1674 -2562
rect 1668 -2574 1674 -2568
rect 1668 -2580 1674 -2574
rect 1668 -2586 1674 -2580
rect 1668 -2592 1674 -2586
rect 1668 -2598 1674 -2592
rect 1668 -2604 1674 -2598
rect 1668 -2610 1674 -2604
rect 1668 -2616 1674 -2610
rect 1668 -2622 1674 -2616
rect 1668 -2628 1674 -2622
rect 1668 -2634 1674 -2628
rect 1668 -2640 1674 -2634
rect 1668 -2646 1674 -2640
rect 1668 -2652 1674 -2646
rect 1668 -2658 1674 -2652
rect 1668 -2664 1674 -2658
rect 1668 -2670 1674 -2664
rect 1668 -2676 1674 -2670
rect 1668 -2682 1674 -2676
rect 1668 -2688 1674 -2682
rect 1668 -2694 1674 -2688
rect 1668 -2700 1674 -2694
rect 1668 -2706 1674 -2700
rect 1668 -2784 1674 -2778
rect 1668 -2790 1674 -2784
rect 1668 -2796 1674 -2790
rect 1668 -2802 1674 -2796
rect 1668 -2808 1674 -2802
rect 1668 -2814 1674 -2808
rect 1668 -2820 1674 -2814
rect 1668 -2826 1674 -2820
rect 1668 -2832 1674 -2826
rect 1668 -2838 1674 -2832
rect 1668 -2844 1674 -2838
rect 1668 -2850 1674 -2844
rect 1668 -2856 1674 -2850
rect 1668 -2862 1674 -2856
rect 1668 -2868 1674 -2862
rect 1668 -2874 1674 -2868
rect 1668 -2880 1674 -2874
rect 1668 -2886 1674 -2880
rect 1668 -2892 1674 -2886
rect 1668 -2898 1674 -2892
rect 1668 -2904 1674 -2898
rect 1668 -2910 1674 -2904
rect 1668 -2916 1674 -2910
rect 1668 -2922 1674 -2916
rect 1668 -2928 1674 -2922
rect 1668 -2934 1674 -2928
rect 1668 -2940 1674 -2934
rect 1668 -2946 1674 -2940
rect 1668 -2952 1674 -2946
rect 1668 -2958 1674 -2952
rect 1668 -2964 1674 -2958
rect 1668 -2970 1674 -2964
rect 1668 -2976 1674 -2970
rect 1668 -2982 1674 -2976
rect 1668 -2988 1674 -2982
rect 1668 -2994 1674 -2988
rect 1668 -3000 1674 -2994
rect 1668 -3006 1674 -3000
rect 1668 -3012 1674 -3006
rect 1668 -3018 1674 -3012
rect 1668 -3024 1674 -3018
rect 1668 -3030 1674 -3024
rect 1668 -3036 1674 -3030
rect 1668 -3042 1674 -3036
rect 1668 -3048 1674 -3042
rect 1668 -3054 1674 -3048
rect 1668 -3060 1674 -3054
rect 1668 -3066 1674 -3060
rect 1668 -3072 1674 -3066
rect 1668 -3078 1674 -3072
rect 1668 -3084 1674 -3078
rect 1668 -3090 1674 -3084
rect 1668 -3096 1674 -3090
rect 1668 -3102 1674 -3096
rect 1668 -3108 1674 -3102
rect 1668 -3114 1674 -3108
rect 1668 -3120 1674 -3114
rect 1668 -3126 1674 -3120
rect 1668 -3132 1674 -3126
rect 1668 -3138 1674 -3132
rect 1668 -3144 1674 -3138
rect 1668 -3150 1674 -3144
rect 1668 -3156 1674 -3150
rect 1668 -3162 1674 -3156
rect 1668 -3168 1674 -3162
rect 1668 -3174 1674 -3168
rect 1668 -3180 1674 -3174
rect 1668 -3186 1674 -3180
rect 1668 -3192 1674 -3186
rect 1668 -3198 1674 -3192
rect 1668 -3204 1674 -3198
rect 1668 -3210 1674 -3204
rect 1668 -3216 1674 -3210
rect 1668 -3222 1674 -3216
rect 1668 -3228 1674 -3222
rect 1668 -3234 1674 -3228
rect 1668 -3276 1674 -3270
rect 1668 -3282 1674 -3276
rect 1668 -3288 1674 -3282
rect 1668 -3294 1674 -3288
rect 1668 -3300 1674 -3294
rect 1668 -3306 1674 -3300
rect 1668 -3312 1674 -3306
rect 1668 -3318 1674 -3312
rect 1668 -3324 1674 -3318
rect 1668 -3330 1674 -3324
rect 1668 -3336 1674 -3330
rect 1668 -3342 1674 -3336
rect 1668 -3348 1674 -3342
rect 1668 -3354 1674 -3348
rect 1668 -3360 1674 -3354
rect 1668 -3366 1674 -3360
rect 1668 -3372 1674 -3366
rect 1668 -3378 1674 -3372
rect 1668 -3384 1674 -3378
rect 1668 -3390 1674 -3384
rect 1668 -3396 1674 -3390
rect 1668 -3402 1674 -3396
rect 1668 -3408 1674 -3402
rect 1668 -3414 1674 -3408
rect 1668 -3420 1674 -3414
rect 1668 -3426 1674 -3420
rect 1668 -3432 1674 -3426
rect 1674 -900 1680 -894
rect 1674 -906 1680 -900
rect 1674 -912 1680 -906
rect 1674 -918 1680 -912
rect 1674 -924 1680 -918
rect 1674 -930 1680 -924
rect 1674 -936 1680 -930
rect 1674 -942 1680 -936
rect 1674 -948 1680 -942
rect 1674 -954 1680 -948
rect 1674 -960 1680 -954
rect 1674 -966 1680 -960
rect 1674 -972 1680 -966
rect 1674 -978 1680 -972
rect 1674 -984 1680 -978
rect 1674 -990 1680 -984
rect 1674 -996 1680 -990
rect 1674 -1002 1680 -996
rect 1674 -1008 1680 -1002
rect 1674 -1014 1680 -1008
rect 1674 -1020 1680 -1014
rect 1674 -1026 1680 -1020
rect 1674 -1032 1680 -1026
rect 1674 -1038 1680 -1032
rect 1674 -1044 1680 -1038
rect 1674 -1050 1680 -1044
rect 1674 -1056 1680 -1050
rect 1674 -1062 1680 -1056
rect 1674 -1068 1680 -1062
rect 1674 -1074 1680 -1068
rect 1674 -1080 1680 -1074
rect 1674 -1086 1680 -1080
rect 1674 -1092 1680 -1086
rect 1674 -1098 1680 -1092
rect 1674 -1104 1680 -1098
rect 1674 -1110 1680 -1104
rect 1674 -1116 1680 -1110
rect 1674 -1122 1680 -1116
rect 1674 -1128 1680 -1122
rect 1674 -1134 1680 -1128
rect 1674 -1140 1680 -1134
rect 1674 -1146 1680 -1140
rect 1674 -1152 1680 -1146
rect 1674 -1158 1680 -1152
rect 1674 -1164 1680 -1158
rect 1674 -1170 1680 -1164
rect 1674 -1176 1680 -1170
rect 1674 -1182 1680 -1176
rect 1674 -1188 1680 -1182
rect 1674 -1194 1680 -1188
rect 1674 -1200 1680 -1194
rect 1674 -1206 1680 -1200
rect 1674 -1212 1680 -1206
rect 1674 -1218 1680 -1212
rect 1674 -1224 1680 -1218
rect 1674 -1230 1680 -1224
rect 1674 -1236 1680 -1230
rect 1674 -1242 1680 -1236
rect 1674 -1248 1680 -1242
rect 1674 -1254 1680 -1248
rect 1674 -1260 1680 -1254
rect 1674 -1266 1680 -1260
rect 1674 -1272 1680 -1266
rect 1674 -1278 1680 -1272
rect 1674 -1284 1680 -1278
rect 1674 -1290 1680 -1284
rect 1674 -1296 1680 -1290
rect 1674 -1302 1680 -1296
rect 1674 -1308 1680 -1302
rect 1674 -1314 1680 -1308
rect 1674 -1320 1680 -1314
rect 1674 -1326 1680 -1320
rect 1674 -1332 1680 -1326
rect 1674 -1338 1680 -1332
rect 1674 -1344 1680 -1338
rect 1674 -1350 1680 -1344
rect 1674 -1356 1680 -1350
rect 1674 -1362 1680 -1356
rect 1674 -1368 1680 -1362
rect 1674 -1374 1680 -1368
rect 1674 -1380 1680 -1374
rect 1674 -1386 1680 -1380
rect 1674 -1392 1680 -1386
rect 1674 -1398 1680 -1392
rect 1674 -1404 1680 -1398
rect 1674 -1410 1680 -1404
rect 1674 -1416 1680 -1410
rect 1674 -1422 1680 -1416
rect 1674 -1428 1680 -1422
rect 1674 -1434 1680 -1428
rect 1674 -1440 1680 -1434
rect 1674 -1446 1680 -1440
rect 1674 -1452 1680 -1446
rect 1674 -1458 1680 -1452
rect 1674 -1464 1680 -1458
rect 1674 -1470 1680 -1464
rect 1674 -1476 1680 -1470
rect 1674 -1482 1680 -1476
rect 1674 -1488 1680 -1482
rect 1674 -1494 1680 -1488
rect 1674 -1500 1680 -1494
rect 1674 -1506 1680 -1500
rect 1674 -1512 1680 -1506
rect 1674 -1518 1680 -1512
rect 1674 -1524 1680 -1518
rect 1674 -1530 1680 -1524
rect 1674 -1536 1680 -1530
rect 1674 -1542 1680 -1536
rect 1674 -1548 1680 -1542
rect 1674 -1554 1680 -1548
rect 1674 -1560 1680 -1554
rect 1674 -1566 1680 -1560
rect 1674 -1572 1680 -1566
rect 1674 -1578 1680 -1572
rect 1674 -1584 1680 -1578
rect 1674 -1590 1680 -1584
rect 1674 -1596 1680 -1590
rect 1674 -1602 1680 -1596
rect 1674 -1608 1680 -1602
rect 1674 -1614 1680 -1608
rect 1674 -1620 1680 -1614
rect 1674 -1626 1680 -1620
rect 1674 -1632 1680 -1626
rect 1674 -1638 1680 -1632
rect 1674 -1644 1680 -1638
rect 1674 -1650 1680 -1644
rect 1674 -1656 1680 -1650
rect 1674 -1662 1680 -1656
rect 1674 -1668 1680 -1662
rect 1674 -1674 1680 -1668
rect 1674 -1680 1680 -1674
rect 1674 -1686 1680 -1680
rect 1674 -1692 1680 -1686
rect 1674 -1698 1680 -1692
rect 1674 -1704 1680 -1698
rect 1674 -1710 1680 -1704
rect 1674 -1716 1680 -1710
rect 1674 -1722 1680 -1716
rect 1674 -1728 1680 -1722
rect 1674 -1734 1680 -1728
rect 1674 -1740 1680 -1734
rect 1674 -1746 1680 -1740
rect 1674 -1752 1680 -1746
rect 1674 -1758 1680 -1752
rect 1674 -1764 1680 -1758
rect 1674 -1770 1680 -1764
rect 1674 -1776 1680 -1770
rect 1674 -1782 1680 -1776
rect 1674 -1788 1680 -1782
rect 1674 -1794 1680 -1788
rect 1674 -1800 1680 -1794
rect 1674 -1806 1680 -1800
rect 1674 -1812 1680 -1806
rect 1674 -1818 1680 -1812
rect 1674 -1824 1680 -1818
rect 1674 -1830 1680 -1824
rect 1674 -1836 1680 -1830
rect 1674 -1842 1680 -1836
rect 1674 -1848 1680 -1842
rect 1674 -1854 1680 -1848
rect 1674 -1860 1680 -1854
rect 1674 -1866 1680 -1860
rect 1674 -1872 1680 -1866
rect 1674 -1878 1680 -1872
rect 1674 -1884 1680 -1878
rect 1674 -1890 1680 -1884
rect 1674 -1896 1680 -1890
rect 1674 -1902 1680 -1896
rect 1674 -1908 1680 -1902
rect 1674 -1914 1680 -1908
rect 1674 -1920 1680 -1914
rect 1674 -1926 1680 -1920
rect 1674 -1932 1680 -1926
rect 1674 -1938 1680 -1932
rect 1674 -1944 1680 -1938
rect 1674 -1950 1680 -1944
rect 1674 -1956 1680 -1950
rect 1674 -1962 1680 -1956
rect 1674 -1968 1680 -1962
rect 1674 -1974 1680 -1968
rect 1674 -1980 1680 -1974
rect 1674 -2058 1680 -2052
rect 1674 -2064 1680 -2058
rect 1674 -2070 1680 -2064
rect 1674 -2076 1680 -2070
rect 1674 -2082 1680 -2076
rect 1674 -2088 1680 -2082
rect 1674 -2094 1680 -2088
rect 1674 -2100 1680 -2094
rect 1674 -2106 1680 -2100
rect 1674 -2112 1680 -2106
rect 1674 -2118 1680 -2112
rect 1674 -2124 1680 -2118
rect 1674 -2130 1680 -2124
rect 1674 -2136 1680 -2130
rect 1674 -2142 1680 -2136
rect 1674 -2148 1680 -2142
rect 1674 -2154 1680 -2148
rect 1674 -2160 1680 -2154
rect 1674 -2166 1680 -2160
rect 1674 -2172 1680 -2166
rect 1674 -2178 1680 -2172
rect 1674 -2184 1680 -2178
rect 1674 -2190 1680 -2184
rect 1674 -2196 1680 -2190
rect 1674 -2202 1680 -2196
rect 1674 -2208 1680 -2202
rect 1674 -2214 1680 -2208
rect 1674 -2220 1680 -2214
rect 1674 -2226 1680 -2220
rect 1674 -2232 1680 -2226
rect 1674 -2238 1680 -2232
rect 1674 -2244 1680 -2238
rect 1674 -2250 1680 -2244
rect 1674 -2256 1680 -2250
rect 1674 -2262 1680 -2256
rect 1674 -2268 1680 -2262
rect 1674 -2274 1680 -2268
rect 1674 -2280 1680 -2274
rect 1674 -2286 1680 -2280
rect 1674 -2292 1680 -2286
rect 1674 -2298 1680 -2292
rect 1674 -2304 1680 -2298
rect 1674 -2310 1680 -2304
rect 1674 -2316 1680 -2310
rect 1674 -2322 1680 -2316
rect 1674 -2328 1680 -2322
rect 1674 -2334 1680 -2328
rect 1674 -2340 1680 -2334
rect 1674 -2346 1680 -2340
rect 1674 -2352 1680 -2346
rect 1674 -2358 1680 -2352
rect 1674 -2364 1680 -2358
rect 1674 -2370 1680 -2364
rect 1674 -2376 1680 -2370
rect 1674 -2382 1680 -2376
rect 1674 -2388 1680 -2382
rect 1674 -2394 1680 -2388
rect 1674 -2400 1680 -2394
rect 1674 -2406 1680 -2400
rect 1674 -2412 1680 -2406
rect 1674 -2418 1680 -2412
rect 1674 -2424 1680 -2418
rect 1674 -2430 1680 -2424
rect 1674 -2436 1680 -2430
rect 1674 -2442 1680 -2436
rect 1674 -2448 1680 -2442
rect 1674 -2454 1680 -2448
rect 1674 -2460 1680 -2454
rect 1674 -2466 1680 -2460
rect 1674 -2472 1680 -2466
rect 1674 -2478 1680 -2472
rect 1674 -2484 1680 -2478
rect 1674 -2490 1680 -2484
rect 1674 -2496 1680 -2490
rect 1674 -2502 1680 -2496
rect 1674 -2508 1680 -2502
rect 1674 -2514 1680 -2508
rect 1674 -2520 1680 -2514
rect 1674 -2526 1680 -2520
rect 1674 -2532 1680 -2526
rect 1674 -2538 1680 -2532
rect 1674 -2544 1680 -2538
rect 1674 -2550 1680 -2544
rect 1674 -2556 1680 -2550
rect 1674 -2562 1680 -2556
rect 1674 -2568 1680 -2562
rect 1674 -2574 1680 -2568
rect 1674 -2580 1680 -2574
rect 1674 -2586 1680 -2580
rect 1674 -2592 1680 -2586
rect 1674 -2598 1680 -2592
rect 1674 -2604 1680 -2598
rect 1674 -2610 1680 -2604
rect 1674 -2616 1680 -2610
rect 1674 -2622 1680 -2616
rect 1674 -2628 1680 -2622
rect 1674 -2634 1680 -2628
rect 1674 -2640 1680 -2634
rect 1674 -2646 1680 -2640
rect 1674 -2652 1680 -2646
rect 1674 -2658 1680 -2652
rect 1674 -2664 1680 -2658
rect 1674 -2670 1680 -2664
rect 1674 -2676 1680 -2670
rect 1674 -2682 1680 -2676
rect 1674 -2688 1680 -2682
rect 1674 -2694 1680 -2688
rect 1674 -2700 1680 -2694
rect 1674 -2778 1680 -2772
rect 1674 -2784 1680 -2778
rect 1674 -2790 1680 -2784
rect 1674 -2796 1680 -2790
rect 1674 -2802 1680 -2796
rect 1674 -2808 1680 -2802
rect 1674 -2814 1680 -2808
rect 1674 -2820 1680 -2814
rect 1674 -2826 1680 -2820
rect 1674 -2832 1680 -2826
rect 1674 -2838 1680 -2832
rect 1674 -2844 1680 -2838
rect 1674 -2850 1680 -2844
rect 1674 -2856 1680 -2850
rect 1674 -2862 1680 -2856
rect 1674 -2868 1680 -2862
rect 1674 -2874 1680 -2868
rect 1674 -2880 1680 -2874
rect 1674 -2886 1680 -2880
rect 1674 -2892 1680 -2886
rect 1674 -2898 1680 -2892
rect 1674 -2904 1680 -2898
rect 1674 -2910 1680 -2904
rect 1674 -2916 1680 -2910
rect 1674 -2922 1680 -2916
rect 1674 -2928 1680 -2922
rect 1674 -2934 1680 -2928
rect 1674 -2940 1680 -2934
rect 1674 -2946 1680 -2940
rect 1674 -2952 1680 -2946
rect 1674 -2958 1680 -2952
rect 1674 -2964 1680 -2958
rect 1674 -2970 1680 -2964
rect 1674 -2976 1680 -2970
rect 1674 -2982 1680 -2976
rect 1674 -2988 1680 -2982
rect 1674 -2994 1680 -2988
rect 1674 -3000 1680 -2994
rect 1674 -3006 1680 -3000
rect 1674 -3012 1680 -3006
rect 1674 -3018 1680 -3012
rect 1674 -3024 1680 -3018
rect 1674 -3030 1680 -3024
rect 1674 -3036 1680 -3030
rect 1674 -3042 1680 -3036
rect 1674 -3048 1680 -3042
rect 1674 -3054 1680 -3048
rect 1674 -3060 1680 -3054
rect 1674 -3066 1680 -3060
rect 1674 -3072 1680 -3066
rect 1674 -3078 1680 -3072
rect 1674 -3084 1680 -3078
rect 1674 -3090 1680 -3084
rect 1674 -3096 1680 -3090
rect 1674 -3102 1680 -3096
rect 1674 -3108 1680 -3102
rect 1674 -3114 1680 -3108
rect 1674 -3120 1680 -3114
rect 1674 -3126 1680 -3120
rect 1674 -3132 1680 -3126
rect 1674 -3138 1680 -3132
rect 1674 -3144 1680 -3138
rect 1674 -3150 1680 -3144
rect 1674 -3156 1680 -3150
rect 1674 -3162 1680 -3156
rect 1674 -3168 1680 -3162
rect 1674 -3174 1680 -3168
rect 1674 -3180 1680 -3174
rect 1674 -3186 1680 -3180
rect 1674 -3192 1680 -3186
rect 1674 -3198 1680 -3192
rect 1674 -3204 1680 -3198
rect 1674 -3210 1680 -3204
rect 1674 -3216 1680 -3210
rect 1674 -3222 1680 -3216
rect 1674 -3228 1680 -3222
rect 1674 -3234 1680 -3228
rect 1674 -3276 1680 -3270
rect 1674 -3282 1680 -3276
rect 1674 -3288 1680 -3282
rect 1674 -3294 1680 -3288
rect 1674 -3300 1680 -3294
rect 1674 -3306 1680 -3300
rect 1674 -3312 1680 -3306
rect 1674 -3318 1680 -3312
rect 1674 -3324 1680 -3318
rect 1674 -3330 1680 -3324
rect 1674 -3336 1680 -3330
rect 1674 -3342 1680 -3336
rect 1674 -3348 1680 -3342
rect 1674 -3354 1680 -3348
rect 1674 -3360 1680 -3354
rect 1674 -3366 1680 -3360
rect 1674 -3372 1680 -3366
rect 1674 -3378 1680 -3372
rect 1674 -3384 1680 -3378
rect 1674 -3390 1680 -3384
rect 1674 -3396 1680 -3390
rect 1674 -3402 1680 -3396
rect 1674 -3408 1680 -3402
rect 1674 -3414 1680 -3408
rect 1674 -3420 1680 -3414
rect 1674 -3426 1680 -3420
rect 1674 -3432 1680 -3426
rect 1680 -894 1686 -888
rect 1680 -900 1686 -894
rect 1680 -906 1686 -900
rect 1680 -912 1686 -906
rect 1680 -918 1686 -912
rect 1680 -924 1686 -918
rect 1680 -930 1686 -924
rect 1680 -936 1686 -930
rect 1680 -942 1686 -936
rect 1680 -948 1686 -942
rect 1680 -954 1686 -948
rect 1680 -960 1686 -954
rect 1680 -966 1686 -960
rect 1680 -972 1686 -966
rect 1680 -978 1686 -972
rect 1680 -984 1686 -978
rect 1680 -990 1686 -984
rect 1680 -996 1686 -990
rect 1680 -1002 1686 -996
rect 1680 -1008 1686 -1002
rect 1680 -1014 1686 -1008
rect 1680 -1020 1686 -1014
rect 1680 -1026 1686 -1020
rect 1680 -1032 1686 -1026
rect 1680 -1038 1686 -1032
rect 1680 -1044 1686 -1038
rect 1680 -1050 1686 -1044
rect 1680 -1056 1686 -1050
rect 1680 -1062 1686 -1056
rect 1680 -1068 1686 -1062
rect 1680 -1074 1686 -1068
rect 1680 -1080 1686 -1074
rect 1680 -1086 1686 -1080
rect 1680 -1092 1686 -1086
rect 1680 -1098 1686 -1092
rect 1680 -1104 1686 -1098
rect 1680 -1110 1686 -1104
rect 1680 -1116 1686 -1110
rect 1680 -1122 1686 -1116
rect 1680 -1128 1686 -1122
rect 1680 -1134 1686 -1128
rect 1680 -1140 1686 -1134
rect 1680 -1146 1686 -1140
rect 1680 -1152 1686 -1146
rect 1680 -1158 1686 -1152
rect 1680 -1164 1686 -1158
rect 1680 -1170 1686 -1164
rect 1680 -1176 1686 -1170
rect 1680 -1182 1686 -1176
rect 1680 -1188 1686 -1182
rect 1680 -1194 1686 -1188
rect 1680 -1200 1686 -1194
rect 1680 -1206 1686 -1200
rect 1680 -1212 1686 -1206
rect 1680 -1218 1686 -1212
rect 1680 -1224 1686 -1218
rect 1680 -1230 1686 -1224
rect 1680 -1236 1686 -1230
rect 1680 -1242 1686 -1236
rect 1680 -1248 1686 -1242
rect 1680 -1254 1686 -1248
rect 1680 -1260 1686 -1254
rect 1680 -1266 1686 -1260
rect 1680 -1272 1686 -1266
rect 1680 -1278 1686 -1272
rect 1680 -1284 1686 -1278
rect 1680 -1290 1686 -1284
rect 1680 -1296 1686 -1290
rect 1680 -1302 1686 -1296
rect 1680 -1308 1686 -1302
rect 1680 -1314 1686 -1308
rect 1680 -1320 1686 -1314
rect 1680 -1326 1686 -1320
rect 1680 -1332 1686 -1326
rect 1680 -1338 1686 -1332
rect 1680 -1344 1686 -1338
rect 1680 -1350 1686 -1344
rect 1680 -1356 1686 -1350
rect 1680 -1362 1686 -1356
rect 1680 -1368 1686 -1362
rect 1680 -1374 1686 -1368
rect 1680 -1380 1686 -1374
rect 1680 -1386 1686 -1380
rect 1680 -1392 1686 -1386
rect 1680 -1398 1686 -1392
rect 1680 -1404 1686 -1398
rect 1680 -1410 1686 -1404
rect 1680 -1416 1686 -1410
rect 1680 -1422 1686 -1416
rect 1680 -1428 1686 -1422
rect 1680 -1434 1686 -1428
rect 1680 -1440 1686 -1434
rect 1680 -1446 1686 -1440
rect 1680 -1452 1686 -1446
rect 1680 -1458 1686 -1452
rect 1680 -1464 1686 -1458
rect 1680 -1470 1686 -1464
rect 1680 -1476 1686 -1470
rect 1680 -1482 1686 -1476
rect 1680 -1488 1686 -1482
rect 1680 -1494 1686 -1488
rect 1680 -1500 1686 -1494
rect 1680 -1506 1686 -1500
rect 1680 -1512 1686 -1506
rect 1680 -1518 1686 -1512
rect 1680 -1524 1686 -1518
rect 1680 -1530 1686 -1524
rect 1680 -1536 1686 -1530
rect 1680 -1542 1686 -1536
rect 1680 -1548 1686 -1542
rect 1680 -1554 1686 -1548
rect 1680 -1560 1686 -1554
rect 1680 -1566 1686 -1560
rect 1680 -1572 1686 -1566
rect 1680 -1578 1686 -1572
rect 1680 -1584 1686 -1578
rect 1680 -1590 1686 -1584
rect 1680 -1596 1686 -1590
rect 1680 -1602 1686 -1596
rect 1680 -1608 1686 -1602
rect 1680 -1614 1686 -1608
rect 1680 -1620 1686 -1614
rect 1680 -1626 1686 -1620
rect 1680 -1632 1686 -1626
rect 1680 -1638 1686 -1632
rect 1680 -1644 1686 -1638
rect 1680 -1650 1686 -1644
rect 1680 -1656 1686 -1650
rect 1680 -1662 1686 -1656
rect 1680 -1668 1686 -1662
rect 1680 -1674 1686 -1668
rect 1680 -1680 1686 -1674
rect 1680 -1686 1686 -1680
rect 1680 -1692 1686 -1686
rect 1680 -1698 1686 -1692
rect 1680 -1704 1686 -1698
rect 1680 -1710 1686 -1704
rect 1680 -1716 1686 -1710
rect 1680 -1722 1686 -1716
rect 1680 -1728 1686 -1722
rect 1680 -1734 1686 -1728
rect 1680 -1740 1686 -1734
rect 1680 -1746 1686 -1740
rect 1680 -1752 1686 -1746
rect 1680 -1758 1686 -1752
rect 1680 -1764 1686 -1758
rect 1680 -1770 1686 -1764
rect 1680 -1776 1686 -1770
rect 1680 -1782 1686 -1776
rect 1680 -1788 1686 -1782
rect 1680 -1794 1686 -1788
rect 1680 -1800 1686 -1794
rect 1680 -1806 1686 -1800
rect 1680 -1812 1686 -1806
rect 1680 -1818 1686 -1812
rect 1680 -1824 1686 -1818
rect 1680 -1830 1686 -1824
rect 1680 -1836 1686 -1830
rect 1680 -1842 1686 -1836
rect 1680 -1848 1686 -1842
rect 1680 -1854 1686 -1848
rect 1680 -1860 1686 -1854
rect 1680 -1866 1686 -1860
rect 1680 -1872 1686 -1866
rect 1680 -1878 1686 -1872
rect 1680 -1884 1686 -1878
rect 1680 -1890 1686 -1884
rect 1680 -1896 1686 -1890
rect 1680 -1902 1686 -1896
rect 1680 -1908 1686 -1902
rect 1680 -1914 1686 -1908
rect 1680 -1920 1686 -1914
rect 1680 -1926 1686 -1920
rect 1680 -1932 1686 -1926
rect 1680 -1938 1686 -1932
rect 1680 -1944 1686 -1938
rect 1680 -1950 1686 -1944
rect 1680 -1956 1686 -1950
rect 1680 -1962 1686 -1956
rect 1680 -1968 1686 -1962
rect 1680 -1974 1686 -1968
rect 1680 -2052 1686 -2046
rect 1680 -2058 1686 -2052
rect 1680 -2064 1686 -2058
rect 1680 -2070 1686 -2064
rect 1680 -2076 1686 -2070
rect 1680 -2082 1686 -2076
rect 1680 -2088 1686 -2082
rect 1680 -2094 1686 -2088
rect 1680 -2100 1686 -2094
rect 1680 -2106 1686 -2100
rect 1680 -2112 1686 -2106
rect 1680 -2118 1686 -2112
rect 1680 -2124 1686 -2118
rect 1680 -2130 1686 -2124
rect 1680 -2136 1686 -2130
rect 1680 -2142 1686 -2136
rect 1680 -2148 1686 -2142
rect 1680 -2154 1686 -2148
rect 1680 -2160 1686 -2154
rect 1680 -2166 1686 -2160
rect 1680 -2172 1686 -2166
rect 1680 -2178 1686 -2172
rect 1680 -2184 1686 -2178
rect 1680 -2190 1686 -2184
rect 1680 -2196 1686 -2190
rect 1680 -2202 1686 -2196
rect 1680 -2208 1686 -2202
rect 1680 -2214 1686 -2208
rect 1680 -2220 1686 -2214
rect 1680 -2226 1686 -2220
rect 1680 -2232 1686 -2226
rect 1680 -2238 1686 -2232
rect 1680 -2244 1686 -2238
rect 1680 -2250 1686 -2244
rect 1680 -2256 1686 -2250
rect 1680 -2262 1686 -2256
rect 1680 -2268 1686 -2262
rect 1680 -2274 1686 -2268
rect 1680 -2280 1686 -2274
rect 1680 -2286 1686 -2280
rect 1680 -2292 1686 -2286
rect 1680 -2298 1686 -2292
rect 1680 -2304 1686 -2298
rect 1680 -2310 1686 -2304
rect 1680 -2316 1686 -2310
rect 1680 -2322 1686 -2316
rect 1680 -2328 1686 -2322
rect 1680 -2334 1686 -2328
rect 1680 -2340 1686 -2334
rect 1680 -2346 1686 -2340
rect 1680 -2352 1686 -2346
rect 1680 -2358 1686 -2352
rect 1680 -2364 1686 -2358
rect 1680 -2370 1686 -2364
rect 1680 -2376 1686 -2370
rect 1680 -2382 1686 -2376
rect 1680 -2388 1686 -2382
rect 1680 -2394 1686 -2388
rect 1680 -2400 1686 -2394
rect 1680 -2406 1686 -2400
rect 1680 -2412 1686 -2406
rect 1680 -2418 1686 -2412
rect 1680 -2424 1686 -2418
rect 1680 -2430 1686 -2424
rect 1680 -2436 1686 -2430
rect 1680 -2442 1686 -2436
rect 1680 -2448 1686 -2442
rect 1680 -2454 1686 -2448
rect 1680 -2460 1686 -2454
rect 1680 -2466 1686 -2460
rect 1680 -2472 1686 -2466
rect 1680 -2478 1686 -2472
rect 1680 -2484 1686 -2478
rect 1680 -2490 1686 -2484
rect 1680 -2496 1686 -2490
rect 1680 -2502 1686 -2496
rect 1680 -2508 1686 -2502
rect 1680 -2514 1686 -2508
rect 1680 -2520 1686 -2514
rect 1680 -2526 1686 -2520
rect 1680 -2532 1686 -2526
rect 1680 -2538 1686 -2532
rect 1680 -2544 1686 -2538
rect 1680 -2550 1686 -2544
rect 1680 -2556 1686 -2550
rect 1680 -2562 1686 -2556
rect 1680 -2568 1686 -2562
rect 1680 -2574 1686 -2568
rect 1680 -2580 1686 -2574
rect 1680 -2586 1686 -2580
rect 1680 -2592 1686 -2586
rect 1680 -2598 1686 -2592
rect 1680 -2604 1686 -2598
rect 1680 -2610 1686 -2604
rect 1680 -2616 1686 -2610
rect 1680 -2622 1686 -2616
rect 1680 -2628 1686 -2622
rect 1680 -2634 1686 -2628
rect 1680 -2640 1686 -2634
rect 1680 -2646 1686 -2640
rect 1680 -2652 1686 -2646
rect 1680 -2658 1686 -2652
rect 1680 -2664 1686 -2658
rect 1680 -2670 1686 -2664
rect 1680 -2676 1686 -2670
rect 1680 -2682 1686 -2676
rect 1680 -2688 1686 -2682
rect 1680 -2694 1686 -2688
rect 1680 -2700 1686 -2694
rect 1680 -2778 1686 -2772
rect 1680 -2784 1686 -2778
rect 1680 -2790 1686 -2784
rect 1680 -2796 1686 -2790
rect 1680 -2802 1686 -2796
rect 1680 -2808 1686 -2802
rect 1680 -2814 1686 -2808
rect 1680 -2820 1686 -2814
rect 1680 -2826 1686 -2820
rect 1680 -2832 1686 -2826
rect 1680 -2838 1686 -2832
rect 1680 -2844 1686 -2838
rect 1680 -2850 1686 -2844
rect 1680 -2856 1686 -2850
rect 1680 -2862 1686 -2856
rect 1680 -2868 1686 -2862
rect 1680 -2874 1686 -2868
rect 1680 -2880 1686 -2874
rect 1680 -2886 1686 -2880
rect 1680 -2892 1686 -2886
rect 1680 -2898 1686 -2892
rect 1680 -2904 1686 -2898
rect 1680 -2910 1686 -2904
rect 1680 -2916 1686 -2910
rect 1680 -2922 1686 -2916
rect 1680 -2928 1686 -2922
rect 1680 -2934 1686 -2928
rect 1680 -2940 1686 -2934
rect 1680 -2946 1686 -2940
rect 1680 -2952 1686 -2946
rect 1680 -2958 1686 -2952
rect 1680 -2964 1686 -2958
rect 1680 -2970 1686 -2964
rect 1680 -2976 1686 -2970
rect 1680 -2982 1686 -2976
rect 1680 -2988 1686 -2982
rect 1680 -2994 1686 -2988
rect 1680 -3000 1686 -2994
rect 1680 -3006 1686 -3000
rect 1680 -3012 1686 -3006
rect 1680 -3018 1686 -3012
rect 1680 -3024 1686 -3018
rect 1680 -3030 1686 -3024
rect 1680 -3036 1686 -3030
rect 1680 -3042 1686 -3036
rect 1680 -3048 1686 -3042
rect 1680 -3054 1686 -3048
rect 1680 -3060 1686 -3054
rect 1680 -3066 1686 -3060
rect 1680 -3072 1686 -3066
rect 1680 -3078 1686 -3072
rect 1680 -3084 1686 -3078
rect 1680 -3090 1686 -3084
rect 1680 -3096 1686 -3090
rect 1680 -3102 1686 -3096
rect 1680 -3108 1686 -3102
rect 1680 -3114 1686 -3108
rect 1680 -3120 1686 -3114
rect 1680 -3126 1686 -3120
rect 1680 -3132 1686 -3126
rect 1680 -3138 1686 -3132
rect 1680 -3144 1686 -3138
rect 1680 -3150 1686 -3144
rect 1680 -3156 1686 -3150
rect 1680 -3162 1686 -3156
rect 1680 -3168 1686 -3162
rect 1680 -3174 1686 -3168
rect 1680 -3180 1686 -3174
rect 1680 -3186 1686 -3180
rect 1680 -3192 1686 -3186
rect 1680 -3198 1686 -3192
rect 1680 -3204 1686 -3198
rect 1680 -3210 1686 -3204
rect 1680 -3216 1686 -3210
rect 1680 -3222 1686 -3216
rect 1680 -3228 1686 -3222
rect 1680 -3276 1686 -3270
rect 1680 -3282 1686 -3276
rect 1680 -3288 1686 -3282
rect 1680 -3294 1686 -3288
rect 1680 -3300 1686 -3294
rect 1680 -3306 1686 -3300
rect 1680 -3312 1686 -3306
rect 1680 -3318 1686 -3312
rect 1680 -3324 1686 -3318
rect 1680 -3330 1686 -3324
rect 1680 -3336 1686 -3330
rect 1680 -3342 1686 -3336
rect 1680 -3348 1686 -3342
rect 1680 -3354 1686 -3348
rect 1680 -3360 1686 -3354
rect 1680 -3366 1686 -3360
rect 1680 -3372 1686 -3366
rect 1680 -3378 1686 -3372
rect 1680 -3384 1686 -3378
rect 1680 -3390 1686 -3384
rect 1680 -3396 1686 -3390
rect 1680 -3402 1686 -3396
rect 1680 -3408 1686 -3402
rect 1680 -3414 1686 -3408
rect 1680 -3420 1686 -3414
rect 1680 -3426 1686 -3420
rect 1686 -882 1692 -876
rect 1686 -888 1692 -882
rect 1686 -894 1692 -888
rect 1686 -900 1692 -894
rect 1686 -906 1692 -900
rect 1686 -912 1692 -906
rect 1686 -918 1692 -912
rect 1686 -924 1692 -918
rect 1686 -930 1692 -924
rect 1686 -936 1692 -930
rect 1686 -942 1692 -936
rect 1686 -948 1692 -942
rect 1686 -954 1692 -948
rect 1686 -960 1692 -954
rect 1686 -966 1692 -960
rect 1686 -972 1692 -966
rect 1686 -978 1692 -972
rect 1686 -984 1692 -978
rect 1686 -990 1692 -984
rect 1686 -996 1692 -990
rect 1686 -1002 1692 -996
rect 1686 -1008 1692 -1002
rect 1686 -1014 1692 -1008
rect 1686 -1020 1692 -1014
rect 1686 -1026 1692 -1020
rect 1686 -1032 1692 -1026
rect 1686 -1038 1692 -1032
rect 1686 -1044 1692 -1038
rect 1686 -1050 1692 -1044
rect 1686 -1056 1692 -1050
rect 1686 -1062 1692 -1056
rect 1686 -1068 1692 -1062
rect 1686 -1074 1692 -1068
rect 1686 -1080 1692 -1074
rect 1686 -1086 1692 -1080
rect 1686 -1092 1692 -1086
rect 1686 -1098 1692 -1092
rect 1686 -1104 1692 -1098
rect 1686 -1110 1692 -1104
rect 1686 -1116 1692 -1110
rect 1686 -1122 1692 -1116
rect 1686 -1128 1692 -1122
rect 1686 -1134 1692 -1128
rect 1686 -1140 1692 -1134
rect 1686 -1146 1692 -1140
rect 1686 -1152 1692 -1146
rect 1686 -1158 1692 -1152
rect 1686 -1164 1692 -1158
rect 1686 -1170 1692 -1164
rect 1686 -1176 1692 -1170
rect 1686 -1182 1692 -1176
rect 1686 -1188 1692 -1182
rect 1686 -1194 1692 -1188
rect 1686 -1200 1692 -1194
rect 1686 -1206 1692 -1200
rect 1686 -1212 1692 -1206
rect 1686 -1218 1692 -1212
rect 1686 -1224 1692 -1218
rect 1686 -1230 1692 -1224
rect 1686 -1236 1692 -1230
rect 1686 -1242 1692 -1236
rect 1686 -1248 1692 -1242
rect 1686 -1254 1692 -1248
rect 1686 -1260 1692 -1254
rect 1686 -1266 1692 -1260
rect 1686 -1272 1692 -1266
rect 1686 -1278 1692 -1272
rect 1686 -1284 1692 -1278
rect 1686 -1290 1692 -1284
rect 1686 -1296 1692 -1290
rect 1686 -1302 1692 -1296
rect 1686 -1308 1692 -1302
rect 1686 -1314 1692 -1308
rect 1686 -1320 1692 -1314
rect 1686 -1326 1692 -1320
rect 1686 -1332 1692 -1326
rect 1686 -1338 1692 -1332
rect 1686 -1344 1692 -1338
rect 1686 -1350 1692 -1344
rect 1686 -1356 1692 -1350
rect 1686 -1362 1692 -1356
rect 1686 -1368 1692 -1362
rect 1686 -1374 1692 -1368
rect 1686 -1380 1692 -1374
rect 1686 -1386 1692 -1380
rect 1686 -1392 1692 -1386
rect 1686 -1398 1692 -1392
rect 1686 -1404 1692 -1398
rect 1686 -1410 1692 -1404
rect 1686 -1416 1692 -1410
rect 1686 -1422 1692 -1416
rect 1686 -1428 1692 -1422
rect 1686 -1434 1692 -1428
rect 1686 -1440 1692 -1434
rect 1686 -1446 1692 -1440
rect 1686 -1452 1692 -1446
rect 1686 -1458 1692 -1452
rect 1686 -1464 1692 -1458
rect 1686 -1470 1692 -1464
rect 1686 -1476 1692 -1470
rect 1686 -1482 1692 -1476
rect 1686 -1488 1692 -1482
rect 1686 -1494 1692 -1488
rect 1686 -1500 1692 -1494
rect 1686 -1506 1692 -1500
rect 1686 -1512 1692 -1506
rect 1686 -1518 1692 -1512
rect 1686 -1524 1692 -1518
rect 1686 -1530 1692 -1524
rect 1686 -1536 1692 -1530
rect 1686 -1542 1692 -1536
rect 1686 -1548 1692 -1542
rect 1686 -1554 1692 -1548
rect 1686 -1560 1692 -1554
rect 1686 -1566 1692 -1560
rect 1686 -1572 1692 -1566
rect 1686 -1578 1692 -1572
rect 1686 -1584 1692 -1578
rect 1686 -1590 1692 -1584
rect 1686 -1596 1692 -1590
rect 1686 -1602 1692 -1596
rect 1686 -1608 1692 -1602
rect 1686 -1614 1692 -1608
rect 1686 -1620 1692 -1614
rect 1686 -1626 1692 -1620
rect 1686 -1632 1692 -1626
rect 1686 -1638 1692 -1632
rect 1686 -1644 1692 -1638
rect 1686 -1650 1692 -1644
rect 1686 -1656 1692 -1650
rect 1686 -1662 1692 -1656
rect 1686 -1668 1692 -1662
rect 1686 -1674 1692 -1668
rect 1686 -1680 1692 -1674
rect 1686 -1686 1692 -1680
rect 1686 -1692 1692 -1686
rect 1686 -1698 1692 -1692
rect 1686 -1704 1692 -1698
rect 1686 -1710 1692 -1704
rect 1686 -1716 1692 -1710
rect 1686 -1722 1692 -1716
rect 1686 -1728 1692 -1722
rect 1686 -1734 1692 -1728
rect 1686 -1740 1692 -1734
rect 1686 -1746 1692 -1740
rect 1686 -1752 1692 -1746
rect 1686 -1758 1692 -1752
rect 1686 -1764 1692 -1758
rect 1686 -1770 1692 -1764
rect 1686 -1776 1692 -1770
rect 1686 -1782 1692 -1776
rect 1686 -1788 1692 -1782
rect 1686 -1794 1692 -1788
rect 1686 -1800 1692 -1794
rect 1686 -1806 1692 -1800
rect 1686 -1812 1692 -1806
rect 1686 -1818 1692 -1812
rect 1686 -1824 1692 -1818
rect 1686 -1830 1692 -1824
rect 1686 -1836 1692 -1830
rect 1686 -1842 1692 -1836
rect 1686 -1848 1692 -1842
rect 1686 -1854 1692 -1848
rect 1686 -1860 1692 -1854
rect 1686 -1866 1692 -1860
rect 1686 -1872 1692 -1866
rect 1686 -1878 1692 -1872
rect 1686 -1884 1692 -1878
rect 1686 -1890 1692 -1884
rect 1686 -1896 1692 -1890
rect 1686 -1902 1692 -1896
rect 1686 -1908 1692 -1902
rect 1686 -1914 1692 -1908
rect 1686 -1920 1692 -1914
rect 1686 -1926 1692 -1920
rect 1686 -1932 1692 -1926
rect 1686 -1938 1692 -1932
rect 1686 -1944 1692 -1938
rect 1686 -1950 1692 -1944
rect 1686 -1956 1692 -1950
rect 1686 -1962 1692 -1956
rect 1686 -1968 1692 -1962
rect 1686 -2046 1692 -2040
rect 1686 -2052 1692 -2046
rect 1686 -2058 1692 -2052
rect 1686 -2064 1692 -2058
rect 1686 -2070 1692 -2064
rect 1686 -2076 1692 -2070
rect 1686 -2082 1692 -2076
rect 1686 -2088 1692 -2082
rect 1686 -2094 1692 -2088
rect 1686 -2100 1692 -2094
rect 1686 -2106 1692 -2100
rect 1686 -2112 1692 -2106
rect 1686 -2118 1692 -2112
rect 1686 -2124 1692 -2118
rect 1686 -2130 1692 -2124
rect 1686 -2136 1692 -2130
rect 1686 -2142 1692 -2136
rect 1686 -2148 1692 -2142
rect 1686 -2154 1692 -2148
rect 1686 -2160 1692 -2154
rect 1686 -2166 1692 -2160
rect 1686 -2172 1692 -2166
rect 1686 -2178 1692 -2172
rect 1686 -2184 1692 -2178
rect 1686 -2190 1692 -2184
rect 1686 -2196 1692 -2190
rect 1686 -2202 1692 -2196
rect 1686 -2208 1692 -2202
rect 1686 -2214 1692 -2208
rect 1686 -2220 1692 -2214
rect 1686 -2226 1692 -2220
rect 1686 -2232 1692 -2226
rect 1686 -2238 1692 -2232
rect 1686 -2244 1692 -2238
rect 1686 -2250 1692 -2244
rect 1686 -2256 1692 -2250
rect 1686 -2262 1692 -2256
rect 1686 -2268 1692 -2262
rect 1686 -2274 1692 -2268
rect 1686 -2280 1692 -2274
rect 1686 -2286 1692 -2280
rect 1686 -2292 1692 -2286
rect 1686 -2298 1692 -2292
rect 1686 -2304 1692 -2298
rect 1686 -2310 1692 -2304
rect 1686 -2316 1692 -2310
rect 1686 -2322 1692 -2316
rect 1686 -2328 1692 -2322
rect 1686 -2334 1692 -2328
rect 1686 -2340 1692 -2334
rect 1686 -2346 1692 -2340
rect 1686 -2352 1692 -2346
rect 1686 -2358 1692 -2352
rect 1686 -2364 1692 -2358
rect 1686 -2370 1692 -2364
rect 1686 -2376 1692 -2370
rect 1686 -2382 1692 -2376
rect 1686 -2388 1692 -2382
rect 1686 -2394 1692 -2388
rect 1686 -2400 1692 -2394
rect 1686 -2406 1692 -2400
rect 1686 -2412 1692 -2406
rect 1686 -2418 1692 -2412
rect 1686 -2424 1692 -2418
rect 1686 -2430 1692 -2424
rect 1686 -2436 1692 -2430
rect 1686 -2442 1692 -2436
rect 1686 -2448 1692 -2442
rect 1686 -2454 1692 -2448
rect 1686 -2460 1692 -2454
rect 1686 -2466 1692 -2460
rect 1686 -2472 1692 -2466
rect 1686 -2478 1692 -2472
rect 1686 -2484 1692 -2478
rect 1686 -2490 1692 -2484
rect 1686 -2496 1692 -2490
rect 1686 -2502 1692 -2496
rect 1686 -2508 1692 -2502
rect 1686 -2514 1692 -2508
rect 1686 -2520 1692 -2514
rect 1686 -2526 1692 -2520
rect 1686 -2532 1692 -2526
rect 1686 -2538 1692 -2532
rect 1686 -2544 1692 -2538
rect 1686 -2550 1692 -2544
rect 1686 -2556 1692 -2550
rect 1686 -2562 1692 -2556
rect 1686 -2568 1692 -2562
rect 1686 -2574 1692 -2568
rect 1686 -2580 1692 -2574
rect 1686 -2586 1692 -2580
rect 1686 -2592 1692 -2586
rect 1686 -2598 1692 -2592
rect 1686 -2604 1692 -2598
rect 1686 -2610 1692 -2604
rect 1686 -2616 1692 -2610
rect 1686 -2622 1692 -2616
rect 1686 -2628 1692 -2622
rect 1686 -2634 1692 -2628
rect 1686 -2640 1692 -2634
rect 1686 -2646 1692 -2640
rect 1686 -2652 1692 -2646
rect 1686 -2658 1692 -2652
rect 1686 -2664 1692 -2658
rect 1686 -2670 1692 -2664
rect 1686 -2676 1692 -2670
rect 1686 -2682 1692 -2676
rect 1686 -2688 1692 -2682
rect 1686 -2694 1692 -2688
rect 1686 -2772 1692 -2766
rect 1686 -2778 1692 -2772
rect 1686 -2784 1692 -2778
rect 1686 -2790 1692 -2784
rect 1686 -2796 1692 -2790
rect 1686 -2802 1692 -2796
rect 1686 -2808 1692 -2802
rect 1686 -2814 1692 -2808
rect 1686 -2820 1692 -2814
rect 1686 -2826 1692 -2820
rect 1686 -2832 1692 -2826
rect 1686 -2838 1692 -2832
rect 1686 -2844 1692 -2838
rect 1686 -2850 1692 -2844
rect 1686 -2856 1692 -2850
rect 1686 -2862 1692 -2856
rect 1686 -2868 1692 -2862
rect 1686 -2874 1692 -2868
rect 1686 -2880 1692 -2874
rect 1686 -2886 1692 -2880
rect 1686 -2892 1692 -2886
rect 1686 -2898 1692 -2892
rect 1686 -2904 1692 -2898
rect 1686 -2910 1692 -2904
rect 1686 -2916 1692 -2910
rect 1686 -2922 1692 -2916
rect 1686 -2928 1692 -2922
rect 1686 -2934 1692 -2928
rect 1686 -2940 1692 -2934
rect 1686 -2946 1692 -2940
rect 1686 -2952 1692 -2946
rect 1686 -2958 1692 -2952
rect 1686 -2964 1692 -2958
rect 1686 -2970 1692 -2964
rect 1686 -2976 1692 -2970
rect 1686 -2982 1692 -2976
rect 1686 -2988 1692 -2982
rect 1686 -2994 1692 -2988
rect 1686 -3000 1692 -2994
rect 1686 -3006 1692 -3000
rect 1686 -3012 1692 -3006
rect 1686 -3018 1692 -3012
rect 1686 -3024 1692 -3018
rect 1686 -3030 1692 -3024
rect 1686 -3036 1692 -3030
rect 1686 -3042 1692 -3036
rect 1686 -3048 1692 -3042
rect 1686 -3054 1692 -3048
rect 1686 -3060 1692 -3054
rect 1686 -3066 1692 -3060
rect 1686 -3072 1692 -3066
rect 1686 -3078 1692 -3072
rect 1686 -3084 1692 -3078
rect 1686 -3090 1692 -3084
rect 1686 -3096 1692 -3090
rect 1686 -3102 1692 -3096
rect 1686 -3108 1692 -3102
rect 1686 -3114 1692 -3108
rect 1686 -3120 1692 -3114
rect 1686 -3126 1692 -3120
rect 1686 -3132 1692 -3126
rect 1686 -3138 1692 -3132
rect 1686 -3144 1692 -3138
rect 1686 -3150 1692 -3144
rect 1686 -3156 1692 -3150
rect 1686 -3162 1692 -3156
rect 1686 -3168 1692 -3162
rect 1686 -3174 1692 -3168
rect 1686 -3180 1692 -3174
rect 1686 -3186 1692 -3180
rect 1686 -3192 1692 -3186
rect 1686 -3198 1692 -3192
rect 1686 -3204 1692 -3198
rect 1686 -3210 1692 -3204
rect 1686 -3216 1692 -3210
rect 1686 -3222 1692 -3216
rect 1686 -3228 1692 -3222
rect 1686 -3276 1692 -3270
rect 1686 -3282 1692 -3276
rect 1686 -3288 1692 -3282
rect 1686 -3294 1692 -3288
rect 1686 -3300 1692 -3294
rect 1686 -3306 1692 -3300
rect 1686 -3312 1692 -3306
rect 1686 -3318 1692 -3312
rect 1686 -3324 1692 -3318
rect 1686 -3330 1692 -3324
rect 1686 -3336 1692 -3330
rect 1686 -3342 1692 -3336
rect 1686 -3348 1692 -3342
rect 1686 -3354 1692 -3348
rect 1686 -3360 1692 -3354
rect 1686 -3366 1692 -3360
rect 1686 -3372 1692 -3366
rect 1686 -3378 1692 -3372
rect 1686 -3384 1692 -3378
rect 1686 -3390 1692 -3384
rect 1686 -3396 1692 -3390
rect 1686 -3402 1692 -3396
rect 1686 -3408 1692 -3402
rect 1686 -3414 1692 -3408
rect 1686 -3420 1692 -3414
rect 1686 -3426 1692 -3420
rect 1692 -876 1698 -870
rect 1692 -882 1698 -876
rect 1692 -888 1698 -882
rect 1692 -894 1698 -888
rect 1692 -900 1698 -894
rect 1692 -906 1698 -900
rect 1692 -912 1698 -906
rect 1692 -918 1698 -912
rect 1692 -924 1698 -918
rect 1692 -930 1698 -924
rect 1692 -936 1698 -930
rect 1692 -942 1698 -936
rect 1692 -948 1698 -942
rect 1692 -954 1698 -948
rect 1692 -960 1698 -954
rect 1692 -966 1698 -960
rect 1692 -972 1698 -966
rect 1692 -978 1698 -972
rect 1692 -984 1698 -978
rect 1692 -990 1698 -984
rect 1692 -996 1698 -990
rect 1692 -1002 1698 -996
rect 1692 -1008 1698 -1002
rect 1692 -1014 1698 -1008
rect 1692 -1020 1698 -1014
rect 1692 -1026 1698 -1020
rect 1692 -1032 1698 -1026
rect 1692 -1038 1698 -1032
rect 1692 -1044 1698 -1038
rect 1692 -1050 1698 -1044
rect 1692 -1056 1698 -1050
rect 1692 -1062 1698 -1056
rect 1692 -1068 1698 -1062
rect 1692 -1074 1698 -1068
rect 1692 -1080 1698 -1074
rect 1692 -1086 1698 -1080
rect 1692 -1092 1698 -1086
rect 1692 -1098 1698 -1092
rect 1692 -1104 1698 -1098
rect 1692 -1110 1698 -1104
rect 1692 -1116 1698 -1110
rect 1692 -1122 1698 -1116
rect 1692 -1128 1698 -1122
rect 1692 -1134 1698 -1128
rect 1692 -1140 1698 -1134
rect 1692 -1146 1698 -1140
rect 1692 -1152 1698 -1146
rect 1692 -1158 1698 -1152
rect 1692 -1164 1698 -1158
rect 1692 -1170 1698 -1164
rect 1692 -1176 1698 -1170
rect 1692 -1182 1698 -1176
rect 1692 -1188 1698 -1182
rect 1692 -1194 1698 -1188
rect 1692 -1200 1698 -1194
rect 1692 -1206 1698 -1200
rect 1692 -1212 1698 -1206
rect 1692 -1218 1698 -1212
rect 1692 -1224 1698 -1218
rect 1692 -1230 1698 -1224
rect 1692 -1236 1698 -1230
rect 1692 -1242 1698 -1236
rect 1692 -1248 1698 -1242
rect 1692 -1254 1698 -1248
rect 1692 -1260 1698 -1254
rect 1692 -1266 1698 -1260
rect 1692 -1272 1698 -1266
rect 1692 -1278 1698 -1272
rect 1692 -1284 1698 -1278
rect 1692 -1290 1698 -1284
rect 1692 -1296 1698 -1290
rect 1692 -1302 1698 -1296
rect 1692 -1308 1698 -1302
rect 1692 -1314 1698 -1308
rect 1692 -1320 1698 -1314
rect 1692 -1326 1698 -1320
rect 1692 -1332 1698 -1326
rect 1692 -1338 1698 -1332
rect 1692 -1344 1698 -1338
rect 1692 -1350 1698 -1344
rect 1692 -1356 1698 -1350
rect 1692 -1362 1698 -1356
rect 1692 -1368 1698 -1362
rect 1692 -1374 1698 -1368
rect 1692 -1380 1698 -1374
rect 1692 -1386 1698 -1380
rect 1692 -1392 1698 -1386
rect 1692 -1398 1698 -1392
rect 1692 -1404 1698 -1398
rect 1692 -1410 1698 -1404
rect 1692 -1416 1698 -1410
rect 1692 -1422 1698 -1416
rect 1692 -1428 1698 -1422
rect 1692 -1434 1698 -1428
rect 1692 -1440 1698 -1434
rect 1692 -1446 1698 -1440
rect 1692 -1452 1698 -1446
rect 1692 -1458 1698 -1452
rect 1692 -1464 1698 -1458
rect 1692 -1470 1698 -1464
rect 1692 -1476 1698 -1470
rect 1692 -1482 1698 -1476
rect 1692 -1488 1698 -1482
rect 1692 -1494 1698 -1488
rect 1692 -1500 1698 -1494
rect 1692 -1506 1698 -1500
rect 1692 -1512 1698 -1506
rect 1692 -1518 1698 -1512
rect 1692 -1524 1698 -1518
rect 1692 -1530 1698 -1524
rect 1692 -1536 1698 -1530
rect 1692 -1542 1698 -1536
rect 1692 -1548 1698 -1542
rect 1692 -1554 1698 -1548
rect 1692 -1560 1698 -1554
rect 1692 -1566 1698 -1560
rect 1692 -1572 1698 -1566
rect 1692 -1578 1698 -1572
rect 1692 -1584 1698 -1578
rect 1692 -1590 1698 -1584
rect 1692 -1596 1698 -1590
rect 1692 -1602 1698 -1596
rect 1692 -1608 1698 -1602
rect 1692 -1614 1698 -1608
rect 1692 -1620 1698 -1614
rect 1692 -1626 1698 -1620
rect 1692 -1632 1698 -1626
rect 1692 -1638 1698 -1632
rect 1692 -1644 1698 -1638
rect 1692 -1650 1698 -1644
rect 1692 -1656 1698 -1650
rect 1692 -1662 1698 -1656
rect 1692 -1668 1698 -1662
rect 1692 -1674 1698 -1668
rect 1692 -1680 1698 -1674
rect 1692 -1686 1698 -1680
rect 1692 -1692 1698 -1686
rect 1692 -1698 1698 -1692
rect 1692 -1704 1698 -1698
rect 1692 -1710 1698 -1704
rect 1692 -1716 1698 -1710
rect 1692 -1722 1698 -1716
rect 1692 -1728 1698 -1722
rect 1692 -1734 1698 -1728
rect 1692 -1740 1698 -1734
rect 1692 -1746 1698 -1740
rect 1692 -1752 1698 -1746
rect 1692 -1758 1698 -1752
rect 1692 -1764 1698 -1758
rect 1692 -1770 1698 -1764
rect 1692 -1776 1698 -1770
rect 1692 -1782 1698 -1776
rect 1692 -1788 1698 -1782
rect 1692 -1794 1698 -1788
rect 1692 -1800 1698 -1794
rect 1692 -1806 1698 -1800
rect 1692 -1812 1698 -1806
rect 1692 -1818 1698 -1812
rect 1692 -1824 1698 -1818
rect 1692 -1830 1698 -1824
rect 1692 -1836 1698 -1830
rect 1692 -1842 1698 -1836
rect 1692 -1848 1698 -1842
rect 1692 -1854 1698 -1848
rect 1692 -1860 1698 -1854
rect 1692 -1866 1698 -1860
rect 1692 -1872 1698 -1866
rect 1692 -1878 1698 -1872
rect 1692 -1884 1698 -1878
rect 1692 -1890 1698 -1884
rect 1692 -1896 1698 -1890
rect 1692 -1902 1698 -1896
rect 1692 -1908 1698 -1902
rect 1692 -1914 1698 -1908
rect 1692 -1920 1698 -1914
rect 1692 -1926 1698 -1920
rect 1692 -1932 1698 -1926
rect 1692 -1938 1698 -1932
rect 1692 -1944 1698 -1938
rect 1692 -1950 1698 -1944
rect 1692 -1956 1698 -1950
rect 1692 -1962 1698 -1956
rect 1692 -2040 1698 -2034
rect 1692 -2046 1698 -2040
rect 1692 -2052 1698 -2046
rect 1692 -2058 1698 -2052
rect 1692 -2064 1698 -2058
rect 1692 -2070 1698 -2064
rect 1692 -2076 1698 -2070
rect 1692 -2082 1698 -2076
rect 1692 -2088 1698 -2082
rect 1692 -2094 1698 -2088
rect 1692 -2100 1698 -2094
rect 1692 -2106 1698 -2100
rect 1692 -2112 1698 -2106
rect 1692 -2118 1698 -2112
rect 1692 -2124 1698 -2118
rect 1692 -2130 1698 -2124
rect 1692 -2136 1698 -2130
rect 1692 -2142 1698 -2136
rect 1692 -2148 1698 -2142
rect 1692 -2154 1698 -2148
rect 1692 -2160 1698 -2154
rect 1692 -2166 1698 -2160
rect 1692 -2172 1698 -2166
rect 1692 -2178 1698 -2172
rect 1692 -2184 1698 -2178
rect 1692 -2190 1698 -2184
rect 1692 -2196 1698 -2190
rect 1692 -2202 1698 -2196
rect 1692 -2208 1698 -2202
rect 1692 -2214 1698 -2208
rect 1692 -2220 1698 -2214
rect 1692 -2226 1698 -2220
rect 1692 -2232 1698 -2226
rect 1692 -2238 1698 -2232
rect 1692 -2244 1698 -2238
rect 1692 -2250 1698 -2244
rect 1692 -2256 1698 -2250
rect 1692 -2262 1698 -2256
rect 1692 -2268 1698 -2262
rect 1692 -2274 1698 -2268
rect 1692 -2280 1698 -2274
rect 1692 -2286 1698 -2280
rect 1692 -2292 1698 -2286
rect 1692 -2298 1698 -2292
rect 1692 -2304 1698 -2298
rect 1692 -2310 1698 -2304
rect 1692 -2316 1698 -2310
rect 1692 -2322 1698 -2316
rect 1692 -2328 1698 -2322
rect 1692 -2334 1698 -2328
rect 1692 -2340 1698 -2334
rect 1692 -2346 1698 -2340
rect 1692 -2352 1698 -2346
rect 1692 -2358 1698 -2352
rect 1692 -2364 1698 -2358
rect 1692 -2370 1698 -2364
rect 1692 -2376 1698 -2370
rect 1692 -2382 1698 -2376
rect 1692 -2388 1698 -2382
rect 1692 -2394 1698 -2388
rect 1692 -2400 1698 -2394
rect 1692 -2406 1698 -2400
rect 1692 -2412 1698 -2406
rect 1692 -2418 1698 -2412
rect 1692 -2424 1698 -2418
rect 1692 -2430 1698 -2424
rect 1692 -2436 1698 -2430
rect 1692 -2442 1698 -2436
rect 1692 -2448 1698 -2442
rect 1692 -2454 1698 -2448
rect 1692 -2460 1698 -2454
rect 1692 -2466 1698 -2460
rect 1692 -2472 1698 -2466
rect 1692 -2478 1698 -2472
rect 1692 -2484 1698 -2478
rect 1692 -2490 1698 -2484
rect 1692 -2496 1698 -2490
rect 1692 -2502 1698 -2496
rect 1692 -2508 1698 -2502
rect 1692 -2514 1698 -2508
rect 1692 -2520 1698 -2514
rect 1692 -2526 1698 -2520
rect 1692 -2532 1698 -2526
rect 1692 -2538 1698 -2532
rect 1692 -2544 1698 -2538
rect 1692 -2550 1698 -2544
rect 1692 -2556 1698 -2550
rect 1692 -2562 1698 -2556
rect 1692 -2568 1698 -2562
rect 1692 -2574 1698 -2568
rect 1692 -2580 1698 -2574
rect 1692 -2586 1698 -2580
rect 1692 -2592 1698 -2586
rect 1692 -2598 1698 -2592
rect 1692 -2604 1698 -2598
rect 1692 -2610 1698 -2604
rect 1692 -2616 1698 -2610
rect 1692 -2622 1698 -2616
rect 1692 -2628 1698 -2622
rect 1692 -2634 1698 -2628
rect 1692 -2640 1698 -2634
rect 1692 -2646 1698 -2640
rect 1692 -2652 1698 -2646
rect 1692 -2658 1698 -2652
rect 1692 -2664 1698 -2658
rect 1692 -2670 1698 -2664
rect 1692 -2676 1698 -2670
rect 1692 -2682 1698 -2676
rect 1692 -2688 1698 -2682
rect 1692 -2694 1698 -2688
rect 1692 -2772 1698 -2766
rect 1692 -2778 1698 -2772
rect 1692 -2784 1698 -2778
rect 1692 -2790 1698 -2784
rect 1692 -2796 1698 -2790
rect 1692 -2802 1698 -2796
rect 1692 -2808 1698 -2802
rect 1692 -2814 1698 -2808
rect 1692 -2820 1698 -2814
rect 1692 -2826 1698 -2820
rect 1692 -2832 1698 -2826
rect 1692 -2838 1698 -2832
rect 1692 -2844 1698 -2838
rect 1692 -2850 1698 -2844
rect 1692 -2856 1698 -2850
rect 1692 -2862 1698 -2856
rect 1692 -2868 1698 -2862
rect 1692 -2874 1698 -2868
rect 1692 -2880 1698 -2874
rect 1692 -2886 1698 -2880
rect 1692 -2892 1698 -2886
rect 1692 -2898 1698 -2892
rect 1692 -2904 1698 -2898
rect 1692 -2910 1698 -2904
rect 1692 -2916 1698 -2910
rect 1692 -2922 1698 -2916
rect 1692 -2928 1698 -2922
rect 1692 -2934 1698 -2928
rect 1692 -2940 1698 -2934
rect 1692 -2946 1698 -2940
rect 1692 -2952 1698 -2946
rect 1692 -2958 1698 -2952
rect 1692 -2964 1698 -2958
rect 1692 -2970 1698 -2964
rect 1692 -2976 1698 -2970
rect 1692 -2982 1698 -2976
rect 1692 -2988 1698 -2982
rect 1692 -2994 1698 -2988
rect 1692 -3000 1698 -2994
rect 1692 -3006 1698 -3000
rect 1692 -3012 1698 -3006
rect 1692 -3018 1698 -3012
rect 1692 -3024 1698 -3018
rect 1692 -3030 1698 -3024
rect 1692 -3036 1698 -3030
rect 1692 -3042 1698 -3036
rect 1692 -3048 1698 -3042
rect 1692 -3054 1698 -3048
rect 1692 -3060 1698 -3054
rect 1692 -3066 1698 -3060
rect 1692 -3072 1698 -3066
rect 1692 -3078 1698 -3072
rect 1692 -3084 1698 -3078
rect 1692 -3090 1698 -3084
rect 1692 -3096 1698 -3090
rect 1692 -3102 1698 -3096
rect 1692 -3108 1698 -3102
rect 1692 -3114 1698 -3108
rect 1692 -3120 1698 -3114
rect 1692 -3126 1698 -3120
rect 1692 -3132 1698 -3126
rect 1692 -3138 1698 -3132
rect 1692 -3144 1698 -3138
rect 1692 -3150 1698 -3144
rect 1692 -3156 1698 -3150
rect 1692 -3162 1698 -3156
rect 1692 -3168 1698 -3162
rect 1692 -3174 1698 -3168
rect 1692 -3180 1698 -3174
rect 1692 -3186 1698 -3180
rect 1692 -3192 1698 -3186
rect 1692 -3198 1698 -3192
rect 1692 -3204 1698 -3198
rect 1692 -3210 1698 -3204
rect 1692 -3216 1698 -3210
rect 1692 -3222 1698 -3216
rect 1692 -3228 1698 -3222
rect 1692 -3276 1698 -3270
rect 1692 -3282 1698 -3276
rect 1692 -3288 1698 -3282
rect 1692 -3294 1698 -3288
rect 1692 -3300 1698 -3294
rect 1692 -3306 1698 -3300
rect 1692 -3312 1698 -3306
rect 1692 -3318 1698 -3312
rect 1692 -3324 1698 -3318
rect 1692 -3330 1698 -3324
rect 1692 -3336 1698 -3330
rect 1692 -3342 1698 -3336
rect 1692 -3348 1698 -3342
rect 1692 -3354 1698 -3348
rect 1692 -3360 1698 -3354
rect 1692 -3366 1698 -3360
rect 1692 -3372 1698 -3366
rect 1692 -3378 1698 -3372
rect 1692 -3384 1698 -3378
rect 1692 -3390 1698 -3384
rect 1692 -3396 1698 -3390
rect 1692 -3402 1698 -3396
rect 1692 -3408 1698 -3402
rect 1692 -3414 1698 -3408
rect 1692 -3420 1698 -3414
rect 1692 -3426 1698 -3420
rect 1698 -864 1704 -858
rect 1698 -870 1704 -864
rect 1698 -876 1704 -870
rect 1698 -882 1704 -876
rect 1698 -888 1704 -882
rect 1698 -894 1704 -888
rect 1698 -900 1704 -894
rect 1698 -906 1704 -900
rect 1698 -912 1704 -906
rect 1698 -918 1704 -912
rect 1698 -924 1704 -918
rect 1698 -930 1704 -924
rect 1698 -936 1704 -930
rect 1698 -942 1704 -936
rect 1698 -948 1704 -942
rect 1698 -954 1704 -948
rect 1698 -960 1704 -954
rect 1698 -966 1704 -960
rect 1698 -972 1704 -966
rect 1698 -978 1704 -972
rect 1698 -984 1704 -978
rect 1698 -990 1704 -984
rect 1698 -996 1704 -990
rect 1698 -1002 1704 -996
rect 1698 -1008 1704 -1002
rect 1698 -1014 1704 -1008
rect 1698 -1020 1704 -1014
rect 1698 -1026 1704 -1020
rect 1698 -1032 1704 -1026
rect 1698 -1038 1704 -1032
rect 1698 -1044 1704 -1038
rect 1698 -1050 1704 -1044
rect 1698 -1056 1704 -1050
rect 1698 -1062 1704 -1056
rect 1698 -1068 1704 -1062
rect 1698 -1074 1704 -1068
rect 1698 -1080 1704 -1074
rect 1698 -1086 1704 -1080
rect 1698 -1092 1704 -1086
rect 1698 -1098 1704 -1092
rect 1698 -1104 1704 -1098
rect 1698 -1110 1704 -1104
rect 1698 -1116 1704 -1110
rect 1698 -1122 1704 -1116
rect 1698 -1128 1704 -1122
rect 1698 -1134 1704 -1128
rect 1698 -1140 1704 -1134
rect 1698 -1146 1704 -1140
rect 1698 -1152 1704 -1146
rect 1698 -1158 1704 -1152
rect 1698 -1164 1704 -1158
rect 1698 -1170 1704 -1164
rect 1698 -1176 1704 -1170
rect 1698 -1182 1704 -1176
rect 1698 -1188 1704 -1182
rect 1698 -1194 1704 -1188
rect 1698 -1200 1704 -1194
rect 1698 -1206 1704 -1200
rect 1698 -1212 1704 -1206
rect 1698 -1218 1704 -1212
rect 1698 -1224 1704 -1218
rect 1698 -1230 1704 -1224
rect 1698 -1236 1704 -1230
rect 1698 -1242 1704 -1236
rect 1698 -1248 1704 -1242
rect 1698 -1254 1704 -1248
rect 1698 -1260 1704 -1254
rect 1698 -1266 1704 -1260
rect 1698 -1272 1704 -1266
rect 1698 -1278 1704 -1272
rect 1698 -1284 1704 -1278
rect 1698 -1290 1704 -1284
rect 1698 -1296 1704 -1290
rect 1698 -1302 1704 -1296
rect 1698 -1308 1704 -1302
rect 1698 -1314 1704 -1308
rect 1698 -1320 1704 -1314
rect 1698 -1326 1704 -1320
rect 1698 -1332 1704 -1326
rect 1698 -1338 1704 -1332
rect 1698 -1344 1704 -1338
rect 1698 -1350 1704 -1344
rect 1698 -1356 1704 -1350
rect 1698 -1362 1704 -1356
rect 1698 -1368 1704 -1362
rect 1698 -1374 1704 -1368
rect 1698 -1380 1704 -1374
rect 1698 -1386 1704 -1380
rect 1698 -1392 1704 -1386
rect 1698 -1398 1704 -1392
rect 1698 -1404 1704 -1398
rect 1698 -1410 1704 -1404
rect 1698 -1416 1704 -1410
rect 1698 -1422 1704 -1416
rect 1698 -1428 1704 -1422
rect 1698 -1434 1704 -1428
rect 1698 -1440 1704 -1434
rect 1698 -1446 1704 -1440
rect 1698 -1452 1704 -1446
rect 1698 -1458 1704 -1452
rect 1698 -1464 1704 -1458
rect 1698 -1470 1704 -1464
rect 1698 -1476 1704 -1470
rect 1698 -1482 1704 -1476
rect 1698 -1488 1704 -1482
rect 1698 -1494 1704 -1488
rect 1698 -1500 1704 -1494
rect 1698 -1506 1704 -1500
rect 1698 -1512 1704 -1506
rect 1698 -1518 1704 -1512
rect 1698 -1524 1704 -1518
rect 1698 -1530 1704 -1524
rect 1698 -1536 1704 -1530
rect 1698 -1542 1704 -1536
rect 1698 -1548 1704 -1542
rect 1698 -1554 1704 -1548
rect 1698 -1560 1704 -1554
rect 1698 -1566 1704 -1560
rect 1698 -1572 1704 -1566
rect 1698 -1578 1704 -1572
rect 1698 -1584 1704 -1578
rect 1698 -1590 1704 -1584
rect 1698 -1596 1704 -1590
rect 1698 -1602 1704 -1596
rect 1698 -1608 1704 -1602
rect 1698 -1614 1704 -1608
rect 1698 -1620 1704 -1614
rect 1698 -1626 1704 -1620
rect 1698 -1632 1704 -1626
rect 1698 -1638 1704 -1632
rect 1698 -1644 1704 -1638
rect 1698 -1650 1704 -1644
rect 1698 -1656 1704 -1650
rect 1698 -1662 1704 -1656
rect 1698 -1668 1704 -1662
rect 1698 -1674 1704 -1668
rect 1698 -1680 1704 -1674
rect 1698 -1686 1704 -1680
rect 1698 -1692 1704 -1686
rect 1698 -1698 1704 -1692
rect 1698 -1704 1704 -1698
rect 1698 -1710 1704 -1704
rect 1698 -1716 1704 -1710
rect 1698 -1722 1704 -1716
rect 1698 -1728 1704 -1722
rect 1698 -1734 1704 -1728
rect 1698 -1740 1704 -1734
rect 1698 -1746 1704 -1740
rect 1698 -1752 1704 -1746
rect 1698 -1758 1704 -1752
rect 1698 -1764 1704 -1758
rect 1698 -1770 1704 -1764
rect 1698 -1776 1704 -1770
rect 1698 -1782 1704 -1776
rect 1698 -1788 1704 -1782
rect 1698 -1794 1704 -1788
rect 1698 -1800 1704 -1794
rect 1698 -1806 1704 -1800
rect 1698 -1812 1704 -1806
rect 1698 -1818 1704 -1812
rect 1698 -1824 1704 -1818
rect 1698 -1830 1704 -1824
rect 1698 -1836 1704 -1830
rect 1698 -1842 1704 -1836
rect 1698 -1848 1704 -1842
rect 1698 -1854 1704 -1848
rect 1698 -1860 1704 -1854
rect 1698 -1866 1704 -1860
rect 1698 -1872 1704 -1866
rect 1698 -1878 1704 -1872
rect 1698 -1884 1704 -1878
rect 1698 -1890 1704 -1884
rect 1698 -1896 1704 -1890
rect 1698 -1902 1704 -1896
rect 1698 -1908 1704 -1902
rect 1698 -1914 1704 -1908
rect 1698 -1920 1704 -1914
rect 1698 -1926 1704 -1920
rect 1698 -1932 1704 -1926
rect 1698 -1938 1704 -1932
rect 1698 -1944 1704 -1938
rect 1698 -1950 1704 -1944
rect 1698 -1956 1704 -1950
rect 1698 -2034 1704 -2028
rect 1698 -2040 1704 -2034
rect 1698 -2046 1704 -2040
rect 1698 -2052 1704 -2046
rect 1698 -2058 1704 -2052
rect 1698 -2064 1704 -2058
rect 1698 -2070 1704 -2064
rect 1698 -2076 1704 -2070
rect 1698 -2082 1704 -2076
rect 1698 -2088 1704 -2082
rect 1698 -2094 1704 -2088
rect 1698 -2100 1704 -2094
rect 1698 -2106 1704 -2100
rect 1698 -2112 1704 -2106
rect 1698 -2118 1704 -2112
rect 1698 -2124 1704 -2118
rect 1698 -2130 1704 -2124
rect 1698 -2136 1704 -2130
rect 1698 -2142 1704 -2136
rect 1698 -2148 1704 -2142
rect 1698 -2154 1704 -2148
rect 1698 -2160 1704 -2154
rect 1698 -2166 1704 -2160
rect 1698 -2172 1704 -2166
rect 1698 -2178 1704 -2172
rect 1698 -2184 1704 -2178
rect 1698 -2190 1704 -2184
rect 1698 -2196 1704 -2190
rect 1698 -2202 1704 -2196
rect 1698 -2208 1704 -2202
rect 1698 -2214 1704 -2208
rect 1698 -2220 1704 -2214
rect 1698 -2226 1704 -2220
rect 1698 -2232 1704 -2226
rect 1698 -2238 1704 -2232
rect 1698 -2244 1704 -2238
rect 1698 -2250 1704 -2244
rect 1698 -2256 1704 -2250
rect 1698 -2262 1704 -2256
rect 1698 -2268 1704 -2262
rect 1698 -2274 1704 -2268
rect 1698 -2280 1704 -2274
rect 1698 -2286 1704 -2280
rect 1698 -2292 1704 -2286
rect 1698 -2298 1704 -2292
rect 1698 -2304 1704 -2298
rect 1698 -2310 1704 -2304
rect 1698 -2316 1704 -2310
rect 1698 -2322 1704 -2316
rect 1698 -2328 1704 -2322
rect 1698 -2334 1704 -2328
rect 1698 -2340 1704 -2334
rect 1698 -2346 1704 -2340
rect 1698 -2352 1704 -2346
rect 1698 -2358 1704 -2352
rect 1698 -2364 1704 -2358
rect 1698 -2370 1704 -2364
rect 1698 -2376 1704 -2370
rect 1698 -2382 1704 -2376
rect 1698 -2388 1704 -2382
rect 1698 -2394 1704 -2388
rect 1698 -2400 1704 -2394
rect 1698 -2406 1704 -2400
rect 1698 -2412 1704 -2406
rect 1698 -2418 1704 -2412
rect 1698 -2424 1704 -2418
rect 1698 -2430 1704 -2424
rect 1698 -2436 1704 -2430
rect 1698 -2442 1704 -2436
rect 1698 -2448 1704 -2442
rect 1698 -2454 1704 -2448
rect 1698 -2460 1704 -2454
rect 1698 -2466 1704 -2460
rect 1698 -2472 1704 -2466
rect 1698 -2478 1704 -2472
rect 1698 -2484 1704 -2478
rect 1698 -2490 1704 -2484
rect 1698 -2496 1704 -2490
rect 1698 -2502 1704 -2496
rect 1698 -2508 1704 -2502
rect 1698 -2514 1704 -2508
rect 1698 -2520 1704 -2514
rect 1698 -2526 1704 -2520
rect 1698 -2532 1704 -2526
rect 1698 -2538 1704 -2532
rect 1698 -2544 1704 -2538
rect 1698 -2550 1704 -2544
rect 1698 -2556 1704 -2550
rect 1698 -2562 1704 -2556
rect 1698 -2568 1704 -2562
rect 1698 -2574 1704 -2568
rect 1698 -2580 1704 -2574
rect 1698 -2586 1704 -2580
rect 1698 -2592 1704 -2586
rect 1698 -2598 1704 -2592
rect 1698 -2604 1704 -2598
rect 1698 -2610 1704 -2604
rect 1698 -2616 1704 -2610
rect 1698 -2622 1704 -2616
rect 1698 -2628 1704 -2622
rect 1698 -2634 1704 -2628
rect 1698 -2640 1704 -2634
rect 1698 -2646 1704 -2640
rect 1698 -2652 1704 -2646
rect 1698 -2658 1704 -2652
rect 1698 -2664 1704 -2658
rect 1698 -2670 1704 -2664
rect 1698 -2676 1704 -2670
rect 1698 -2682 1704 -2676
rect 1698 -2688 1704 -2682
rect 1698 -2766 1704 -2760
rect 1698 -2772 1704 -2766
rect 1698 -2778 1704 -2772
rect 1698 -2784 1704 -2778
rect 1698 -2790 1704 -2784
rect 1698 -2796 1704 -2790
rect 1698 -2802 1704 -2796
rect 1698 -2808 1704 -2802
rect 1698 -2814 1704 -2808
rect 1698 -2820 1704 -2814
rect 1698 -2826 1704 -2820
rect 1698 -2832 1704 -2826
rect 1698 -2838 1704 -2832
rect 1698 -2844 1704 -2838
rect 1698 -2850 1704 -2844
rect 1698 -2856 1704 -2850
rect 1698 -2862 1704 -2856
rect 1698 -2868 1704 -2862
rect 1698 -2874 1704 -2868
rect 1698 -2880 1704 -2874
rect 1698 -2886 1704 -2880
rect 1698 -2892 1704 -2886
rect 1698 -2898 1704 -2892
rect 1698 -2904 1704 -2898
rect 1698 -2910 1704 -2904
rect 1698 -2916 1704 -2910
rect 1698 -2922 1704 -2916
rect 1698 -2928 1704 -2922
rect 1698 -2934 1704 -2928
rect 1698 -2940 1704 -2934
rect 1698 -2946 1704 -2940
rect 1698 -2952 1704 -2946
rect 1698 -2958 1704 -2952
rect 1698 -2964 1704 -2958
rect 1698 -2970 1704 -2964
rect 1698 -2976 1704 -2970
rect 1698 -2982 1704 -2976
rect 1698 -2988 1704 -2982
rect 1698 -2994 1704 -2988
rect 1698 -3000 1704 -2994
rect 1698 -3006 1704 -3000
rect 1698 -3012 1704 -3006
rect 1698 -3018 1704 -3012
rect 1698 -3024 1704 -3018
rect 1698 -3030 1704 -3024
rect 1698 -3036 1704 -3030
rect 1698 -3042 1704 -3036
rect 1698 -3048 1704 -3042
rect 1698 -3054 1704 -3048
rect 1698 -3060 1704 -3054
rect 1698 -3066 1704 -3060
rect 1698 -3072 1704 -3066
rect 1698 -3078 1704 -3072
rect 1698 -3084 1704 -3078
rect 1698 -3090 1704 -3084
rect 1698 -3096 1704 -3090
rect 1698 -3102 1704 -3096
rect 1698 -3108 1704 -3102
rect 1698 -3114 1704 -3108
rect 1698 -3120 1704 -3114
rect 1698 -3126 1704 -3120
rect 1698 -3132 1704 -3126
rect 1698 -3138 1704 -3132
rect 1698 -3144 1704 -3138
rect 1698 -3150 1704 -3144
rect 1698 -3156 1704 -3150
rect 1698 -3162 1704 -3156
rect 1698 -3168 1704 -3162
rect 1698 -3174 1704 -3168
rect 1698 -3180 1704 -3174
rect 1698 -3186 1704 -3180
rect 1698 -3192 1704 -3186
rect 1698 -3198 1704 -3192
rect 1698 -3204 1704 -3198
rect 1698 -3210 1704 -3204
rect 1698 -3216 1704 -3210
rect 1698 -3222 1704 -3216
rect 1698 -3270 1704 -3264
rect 1698 -3276 1704 -3270
rect 1698 -3282 1704 -3276
rect 1698 -3288 1704 -3282
rect 1698 -3294 1704 -3288
rect 1698 -3300 1704 -3294
rect 1698 -3306 1704 -3300
rect 1698 -3312 1704 -3306
rect 1698 -3318 1704 -3312
rect 1698 -3324 1704 -3318
rect 1698 -3330 1704 -3324
rect 1698 -3336 1704 -3330
rect 1698 -3342 1704 -3336
rect 1698 -3348 1704 -3342
rect 1698 -3354 1704 -3348
rect 1698 -3360 1704 -3354
rect 1698 -3366 1704 -3360
rect 1698 -3372 1704 -3366
rect 1698 -3378 1704 -3372
rect 1698 -3384 1704 -3378
rect 1698 -3390 1704 -3384
rect 1698 -3396 1704 -3390
rect 1698 -3402 1704 -3396
rect 1698 -3408 1704 -3402
rect 1698 -3414 1704 -3408
rect 1698 -3420 1704 -3414
rect 1704 -858 1710 -852
rect 1704 -864 1710 -858
rect 1704 -870 1710 -864
rect 1704 -876 1710 -870
rect 1704 -882 1710 -876
rect 1704 -888 1710 -882
rect 1704 -894 1710 -888
rect 1704 -900 1710 -894
rect 1704 -906 1710 -900
rect 1704 -912 1710 -906
rect 1704 -918 1710 -912
rect 1704 -924 1710 -918
rect 1704 -930 1710 -924
rect 1704 -936 1710 -930
rect 1704 -942 1710 -936
rect 1704 -948 1710 -942
rect 1704 -954 1710 -948
rect 1704 -960 1710 -954
rect 1704 -966 1710 -960
rect 1704 -972 1710 -966
rect 1704 -978 1710 -972
rect 1704 -984 1710 -978
rect 1704 -990 1710 -984
rect 1704 -996 1710 -990
rect 1704 -1002 1710 -996
rect 1704 -1008 1710 -1002
rect 1704 -1014 1710 -1008
rect 1704 -1020 1710 -1014
rect 1704 -1026 1710 -1020
rect 1704 -1032 1710 -1026
rect 1704 -1038 1710 -1032
rect 1704 -1044 1710 -1038
rect 1704 -1050 1710 -1044
rect 1704 -1056 1710 -1050
rect 1704 -1062 1710 -1056
rect 1704 -1068 1710 -1062
rect 1704 -1074 1710 -1068
rect 1704 -1080 1710 -1074
rect 1704 -1086 1710 -1080
rect 1704 -1092 1710 -1086
rect 1704 -1098 1710 -1092
rect 1704 -1104 1710 -1098
rect 1704 -1110 1710 -1104
rect 1704 -1116 1710 -1110
rect 1704 -1122 1710 -1116
rect 1704 -1128 1710 -1122
rect 1704 -1134 1710 -1128
rect 1704 -1140 1710 -1134
rect 1704 -1146 1710 -1140
rect 1704 -1152 1710 -1146
rect 1704 -1158 1710 -1152
rect 1704 -1164 1710 -1158
rect 1704 -1170 1710 -1164
rect 1704 -1176 1710 -1170
rect 1704 -1182 1710 -1176
rect 1704 -1188 1710 -1182
rect 1704 -1194 1710 -1188
rect 1704 -1200 1710 -1194
rect 1704 -1206 1710 -1200
rect 1704 -1212 1710 -1206
rect 1704 -1218 1710 -1212
rect 1704 -1224 1710 -1218
rect 1704 -1230 1710 -1224
rect 1704 -1236 1710 -1230
rect 1704 -1242 1710 -1236
rect 1704 -1248 1710 -1242
rect 1704 -1254 1710 -1248
rect 1704 -1260 1710 -1254
rect 1704 -1266 1710 -1260
rect 1704 -1272 1710 -1266
rect 1704 -1278 1710 -1272
rect 1704 -1284 1710 -1278
rect 1704 -1290 1710 -1284
rect 1704 -1296 1710 -1290
rect 1704 -1302 1710 -1296
rect 1704 -1308 1710 -1302
rect 1704 -1314 1710 -1308
rect 1704 -1320 1710 -1314
rect 1704 -1326 1710 -1320
rect 1704 -1332 1710 -1326
rect 1704 -1338 1710 -1332
rect 1704 -1344 1710 -1338
rect 1704 -1350 1710 -1344
rect 1704 -1356 1710 -1350
rect 1704 -1362 1710 -1356
rect 1704 -1368 1710 -1362
rect 1704 -1374 1710 -1368
rect 1704 -1380 1710 -1374
rect 1704 -1386 1710 -1380
rect 1704 -1392 1710 -1386
rect 1704 -1398 1710 -1392
rect 1704 -1404 1710 -1398
rect 1704 -1410 1710 -1404
rect 1704 -1416 1710 -1410
rect 1704 -1422 1710 -1416
rect 1704 -1428 1710 -1422
rect 1704 -1434 1710 -1428
rect 1704 -1440 1710 -1434
rect 1704 -1446 1710 -1440
rect 1704 -1452 1710 -1446
rect 1704 -1458 1710 -1452
rect 1704 -1464 1710 -1458
rect 1704 -1470 1710 -1464
rect 1704 -1476 1710 -1470
rect 1704 -1482 1710 -1476
rect 1704 -1488 1710 -1482
rect 1704 -1494 1710 -1488
rect 1704 -1500 1710 -1494
rect 1704 -1506 1710 -1500
rect 1704 -1512 1710 -1506
rect 1704 -1518 1710 -1512
rect 1704 -1524 1710 -1518
rect 1704 -1530 1710 -1524
rect 1704 -1536 1710 -1530
rect 1704 -1542 1710 -1536
rect 1704 -1548 1710 -1542
rect 1704 -1554 1710 -1548
rect 1704 -1560 1710 -1554
rect 1704 -1566 1710 -1560
rect 1704 -1572 1710 -1566
rect 1704 -1578 1710 -1572
rect 1704 -1584 1710 -1578
rect 1704 -1590 1710 -1584
rect 1704 -1596 1710 -1590
rect 1704 -1602 1710 -1596
rect 1704 -1608 1710 -1602
rect 1704 -1614 1710 -1608
rect 1704 -1620 1710 -1614
rect 1704 -1626 1710 -1620
rect 1704 -1632 1710 -1626
rect 1704 -1638 1710 -1632
rect 1704 -1644 1710 -1638
rect 1704 -1650 1710 -1644
rect 1704 -1656 1710 -1650
rect 1704 -1662 1710 -1656
rect 1704 -1668 1710 -1662
rect 1704 -1674 1710 -1668
rect 1704 -1680 1710 -1674
rect 1704 -1686 1710 -1680
rect 1704 -1692 1710 -1686
rect 1704 -1698 1710 -1692
rect 1704 -1704 1710 -1698
rect 1704 -1710 1710 -1704
rect 1704 -1716 1710 -1710
rect 1704 -1722 1710 -1716
rect 1704 -1728 1710 -1722
rect 1704 -1734 1710 -1728
rect 1704 -1740 1710 -1734
rect 1704 -1746 1710 -1740
rect 1704 -1752 1710 -1746
rect 1704 -1758 1710 -1752
rect 1704 -1764 1710 -1758
rect 1704 -1770 1710 -1764
rect 1704 -1776 1710 -1770
rect 1704 -1782 1710 -1776
rect 1704 -1788 1710 -1782
rect 1704 -1794 1710 -1788
rect 1704 -1800 1710 -1794
rect 1704 -1806 1710 -1800
rect 1704 -1812 1710 -1806
rect 1704 -1818 1710 -1812
rect 1704 -1824 1710 -1818
rect 1704 -1830 1710 -1824
rect 1704 -1836 1710 -1830
rect 1704 -1842 1710 -1836
rect 1704 -1848 1710 -1842
rect 1704 -1854 1710 -1848
rect 1704 -1860 1710 -1854
rect 1704 -1866 1710 -1860
rect 1704 -1872 1710 -1866
rect 1704 -1878 1710 -1872
rect 1704 -1884 1710 -1878
rect 1704 -1890 1710 -1884
rect 1704 -1896 1710 -1890
rect 1704 -1902 1710 -1896
rect 1704 -1908 1710 -1902
rect 1704 -1914 1710 -1908
rect 1704 -1920 1710 -1914
rect 1704 -1926 1710 -1920
rect 1704 -1932 1710 -1926
rect 1704 -1938 1710 -1932
rect 1704 -1944 1710 -1938
rect 1704 -1950 1710 -1944
rect 1704 -2028 1710 -2022
rect 1704 -2034 1710 -2028
rect 1704 -2040 1710 -2034
rect 1704 -2046 1710 -2040
rect 1704 -2052 1710 -2046
rect 1704 -2058 1710 -2052
rect 1704 -2064 1710 -2058
rect 1704 -2070 1710 -2064
rect 1704 -2076 1710 -2070
rect 1704 -2082 1710 -2076
rect 1704 -2088 1710 -2082
rect 1704 -2094 1710 -2088
rect 1704 -2100 1710 -2094
rect 1704 -2106 1710 -2100
rect 1704 -2112 1710 -2106
rect 1704 -2118 1710 -2112
rect 1704 -2124 1710 -2118
rect 1704 -2130 1710 -2124
rect 1704 -2136 1710 -2130
rect 1704 -2142 1710 -2136
rect 1704 -2148 1710 -2142
rect 1704 -2154 1710 -2148
rect 1704 -2160 1710 -2154
rect 1704 -2166 1710 -2160
rect 1704 -2172 1710 -2166
rect 1704 -2178 1710 -2172
rect 1704 -2184 1710 -2178
rect 1704 -2190 1710 -2184
rect 1704 -2196 1710 -2190
rect 1704 -2202 1710 -2196
rect 1704 -2208 1710 -2202
rect 1704 -2214 1710 -2208
rect 1704 -2220 1710 -2214
rect 1704 -2226 1710 -2220
rect 1704 -2232 1710 -2226
rect 1704 -2238 1710 -2232
rect 1704 -2244 1710 -2238
rect 1704 -2250 1710 -2244
rect 1704 -2256 1710 -2250
rect 1704 -2262 1710 -2256
rect 1704 -2268 1710 -2262
rect 1704 -2274 1710 -2268
rect 1704 -2280 1710 -2274
rect 1704 -2286 1710 -2280
rect 1704 -2292 1710 -2286
rect 1704 -2298 1710 -2292
rect 1704 -2304 1710 -2298
rect 1704 -2310 1710 -2304
rect 1704 -2316 1710 -2310
rect 1704 -2322 1710 -2316
rect 1704 -2328 1710 -2322
rect 1704 -2334 1710 -2328
rect 1704 -2340 1710 -2334
rect 1704 -2346 1710 -2340
rect 1704 -2352 1710 -2346
rect 1704 -2358 1710 -2352
rect 1704 -2364 1710 -2358
rect 1704 -2370 1710 -2364
rect 1704 -2376 1710 -2370
rect 1704 -2382 1710 -2376
rect 1704 -2388 1710 -2382
rect 1704 -2394 1710 -2388
rect 1704 -2400 1710 -2394
rect 1704 -2406 1710 -2400
rect 1704 -2412 1710 -2406
rect 1704 -2418 1710 -2412
rect 1704 -2424 1710 -2418
rect 1704 -2430 1710 -2424
rect 1704 -2436 1710 -2430
rect 1704 -2442 1710 -2436
rect 1704 -2448 1710 -2442
rect 1704 -2454 1710 -2448
rect 1704 -2460 1710 -2454
rect 1704 -2466 1710 -2460
rect 1704 -2472 1710 -2466
rect 1704 -2478 1710 -2472
rect 1704 -2484 1710 -2478
rect 1704 -2490 1710 -2484
rect 1704 -2496 1710 -2490
rect 1704 -2502 1710 -2496
rect 1704 -2508 1710 -2502
rect 1704 -2514 1710 -2508
rect 1704 -2520 1710 -2514
rect 1704 -2526 1710 -2520
rect 1704 -2532 1710 -2526
rect 1704 -2538 1710 -2532
rect 1704 -2544 1710 -2538
rect 1704 -2550 1710 -2544
rect 1704 -2556 1710 -2550
rect 1704 -2562 1710 -2556
rect 1704 -2568 1710 -2562
rect 1704 -2574 1710 -2568
rect 1704 -2580 1710 -2574
rect 1704 -2586 1710 -2580
rect 1704 -2592 1710 -2586
rect 1704 -2598 1710 -2592
rect 1704 -2604 1710 -2598
rect 1704 -2610 1710 -2604
rect 1704 -2616 1710 -2610
rect 1704 -2622 1710 -2616
rect 1704 -2628 1710 -2622
rect 1704 -2634 1710 -2628
rect 1704 -2640 1710 -2634
rect 1704 -2646 1710 -2640
rect 1704 -2652 1710 -2646
rect 1704 -2658 1710 -2652
rect 1704 -2664 1710 -2658
rect 1704 -2670 1710 -2664
rect 1704 -2676 1710 -2670
rect 1704 -2682 1710 -2676
rect 1704 -2688 1710 -2682
rect 1704 -2760 1710 -2754
rect 1704 -2766 1710 -2760
rect 1704 -2772 1710 -2766
rect 1704 -2778 1710 -2772
rect 1704 -2784 1710 -2778
rect 1704 -2790 1710 -2784
rect 1704 -2796 1710 -2790
rect 1704 -2802 1710 -2796
rect 1704 -2808 1710 -2802
rect 1704 -2814 1710 -2808
rect 1704 -2820 1710 -2814
rect 1704 -2826 1710 -2820
rect 1704 -2832 1710 -2826
rect 1704 -2838 1710 -2832
rect 1704 -2844 1710 -2838
rect 1704 -2850 1710 -2844
rect 1704 -2856 1710 -2850
rect 1704 -2862 1710 -2856
rect 1704 -2868 1710 -2862
rect 1704 -2874 1710 -2868
rect 1704 -2880 1710 -2874
rect 1704 -2886 1710 -2880
rect 1704 -2892 1710 -2886
rect 1704 -2898 1710 -2892
rect 1704 -2904 1710 -2898
rect 1704 -2910 1710 -2904
rect 1704 -2916 1710 -2910
rect 1704 -2922 1710 -2916
rect 1704 -2928 1710 -2922
rect 1704 -2934 1710 -2928
rect 1704 -2940 1710 -2934
rect 1704 -2946 1710 -2940
rect 1704 -2952 1710 -2946
rect 1704 -2958 1710 -2952
rect 1704 -2964 1710 -2958
rect 1704 -2970 1710 -2964
rect 1704 -2976 1710 -2970
rect 1704 -2982 1710 -2976
rect 1704 -2988 1710 -2982
rect 1704 -2994 1710 -2988
rect 1704 -3000 1710 -2994
rect 1704 -3006 1710 -3000
rect 1704 -3012 1710 -3006
rect 1704 -3018 1710 -3012
rect 1704 -3024 1710 -3018
rect 1704 -3030 1710 -3024
rect 1704 -3036 1710 -3030
rect 1704 -3042 1710 -3036
rect 1704 -3048 1710 -3042
rect 1704 -3054 1710 -3048
rect 1704 -3060 1710 -3054
rect 1704 -3066 1710 -3060
rect 1704 -3072 1710 -3066
rect 1704 -3078 1710 -3072
rect 1704 -3084 1710 -3078
rect 1704 -3090 1710 -3084
rect 1704 -3096 1710 -3090
rect 1704 -3102 1710 -3096
rect 1704 -3108 1710 -3102
rect 1704 -3114 1710 -3108
rect 1704 -3120 1710 -3114
rect 1704 -3126 1710 -3120
rect 1704 -3132 1710 -3126
rect 1704 -3138 1710 -3132
rect 1704 -3144 1710 -3138
rect 1704 -3150 1710 -3144
rect 1704 -3156 1710 -3150
rect 1704 -3162 1710 -3156
rect 1704 -3168 1710 -3162
rect 1704 -3174 1710 -3168
rect 1704 -3180 1710 -3174
rect 1704 -3186 1710 -3180
rect 1704 -3192 1710 -3186
rect 1704 -3198 1710 -3192
rect 1704 -3204 1710 -3198
rect 1704 -3210 1710 -3204
rect 1704 -3216 1710 -3210
rect 1704 -3222 1710 -3216
rect 1704 -3270 1710 -3264
rect 1704 -3276 1710 -3270
rect 1704 -3282 1710 -3276
rect 1704 -3288 1710 -3282
rect 1704 -3294 1710 -3288
rect 1704 -3300 1710 -3294
rect 1704 -3306 1710 -3300
rect 1704 -3312 1710 -3306
rect 1704 -3318 1710 -3312
rect 1704 -3324 1710 -3318
rect 1704 -3330 1710 -3324
rect 1704 -3336 1710 -3330
rect 1704 -3342 1710 -3336
rect 1704 -3348 1710 -3342
rect 1704 -3354 1710 -3348
rect 1704 -3360 1710 -3354
rect 1704 -3366 1710 -3360
rect 1704 -3372 1710 -3366
rect 1704 -3378 1710 -3372
rect 1704 -3384 1710 -3378
rect 1704 -3390 1710 -3384
rect 1704 -3396 1710 -3390
rect 1704 -3402 1710 -3396
rect 1704 -3408 1710 -3402
rect 1704 -3414 1710 -3408
rect 1704 -3420 1710 -3414
rect 1710 -846 1716 -840
rect 1710 -852 1716 -846
rect 1710 -858 1716 -852
rect 1710 -864 1716 -858
rect 1710 -870 1716 -864
rect 1710 -876 1716 -870
rect 1710 -882 1716 -876
rect 1710 -888 1716 -882
rect 1710 -894 1716 -888
rect 1710 -900 1716 -894
rect 1710 -906 1716 -900
rect 1710 -912 1716 -906
rect 1710 -918 1716 -912
rect 1710 -924 1716 -918
rect 1710 -930 1716 -924
rect 1710 -936 1716 -930
rect 1710 -942 1716 -936
rect 1710 -948 1716 -942
rect 1710 -954 1716 -948
rect 1710 -960 1716 -954
rect 1710 -966 1716 -960
rect 1710 -972 1716 -966
rect 1710 -978 1716 -972
rect 1710 -984 1716 -978
rect 1710 -990 1716 -984
rect 1710 -996 1716 -990
rect 1710 -1002 1716 -996
rect 1710 -1008 1716 -1002
rect 1710 -1014 1716 -1008
rect 1710 -1020 1716 -1014
rect 1710 -1026 1716 -1020
rect 1710 -1032 1716 -1026
rect 1710 -1038 1716 -1032
rect 1710 -1044 1716 -1038
rect 1710 -1050 1716 -1044
rect 1710 -1056 1716 -1050
rect 1710 -1062 1716 -1056
rect 1710 -1068 1716 -1062
rect 1710 -1074 1716 -1068
rect 1710 -1080 1716 -1074
rect 1710 -1086 1716 -1080
rect 1710 -1092 1716 -1086
rect 1710 -1098 1716 -1092
rect 1710 -1104 1716 -1098
rect 1710 -1110 1716 -1104
rect 1710 -1116 1716 -1110
rect 1710 -1122 1716 -1116
rect 1710 -1128 1716 -1122
rect 1710 -1134 1716 -1128
rect 1710 -1140 1716 -1134
rect 1710 -1146 1716 -1140
rect 1710 -1152 1716 -1146
rect 1710 -1158 1716 -1152
rect 1710 -1164 1716 -1158
rect 1710 -1170 1716 -1164
rect 1710 -1176 1716 -1170
rect 1710 -1182 1716 -1176
rect 1710 -1188 1716 -1182
rect 1710 -1194 1716 -1188
rect 1710 -1200 1716 -1194
rect 1710 -1206 1716 -1200
rect 1710 -1212 1716 -1206
rect 1710 -1218 1716 -1212
rect 1710 -1224 1716 -1218
rect 1710 -1230 1716 -1224
rect 1710 -1236 1716 -1230
rect 1710 -1242 1716 -1236
rect 1710 -1248 1716 -1242
rect 1710 -1254 1716 -1248
rect 1710 -1260 1716 -1254
rect 1710 -1266 1716 -1260
rect 1710 -1272 1716 -1266
rect 1710 -1278 1716 -1272
rect 1710 -1284 1716 -1278
rect 1710 -1290 1716 -1284
rect 1710 -1296 1716 -1290
rect 1710 -1302 1716 -1296
rect 1710 -1308 1716 -1302
rect 1710 -1314 1716 -1308
rect 1710 -1320 1716 -1314
rect 1710 -1326 1716 -1320
rect 1710 -1332 1716 -1326
rect 1710 -1338 1716 -1332
rect 1710 -1344 1716 -1338
rect 1710 -1350 1716 -1344
rect 1710 -1356 1716 -1350
rect 1710 -1362 1716 -1356
rect 1710 -1368 1716 -1362
rect 1710 -1374 1716 -1368
rect 1710 -1380 1716 -1374
rect 1710 -1386 1716 -1380
rect 1710 -1392 1716 -1386
rect 1710 -1398 1716 -1392
rect 1710 -1404 1716 -1398
rect 1710 -1410 1716 -1404
rect 1710 -1416 1716 -1410
rect 1710 -1422 1716 -1416
rect 1710 -1428 1716 -1422
rect 1710 -1434 1716 -1428
rect 1710 -1440 1716 -1434
rect 1710 -1446 1716 -1440
rect 1710 -1452 1716 -1446
rect 1710 -1458 1716 -1452
rect 1710 -1464 1716 -1458
rect 1710 -1470 1716 -1464
rect 1710 -1476 1716 -1470
rect 1710 -1482 1716 -1476
rect 1710 -1488 1716 -1482
rect 1710 -1494 1716 -1488
rect 1710 -1500 1716 -1494
rect 1710 -1506 1716 -1500
rect 1710 -1512 1716 -1506
rect 1710 -1518 1716 -1512
rect 1710 -1524 1716 -1518
rect 1710 -1530 1716 -1524
rect 1710 -1536 1716 -1530
rect 1710 -1542 1716 -1536
rect 1710 -1548 1716 -1542
rect 1710 -1554 1716 -1548
rect 1710 -1560 1716 -1554
rect 1710 -1566 1716 -1560
rect 1710 -1572 1716 -1566
rect 1710 -1578 1716 -1572
rect 1710 -1584 1716 -1578
rect 1710 -1590 1716 -1584
rect 1710 -1596 1716 -1590
rect 1710 -1602 1716 -1596
rect 1710 -1608 1716 -1602
rect 1710 -1614 1716 -1608
rect 1710 -1620 1716 -1614
rect 1710 -1626 1716 -1620
rect 1710 -1632 1716 -1626
rect 1710 -1638 1716 -1632
rect 1710 -1644 1716 -1638
rect 1710 -1650 1716 -1644
rect 1710 -1656 1716 -1650
rect 1710 -1662 1716 -1656
rect 1710 -1668 1716 -1662
rect 1710 -1674 1716 -1668
rect 1710 -1680 1716 -1674
rect 1710 -1686 1716 -1680
rect 1710 -1692 1716 -1686
rect 1710 -1698 1716 -1692
rect 1710 -1704 1716 -1698
rect 1710 -1710 1716 -1704
rect 1710 -1716 1716 -1710
rect 1710 -1722 1716 -1716
rect 1710 -1728 1716 -1722
rect 1710 -1734 1716 -1728
rect 1710 -1740 1716 -1734
rect 1710 -1746 1716 -1740
rect 1710 -1752 1716 -1746
rect 1710 -1758 1716 -1752
rect 1710 -1764 1716 -1758
rect 1710 -1770 1716 -1764
rect 1710 -1776 1716 -1770
rect 1710 -1782 1716 -1776
rect 1710 -1788 1716 -1782
rect 1710 -1794 1716 -1788
rect 1710 -1800 1716 -1794
rect 1710 -1806 1716 -1800
rect 1710 -1812 1716 -1806
rect 1710 -1818 1716 -1812
rect 1710 -1824 1716 -1818
rect 1710 -1830 1716 -1824
rect 1710 -1836 1716 -1830
rect 1710 -1842 1716 -1836
rect 1710 -1848 1716 -1842
rect 1710 -1854 1716 -1848
rect 1710 -1860 1716 -1854
rect 1710 -1866 1716 -1860
rect 1710 -1872 1716 -1866
rect 1710 -1878 1716 -1872
rect 1710 -1884 1716 -1878
rect 1710 -1890 1716 -1884
rect 1710 -1896 1716 -1890
rect 1710 -1902 1716 -1896
rect 1710 -1908 1716 -1902
rect 1710 -1914 1716 -1908
rect 1710 -1920 1716 -1914
rect 1710 -1926 1716 -1920
rect 1710 -1932 1716 -1926
rect 1710 -1938 1716 -1932
rect 1710 -1944 1716 -1938
rect 1710 -2022 1716 -2016
rect 1710 -2028 1716 -2022
rect 1710 -2034 1716 -2028
rect 1710 -2040 1716 -2034
rect 1710 -2046 1716 -2040
rect 1710 -2052 1716 -2046
rect 1710 -2058 1716 -2052
rect 1710 -2064 1716 -2058
rect 1710 -2070 1716 -2064
rect 1710 -2076 1716 -2070
rect 1710 -2082 1716 -2076
rect 1710 -2088 1716 -2082
rect 1710 -2094 1716 -2088
rect 1710 -2100 1716 -2094
rect 1710 -2106 1716 -2100
rect 1710 -2112 1716 -2106
rect 1710 -2118 1716 -2112
rect 1710 -2124 1716 -2118
rect 1710 -2130 1716 -2124
rect 1710 -2136 1716 -2130
rect 1710 -2142 1716 -2136
rect 1710 -2148 1716 -2142
rect 1710 -2154 1716 -2148
rect 1710 -2160 1716 -2154
rect 1710 -2166 1716 -2160
rect 1710 -2172 1716 -2166
rect 1710 -2178 1716 -2172
rect 1710 -2184 1716 -2178
rect 1710 -2190 1716 -2184
rect 1710 -2196 1716 -2190
rect 1710 -2202 1716 -2196
rect 1710 -2208 1716 -2202
rect 1710 -2214 1716 -2208
rect 1710 -2220 1716 -2214
rect 1710 -2226 1716 -2220
rect 1710 -2232 1716 -2226
rect 1710 -2238 1716 -2232
rect 1710 -2244 1716 -2238
rect 1710 -2250 1716 -2244
rect 1710 -2256 1716 -2250
rect 1710 -2262 1716 -2256
rect 1710 -2268 1716 -2262
rect 1710 -2274 1716 -2268
rect 1710 -2280 1716 -2274
rect 1710 -2286 1716 -2280
rect 1710 -2292 1716 -2286
rect 1710 -2298 1716 -2292
rect 1710 -2304 1716 -2298
rect 1710 -2310 1716 -2304
rect 1710 -2316 1716 -2310
rect 1710 -2322 1716 -2316
rect 1710 -2328 1716 -2322
rect 1710 -2334 1716 -2328
rect 1710 -2340 1716 -2334
rect 1710 -2346 1716 -2340
rect 1710 -2352 1716 -2346
rect 1710 -2358 1716 -2352
rect 1710 -2364 1716 -2358
rect 1710 -2370 1716 -2364
rect 1710 -2376 1716 -2370
rect 1710 -2382 1716 -2376
rect 1710 -2388 1716 -2382
rect 1710 -2394 1716 -2388
rect 1710 -2400 1716 -2394
rect 1710 -2406 1716 -2400
rect 1710 -2412 1716 -2406
rect 1710 -2418 1716 -2412
rect 1710 -2424 1716 -2418
rect 1710 -2430 1716 -2424
rect 1710 -2436 1716 -2430
rect 1710 -2442 1716 -2436
rect 1710 -2448 1716 -2442
rect 1710 -2454 1716 -2448
rect 1710 -2460 1716 -2454
rect 1710 -2466 1716 -2460
rect 1710 -2472 1716 -2466
rect 1710 -2478 1716 -2472
rect 1710 -2484 1716 -2478
rect 1710 -2490 1716 -2484
rect 1710 -2496 1716 -2490
rect 1710 -2502 1716 -2496
rect 1710 -2508 1716 -2502
rect 1710 -2514 1716 -2508
rect 1710 -2520 1716 -2514
rect 1710 -2526 1716 -2520
rect 1710 -2532 1716 -2526
rect 1710 -2538 1716 -2532
rect 1710 -2544 1716 -2538
rect 1710 -2550 1716 -2544
rect 1710 -2556 1716 -2550
rect 1710 -2562 1716 -2556
rect 1710 -2568 1716 -2562
rect 1710 -2574 1716 -2568
rect 1710 -2580 1716 -2574
rect 1710 -2586 1716 -2580
rect 1710 -2592 1716 -2586
rect 1710 -2598 1716 -2592
rect 1710 -2604 1716 -2598
rect 1710 -2610 1716 -2604
rect 1710 -2616 1716 -2610
rect 1710 -2622 1716 -2616
rect 1710 -2628 1716 -2622
rect 1710 -2634 1716 -2628
rect 1710 -2640 1716 -2634
rect 1710 -2646 1716 -2640
rect 1710 -2652 1716 -2646
rect 1710 -2658 1716 -2652
rect 1710 -2664 1716 -2658
rect 1710 -2670 1716 -2664
rect 1710 -2676 1716 -2670
rect 1710 -2682 1716 -2676
rect 1710 -2760 1716 -2754
rect 1710 -2766 1716 -2760
rect 1710 -2772 1716 -2766
rect 1710 -2778 1716 -2772
rect 1710 -2784 1716 -2778
rect 1710 -2790 1716 -2784
rect 1710 -2796 1716 -2790
rect 1710 -2802 1716 -2796
rect 1710 -2808 1716 -2802
rect 1710 -2814 1716 -2808
rect 1710 -2820 1716 -2814
rect 1710 -2826 1716 -2820
rect 1710 -2832 1716 -2826
rect 1710 -2838 1716 -2832
rect 1710 -2844 1716 -2838
rect 1710 -2850 1716 -2844
rect 1710 -2856 1716 -2850
rect 1710 -2862 1716 -2856
rect 1710 -2868 1716 -2862
rect 1710 -2874 1716 -2868
rect 1710 -2880 1716 -2874
rect 1710 -2886 1716 -2880
rect 1710 -2892 1716 -2886
rect 1710 -2898 1716 -2892
rect 1710 -2904 1716 -2898
rect 1710 -2910 1716 -2904
rect 1710 -2916 1716 -2910
rect 1710 -2922 1716 -2916
rect 1710 -2928 1716 -2922
rect 1710 -2934 1716 -2928
rect 1710 -2940 1716 -2934
rect 1710 -2946 1716 -2940
rect 1710 -2952 1716 -2946
rect 1710 -2958 1716 -2952
rect 1710 -2964 1716 -2958
rect 1710 -2970 1716 -2964
rect 1710 -2976 1716 -2970
rect 1710 -2982 1716 -2976
rect 1710 -2988 1716 -2982
rect 1710 -2994 1716 -2988
rect 1710 -3000 1716 -2994
rect 1710 -3006 1716 -3000
rect 1710 -3012 1716 -3006
rect 1710 -3018 1716 -3012
rect 1710 -3024 1716 -3018
rect 1710 -3030 1716 -3024
rect 1710 -3036 1716 -3030
rect 1710 -3042 1716 -3036
rect 1710 -3048 1716 -3042
rect 1710 -3054 1716 -3048
rect 1710 -3060 1716 -3054
rect 1710 -3066 1716 -3060
rect 1710 -3072 1716 -3066
rect 1710 -3078 1716 -3072
rect 1710 -3084 1716 -3078
rect 1710 -3090 1716 -3084
rect 1710 -3096 1716 -3090
rect 1710 -3102 1716 -3096
rect 1710 -3108 1716 -3102
rect 1710 -3114 1716 -3108
rect 1710 -3120 1716 -3114
rect 1710 -3126 1716 -3120
rect 1710 -3132 1716 -3126
rect 1710 -3138 1716 -3132
rect 1710 -3144 1716 -3138
rect 1710 -3150 1716 -3144
rect 1710 -3156 1716 -3150
rect 1710 -3162 1716 -3156
rect 1710 -3168 1716 -3162
rect 1710 -3174 1716 -3168
rect 1710 -3180 1716 -3174
rect 1710 -3186 1716 -3180
rect 1710 -3192 1716 -3186
rect 1710 -3198 1716 -3192
rect 1710 -3204 1716 -3198
rect 1710 -3210 1716 -3204
rect 1710 -3216 1716 -3210
rect 1710 -3270 1716 -3264
rect 1710 -3276 1716 -3270
rect 1710 -3282 1716 -3276
rect 1710 -3288 1716 -3282
rect 1710 -3294 1716 -3288
rect 1710 -3300 1716 -3294
rect 1710 -3306 1716 -3300
rect 1710 -3312 1716 -3306
rect 1710 -3318 1716 -3312
rect 1710 -3324 1716 -3318
rect 1710 -3330 1716 -3324
rect 1710 -3336 1716 -3330
rect 1710 -3342 1716 -3336
rect 1710 -3348 1716 -3342
rect 1710 -3354 1716 -3348
rect 1710 -3360 1716 -3354
rect 1710 -3366 1716 -3360
rect 1710 -3372 1716 -3366
rect 1710 -3378 1716 -3372
rect 1710 -3384 1716 -3378
rect 1710 -3390 1716 -3384
rect 1710 -3396 1716 -3390
rect 1710 -3402 1716 -3396
rect 1710 -3408 1716 -3402
rect 1710 -3414 1716 -3408
rect 1716 -840 1722 -834
rect 1716 -846 1722 -840
rect 1716 -852 1722 -846
rect 1716 -858 1722 -852
rect 1716 -864 1722 -858
rect 1716 -870 1722 -864
rect 1716 -876 1722 -870
rect 1716 -882 1722 -876
rect 1716 -888 1722 -882
rect 1716 -894 1722 -888
rect 1716 -900 1722 -894
rect 1716 -906 1722 -900
rect 1716 -912 1722 -906
rect 1716 -918 1722 -912
rect 1716 -924 1722 -918
rect 1716 -930 1722 -924
rect 1716 -936 1722 -930
rect 1716 -942 1722 -936
rect 1716 -948 1722 -942
rect 1716 -954 1722 -948
rect 1716 -960 1722 -954
rect 1716 -966 1722 -960
rect 1716 -972 1722 -966
rect 1716 -978 1722 -972
rect 1716 -984 1722 -978
rect 1716 -990 1722 -984
rect 1716 -996 1722 -990
rect 1716 -1002 1722 -996
rect 1716 -1008 1722 -1002
rect 1716 -1014 1722 -1008
rect 1716 -1020 1722 -1014
rect 1716 -1026 1722 -1020
rect 1716 -1032 1722 -1026
rect 1716 -1038 1722 -1032
rect 1716 -1044 1722 -1038
rect 1716 -1050 1722 -1044
rect 1716 -1056 1722 -1050
rect 1716 -1062 1722 -1056
rect 1716 -1068 1722 -1062
rect 1716 -1074 1722 -1068
rect 1716 -1080 1722 -1074
rect 1716 -1086 1722 -1080
rect 1716 -1092 1722 -1086
rect 1716 -1098 1722 -1092
rect 1716 -1104 1722 -1098
rect 1716 -1110 1722 -1104
rect 1716 -1116 1722 -1110
rect 1716 -1122 1722 -1116
rect 1716 -1128 1722 -1122
rect 1716 -1134 1722 -1128
rect 1716 -1140 1722 -1134
rect 1716 -1146 1722 -1140
rect 1716 -1152 1722 -1146
rect 1716 -1158 1722 -1152
rect 1716 -1164 1722 -1158
rect 1716 -1170 1722 -1164
rect 1716 -1176 1722 -1170
rect 1716 -1182 1722 -1176
rect 1716 -1188 1722 -1182
rect 1716 -1194 1722 -1188
rect 1716 -1200 1722 -1194
rect 1716 -1206 1722 -1200
rect 1716 -1212 1722 -1206
rect 1716 -1218 1722 -1212
rect 1716 -1224 1722 -1218
rect 1716 -1230 1722 -1224
rect 1716 -1236 1722 -1230
rect 1716 -1242 1722 -1236
rect 1716 -1248 1722 -1242
rect 1716 -1254 1722 -1248
rect 1716 -1260 1722 -1254
rect 1716 -1266 1722 -1260
rect 1716 -1272 1722 -1266
rect 1716 -1278 1722 -1272
rect 1716 -1284 1722 -1278
rect 1716 -1290 1722 -1284
rect 1716 -1296 1722 -1290
rect 1716 -1302 1722 -1296
rect 1716 -1308 1722 -1302
rect 1716 -1314 1722 -1308
rect 1716 -1320 1722 -1314
rect 1716 -1326 1722 -1320
rect 1716 -1332 1722 -1326
rect 1716 -1338 1722 -1332
rect 1716 -1344 1722 -1338
rect 1716 -1350 1722 -1344
rect 1716 -1356 1722 -1350
rect 1716 -1362 1722 -1356
rect 1716 -1368 1722 -1362
rect 1716 -1374 1722 -1368
rect 1716 -1380 1722 -1374
rect 1716 -1386 1722 -1380
rect 1716 -1392 1722 -1386
rect 1716 -1398 1722 -1392
rect 1716 -1404 1722 -1398
rect 1716 -1410 1722 -1404
rect 1716 -1416 1722 -1410
rect 1716 -1422 1722 -1416
rect 1716 -1428 1722 -1422
rect 1716 -1434 1722 -1428
rect 1716 -1440 1722 -1434
rect 1716 -1446 1722 -1440
rect 1716 -1452 1722 -1446
rect 1716 -1458 1722 -1452
rect 1716 -1464 1722 -1458
rect 1716 -1470 1722 -1464
rect 1716 -1476 1722 -1470
rect 1716 -1482 1722 -1476
rect 1716 -1488 1722 -1482
rect 1716 -1494 1722 -1488
rect 1716 -1500 1722 -1494
rect 1716 -1506 1722 -1500
rect 1716 -1512 1722 -1506
rect 1716 -1518 1722 -1512
rect 1716 -1524 1722 -1518
rect 1716 -1530 1722 -1524
rect 1716 -1536 1722 -1530
rect 1716 -1542 1722 -1536
rect 1716 -1548 1722 -1542
rect 1716 -1554 1722 -1548
rect 1716 -1560 1722 -1554
rect 1716 -1566 1722 -1560
rect 1716 -1572 1722 -1566
rect 1716 -1578 1722 -1572
rect 1716 -1584 1722 -1578
rect 1716 -1590 1722 -1584
rect 1716 -1596 1722 -1590
rect 1716 -1602 1722 -1596
rect 1716 -1608 1722 -1602
rect 1716 -1614 1722 -1608
rect 1716 -1620 1722 -1614
rect 1716 -1626 1722 -1620
rect 1716 -1632 1722 -1626
rect 1716 -1638 1722 -1632
rect 1716 -1644 1722 -1638
rect 1716 -1650 1722 -1644
rect 1716 -1656 1722 -1650
rect 1716 -1662 1722 -1656
rect 1716 -1668 1722 -1662
rect 1716 -1674 1722 -1668
rect 1716 -1680 1722 -1674
rect 1716 -1686 1722 -1680
rect 1716 -1692 1722 -1686
rect 1716 -1698 1722 -1692
rect 1716 -1704 1722 -1698
rect 1716 -1710 1722 -1704
rect 1716 -1716 1722 -1710
rect 1716 -1722 1722 -1716
rect 1716 -1728 1722 -1722
rect 1716 -1734 1722 -1728
rect 1716 -1740 1722 -1734
rect 1716 -1746 1722 -1740
rect 1716 -1752 1722 -1746
rect 1716 -1758 1722 -1752
rect 1716 -1764 1722 -1758
rect 1716 -1770 1722 -1764
rect 1716 -1776 1722 -1770
rect 1716 -1782 1722 -1776
rect 1716 -1788 1722 -1782
rect 1716 -1794 1722 -1788
rect 1716 -1800 1722 -1794
rect 1716 -1806 1722 -1800
rect 1716 -1812 1722 -1806
rect 1716 -1818 1722 -1812
rect 1716 -1824 1722 -1818
rect 1716 -1830 1722 -1824
rect 1716 -1836 1722 -1830
rect 1716 -1842 1722 -1836
rect 1716 -1848 1722 -1842
rect 1716 -1854 1722 -1848
rect 1716 -1860 1722 -1854
rect 1716 -1866 1722 -1860
rect 1716 -1872 1722 -1866
rect 1716 -1878 1722 -1872
rect 1716 -1884 1722 -1878
rect 1716 -1890 1722 -1884
rect 1716 -1896 1722 -1890
rect 1716 -1902 1722 -1896
rect 1716 -1908 1722 -1902
rect 1716 -1914 1722 -1908
rect 1716 -1920 1722 -1914
rect 1716 -1926 1722 -1920
rect 1716 -1932 1722 -1926
rect 1716 -1938 1722 -1932
rect 1716 -2016 1722 -2010
rect 1716 -2022 1722 -2016
rect 1716 -2028 1722 -2022
rect 1716 -2034 1722 -2028
rect 1716 -2040 1722 -2034
rect 1716 -2046 1722 -2040
rect 1716 -2052 1722 -2046
rect 1716 -2058 1722 -2052
rect 1716 -2064 1722 -2058
rect 1716 -2070 1722 -2064
rect 1716 -2076 1722 -2070
rect 1716 -2082 1722 -2076
rect 1716 -2088 1722 -2082
rect 1716 -2094 1722 -2088
rect 1716 -2100 1722 -2094
rect 1716 -2106 1722 -2100
rect 1716 -2112 1722 -2106
rect 1716 -2118 1722 -2112
rect 1716 -2124 1722 -2118
rect 1716 -2130 1722 -2124
rect 1716 -2136 1722 -2130
rect 1716 -2142 1722 -2136
rect 1716 -2148 1722 -2142
rect 1716 -2154 1722 -2148
rect 1716 -2160 1722 -2154
rect 1716 -2166 1722 -2160
rect 1716 -2172 1722 -2166
rect 1716 -2178 1722 -2172
rect 1716 -2184 1722 -2178
rect 1716 -2190 1722 -2184
rect 1716 -2196 1722 -2190
rect 1716 -2202 1722 -2196
rect 1716 -2208 1722 -2202
rect 1716 -2214 1722 -2208
rect 1716 -2220 1722 -2214
rect 1716 -2226 1722 -2220
rect 1716 -2232 1722 -2226
rect 1716 -2238 1722 -2232
rect 1716 -2244 1722 -2238
rect 1716 -2250 1722 -2244
rect 1716 -2256 1722 -2250
rect 1716 -2262 1722 -2256
rect 1716 -2268 1722 -2262
rect 1716 -2274 1722 -2268
rect 1716 -2280 1722 -2274
rect 1716 -2286 1722 -2280
rect 1716 -2292 1722 -2286
rect 1716 -2298 1722 -2292
rect 1716 -2304 1722 -2298
rect 1716 -2310 1722 -2304
rect 1716 -2316 1722 -2310
rect 1716 -2322 1722 -2316
rect 1716 -2328 1722 -2322
rect 1716 -2334 1722 -2328
rect 1716 -2340 1722 -2334
rect 1716 -2346 1722 -2340
rect 1716 -2352 1722 -2346
rect 1716 -2358 1722 -2352
rect 1716 -2364 1722 -2358
rect 1716 -2370 1722 -2364
rect 1716 -2376 1722 -2370
rect 1716 -2382 1722 -2376
rect 1716 -2388 1722 -2382
rect 1716 -2394 1722 -2388
rect 1716 -2400 1722 -2394
rect 1716 -2406 1722 -2400
rect 1716 -2412 1722 -2406
rect 1716 -2418 1722 -2412
rect 1716 -2424 1722 -2418
rect 1716 -2430 1722 -2424
rect 1716 -2436 1722 -2430
rect 1716 -2442 1722 -2436
rect 1716 -2448 1722 -2442
rect 1716 -2454 1722 -2448
rect 1716 -2460 1722 -2454
rect 1716 -2466 1722 -2460
rect 1716 -2472 1722 -2466
rect 1716 -2478 1722 -2472
rect 1716 -2484 1722 -2478
rect 1716 -2490 1722 -2484
rect 1716 -2496 1722 -2490
rect 1716 -2502 1722 -2496
rect 1716 -2508 1722 -2502
rect 1716 -2514 1722 -2508
rect 1716 -2520 1722 -2514
rect 1716 -2526 1722 -2520
rect 1716 -2532 1722 -2526
rect 1716 -2538 1722 -2532
rect 1716 -2544 1722 -2538
rect 1716 -2550 1722 -2544
rect 1716 -2556 1722 -2550
rect 1716 -2562 1722 -2556
rect 1716 -2568 1722 -2562
rect 1716 -2574 1722 -2568
rect 1716 -2580 1722 -2574
rect 1716 -2586 1722 -2580
rect 1716 -2592 1722 -2586
rect 1716 -2598 1722 -2592
rect 1716 -2604 1722 -2598
rect 1716 -2610 1722 -2604
rect 1716 -2616 1722 -2610
rect 1716 -2622 1722 -2616
rect 1716 -2628 1722 -2622
rect 1716 -2634 1722 -2628
rect 1716 -2640 1722 -2634
rect 1716 -2646 1722 -2640
rect 1716 -2652 1722 -2646
rect 1716 -2658 1722 -2652
rect 1716 -2664 1722 -2658
rect 1716 -2670 1722 -2664
rect 1716 -2676 1722 -2670
rect 1716 -2754 1722 -2748
rect 1716 -2760 1722 -2754
rect 1716 -2766 1722 -2760
rect 1716 -2772 1722 -2766
rect 1716 -2778 1722 -2772
rect 1716 -2784 1722 -2778
rect 1716 -2790 1722 -2784
rect 1716 -2796 1722 -2790
rect 1716 -2802 1722 -2796
rect 1716 -2808 1722 -2802
rect 1716 -2814 1722 -2808
rect 1716 -2820 1722 -2814
rect 1716 -2826 1722 -2820
rect 1716 -2832 1722 -2826
rect 1716 -2838 1722 -2832
rect 1716 -2844 1722 -2838
rect 1716 -2850 1722 -2844
rect 1716 -2856 1722 -2850
rect 1716 -2862 1722 -2856
rect 1716 -2868 1722 -2862
rect 1716 -2874 1722 -2868
rect 1716 -2880 1722 -2874
rect 1716 -2886 1722 -2880
rect 1716 -2892 1722 -2886
rect 1716 -2898 1722 -2892
rect 1716 -2904 1722 -2898
rect 1716 -2910 1722 -2904
rect 1716 -2916 1722 -2910
rect 1716 -2922 1722 -2916
rect 1716 -2928 1722 -2922
rect 1716 -2934 1722 -2928
rect 1716 -2940 1722 -2934
rect 1716 -2946 1722 -2940
rect 1716 -2952 1722 -2946
rect 1716 -2958 1722 -2952
rect 1716 -2964 1722 -2958
rect 1716 -2970 1722 -2964
rect 1716 -2976 1722 -2970
rect 1716 -2982 1722 -2976
rect 1716 -2988 1722 -2982
rect 1716 -2994 1722 -2988
rect 1716 -3000 1722 -2994
rect 1716 -3006 1722 -3000
rect 1716 -3012 1722 -3006
rect 1716 -3018 1722 -3012
rect 1716 -3024 1722 -3018
rect 1716 -3030 1722 -3024
rect 1716 -3036 1722 -3030
rect 1716 -3042 1722 -3036
rect 1716 -3048 1722 -3042
rect 1716 -3054 1722 -3048
rect 1716 -3060 1722 -3054
rect 1716 -3066 1722 -3060
rect 1716 -3072 1722 -3066
rect 1716 -3078 1722 -3072
rect 1716 -3084 1722 -3078
rect 1716 -3090 1722 -3084
rect 1716 -3096 1722 -3090
rect 1716 -3102 1722 -3096
rect 1716 -3108 1722 -3102
rect 1716 -3114 1722 -3108
rect 1716 -3120 1722 -3114
rect 1716 -3126 1722 -3120
rect 1716 -3132 1722 -3126
rect 1716 -3138 1722 -3132
rect 1716 -3144 1722 -3138
rect 1716 -3150 1722 -3144
rect 1716 -3156 1722 -3150
rect 1716 -3162 1722 -3156
rect 1716 -3168 1722 -3162
rect 1716 -3174 1722 -3168
rect 1716 -3180 1722 -3174
rect 1716 -3186 1722 -3180
rect 1716 -3192 1722 -3186
rect 1716 -3198 1722 -3192
rect 1716 -3204 1722 -3198
rect 1716 -3210 1722 -3204
rect 1716 -3216 1722 -3210
rect 1716 -3264 1722 -3258
rect 1716 -3270 1722 -3264
rect 1716 -3276 1722 -3270
rect 1716 -3282 1722 -3276
rect 1716 -3288 1722 -3282
rect 1716 -3294 1722 -3288
rect 1716 -3300 1722 -3294
rect 1716 -3306 1722 -3300
rect 1716 -3312 1722 -3306
rect 1716 -3318 1722 -3312
rect 1716 -3324 1722 -3318
rect 1716 -3330 1722 -3324
rect 1716 -3336 1722 -3330
rect 1716 -3342 1722 -3336
rect 1716 -3348 1722 -3342
rect 1716 -3354 1722 -3348
rect 1716 -3360 1722 -3354
rect 1716 -3366 1722 -3360
rect 1716 -3372 1722 -3366
rect 1716 -3378 1722 -3372
rect 1716 -3384 1722 -3378
rect 1716 -3390 1722 -3384
rect 1716 -3396 1722 -3390
rect 1716 -3402 1722 -3396
rect 1716 -3408 1722 -3402
rect 1716 -3414 1722 -3408
rect 1722 -834 1728 -828
rect 1722 -840 1728 -834
rect 1722 -846 1728 -840
rect 1722 -852 1728 -846
rect 1722 -858 1728 -852
rect 1722 -864 1728 -858
rect 1722 -870 1728 -864
rect 1722 -876 1728 -870
rect 1722 -882 1728 -876
rect 1722 -888 1728 -882
rect 1722 -894 1728 -888
rect 1722 -900 1728 -894
rect 1722 -906 1728 -900
rect 1722 -912 1728 -906
rect 1722 -918 1728 -912
rect 1722 -924 1728 -918
rect 1722 -930 1728 -924
rect 1722 -936 1728 -930
rect 1722 -942 1728 -936
rect 1722 -948 1728 -942
rect 1722 -954 1728 -948
rect 1722 -960 1728 -954
rect 1722 -966 1728 -960
rect 1722 -972 1728 -966
rect 1722 -978 1728 -972
rect 1722 -984 1728 -978
rect 1722 -990 1728 -984
rect 1722 -996 1728 -990
rect 1722 -1002 1728 -996
rect 1722 -1008 1728 -1002
rect 1722 -1014 1728 -1008
rect 1722 -1020 1728 -1014
rect 1722 -1026 1728 -1020
rect 1722 -1032 1728 -1026
rect 1722 -1038 1728 -1032
rect 1722 -1044 1728 -1038
rect 1722 -1050 1728 -1044
rect 1722 -1056 1728 -1050
rect 1722 -1062 1728 -1056
rect 1722 -1068 1728 -1062
rect 1722 -1074 1728 -1068
rect 1722 -1080 1728 -1074
rect 1722 -1086 1728 -1080
rect 1722 -1092 1728 -1086
rect 1722 -1098 1728 -1092
rect 1722 -1104 1728 -1098
rect 1722 -1110 1728 -1104
rect 1722 -1116 1728 -1110
rect 1722 -1122 1728 -1116
rect 1722 -1128 1728 -1122
rect 1722 -1134 1728 -1128
rect 1722 -1140 1728 -1134
rect 1722 -1146 1728 -1140
rect 1722 -1152 1728 -1146
rect 1722 -1158 1728 -1152
rect 1722 -1164 1728 -1158
rect 1722 -1170 1728 -1164
rect 1722 -1176 1728 -1170
rect 1722 -1182 1728 -1176
rect 1722 -1188 1728 -1182
rect 1722 -1194 1728 -1188
rect 1722 -1200 1728 -1194
rect 1722 -1206 1728 -1200
rect 1722 -1212 1728 -1206
rect 1722 -1218 1728 -1212
rect 1722 -1224 1728 -1218
rect 1722 -1230 1728 -1224
rect 1722 -1236 1728 -1230
rect 1722 -1242 1728 -1236
rect 1722 -1248 1728 -1242
rect 1722 -1254 1728 -1248
rect 1722 -1260 1728 -1254
rect 1722 -1266 1728 -1260
rect 1722 -1272 1728 -1266
rect 1722 -1278 1728 -1272
rect 1722 -1284 1728 -1278
rect 1722 -1290 1728 -1284
rect 1722 -1296 1728 -1290
rect 1722 -1302 1728 -1296
rect 1722 -1308 1728 -1302
rect 1722 -1314 1728 -1308
rect 1722 -1320 1728 -1314
rect 1722 -1326 1728 -1320
rect 1722 -1332 1728 -1326
rect 1722 -1338 1728 -1332
rect 1722 -1344 1728 -1338
rect 1722 -1350 1728 -1344
rect 1722 -1356 1728 -1350
rect 1722 -1362 1728 -1356
rect 1722 -1368 1728 -1362
rect 1722 -1374 1728 -1368
rect 1722 -1380 1728 -1374
rect 1722 -1386 1728 -1380
rect 1722 -1392 1728 -1386
rect 1722 -1398 1728 -1392
rect 1722 -1404 1728 -1398
rect 1722 -1410 1728 -1404
rect 1722 -1416 1728 -1410
rect 1722 -1422 1728 -1416
rect 1722 -1428 1728 -1422
rect 1722 -1434 1728 -1428
rect 1722 -1440 1728 -1434
rect 1722 -1446 1728 -1440
rect 1722 -1452 1728 -1446
rect 1722 -1458 1728 -1452
rect 1722 -1464 1728 -1458
rect 1722 -1470 1728 -1464
rect 1722 -1476 1728 -1470
rect 1722 -1482 1728 -1476
rect 1722 -1488 1728 -1482
rect 1722 -1494 1728 -1488
rect 1722 -1500 1728 -1494
rect 1722 -1506 1728 -1500
rect 1722 -1512 1728 -1506
rect 1722 -1518 1728 -1512
rect 1722 -1524 1728 -1518
rect 1722 -1530 1728 -1524
rect 1722 -1536 1728 -1530
rect 1722 -1542 1728 -1536
rect 1722 -1548 1728 -1542
rect 1722 -1554 1728 -1548
rect 1722 -1560 1728 -1554
rect 1722 -1566 1728 -1560
rect 1722 -1572 1728 -1566
rect 1722 -1578 1728 -1572
rect 1722 -1584 1728 -1578
rect 1722 -1590 1728 -1584
rect 1722 -1596 1728 -1590
rect 1722 -1602 1728 -1596
rect 1722 -1608 1728 -1602
rect 1722 -1614 1728 -1608
rect 1722 -1620 1728 -1614
rect 1722 -1626 1728 -1620
rect 1722 -1632 1728 -1626
rect 1722 -1638 1728 -1632
rect 1722 -1644 1728 -1638
rect 1722 -1650 1728 -1644
rect 1722 -1656 1728 -1650
rect 1722 -1662 1728 -1656
rect 1722 -1668 1728 -1662
rect 1722 -1674 1728 -1668
rect 1722 -1680 1728 -1674
rect 1722 -1686 1728 -1680
rect 1722 -1692 1728 -1686
rect 1722 -1698 1728 -1692
rect 1722 -1704 1728 -1698
rect 1722 -1710 1728 -1704
rect 1722 -1716 1728 -1710
rect 1722 -1722 1728 -1716
rect 1722 -1728 1728 -1722
rect 1722 -1734 1728 -1728
rect 1722 -1740 1728 -1734
rect 1722 -1746 1728 -1740
rect 1722 -1752 1728 -1746
rect 1722 -1758 1728 -1752
rect 1722 -1764 1728 -1758
rect 1722 -1770 1728 -1764
rect 1722 -1776 1728 -1770
rect 1722 -1782 1728 -1776
rect 1722 -1788 1728 -1782
rect 1722 -1794 1728 -1788
rect 1722 -1800 1728 -1794
rect 1722 -1806 1728 -1800
rect 1722 -1812 1728 -1806
rect 1722 -1818 1728 -1812
rect 1722 -1824 1728 -1818
rect 1722 -1830 1728 -1824
rect 1722 -1836 1728 -1830
rect 1722 -1842 1728 -1836
rect 1722 -1848 1728 -1842
rect 1722 -1854 1728 -1848
rect 1722 -1860 1728 -1854
rect 1722 -1866 1728 -1860
rect 1722 -1872 1728 -1866
rect 1722 -1878 1728 -1872
rect 1722 -1884 1728 -1878
rect 1722 -1890 1728 -1884
rect 1722 -1896 1728 -1890
rect 1722 -1902 1728 -1896
rect 1722 -1908 1728 -1902
rect 1722 -1914 1728 -1908
rect 1722 -1920 1728 -1914
rect 1722 -1926 1728 -1920
rect 1722 -1932 1728 -1926
rect 1722 -2010 1728 -2004
rect 1722 -2016 1728 -2010
rect 1722 -2022 1728 -2016
rect 1722 -2028 1728 -2022
rect 1722 -2034 1728 -2028
rect 1722 -2040 1728 -2034
rect 1722 -2046 1728 -2040
rect 1722 -2052 1728 -2046
rect 1722 -2058 1728 -2052
rect 1722 -2064 1728 -2058
rect 1722 -2070 1728 -2064
rect 1722 -2076 1728 -2070
rect 1722 -2082 1728 -2076
rect 1722 -2088 1728 -2082
rect 1722 -2094 1728 -2088
rect 1722 -2100 1728 -2094
rect 1722 -2106 1728 -2100
rect 1722 -2112 1728 -2106
rect 1722 -2118 1728 -2112
rect 1722 -2124 1728 -2118
rect 1722 -2130 1728 -2124
rect 1722 -2136 1728 -2130
rect 1722 -2142 1728 -2136
rect 1722 -2148 1728 -2142
rect 1722 -2154 1728 -2148
rect 1722 -2160 1728 -2154
rect 1722 -2166 1728 -2160
rect 1722 -2172 1728 -2166
rect 1722 -2178 1728 -2172
rect 1722 -2184 1728 -2178
rect 1722 -2190 1728 -2184
rect 1722 -2196 1728 -2190
rect 1722 -2202 1728 -2196
rect 1722 -2208 1728 -2202
rect 1722 -2214 1728 -2208
rect 1722 -2220 1728 -2214
rect 1722 -2226 1728 -2220
rect 1722 -2232 1728 -2226
rect 1722 -2238 1728 -2232
rect 1722 -2244 1728 -2238
rect 1722 -2250 1728 -2244
rect 1722 -2256 1728 -2250
rect 1722 -2262 1728 -2256
rect 1722 -2268 1728 -2262
rect 1722 -2274 1728 -2268
rect 1722 -2280 1728 -2274
rect 1722 -2286 1728 -2280
rect 1722 -2292 1728 -2286
rect 1722 -2298 1728 -2292
rect 1722 -2304 1728 -2298
rect 1722 -2310 1728 -2304
rect 1722 -2316 1728 -2310
rect 1722 -2322 1728 -2316
rect 1722 -2328 1728 -2322
rect 1722 -2334 1728 -2328
rect 1722 -2340 1728 -2334
rect 1722 -2346 1728 -2340
rect 1722 -2352 1728 -2346
rect 1722 -2358 1728 -2352
rect 1722 -2364 1728 -2358
rect 1722 -2370 1728 -2364
rect 1722 -2376 1728 -2370
rect 1722 -2382 1728 -2376
rect 1722 -2388 1728 -2382
rect 1722 -2394 1728 -2388
rect 1722 -2400 1728 -2394
rect 1722 -2406 1728 -2400
rect 1722 -2412 1728 -2406
rect 1722 -2418 1728 -2412
rect 1722 -2424 1728 -2418
rect 1722 -2430 1728 -2424
rect 1722 -2436 1728 -2430
rect 1722 -2442 1728 -2436
rect 1722 -2448 1728 -2442
rect 1722 -2454 1728 -2448
rect 1722 -2460 1728 -2454
rect 1722 -2466 1728 -2460
rect 1722 -2472 1728 -2466
rect 1722 -2478 1728 -2472
rect 1722 -2484 1728 -2478
rect 1722 -2490 1728 -2484
rect 1722 -2496 1728 -2490
rect 1722 -2502 1728 -2496
rect 1722 -2508 1728 -2502
rect 1722 -2514 1728 -2508
rect 1722 -2520 1728 -2514
rect 1722 -2526 1728 -2520
rect 1722 -2532 1728 -2526
rect 1722 -2538 1728 -2532
rect 1722 -2544 1728 -2538
rect 1722 -2550 1728 -2544
rect 1722 -2556 1728 -2550
rect 1722 -2562 1728 -2556
rect 1722 -2568 1728 -2562
rect 1722 -2574 1728 -2568
rect 1722 -2580 1728 -2574
rect 1722 -2586 1728 -2580
rect 1722 -2592 1728 -2586
rect 1722 -2598 1728 -2592
rect 1722 -2604 1728 -2598
rect 1722 -2610 1728 -2604
rect 1722 -2616 1728 -2610
rect 1722 -2622 1728 -2616
rect 1722 -2628 1728 -2622
rect 1722 -2634 1728 -2628
rect 1722 -2640 1728 -2634
rect 1722 -2646 1728 -2640
rect 1722 -2652 1728 -2646
rect 1722 -2658 1728 -2652
rect 1722 -2664 1728 -2658
rect 1722 -2670 1728 -2664
rect 1722 -2676 1728 -2670
rect 1722 -2748 1728 -2742
rect 1722 -2754 1728 -2748
rect 1722 -2760 1728 -2754
rect 1722 -2766 1728 -2760
rect 1722 -2772 1728 -2766
rect 1722 -2778 1728 -2772
rect 1722 -2784 1728 -2778
rect 1722 -2790 1728 -2784
rect 1722 -2796 1728 -2790
rect 1722 -2802 1728 -2796
rect 1722 -2808 1728 -2802
rect 1722 -2814 1728 -2808
rect 1722 -2820 1728 -2814
rect 1722 -2826 1728 -2820
rect 1722 -2832 1728 -2826
rect 1722 -2838 1728 -2832
rect 1722 -2844 1728 -2838
rect 1722 -2850 1728 -2844
rect 1722 -2856 1728 -2850
rect 1722 -2862 1728 -2856
rect 1722 -2868 1728 -2862
rect 1722 -2874 1728 -2868
rect 1722 -2880 1728 -2874
rect 1722 -2886 1728 -2880
rect 1722 -2892 1728 -2886
rect 1722 -2898 1728 -2892
rect 1722 -2904 1728 -2898
rect 1722 -2910 1728 -2904
rect 1722 -2916 1728 -2910
rect 1722 -2922 1728 -2916
rect 1722 -2928 1728 -2922
rect 1722 -2934 1728 -2928
rect 1722 -2940 1728 -2934
rect 1722 -2946 1728 -2940
rect 1722 -2952 1728 -2946
rect 1722 -2958 1728 -2952
rect 1722 -2964 1728 -2958
rect 1722 -2970 1728 -2964
rect 1722 -2976 1728 -2970
rect 1722 -2982 1728 -2976
rect 1722 -2988 1728 -2982
rect 1722 -2994 1728 -2988
rect 1722 -3000 1728 -2994
rect 1722 -3006 1728 -3000
rect 1722 -3012 1728 -3006
rect 1722 -3018 1728 -3012
rect 1722 -3024 1728 -3018
rect 1722 -3030 1728 -3024
rect 1722 -3036 1728 -3030
rect 1722 -3042 1728 -3036
rect 1722 -3048 1728 -3042
rect 1722 -3054 1728 -3048
rect 1722 -3060 1728 -3054
rect 1722 -3066 1728 -3060
rect 1722 -3072 1728 -3066
rect 1722 -3078 1728 -3072
rect 1722 -3084 1728 -3078
rect 1722 -3090 1728 -3084
rect 1722 -3096 1728 -3090
rect 1722 -3102 1728 -3096
rect 1722 -3108 1728 -3102
rect 1722 -3114 1728 -3108
rect 1722 -3120 1728 -3114
rect 1722 -3126 1728 -3120
rect 1722 -3132 1728 -3126
rect 1722 -3138 1728 -3132
rect 1722 -3144 1728 -3138
rect 1722 -3150 1728 -3144
rect 1722 -3156 1728 -3150
rect 1722 -3162 1728 -3156
rect 1722 -3168 1728 -3162
rect 1722 -3174 1728 -3168
rect 1722 -3180 1728 -3174
rect 1722 -3186 1728 -3180
rect 1722 -3192 1728 -3186
rect 1722 -3198 1728 -3192
rect 1722 -3204 1728 -3198
rect 1722 -3210 1728 -3204
rect 1722 -3216 1728 -3210
rect 1722 -3264 1728 -3258
rect 1722 -3270 1728 -3264
rect 1722 -3276 1728 -3270
rect 1722 -3282 1728 -3276
rect 1722 -3288 1728 -3282
rect 1722 -3294 1728 -3288
rect 1722 -3300 1728 -3294
rect 1722 -3306 1728 -3300
rect 1722 -3312 1728 -3306
rect 1722 -3318 1728 -3312
rect 1722 -3324 1728 -3318
rect 1722 -3330 1728 -3324
rect 1722 -3336 1728 -3330
rect 1722 -3342 1728 -3336
rect 1722 -3348 1728 -3342
rect 1722 -3354 1728 -3348
rect 1722 -3360 1728 -3354
rect 1722 -3366 1728 -3360
rect 1722 -3372 1728 -3366
rect 1722 -3378 1728 -3372
rect 1722 -3384 1728 -3378
rect 1722 -3390 1728 -3384
rect 1722 -3396 1728 -3390
rect 1722 -3402 1728 -3396
rect 1722 -3408 1728 -3402
rect 1728 -822 1734 -816
rect 1728 -828 1734 -822
rect 1728 -834 1734 -828
rect 1728 -840 1734 -834
rect 1728 -846 1734 -840
rect 1728 -852 1734 -846
rect 1728 -858 1734 -852
rect 1728 -864 1734 -858
rect 1728 -870 1734 -864
rect 1728 -876 1734 -870
rect 1728 -882 1734 -876
rect 1728 -888 1734 -882
rect 1728 -894 1734 -888
rect 1728 -900 1734 -894
rect 1728 -906 1734 -900
rect 1728 -912 1734 -906
rect 1728 -918 1734 -912
rect 1728 -924 1734 -918
rect 1728 -930 1734 -924
rect 1728 -936 1734 -930
rect 1728 -942 1734 -936
rect 1728 -948 1734 -942
rect 1728 -954 1734 -948
rect 1728 -960 1734 -954
rect 1728 -966 1734 -960
rect 1728 -972 1734 -966
rect 1728 -978 1734 -972
rect 1728 -984 1734 -978
rect 1728 -990 1734 -984
rect 1728 -996 1734 -990
rect 1728 -1002 1734 -996
rect 1728 -1008 1734 -1002
rect 1728 -1014 1734 -1008
rect 1728 -1020 1734 -1014
rect 1728 -1026 1734 -1020
rect 1728 -1032 1734 -1026
rect 1728 -1038 1734 -1032
rect 1728 -1044 1734 -1038
rect 1728 -1050 1734 -1044
rect 1728 -1056 1734 -1050
rect 1728 -1062 1734 -1056
rect 1728 -1068 1734 -1062
rect 1728 -1074 1734 -1068
rect 1728 -1080 1734 -1074
rect 1728 -1086 1734 -1080
rect 1728 -1092 1734 -1086
rect 1728 -1098 1734 -1092
rect 1728 -1104 1734 -1098
rect 1728 -1110 1734 -1104
rect 1728 -1116 1734 -1110
rect 1728 -1122 1734 -1116
rect 1728 -1128 1734 -1122
rect 1728 -1134 1734 -1128
rect 1728 -1140 1734 -1134
rect 1728 -1146 1734 -1140
rect 1728 -1152 1734 -1146
rect 1728 -1158 1734 -1152
rect 1728 -1164 1734 -1158
rect 1728 -1170 1734 -1164
rect 1728 -1176 1734 -1170
rect 1728 -1182 1734 -1176
rect 1728 -1188 1734 -1182
rect 1728 -1194 1734 -1188
rect 1728 -1200 1734 -1194
rect 1728 -1206 1734 -1200
rect 1728 -1212 1734 -1206
rect 1728 -1218 1734 -1212
rect 1728 -1224 1734 -1218
rect 1728 -1230 1734 -1224
rect 1728 -1236 1734 -1230
rect 1728 -1242 1734 -1236
rect 1728 -1248 1734 -1242
rect 1728 -1254 1734 -1248
rect 1728 -1260 1734 -1254
rect 1728 -1266 1734 -1260
rect 1728 -1272 1734 -1266
rect 1728 -1278 1734 -1272
rect 1728 -1284 1734 -1278
rect 1728 -1290 1734 -1284
rect 1728 -1296 1734 -1290
rect 1728 -1302 1734 -1296
rect 1728 -1308 1734 -1302
rect 1728 -1314 1734 -1308
rect 1728 -1320 1734 -1314
rect 1728 -1326 1734 -1320
rect 1728 -1332 1734 -1326
rect 1728 -1338 1734 -1332
rect 1728 -1344 1734 -1338
rect 1728 -1350 1734 -1344
rect 1728 -1356 1734 -1350
rect 1728 -1362 1734 -1356
rect 1728 -1368 1734 -1362
rect 1728 -1374 1734 -1368
rect 1728 -1380 1734 -1374
rect 1728 -1386 1734 -1380
rect 1728 -1392 1734 -1386
rect 1728 -1398 1734 -1392
rect 1728 -1404 1734 -1398
rect 1728 -1410 1734 -1404
rect 1728 -1416 1734 -1410
rect 1728 -1422 1734 -1416
rect 1728 -1428 1734 -1422
rect 1728 -1434 1734 -1428
rect 1728 -1440 1734 -1434
rect 1728 -1446 1734 -1440
rect 1728 -1452 1734 -1446
rect 1728 -1458 1734 -1452
rect 1728 -1464 1734 -1458
rect 1728 -1470 1734 -1464
rect 1728 -1476 1734 -1470
rect 1728 -1482 1734 -1476
rect 1728 -1488 1734 -1482
rect 1728 -1494 1734 -1488
rect 1728 -1500 1734 -1494
rect 1728 -1506 1734 -1500
rect 1728 -1512 1734 -1506
rect 1728 -1518 1734 -1512
rect 1728 -1524 1734 -1518
rect 1728 -1530 1734 -1524
rect 1728 -1536 1734 -1530
rect 1728 -1542 1734 -1536
rect 1728 -1548 1734 -1542
rect 1728 -1554 1734 -1548
rect 1728 -1560 1734 -1554
rect 1728 -1566 1734 -1560
rect 1728 -1572 1734 -1566
rect 1728 -1578 1734 -1572
rect 1728 -1584 1734 -1578
rect 1728 -1590 1734 -1584
rect 1728 -1596 1734 -1590
rect 1728 -1602 1734 -1596
rect 1728 -1608 1734 -1602
rect 1728 -1614 1734 -1608
rect 1728 -1620 1734 -1614
rect 1728 -1626 1734 -1620
rect 1728 -1632 1734 -1626
rect 1728 -1638 1734 -1632
rect 1728 -1644 1734 -1638
rect 1728 -1650 1734 -1644
rect 1728 -1656 1734 -1650
rect 1728 -1662 1734 -1656
rect 1728 -1668 1734 -1662
rect 1728 -1674 1734 -1668
rect 1728 -1680 1734 -1674
rect 1728 -1686 1734 -1680
rect 1728 -1692 1734 -1686
rect 1728 -1698 1734 -1692
rect 1728 -1704 1734 -1698
rect 1728 -1710 1734 -1704
rect 1728 -1716 1734 -1710
rect 1728 -1722 1734 -1716
rect 1728 -1728 1734 -1722
rect 1728 -1734 1734 -1728
rect 1728 -1740 1734 -1734
rect 1728 -1746 1734 -1740
rect 1728 -1752 1734 -1746
rect 1728 -1758 1734 -1752
rect 1728 -1764 1734 -1758
rect 1728 -1770 1734 -1764
rect 1728 -1776 1734 -1770
rect 1728 -1782 1734 -1776
rect 1728 -1788 1734 -1782
rect 1728 -1794 1734 -1788
rect 1728 -1800 1734 -1794
rect 1728 -1806 1734 -1800
rect 1728 -1812 1734 -1806
rect 1728 -1818 1734 -1812
rect 1728 -1824 1734 -1818
rect 1728 -1830 1734 -1824
rect 1728 -1836 1734 -1830
rect 1728 -1842 1734 -1836
rect 1728 -1848 1734 -1842
rect 1728 -1854 1734 -1848
rect 1728 -1860 1734 -1854
rect 1728 -1866 1734 -1860
rect 1728 -1872 1734 -1866
rect 1728 -1878 1734 -1872
rect 1728 -1884 1734 -1878
rect 1728 -1890 1734 -1884
rect 1728 -1896 1734 -1890
rect 1728 -1902 1734 -1896
rect 1728 -1908 1734 -1902
rect 1728 -1914 1734 -1908
rect 1728 -1920 1734 -1914
rect 1728 -1926 1734 -1920
rect 1728 -2004 1734 -1998
rect 1728 -2010 1734 -2004
rect 1728 -2016 1734 -2010
rect 1728 -2022 1734 -2016
rect 1728 -2028 1734 -2022
rect 1728 -2034 1734 -2028
rect 1728 -2040 1734 -2034
rect 1728 -2046 1734 -2040
rect 1728 -2052 1734 -2046
rect 1728 -2058 1734 -2052
rect 1728 -2064 1734 -2058
rect 1728 -2070 1734 -2064
rect 1728 -2076 1734 -2070
rect 1728 -2082 1734 -2076
rect 1728 -2088 1734 -2082
rect 1728 -2094 1734 -2088
rect 1728 -2100 1734 -2094
rect 1728 -2106 1734 -2100
rect 1728 -2112 1734 -2106
rect 1728 -2118 1734 -2112
rect 1728 -2124 1734 -2118
rect 1728 -2130 1734 -2124
rect 1728 -2136 1734 -2130
rect 1728 -2142 1734 -2136
rect 1728 -2148 1734 -2142
rect 1728 -2154 1734 -2148
rect 1728 -2160 1734 -2154
rect 1728 -2166 1734 -2160
rect 1728 -2172 1734 -2166
rect 1728 -2178 1734 -2172
rect 1728 -2184 1734 -2178
rect 1728 -2190 1734 -2184
rect 1728 -2196 1734 -2190
rect 1728 -2202 1734 -2196
rect 1728 -2208 1734 -2202
rect 1728 -2214 1734 -2208
rect 1728 -2220 1734 -2214
rect 1728 -2226 1734 -2220
rect 1728 -2232 1734 -2226
rect 1728 -2238 1734 -2232
rect 1728 -2244 1734 -2238
rect 1728 -2250 1734 -2244
rect 1728 -2256 1734 -2250
rect 1728 -2262 1734 -2256
rect 1728 -2268 1734 -2262
rect 1728 -2274 1734 -2268
rect 1728 -2280 1734 -2274
rect 1728 -2286 1734 -2280
rect 1728 -2292 1734 -2286
rect 1728 -2298 1734 -2292
rect 1728 -2304 1734 -2298
rect 1728 -2310 1734 -2304
rect 1728 -2316 1734 -2310
rect 1728 -2322 1734 -2316
rect 1728 -2328 1734 -2322
rect 1728 -2334 1734 -2328
rect 1728 -2340 1734 -2334
rect 1728 -2346 1734 -2340
rect 1728 -2352 1734 -2346
rect 1728 -2358 1734 -2352
rect 1728 -2364 1734 -2358
rect 1728 -2370 1734 -2364
rect 1728 -2376 1734 -2370
rect 1728 -2382 1734 -2376
rect 1728 -2388 1734 -2382
rect 1728 -2394 1734 -2388
rect 1728 -2400 1734 -2394
rect 1728 -2406 1734 -2400
rect 1728 -2412 1734 -2406
rect 1728 -2418 1734 -2412
rect 1728 -2424 1734 -2418
rect 1728 -2430 1734 -2424
rect 1728 -2436 1734 -2430
rect 1728 -2442 1734 -2436
rect 1728 -2448 1734 -2442
rect 1728 -2454 1734 -2448
rect 1728 -2460 1734 -2454
rect 1728 -2466 1734 -2460
rect 1728 -2472 1734 -2466
rect 1728 -2478 1734 -2472
rect 1728 -2484 1734 -2478
rect 1728 -2490 1734 -2484
rect 1728 -2496 1734 -2490
rect 1728 -2502 1734 -2496
rect 1728 -2508 1734 -2502
rect 1728 -2514 1734 -2508
rect 1728 -2520 1734 -2514
rect 1728 -2526 1734 -2520
rect 1728 -2532 1734 -2526
rect 1728 -2538 1734 -2532
rect 1728 -2544 1734 -2538
rect 1728 -2550 1734 -2544
rect 1728 -2556 1734 -2550
rect 1728 -2562 1734 -2556
rect 1728 -2568 1734 -2562
rect 1728 -2574 1734 -2568
rect 1728 -2580 1734 -2574
rect 1728 -2586 1734 -2580
rect 1728 -2592 1734 -2586
rect 1728 -2598 1734 -2592
rect 1728 -2604 1734 -2598
rect 1728 -2610 1734 -2604
rect 1728 -2616 1734 -2610
rect 1728 -2622 1734 -2616
rect 1728 -2628 1734 -2622
rect 1728 -2634 1734 -2628
rect 1728 -2640 1734 -2634
rect 1728 -2646 1734 -2640
rect 1728 -2652 1734 -2646
rect 1728 -2658 1734 -2652
rect 1728 -2664 1734 -2658
rect 1728 -2670 1734 -2664
rect 1728 -2748 1734 -2742
rect 1728 -2754 1734 -2748
rect 1728 -2760 1734 -2754
rect 1728 -2766 1734 -2760
rect 1728 -2772 1734 -2766
rect 1728 -2778 1734 -2772
rect 1728 -2784 1734 -2778
rect 1728 -2790 1734 -2784
rect 1728 -2796 1734 -2790
rect 1728 -2802 1734 -2796
rect 1728 -2808 1734 -2802
rect 1728 -2814 1734 -2808
rect 1728 -2820 1734 -2814
rect 1728 -2826 1734 -2820
rect 1728 -2832 1734 -2826
rect 1728 -2838 1734 -2832
rect 1728 -2844 1734 -2838
rect 1728 -2850 1734 -2844
rect 1728 -2856 1734 -2850
rect 1728 -2862 1734 -2856
rect 1728 -2868 1734 -2862
rect 1728 -2874 1734 -2868
rect 1728 -2880 1734 -2874
rect 1728 -2886 1734 -2880
rect 1728 -2892 1734 -2886
rect 1728 -2898 1734 -2892
rect 1728 -2904 1734 -2898
rect 1728 -2910 1734 -2904
rect 1728 -2916 1734 -2910
rect 1728 -2922 1734 -2916
rect 1728 -2928 1734 -2922
rect 1728 -2934 1734 -2928
rect 1728 -2940 1734 -2934
rect 1728 -2946 1734 -2940
rect 1728 -2952 1734 -2946
rect 1728 -2958 1734 -2952
rect 1728 -2964 1734 -2958
rect 1728 -2970 1734 -2964
rect 1728 -2976 1734 -2970
rect 1728 -2982 1734 -2976
rect 1728 -2988 1734 -2982
rect 1728 -2994 1734 -2988
rect 1728 -3000 1734 -2994
rect 1728 -3006 1734 -3000
rect 1728 -3012 1734 -3006
rect 1728 -3018 1734 -3012
rect 1728 -3024 1734 -3018
rect 1728 -3030 1734 -3024
rect 1728 -3036 1734 -3030
rect 1728 -3042 1734 -3036
rect 1728 -3048 1734 -3042
rect 1728 -3054 1734 -3048
rect 1728 -3060 1734 -3054
rect 1728 -3066 1734 -3060
rect 1728 -3072 1734 -3066
rect 1728 -3078 1734 -3072
rect 1728 -3084 1734 -3078
rect 1728 -3090 1734 -3084
rect 1728 -3096 1734 -3090
rect 1728 -3102 1734 -3096
rect 1728 -3108 1734 -3102
rect 1728 -3114 1734 -3108
rect 1728 -3120 1734 -3114
rect 1728 -3126 1734 -3120
rect 1728 -3132 1734 -3126
rect 1728 -3138 1734 -3132
rect 1728 -3144 1734 -3138
rect 1728 -3150 1734 -3144
rect 1728 -3156 1734 -3150
rect 1728 -3162 1734 -3156
rect 1728 -3168 1734 -3162
rect 1728 -3174 1734 -3168
rect 1728 -3180 1734 -3174
rect 1728 -3186 1734 -3180
rect 1728 -3192 1734 -3186
rect 1728 -3198 1734 -3192
rect 1728 -3204 1734 -3198
rect 1728 -3210 1734 -3204
rect 1728 -3258 1734 -3252
rect 1728 -3264 1734 -3258
rect 1728 -3270 1734 -3264
rect 1728 -3276 1734 -3270
rect 1728 -3282 1734 -3276
rect 1728 -3288 1734 -3282
rect 1728 -3294 1734 -3288
rect 1728 -3300 1734 -3294
rect 1728 -3306 1734 -3300
rect 1728 -3312 1734 -3306
rect 1728 -3318 1734 -3312
rect 1728 -3324 1734 -3318
rect 1728 -3330 1734 -3324
rect 1728 -3336 1734 -3330
rect 1728 -3342 1734 -3336
rect 1728 -3348 1734 -3342
rect 1728 -3354 1734 -3348
rect 1728 -3360 1734 -3354
rect 1728 -3366 1734 -3360
rect 1728 -3372 1734 -3366
rect 1728 -3378 1734 -3372
rect 1728 -3384 1734 -3378
rect 1728 -3390 1734 -3384
rect 1728 -3396 1734 -3390
rect 1728 -3402 1734 -3396
rect 1728 -3408 1734 -3402
rect 1734 -816 1740 -810
rect 1734 -822 1740 -816
rect 1734 -828 1740 -822
rect 1734 -834 1740 -828
rect 1734 -840 1740 -834
rect 1734 -846 1740 -840
rect 1734 -852 1740 -846
rect 1734 -858 1740 -852
rect 1734 -864 1740 -858
rect 1734 -870 1740 -864
rect 1734 -876 1740 -870
rect 1734 -882 1740 -876
rect 1734 -888 1740 -882
rect 1734 -894 1740 -888
rect 1734 -900 1740 -894
rect 1734 -906 1740 -900
rect 1734 -912 1740 -906
rect 1734 -918 1740 -912
rect 1734 -924 1740 -918
rect 1734 -930 1740 -924
rect 1734 -936 1740 -930
rect 1734 -942 1740 -936
rect 1734 -948 1740 -942
rect 1734 -954 1740 -948
rect 1734 -960 1740 -954
rect 1734 -966 1740 -960
rect 1734 -972 1740 -966
rect 1734 -978 1740 -972
rect 1734 -984 1740 -978
rect 1734 -990 1740 -984
rect 1734 -996 1740 -990
rect 1734 -1002 1740 -996
rect 1734 -1008 1740 -1002
rect 1734 -1014 1740 -1008
rect 1734 -1020 1740 -1014
rect 1734 -1026 1740 -1020
rect 1734 -1032 1740 -1026
rect 1734 -1038 1740 -1032
rect 1734 -1044 1740 -1038
rect 1734 -1050 1740 -1044
rect 1734 -1056 1740 -1050
rect 1734 -1062 1740 -1056
rect 1734 -1068 1740 -1062
rect 1734 -1074 1740 -1068
rect 1734 -1080 1740 -1074
rect 1734 -1086 1740 -1080
rect 1734 -1092 1740 -1086
rect 1734 -1098 1740 -1092
rect 1734 -1104 1740 -1098
rect 1734 -1110 1740 -1104
rect 1734 -1116 1740 -1110
rect 1734 -1122 1740 -1116
rect 1734 -1128 1740 -1122
rect 1734 -1134 1740 -1128
rect 1734 -1140 1740 -1134
rect 1734 -1146 1740 -1140
rect 1734 -1152 1740 -1146
rect 1734 -1158 1740 -1152
rect 1734 -1164 1740 -1158
rect 1734 -1170 1740 -1164
rect 1734 -1176 1740 -1170
rect 1734 -1182 1740 -1176
rect 1734 -1188 1740 -1182
rect 1734 -1194 1740 -1188
rect 1734 -1200 1740 -1194
rect 1734 -1206 1740 -1200
rect 1734 -1212 1740 -1206
rect 1734 -1218 1740 -1212
rect 1734 -1224 1740 -1218
rect 1734 -1230 1740 -1224
rect 1734 -1236 1740 -1230
rect 1734 -1242 1740 -1236
rect 1734 -1248 1740 -1242
rect 1734 -1254 1740 -1248
rect 1734 -1260 1740 -1254
rect 1734 -1266 1740 -1260
rect 1734 -1272 1740 -1266
rect 1734 -1278 1740 -1272
rect 1734 -1284 1740 -1278
rect 1734 -1290 1740 -1284
rect 1734 -1296 1740 -1290
rect 1734 -1302 1740 -1296
rect 1734 -1308 1740 -1302
rect 1734 -1314 1740 -1308
rect 1734 -1320 1740 -1314
rect 1734 -1326 1740 -1320
rect 1734 -1332 1740 -1326
rect 1734 -1338 1740 -1332
rect 1734 -1344 1740 -1338
rect 1734 -1350 1740 -1344
rect 1734 -1356 1740 -1350
rect 1734 -1362 1740 -1356
rect 1734 -1368 1740 -1362
rect 1734 -1374 1740 -1368
rect 1734 -1380 1740 -1374
rect 1734 -1386 1740 -1380
rect 1734 -1392 1740 -1386
rect 1734 -1398 1740 -1392
rect 1734 -1404 1740 -1398
rect 1734 -1410 1740 -1404
rect 1734 -1416 1740 -1410
rect 1734 -1422 1740 -1416
rect 1734 -1428 1740 -1422
rect 1734 -1434 1740 -1428
rect 1734 -1440 1740 -1434
rect 1734 -1446 1740 -1440
rect 1734 -1452 1740 -1446
rect 1734 -1458 1740 -1452
rect 1734 -1464 1740 -1458
rect 1734 -1470 1740 -1464
rect 1734 -1476 1740 -1470
rect 1734 -1482 1740 -1476
rect 1734 -1488 1740 -1482
rect 1734 -1494 1740 -1488
rect 1734 -1500 1740 -1494
rect 1734 -1506 1740 -1500
rect 1734 -1512 1740 -1506
rect 1734 -1518 1740 -1512
rect 1734 -1524 1740 -1518
rect 1734 -1530 1740 -1524
rect 1734 -1536 1740 -1530
rect 1734 -1542 1740 -1536
rect 1734 -1548 1740 -1542
rect 1734 -1554 1740 -1548
rect 1734 -1560 1740 -1554
rect 1734 -1566 1740 -1560
rect 1734 -1572 1740 -1566
rect 1734 -1578 1740 -1572
rect 1734 -1584 1740 -1578
rect 1734 -1590 1740 -1584
rect 1734 -1596 1740 -1590
rect 1734 -1602 1740 -1596
rect 1734 -1608 1740 -1602
rect 1734 -1614 1740 -1608
rect 1734 -1620 1740 -1614
rect 1734 -1626 1740 -1620
rect 1734 -1632 1740 -1626
rect 1734 -1638 1740 -1632
rect 1734 -1644 1740 -1638
rect 1734 -1650 1740 -1644
rect 1734 -1656 1740 -1650
rect 1734 -1662 1740 -1656
rect 1734 -1668 1740 -1662
rect 1734 -1674 1740 -1668
rect 1734 -1680 1740 -1674
rect 1734 -1686 1740 -1680
rect 1734 -1692 1740 -1686
rect 1734 -1698 1740 -1692
rect 1734 -1704 1740 -1698
rect 1734 -1710 1740 -1704
rect 1734 -1716 1740 -1710
rect 1734 -1722 1740 -1716
rect 1734 -1728 1740 -1722
rect 1734 -1734 1740 -1728
rect 1734 -1740 1740 -1734
rect 1734 -1746 1740 -1740
rect 1734 -1752 1740 -1746
rect 1734 -1758 1740 -1752
rect 1734 -1764 1740 -1758
rect 1734 -1770 1740 -1764
rect 1734 -1776 1740 -1770
rect 1734 -1782 1740 -1776
rect 1734 -1788 1740 -1782
rect 1734 -1794 1740 -1788
rect 1734 -1800 1740 -1794
rect 1734 -1806 1740 -1800
rect 1734 -1812 1740 -1806
rect 1734 -1818 1740 -1812
rect 1734 -1824 1740 -1818
rect 1734 -1830 1740 -1824
rect 1734 -1836 1740 -1830
rect 1734 -1842 1740 -1836
rect 1734 -1848 1740 -1842
rect 1734 -1854 1740 -1848
rect 1734 -1860 1740 -1854
rect 1734 -1866 1740 -1860
rect 1734 -1872 1740 -1866
rect 1734 -1878 1740 -1872
rect 1734 -1884 1740 -1878
rect 1734 -1890 1740 -1884
rect 1734 -1896 1740 -1890
rect 1734 -1902 1740 -1896
rect 1734 -1908 1740 -1902
rect 1734 -1914 1740 -1908
rect 1734 -1920 1740 -1914
rect 1734 -1992 1740 -1986
rect 1734 -1998 1740 -1992
rect 1734 -2004 1740 -1998
rect 1734 -2010 1740 -2004
rect 1734 -2016 1740 -2010
rect 1734 -2022 1740 -2016
rect 1734 -2028 1740 -2022
rect 1734 -2034 1740 -2028
rect 1734 -2040 1740 -2034
rect 1734 -2046 1740 -2040
rect 1734 -2052 1740 -2046
rect 1734 -2058 1740 -2052
rect 1734 -2064 1740 -2058
rect 1734 -2070 1740 -2064
rect 1734 -2076 1740 -2070
rect 1734 -2082 1740 -2076
rect 1734 -2088 1740 -2082
rect 1734 -2094 1740 -2088
rect 1734 -2100 1740 -2094
rect 1734 -2106 1740 -2100
rect 1734 -2112 1740 -2106
rect 1734 -2118 1740 -2112
rect 1734 -2124 1740 -2118
rect 1734 -2130 1740 -2124
rect 1734 -2136 1740 -2130
rect 1734 -2142 1740 -2136
rect 1734 -2148 1740 -2142
rect 1734 -2154 1740 -2148
rect 1734 -2160 1740 -2154
rect 1734 -2166 1740 -2160
rect 1734 -2172 1740 -2166
rect 1734 -2178 1740 -2172
rect 1734 -2184 1740 -2178
rect 1734 -2190 1740 -2184
rect 1734 -2196 1740 -2190
rect 1734 -2202 1740 -2196
rect 1734 -2208 1740 -2202
rect 1734 -2214 1740 -2208
rect 1734 -2220 1740 -2214
rect 1734 -2226 1740 -2220
rect 1734 -2232 1740 -2226
rect 1734 -2238 1740 -2232
rect 1734 -2244 1740 -2238
rect 1734 -2250 1740 -2244
rect 1734 -2256 1740 -2250
rect 1734 -2262 1740 -2256
rect 1734 -2268 1740 -2262
rect 1734 -2274 1740 -2268
rect 1734 -2280 1740 -2274
rect 1734 -2286 1740 -2280
rect 1734 -2292 1740 -2286
rect 1734 -2298 1740 -2292
rect 1734 -2304 1740 -2298
rect 1734 -2310 1740 -2304
rect 1734 -2316 1740 -2310
rect 1734 -2322 1740 -2316
rect 1734 -2328 1740 -2322
rect 1734 -2334 1740 -2328
rect 1734 -2340 1740 -2334
rect 1734 -2346 1740 -2340
rect 1734 -2352 1740 -2346
rect 1734 -2358 1740 -2352
rect 1734 -2364 1740 -2358
rect 1734 -2370 1740 -2364
rect 1734 -2376 1740 -2370
rect 1734 -2382 1740 -2376
rect 1734 -2388 1740 -2382
rect 1734 -2394 1740 -2388
rect 1734 -2400 1740 -2394
rect 1734 -2406 1740 -2400
rect 1734 -2412 1740 -2406
rect 1734 -2418 1740 -2412
rect 1734 -2424 1740 -2418
rect 1734 -2430 1740 -2424
rect 1734 -2436 1740 -2430
rect 1734 -2442 1740 -2436
rect 1734 -2448 1740 -2442
rect 1734 -2454 1740 -2448
rect 1734 -2460 1740 -2454
rect 1734 -2466 1740 -2460
rect 1734 -2472 1740 -2466
rect 1734 -2478 1740 -2472
rect 1734 -2484 1740 -2478
rect 1734 -2490 1740 -2484
rect 1734 -2496 1740 -2490
rect 1734 -2502 1740 -2496
rect 1734 -2508 1740 -2502
rect 1734 -2514 1740 -2508
rect 1734 -2520 1740 -2514
rect 1734 -2526 1740 -2520
rect 1734 -2532 1740 -2526
rect 1734 -2538 1740 -2532
rect 1734 -2544 1740 -2538
rect 1734 -2550 1740 -2544
rect 1734 -2556 1740 -2550
rect 1734 -2562 1740 -2556
rect 1734 -2568 1740 -2562
rect 1734 -2574 1740 -2568
rect 1734 -2580 1740 -2574
rect 1734 -2586 1740 -2580
rect 1734 -2592 1740 -2586
rect 1734 -2598 1740 -2592
rect 1734 -2604 1740 -2598
rect 1734 -2610 1740 -2604
rect 1734 -2616 1740 -2610
rect 1734 -2622 1740 -2616
rect 1734 -2628 1740 -2622
rect 1734 -2634 1740 -2628
rect 1734 -2640 1740 -2634
rect 1734 -2646 1740 -2640
rect 1734 -2652 1740 -2646
rect 1734 -2658 1740 -2652
rect 1734 -2664 1740 -2658
rect 1734 -2670 1740 -2664
rect 1734 -2742 1740 -2736
rect 1734 -2748 1740 -2742
rect 1734 -2754 1740 -2748
rect 1734 -2760 1740 -2754
rect 1734 -2766 1740 -2760
rect 1734 -2772 1740 -2766
rect 1734 -2778 1740 -2772
rect 1734 -2784 1740 -2778
rect 1734 -2790 1740 -2784
rect 1734 -2796 1740 -2790
rect 1734 -2802 1740 -2796
rect 1734 -2808 1740 -2802
rect 1734 -2814 1740 -2808
rect 1734 -2820 1740 -2814
rect 1734 -2826 1740 -2820
rect 1734 -2832 1740 -2826
rect 1734 -2838 1740 -2832
rect 1734 -2844 1740 -2838
rect 1734 -2850 1740 -2844
rect 1734 -2856 1740 -2850
rect 1734 -2862 1740 -2856
rect 1734 -2868 1740 -2862
rect 1734 -2874 1740 -2868
rect 1734 -2880 1740 -2874
rect 1734 -2886 1740 -2880
rect 1734 -2892 1740 -2886
rect 1734 -2898 1740 -2892
rect 1734 -2904 1740 -2898
rect 1734 -2910 1740 -2904
rect 1734 -2916 1740 -2910
rect 1734 -2922 1740 -2916
rect 1734 -2928 1740 -2922
rect 1734 -2934 1740 -2928
rect 1734 -2940 1740 -2934
rect 1734 -2946 1740 -2940
rect 1734 -2952 1740 -2946
rect 1734 -2958 1740 -2952
rect 1734 -2964 1740 -2958
rect 1734 -2970 1740 -2964
rect 1734 -2976 1740 -2970
rect 1734 -2982 1740 -2976
rect 1734 -2988 1740 -2982
rect 1734 -2994 1740 -2988
rect 1734 -3000 1740 -2994
rect 1734 -3006 1740 -3000
rect 1734 -3012 1740 -3006
rect 1734 -3018 1740 -3012
rect 1734 -3024 1740 -3018
rect 1734 -3030 1740 -3024
rect 1734 -3036 1740 -3030
rect 1734 -3042 1740 -3036
rect 1734 -3048 1740 -3042
rect 1734 -3054 1740 -3048
rect 1734 -3060 1740 -3054
rect 1734 -3066 1740 -3060
rect 1734 -3072 1740 -3066
rect 1734 -3078 1740 -3072
rect 1734 -3084 1740 -3078
rect 1734 -3090 1740 -3084
rect 1734 -3096 1740 -3090
rect 1734 -3102 1740 -3096
rect 1734 -3108 1740 -3102
rect 1734 -3114 1740 -3108
rect 1734 -3120 1740 -3114
rect 1734 -3126 1740 -3120
rect 1734 -3132 1740 -3126
rect 1734 -3138 1740 -3132
rect 1734 -3144 1740 -3138
rect 1734 -3150 1740 -3144
rect 1734 -3156 1740 -3150
rect 1734 -3162 1740 -3156
rect 1734 -3168 1740 -3162
rect 1734 -3174 1740 -3168
rect 1734 -3180 1740 -3174
rect 1734 -3186 1740 -3180
rect 1734 -3192 1740 -3186
rect 1734 -3198 1740 -3192
rect 1734 -3204 1740 -3198
rect 1734 -3210 1740 -3204
rect 1734 -3258 1740 -3252
rect 1734 -3264 1740 -3258
rect 1734 -3270 1740 -3264
rect 1734 -3276 1740 -3270
rect 1734 -3282 1740 -3276
rect 1734 -3288 1740 -3282
rect 1734 -3294 1740 -3288
rect 1734 -3300 1740 -3294
rect 1734 -3306 1740 -3300
rect 1734 -3312 1740 -3306
rect 1734 -3318 1740 -3312
rect 1734 -3324 1740 -3318
rect 1734 -3330 1740 -3324
rect 1734 -3336 1740 -3330
rect 1734 -3342 1740 -3336
rect 1734 -3348 1740 -3342
rect 1734 -3354 1740 -3348
rect 1734 -3360 1740 -3354
rect 1734 -3366 1740 -3360
rect 1734 -3372 1740 -3366
rect 1734 -3378 1740 -3372
rect 1734 -3384 1740 -3378
rect 1734 -3390 1740 -3384
rect 1734 -3396 1740 -3390
rect 1734 -3402 1740 -3396
rect 1740 -804 1746 -798
rect 1740 -810 1746 -804
rect 1740 -816 1746 -810
rect 1740 -822 1746 -816
rect 1740 -828 1746 -822
rect 1740 -834 1746 -828
rect 1740 -840 1746 -834
rect 1740 -846 1746 -840
rect 1740 -852 1746 -846
rect 1740 -858 1746 -852
rect 1740 -864 1746 -858
rect 1740 -870 1746 -864
rect 1740 -876 1746 -870
rect 1740 -882 1746 -876
rect 1740 -888 1746 -882
rect 1740 -894 1746 -888
rect 1740 -900 1746 -894
rect 1740 -906 1746 -900
rect 1740 -912 1746 -906
rect 1740 -918 1746 -912
rect 1740 -924 1746 -918
rect 1740 -930 1746 -924
rect 1740 -936 1746 -930
rect 1740 -942 1746 -936
rect 1740 -948 1746 -942
rect 1740 -954 1746 -948
rect 1740 -960 1746 -954
rect 1740 -966 1746 -960
rect 1740 -972 1746 -966
rect 1740 -978 1746 -972
rect 1740 -984 1746 -978
rect 1740 -990 1746 -984
rect 1740 -996 1746 -990
rect 1740 -1002 1746 -996
rect 1740 -1008 1746 -1002
rect 1740 -1014 1746 -1008
rect 1740 -1020 1746 -1014
rect 1740 -1026 1746 -1020
rect 1740 -1032 1746 -1026
rect 1740 -1038 1746 -1032
rect 1740 -1044 1746 -1038
rect 1740 -1050 1746 -1044
rect 1740 -1056 1746 -1050
rect 1740 -1062 1746 -1056
rect 1740 -1068 1746 -1062
rect 1740 -1074 1746 -1068
rect 1740 -1080 1746 -1074
rect 1740 -1086 1746 -1080
rect 1740 -1092 1746 -1086
rect 1740 -1098 1746 -1092
rect 1740 -1104 1746 -1098
rect 1740 -1110 1746 -1104
rect 1740 -1116 1746 -1110
rect 1740 -1122 1746 -1116
rect 1740 -1128 1746 -1122
rect 1740 -1134 1746 -1128
rect 1740 -1140 1746 -1134
rect 1740 -1146 1746 -1140
rect 1740 -1152 1746 -1146
rect 1740 -1158 1746 -1152
rect 1740 -1164 1746 -1158
rect 1740 -1170 1746 -1164
rect 1740 -1176 1746 -1170
rect 1740 -1182 1746 -1176
rect 1740 -1188 1746 -1182
rect 1740 -1194 1746 -1188
rect 1740 -1200 1746 -1194
rect 1740 -1206 1746 -1200
rect 1740 -1212 1746 -1206
rect 1740 -1218 1746 -1212
rect 1740 -1224 1746 -1218
rect 1740 -1230 1746 -1224
rect 1740 -1236 1746 -1230
rect 1740 -1242 1746 -1236
rect 1740 -1248 1746 -1242
rect 1740 -1254 1746 -1248
rect 1740 -1260 1746 -1254
rect 1740 -1266 1746 -1260
rect 1740 -1272 1746 -1266
rect 1740 -1278 1746 -1272
rect 1740 -1284 1746 -1278
rect 1740 -1290 1746 -1284
rect 1740 -1296 1746 -1290
rect 1740 -1302 1746 -1296
rect 1740 -1308 1746 -1302
rect 1740 -1314 1746 -1308
rect 1740 -1320 1746 -1314
rect 1740 -1326 1746 -1320
rect 1740 -1332 1746 -1326
rect 1740 -1338 1746 -1332
rect 1740 -1344 1746 -1338
rect 1740 -1350 1746 -1344
rect 1740 -1356 1746 -1350
rect 1740 -1362 1746 -1356
rect 1740 -1368 1746 -1362
rect 1740 -1374 1746 -1368
rect 1740 -1380 1746 -1374
rect 1740 -1386 1746 -1380
rect 1740 -1392 1746 -1386
rect 1740 -1398 1746 -1392
rect 1740 -1404 1746 -1398
rect 1740 -1410 1746 -1404
rect 1740 -1416 1746 -1410
rect 1740 -1422 1746 -1416
rect 1740 -1428 1746 -1422
rect 1740 -1434 1746 -1428
rect 1740 -1440 1746 -1434
rect 1740 -1446 1746 -1440
rect 1740 -1452 1746 -1446
rect 1740 -1458 1746 -1452
rect 1740 -1464 1746 -1458
rect 1740 -1470 1746 -1464
rect 1740 -1476 1746 -1470
rect 1740 -1482 1746 -1476
rect 1740 -1488 1746 -1482
rect 1740 -1494 1746 -1488
rect 1740 -1500 1746 -1494
rect 1740 -1506 1746 -1500
rect 1740 -1512 1746 -1506
rect 1740 -1518 1746 -1512
rect 1740 -1524 1746 -1518
rect 1740 -1530 1746 -1524
rect 1740 -1536 1746 -1530
rect 1740 -1542 1746 -1536
rect 1740 -1548 1746 -1542
rect 1740 -1554 1746 -1548
rect 1740 -1560 1746 -1554
rect 1740 -1566 1746 -1560
rect 1740 -1572 1746 -1566
rect 1740 -1578 1746 -1572
rect 1740 -1584 1746 -1578
rect 1740 -1590 1746 -1584
rect 1740 -1596 1746 -1590
rect 1740 -1602 1746 -1596
rect 1740 -1608 1746 -1602
rect 1740 -1614 1746 -1608
rect 1740 -1620 1746 -1614
rect 1740 -1626 1746 -1620
rect 1740 -1632 1746 -1626
rect 1740 -1638 1746 -1632
rect 1740 -1644 1746 -1638
rect 1740 -1650 1746 -1644
rect 1740 -1656 1746 -1650
rect 1740 -1662 1746 -1656
rect 1740 -1668 1746 -1662
rect 1740 -1674 1746 -1668
rect 1740 -1680 1746 -1674
rect 1740 -1686 1746 -1680
rect 1740 -1692 1746 -1686
rect 1740 -1698 1746 -1692
rect 1740 -1704 1746 -1698
rect 1740 -1710 1746 -1704
rect 1740 -1716 1746 -1710
rect 1740 -1722 1746 -1716
rect 1740 -1728 1746 -1722
rect 1740 -1734 1746 -1728
rect 1740 -1740 1746 -1734
rect 1740 -1746 1746 -1740
rect 1740 -1752 1746 -1746
rect 1740 -1758 1746 -1752
rect 1740 -1764 1746 -1758
rect 1740 -1770 1746 -1764
rect 1740 -1776 1746 -1770
rect 1740 -1782 1746 -1776
rect 1740 -1788 1746 -1782
rect 1740 -1794 1746 -1788
rect 1740 -1800 1746 -1794
rect 1740 -1806 1746 -1800
rect 1740 -1812 1746 -1806
rect 1740 -1818 1746 -1812
rect 1740 -1824 1746 -1818
rect 1740 -1830 1746 -1824
rect 1740 -1836 1746 -1830
rect 1740 -1842 1746 -1836
rect 1740 -1848 1746 -1842
rect 1740 -1854 1746 -1848
rect 1740 -1860 1746 -1854
rect 1740 -1866 1746 -1860
rect 1740 -1872 1746 -1866
rect 1740 -1878 1746 -1872
rect 1740 -1884 1746 -1878
rect 1740 -1890 1746 -1884
rect 1740 -1896 1746 -1890
rect 1740 -1902 1746 -1896
rect 1740 -1908 1746 -1902
rect 1740 -1914 1746 -1908
rect 1740 -1986 1746 -1980
rect 1740 -1992 1746 -1986
rect 1740 -1998 1746 -1992
rect 1740 -2004 1746 -1998
rect 1740 -2010 1746 -2004
rect 1740 -2016 1746 -2010
rect 1740 -2022 1746 -2016
rect 1740 -2028 1746 -2022
rect 1740 -2034 1746 -2028
rect 1740 -2040 1746 -2034
rect 1740 -2046 1746 -2040
rect 1740 -2052 1746 -2046
rect 1740 -2058 1746 -2052
rect 1740 -2064 1746 -2058
rect 1740 -2070 1746 -2064
rect 1740 -2076 1746 -2070
rect 1740 -2082 1746 -2076
rect 1740 -2088 1746 -2082
rect 1740 -2094 1746 -2088
rect 1740 -2100 1746 -2094
rect 1740 -2106 1746 -2100
rect 1740 -2112 1746 -2106
rect 1740 -2118 1746 -2112
rect 1740 -2124 1746 -2118
rect 1740 -2130 1746 -2124
rect 1740 -2136 1746 -2130
rect 1740 -2142 1746 -2136
rect 1740 -2148 1746 -2142
rect 1740 -2154 1746 -2148
rect 1740 -2160 1746 -2154
rect 1740 -2166 1746 -2160
rect 1740 -2172 1746 -2166
rect 1740 -2178 1746 -2172
rect 1740 -2184 1746 -2178
rect 1740 -2190 1746 -2184
rect 1740 -2196 1746 -2190
rect 1740 -2202 1746 -2196
rect 1740 -2208 1746 -2202
rect 1740 -2214 1746 -2208
rect 1740 -2220 1746 -2214
rect 1740 -2226 1746 -2220
rect 1740 -2232 1746 -2226
rect 1740 -2238 1746 -2232
rect 1740 -2244 1746 -2238
rect 1740 -2250 1746 -2244
rect 1740 -2256 1746 -2250
rect 1740 -2262 1746 -2256
rect 1740 -2268 1746 -2262
rect 1740 -2274 1746 -2268
rect 1740 -2280 1746 -2274
rect 1740 -2286 1746 -2280
rect 1740 -2292 1746 -2286
rect 1740 -2298 1746 -2292
rect 1740 -2304 1746 -2298
rect 1740 -2310 1746 -2304
rect 1740 -2316 1746 -2310
rect 1740 -2322 1746 -2316
rect 1740 -2328 1746 -2322
rect 1740 -2334 1746 -2328
rect 1740 -2340 1746 -2334
rect 1740 -2346 1746 -2340
rect 1740 -2352 1746 -2346
rect 1740 -2358 1746 -2352
rect 1740 -2364 1746 -2358
rect 1740 -2370 1746 -2364
rect 1740 -2376 1746 -2370
rect 1740 -2382 1746 -2376
rect 1740 -2388 1746 -2382
rect 1740 -2394 1746 -2388
rect 1740 -2400 1746 -2394
rect 1740 -2406 1746 -2400
rect 1740 -2412 1746 -2406
rect 1740 -2418 1746 -2412
rect 1740 -2424 1746 -2418
rect 1740 -2430 1746 -2424
rect 1740 -2436 1746 -2430
rect 1740 -2442 1746 -2436
rect 1740 -2448 1746 -2442
rect 1740 -2454 1746 -2448
rect 1740 -2460 1746 -2454
rect 1740 -2466 1746 -2460
rect 1740 -2472 1746 -2466
rect 1740 -2478 1746 -2472
rect 1740 -2484 1746 -2478
rect 1740 -2490 1746 -2484
rect 1740 -2496 1746 -2490
rect 1740 -2502 1746 -2496
rect 1740 -2508 1746 -2502
rect 1740 -2514 1746 -2508
rect 1740 -2520 1746 -2514
rect 1740 -2526 1746 -2520
rect 1740 -2532 1746 -2526
rect 1740 -2538 1746 -2532
rect 1740 -2544 1746 -2538
rect 1740 -2550 1746 -2544
rect 1740 -2556 1746 -2550
rect 1740 -2562 1746 -2556
rect 1740 -2568 1746 -2562
rect 1740 -2574 1746 -2568
rect 1740 -2580 1746 -2574
rect 1740 -2586 1746 -2580
rect 1740 -2592 1746 -2586
rect 1740 -2598 1746 -2592
rect 1740 -2604 1746 -2598
rect 1740 -2610 1746 -2604
rect 1740 -2616 1746 -2610
rect 1740 -2622 1746 -2616
rect 1740 -2628 1746 -2622
rect 1740 -2634 1746 -2628
rect 1740 -2640 1746 -2634
rect 1740 -2646 1746 -2640
rect 1740 -2652 1746 -2646
rect 1740 -2658 1746 -2652
rect 1740 -2664 1746 -2658
rect 1740 -2742 1746 -2736
rect 1740 -2748 1746 -2742
rect 1740 -2754 1746 -2748
rect 1740 -2760 1746 -2754
rect 1740 -2766 1746 -2760
rect 1740 -2772 1746 -2766
rect 1740 -2778 1746 -2772
rect 1740 -2784 1746 -2778
rect 1740 -2790 1746 -2784
rect 1740 -2796 1746 -2790
rect 1740 -2802 1746 -2796
rect 1740 -2808 1746 -2802
rect 1740 -2814 1746 -2808
rect 1740 -2820 1746 -2814
rect 1740 -2826 1746 -2820
rect 1740 -2832 1746 -2826
rect 1740 -2838 1746 -2832
rect 1740 -2844 1746 -2838
rect 1740 -2850 1746 -2844
rect 1740 -2856 1746 -2850
rect 1740 -2862 1746 -2856
rect 1740 -2868 1746 -2862
rect 1740 -2874 1746 -2868
rect 1740 -2880 1746 -2874
rect 1740 -2886 1746 -2880
rect 1740 -2892 1746 -2886
rect 1740 -2898 1746 -2892
rect 1740 -2904 1746 -2898
rect 1740 -2910 1746 -2904
rect 1740 -2916 1746 -2910
rect 1740 -2922 1746 -2916
rect 1740 -2928 1746 -2922
rect 1740 -2934 1746 -2928
rect 1740 -2940 1746 -2934
rect 1740 -2946 1746 -2940
rect 1740 -2952 1746 -2946
rect 1740 -2958 1746 -2952
rect 1740 -2964 1746 -2958
rect 1740 -2970 1746 -2964
rect 1740 -2976 1746 -2970
rect 1740 -2982 1746 -2976
rect 1740 -2988 1746 -2982
rect 1740 -2994 1746 -2988
rect 1740 -3000 1746 -2994
rect 1740 -3006 1746 -3000
rect 1740 -3012 1746 -3006
rect 1740 -3018 1746 -3012
rect 1740 -3024 1746 -3018
rect 1740 -3030 1746 -3024
rect 1740 -3036 1746 -3030
rect 1740 -3042 1746 -3036
rect 1740 -3048 1746 -3042
rect 1740 -3054 1746 -3048
rect 1740 -3060 1746 -3054
rect 1740 -3066 1746 -3060
rect 1740 -3072 1746 -3066
rect 1740 -3078 1746 -3072
rect 1740 -3084 1746 -3078
rect 1740 -3090 1746 -3084
rect 1740 -3096 1746 -3090
rect 1740 -3102 1746 -3096
rect 1740 -3108 1746 -3102
rect 1740 -3114 1746 -3108
rect 1740 -3120 1746 -3114
rect 1740 -3126 1746 -3120
rect 1740 -3132 1746 -3126
rect 1740 -3138 1746 -3132
rect 1740 -3144 1746 -3138
rect 1740 -3150 1746 -3144
rect 1740 -3156 1746 -3150
rect 1740 -3162 1746 -3156
rect 1740 -3168 1746 -3162
rect 1740 -3174 1746 -3168
rect 1740 -3180 1746 -3174
rect 1740 -3186 1746 -3180
rect 1740 -3192 1746 -3186
rect 1740 -3198 1746 -3192
rect 1740 -3204 1746 -3198
rect 1740 -3258 1746 -3252
rect 1740 -3264 1746 -3258
rect 1740 -3270 1746 -3264
rect 1740 -3276 1746 -3270
rect 1740 -3282 1746 -3276
rect 1740 -3288 1746 -3282
rect 1740 -3294 1746 -3288
rect 1740 -3300 1746 -3294
rect 1740 -3306 1746 -3300
rect 1740 -3312 1746 -3306
rect 1740 -3318 1746 -3312
rect 1740 -3324 1746 -3318
rect 1740 -3330 1746 -3324
rect 1740 -3336 1746 -3330
rect 1740 -3342 1746 -3336
rect 1740 -3348 1746 -3342
rect 1740 -3354 1746 -3348
rect 1740 -3360 1746 -3354
rect 1740 -3366 1746 -3360
rect 1740 -3372 1746 -3366
rect 1740 -3378 1746 -3372
rect 1740 -3384 1746 -3378
rect 1740 -3390 1746 -3384
rect 1740 -3396 1746 -3390
rect 1740 -3402 1746 -3396
rect 1746 -798 1752 -792
rect 1746 -804 1752 -798
rect 1746 -810 1752 -804
rect 1746 -816 1752 -810
rect 1746 -822 1752 -816
rect 1746 -828 1752 -822
rect 1746 -834 1752 -828
rect 1746 -840 1752 -834
rect 1746 -846 1752 -840
rect 1746 -852 1752 -846
rect 1746 -858 1752 -852
rect 1746 -864 1752 -858
rect 1746 -870 1752 -864
rect 1746 -876 1752 -870
rect 1746 -882 1752 -876
rect 1746 -888 1752 -882
rect 1746 -894 1752 -888
rect 1746 -900 1752 -894
rect 1746 -906 1752 -900
rect 1746 -912 1752 -906
rect 1746 -918 1752 -912
rect 1746 -924 1752 -918
rect 1746 -930 1752 -924
rect 1746 -936 1752 -930
rect 1746 -942 1752 -936
rect 1746 -948 1752 -942
rect 1746 -954 1752 -948
rect 1746 -960 1752 -954
rect 1746 -966 1752 -960
rect 1746 -972 1752 -966
rect 1746 -978 1752 -972
rect 1746 -984 1752 -978
rect 1746 -990 1752 -984
rect 1746 -996 1752 -990
rect 1746 -1002 1752 -996
rect 1746 -1008 1752 -1002
rect 1746 -1014 1752 -1008
rect 1746 -1020 1752 -1014
rect 1746 -1026 1752 -1020
rect 1746 -1032 1752 -1026
rect 1746 -1038 1752 -1032
rect 1746 -1044 1752 -1038
rect 1746 -1050 1752 -1044
rect 1746 -1056 1752 -1050
rect 1746 -1062 1752 -1056
rect 1746 -1068 1752 -1062
rect 1746 -1074 1752 -1068
rect 1746 -1080 1752 -1074
rect 1746 -1086 1752 -1080
rect 1746 -1092 1752 -1086
rect 1746 -1098 1752 -1092
rect 1746 -1104 1752 -1098
rect 1746 -1110 1752 -1104
rect 1746 -1116 1752 -1110
rect 1746 -1122 1752 -1116
rect 1746 -1128 1752 -1122
rect 1746 -1134 1752 -1128
rect 1746 -1140 1752 -1134
rect 1746 -1146 1752 -1140
rect 1746 -1152 1752 -1146
rect 1746 -1158 1752 -1152
rect 1746 -1164 1752 -1158
rect 1746 -1170 1752 -1164
rect 1746 -1176 1752 -1170
rect 1746 -1182 1752 -1176
rect 1746 -1188 1752 -1182
rect 1746 -1194 1752 -1188
rect 1746 -1200 1752 -1194
rect 1746 -1206 1752 -1200
rect 1746 -1212 1752 -1206
rect 1746 -1218 1752 -1212
rect 1746 -1224 1752 -1218
rect 1746 -1230 1752 -1224
rect 1746 -1236 1752 -1230
rect 1746 -1242 1752 -1236
rect 1746 -1248 1752 -1242
rect 1746 -1254 1752 -1248
rect 1746 -1260 1752 -1254
rect 1746 -1266 1752 -1260
rect 1746 -1272 1752 -1266
rect 1746 -1278 1752 -1272
rect 1746 -1284 1752 -1278
rect 1746 -1290 1752 -1284
rect 1746 -1296 1752 -1290
rect 1746 -1302 1752 -1296
rect 1746 -1308 1752 -1302
rect 1746 -1314 1752 -1308
rect 1746 -1320 1752 -1314
rect 1746 -1326 1752 -1320
rect 1746 -1332 1752 -1326
rect 1746 -1338 1752 -1332
rect 1746 -1344 1752 -1338
rect 1746 -1350 1752 -1344
rect 1746 -1356 1752 -1350
rect 1746 -1362 1752 -1356
rect 1746 -1368 1752 -1362
rect 1746 -1374 1752 -1368
rect 1746 -1380 1752 -1374
rect 1746 -1386 1752 -1380
rect 1746 -1392 1752 -1386
rect 1746 -1398 1752 -1392
rect 1746 -1404 1752 -1398
rect 1746 -1410 1752 -1404
rect 1746 -1416 1752 -1410
rect 1746 -1422 1752 -1416
rect 1746 -1428 1752 -1422
rect 1746 -1434 1752 -1428
rect 1746 -1440 1752 -1434
rect 1746 -1446 1752 -1440
rect 1746 -1452 1752 -1446
rect 1746 -1458 1752 -1452
rect 1746 -1464 1752 -1458
rect 1746 -1470 1752 -1464
rect 1746 -1476 1752 -1470
rect 1746 -1482 1752 -1476
rect 1746 -1488 1752 -1482
rect 1746 -1494 1752 -1488
rect 1746 -1500 1752 -1494
rect 1746 -1506 1752 -1500
rect 1746 -1512 1752 -1506
rect 1746 -1518 1752 -1512
rect 1746 -1524 1752 -1518
rect 1746 -1530 1752 -1524
rect 1746 -1536 1752 -1530
rect 1746 -1542 1752 -1536
rect 1746 -1548 1752 -1542
rect 1746 -1554 1752 -1548
rect 1746 -1560 1752 -1554
rect 1746 -1566 1752 -1560
rect 1746 -1572 1752 -1566
rect 1746 -1578 1752 -1572
rect 1746 -1584 1752 -1578
rect 1746 -1590 1752 -1584
rect 1746 -1596 1752 -1590
rect 1746 -1602 1752 -1596
rect 1746 -1608 1752 -1602
rect 1746 -1614 1752 -1608
rect 1746 -1620 1752 -1614
rect 1746 -1626 1752 -1620
rect 1746 -1632 1752 -1626
rect 1746 -1638 1752 -1632
rect 1746 -1644 1752 -1638
rect 1746 -1650 1752 -1644
rect 1746 -1656 1752 -1650
rect 1746 -1662 1752 -1656
rect 1746 -1668 1752 -1662
rect 1746 -1674 1752 -1668
rect 1746 -1680 1752 -1674
rect 1746 -1686 1752 -1680
rect 1746 -1692 1752 -1686
rect 1746 -1698 1752 -1692
rect 1746 -1704 1752 -1698
rect 1746 -1710 1752 -1704
rect 1746 -1716 1752 -1710
rect 1746 -1722 1752 -1716
rect 1746 -1728 1752 -1722
rect 1746 -1734 1752 -1728
rect 1746 -1740 1752 -1734
rect 1746 -1746 1752 -1740
rect 1746 -1752 1752 -1746
rect 1746 -1758 1752 -1752
rect 1746 -1764 1752 -1758
rect 1746 -1770 1752 -1764
rect 1746 -1776 1752 -1770
rect 1746 -1782 1752 -1776
rect 1746 -1788 1752 -1782
rect 1746 -1794 1752 -1788
rect 1746 -1800 1752 -1794
rect 1746 -1806 1752 -1800
rect 1746 -1812 1752 -1806
rect 1746 -1818 1752 -1812
rect 1746 -1824 1752 -1818
rect 1746 -1830 1752 -1824
rect 1746 -1836 1752 -1830
rect 1746 -1842 1752 -1836
rect 1746 -1848 1752 -1842
rect 1746 -1854 1752 -1848
rect 1746 -1860 1752 -1854
rect 1746 -1866 1752 -1860
rect 1746 -1872 1752 -1866
rect 1746 -1878 1752 -1872
rect 1746 -1884 1752 -1878
rect 1746 -1890 1752 -1884
rect 1746 -1896 1752 -1890
rect 1746 -1902 1752 -1896
rect 1746 -1908 1752 -1902
rect 1746 -1980 1752 -1974
rect 1746 -1986 1752 -1980
rect 1746 -1992 1752 -1986
rect 1746 -1998 1752 -1992
rect 1746 -2004 1752 -1998
rect 1746 -2010 1752 -2004
rect 1746 -2016 1752 -2010
rect 1746 -2022 1752 -2016
rect 1746 -2028 1752 -2022
rect 1746 -2034 1752 -2028
rect 1746 -2040 1752 -2034
rect 1746 -2046 1752 -2040
rect 1746 -2052 1752 -2046
rect 1746 -2058 1752 -2052
rect 1746 -2064 1752 -2058
rect 1746 -2070 1752 -2064
rect 1746 -2076 1752 -2070
rect 1746 -2082 1752 -2076
rect 1746 -2088 1752 -2082
rect 1746 -2094 1752 -2088
rect 1746 -2100 1752 -2094
rect 1746 -2106 1752 -2100
rect 1746 -2112 1752 -2106
rect 1746 -2118 1752 -2112
rect 1746 -2124 1752 -2118
rect 1746 -2130 1752 -2124
rect 1746 -2136 1752 -2130
rect 1746 -2142 1752 -2136
rect 1746 -2148 1752 -2142
rect 1746 -2154 1752 -2148
rect 1746 -2160 1752 -2154
rect 1746 -2166 1752 -2160
rect 1746 -2172 1752 -2166
rect 1746 -2178 1752 -2172
rect 1746 -2184 1752 -2178
rect 1746 -2190 1752 -2184
rect 1746 -2196 1752 -2190
rect 1746 -2202 1752 -2196
rect 1746 -2208 1752 -2202
rect 1746 -2214 1752 -2208
rect 1746 -2220 1752 -2214
rect 1746 -2226 1752 -2220
rect 1746 -2232 1752 -2226
rect 1746 -2238 1752 -2232
rect 1746 -2244 1752 -2238
rect 1746 -2250 1752 -2244
rect 1746 -2256 1752 -2250
rect 1746 -2262 1752 -2256
rect 1746 -2268 1752 -2262
rect 1746 -2274 1752 -2268
rect 1746 -2280 1752 -2274
rect 1746 -2286 1752 -2280
rect 1746 -2292 1752 -2286
rect 1746 -2298 1752 -2292
rect 1746 -2304 1752 -2298
rect 1746 -2310 1752 -2304
rect 1746 -2316 1752 -2310
rect 1746 -2322 1752 -2316
rect 1746 -2328 1752 -2322
rect 1746 -2334 1752 -2328
rect 1746 -2340 1752 -2334
rect 1746 -2346 1752 -2340
rect 1746 -2352 1752 -2346
rect 1746 -2358 1752 -2352
rect 1746 -2364 1752 -2358
rect 1746 -2370 1752 -2364
rect 1746 -2376 1752 -2370
rect 1746 -2382 1752 -2376
rect 1746 -2388 1752 -2382
rect 1746 -2394 1752 -2388
rect 1746 -2400 1752 -2394
rect 1746 -2406 1752 -2400
rect 1746 -2412 1752 -2406
rect 1746 -2418 1752 -2412
rect 1746 -2424 1752 -2418
rect 1746 -2430 1752 -2424
rect 1746 -2436 1752 -2430
rect 1746 -2442 1752 -2436
rect 1746 -2448 1752 -2442
rect 1746 -2454 1752 -2448
rect 1746 -2460 1752 -2454
rect 1746 -2466 1752 -2460
rect 1746 -2472 1752 -2466
rect 1746 -2478 1752 -2472
rect 1746 -2484 1752 -2478
rect 1746 -2490 1752 -2484
rect 1746 -2496 1752 -2490
rect 1746 -2502 1752 -2496
rect 1746 -2508 1752 -2502
rect 1746 -2514 1752 -2508
rect 1746 -2520 1752 -2514
rect 1746 -2526 1752 -2520
rect 1746 -2532 1752 -2526
rect 1746 -2538 1752 -2532
rect 1746 -2544 1752 -2538
rect 1746 -2550 1752 -2544
rect 1746 -2556 1752 -2550
rect 1746 -2562 1752 -2556
rect 1746 -2568 1752 -2562
rect 1746 -2574 1752 -2568
rect 1746 -2580 1752 -2574
rect 1746 -2586 1752 -2580
rect 1746 -2592 1752 -2586
rect 1746 -2598 1752 -2592
rect 1746 -2604 1752 -2598
rect 1746 -2610 1752 -2604
rect 1746 -2616 1752 -2610
rect 1746 -2622 1752 -2616
rect 1746 -2628 1752 -2622
rect 1746 -2634 1752 -2628
rect 1746 -2640 1752 -2634
rect 1746 -2646 1752 -2640
rect 1746 -2652 1752 -2646
rect 1746 -2658 1752 -2652
rect 1746 -2664 1752 -2658
rect 1746 -2736 1752 -2730
rect 1746 -2742 1752 -2736
rect 1746 -2748 1752 -2742
rect 1746 -2754 1752 -2748
rect 1746 -2760 1752 -2754
rect 1746 -2766 1752 -2760
rect 1746 -2772 1752 -2766
rect 1746 -2778 1752 -2772
rect 1746 -2784 1752 -2778
rect 1746 -2790 1752 -2784
rect 1746 -2796 1752 -2790
rect 1746 -2802 1752 -2796
rect 1746 -2808 1752 -2802
rect 1746 -2814 1752 -2808
rect 1746 -2820 1752 -2814
rect 1746 -2826 1752 -2820
rect 1746 -2832 1752 -2826
rect 1746 -2838 1752 -2832
rect 1746 -2844 1752 -2838
rect 1746 -2850 1752 -2844
rect 1746 -2856 1752 -2850
rect 1746 -2862 1752 -2856
rect 1746 -2868 1752 -2862
rect 1746 -2874 1752 -2868
rect 1746 -2880 1752 -2874
rect 1746 -2886 1752 -2880
rect 1746 -2892 1752 -2886
rect 1746 -2898 1752 -2892
rect 1746 -2904 1752 -2898
rect 1746 -2910 1752 -2904
rect 1746 -2916 1752 -2910
rect 1746 -2922 1752 -2916
rect 1746 -2928 1752 -2922
rect 1746 -2934 1752 -2928
rect 1746 -2940 1752 -2934
rect 1746 -2946 1752 -2940
rect 1746 -2952 1752 -2946
rect 1746 -2958 1752 -2952
rect 1746 -2964 1752 -2958
rect 1746 -2970 1752 -2964
rect 1746 -2976 1752 -2970
rect 1746 -2982 1752 -2976
rect 1746 -2988 1752 -2982
rect 1746 -2994 1752 -2988
rect 1746 -3000 1752 -2994
rect 1746 -3006 1752 -3000
rect 1746 -3012 1752 -3006
rect 1746 -3018 1752 -3012
rect 1746 -3024 1752 -3018
rect 1746 -3030 1752 -3024
rect 1746 -3036 1752 -3030
rect 1746 -3042 1752 -3036
rect 1746 -3048 1752 -3042
rect 1746 -3054 1752 -3048
rect 1746 -3060 1752 -3054
rect 1746 -3066 1752 -3060
rect 1746 -3072 1752 -3066
rect 1746 -3078 1752 -3072
rect 1746 -3084 1752 -3078
rect 1746 -3090 1752 -3084
rect 1746 -3096 1752 -3090
rect 1746 -3102 1752 -3096
rect 1746 -3108 1752 -3102
rect 1746 -3114 1752 -3108
rect 1746 -3120 1752 -3114
rect 1746 -3126 1752 -3120
rect 1746 -3132 1752 -3126
rect 1746 -3138 1752 -3132
rect 1746 -3144 1752 -3138
rect 1746 -3150 1752 -3144
rect 1746 -3156 1752 -3150
rect 1746 -3162 1752 -3156
rect 1746 -3168 1752 -3162
rect 1746 -3174 1752 -3168
rect 1746 -3180 1752 -3174
rect 1746 -3186 1752 -3180
rect 1746 -3192 1752 -3186
rect 1746 -3198 1752 -3192
rect 1746 -3204 1752 -3198
rect 1746 -3252 1752 -3246
rect 1746 -3258 1752 -3252
rect 1746 -3264 1752 -3258
rect 1746 -3270 1752 -3264
rect 1746 -3276 1752 -3270
rect 1746 -3282 1752 -3276
rect 1746 -3288 1752 -3282
rect 1746 -3294 1752 -3288
rect 1746 -3300 1752 -3294
rect 1746 -3306 1752 -3300
rect 1746 -3312 1752 -3306
rect 1746 -3318 1752 -3312
rect 1746 -3324 1752 -3318
rect 1746 -3330 1752 -3324
rect 1746 -3336 1752 -3330
rect 1746 -3342 1752 -3336
rect 1746 -3348 1752 -3342
rect 1746 -3354 1752 -3348
rect 1746 -3360 1752 -3354
rect 1746 -3366 1752 -3360
rect 1746 -3372 1752 -3366
rect 1746 -3378 1752 -3372
rect 1746 -3384 1752 -3378
rect 1746 -3390 1752 -3384
rect 1746 -3396 1752 -3390
rect 1752 -786 1758 -780
rect 1752 -792 1758 -786
rect 1752 -798 1758 -792
rect 1752 -804 1758 -798
rect 1752 -810 1758 -804
rect 1752 -816 1758 -810
rect 1752 -822 1758 -816
rect 1752 -828 1758 -822
rect 1752 -834 1758 -828
rect 1752 -840 1758 -834
rect 1752 -846 1758 -840
rect 1752 -852 1758 -846
rect 1752 -858 1758 -852
rect 1752 -864 1758 -858
rect 1752 -870 1758 -864
rect 1752 -876 1758 -870
rect 1752 -882 1758 -876
rect 1752 -888 1758 -882
rect 1752 -894 1758 -888
rect 1752 -900 1758 -894
rect 1752 -906 1758 -900
rect 1752 -912 1758 -906
rect 1752 -918 1758 -912
rect 1752 -924 1758 -918
rect 1752 -930 1758 -924
rect 1752 -936 1758 -930
rect 1752 -942 1758 -936
rect 1752 -948 1758 -942
rect 1752 -954 1758 -948
rect 1752 -960 1758 -954
rect 1752 -966 1758 -960
rect 1752 -972 1758 -966
rect 1752 -978 1758 -972
rect 1752 -984 1758 -978
rect 1752 -990 1758 -984
rect 1752 -996 1758 -990
rect 1752 -1002 1758 -996
rect 1752 -1008 1758 -1002
rect 1752 -1014 1758 -1008
rect 1752 -1020 1758 -1014
rect 1752 -1026 1758 -1020
rect 1752 -1032 1758 -1026
rect 1752 -1038 1758 -1032
rect 1752 -1044 1758 -1038
rect 1752 -1050 1758 -1044
rect 1752 -1056 1758 -1050
rect 1752 -1062 1758 -1056
rect 1752 -1068 1758 -1062
rect 1752 -1074 1758 -1068
rect 1752 -1080 1758 -1074
rect 1752 -1086 1758 -1080
rect 1752 -1092 1758 -1086
rect 1752 -1098 1758 -1092
rect 1752 -1104 1758 -1098
rect 1752 -1110 1758 -1104
rect 1752 -1116 1758 -1110
rect 1752 -1122 1758 -1116
rect 1752 -1128 1758 -1122
rect 1752 -1134 1758 -1128
rect 1752 -1140 1758 -1134
rect 1752 -1146 1758 -1140
rect 1752 -1152 1758 -1146
rect 1752 -1158 1758 -1152
rect 1752 -1164 1758 -1158
rect 1752 -1170 1758 -1164
rect 1752 -1176 1758 -1170
rect 1752 -1182 1758 -1176
rect 1752 -1188 1758 -1182
rect 1752 -1194 1758 -1188
rect 1752 -1200 1758 -1194
rect 1752 -1206 1758 -1200
rect 1752 -1212 1758 -1206
rect 1752 -1218 1758 -1212
rect 1752 -1224 1758 -1218
rect 1752 -1230 1758 -1224
rect 1752 -1236 1758 -1230
rect 1752 -1242 1758 -1236
rect 1752 -1248 1758 -1242
rect 1752 -1254 1758 -1248
rect 1752 -1260 1758 -1254
rect 1752 -1266 1758 -1260
rect 1752 -1272 1758 -1266
rect 1752 -1278 1758 -1272
rect 1752 -1284 1758 -1278
rect 1752 -1290 1758 -1284
rect 1752 -1296 1758 -1290
rect 1752 -1302 1758 -1296
rect 1752 -1308 1758 -1302
rect 1752 -1314 1758 -1308
rect 1752 -1320 1758 -1314
rect 1752 -1326 1758 -1320
rect 1752 -1332 1758 -1326
rect 1752 -1338 1758 -1332
rect 1752 -1344 1758 -1338
rect 1752 -1350 1758 -1344
rect 1752 -1356 1758 -1350
rect 1752 -1362 1758 -1356
rect 1752 -1368 1758 -1362
rect 1752 -1374 1758 -1368
rect 1752 -1380 1758 -1374
rect 1752 -1386 1758 -1380
rect 1752 -1392 1758 -1386
rect 1752 -1398 1758 -1392
rect 1752 -1404 1758 -1398
rect 1752 -1410 1758 -1404
rect 1752 -1416 1758 -1410
rect 1752 -1422 1758 -1416
rect 1752 -1428 1758 -1422
rect 1752 -1434 1758 -1428
rect 1752 -1440 1758 -1434
rect 1752 -1446 1758 -1440
rect 1752 -1452 1758 -1446
rect 1752 -1458 1758 -1452
rect 1752 -1464 1758 -1458
rect 1752 -1470 1758 -1464
rect 1752 -1476 1758 -1470
rect 1752 -1482 1758 -1476
rect 1752 -1488 1758 -1482
rect 1752 -1494 1758 -1488
rect 1752 -1500 1758 -1494
rect 1752 -1506 1758 -1500
rect 1752 -1512 1758 -1506
rect 1752 -1518 1758 -1512
rect 1752 -1524 1758 -1518
rect 1752 -1530 1758 -1524
rect 1752 -1536 1758 -1530
rect 1752 -1542 1758 -1536
rect 1752 -1548 1758 -1542
rect 1752 -1554 1758 -1548
rect 1752 -1560 1758 -1554
rect 1752 -1566 1758 -1560
rect 1752 -1572 1758 -1566
rect 1752 -1578 1758 -1572
rect 1752 -1584 1758 -1578
rect 1752 -1590 1758 -1584
rect 1752 -1596 1758 -1590
rect 1752 -1602 1758 -1596
rect 1752 -1608 1758 -1602
rect 1752 -1614 1758 -1608
rect 1752 -1620 1758 -1614
rect 1752 -1626 1758 -1620
rect 1752 -1632 1758 -1626
rect 1752 -1638 1758 -1632
rect 1752 -1644 1758 -1638
rect 1752 -1650 1758 -1644
rect 1752 -1656 1758 -1650
rect 1752 -1662 1758 -1656
rect 1752 -1668 1758 -1662
rect 1752 -1674 1758 -1668
rect 1752 -1680 1758 -1674
rect 1752 -1686 1758 -1680
rect 1752 -1692 1758 -1686
rect 1752 -1698 1758 -1692
rect 1752 -1704 1758 -1698
rect 1752 -1710 1758 -1704
rect 1752 -1716 1758 -1710
rect 1752 -1722 1758 -1716
rect 1752 -1728 1758 -1722
rect 1752 -1734 1758 -1728
rect 1752 -1740 1758 -1734
rect 1752 -1746 1758 -1740
rect 1752 -1752 1758 -1746
rect 1752 -1758 1758 -1752
rect 1752 -1764 1758 -1758
rect 1752 -1770 1758 -1764
rect 1752 -1776 1758 -1770
rect 1752 -1782 1758 -1776
rect 1752 -1788 1758 -1782
rect 1752 -1794 1758 -1788
rect 1752 -1800 1758 -1794
rect 1752 -1806 1758 -1800
rect 1752 -1812 1758 -1806
rect 1752 -1818 1758 -1812
rect 1752 -1824 1758 -1818
rect 1752 -1830 1758 -1824
rect 1752 -1836 1758 -1830
rect 1752 -1842 1758 -1836
rect 1752 -1848 1758 -1842
rect 1752 -1854 1758 -1848
rect 1752 -1860 1758 -1854
rect 1752 -1866 1758 -1860
rect 1752 -1872 1758 -1866
rect 1752 -1878 1758 -1872
rect 1752 -1884 1758 -1878
rect 1752 -1890 1758 -1884
rect 1752 -1896 1758 -1890
rect 1752 -1974 1758 -1968
rect 1752 -1980 1758 -1974
rect 1752 -1986 1758 -1980
rect 1752 -1992 1758 -1986
rect 1752 -1998 1758 -1992
rect 1752 -2004 1758 -1998
rect 1752 -2010 1758 -2004
rect 1752 -2016 1758 -2010
rect 1752 -2022 1758 -2016
rect 1752 -2028 1758 -2022
rect 1752 -2034 1758 -2028
rect 1752 -2040 1758 -2034
rect 1752 -2046 1758 -2040
rect 1752 -2052 1758 -2046
rect 1752 -2058 1758 -2052
rect 1752 -2064 1758 -2058
rect 1752 -2070 1758 -2064
rect 1752 -2076 1758 -2070
rect 1752 -2082 1758 -2076
rect 1752 -2088 1758 -2082
rect 1752 -2094 1758 -2088
rect 1752 -2100 1758 -2094
rect 1752 -2106 1758 -2100
rect 1752 -2112 1758 -2106
rect 1752 -2118 1758 -2112
rect 1752 -2124 1758 -2118
rect 1752 -2130 1758 -2124
rect 1752 -2136 1758 -2130
rect 1752 -2142 1758 -2136
rect 1752 -2148 1758 -2142
rect 1752 -2154 1758 -2148
rect 1752 -2160 1758 -2154
rect 1752 -2166 1758 -2160
rect 1752 -2172 1758 -2166
rect 1752 -2178 1758 -2172
rect 1752 -2184 1758 -2178
rect 1752 -2190 1758 -2184
rect 1752 -2196 1758 -2190
rect 1752 -2202 1758 -2196
rect 1752 -2208 1758 -2202
rect 1752 -2214 1758 -2208
rect 1752 -2220 1758 -2214
rect 1752 -2226 1758 -2220
rect 1752 -2232 1758 -2226
rect 1752 -2238 1758 -2232
rect 1752 -2244 1758 -2238
rect 1752 -2250 1758 -2244
rect 1752 -2256 1758 -2250
rect 1752 -2262 1758 -2256
rect 1752 -2268 1758 -2262
rect 1752 -2274 1758 -2268
rect 1752 -2280 1758 -2274
rect 1752 -2286 1758 -2280
rect 1752 -2292 1758 -2286
rect 1752 -2298 1758 -2292
rect 1752 -2304 1758 -2298
rect 1752 -2310 1758 -2304
rect 1752 -2316 1758 -2310
rect 1752 -2322 1758 -2316
rect 1752 -2328 1758 -2322
rect 1752 -2334 1758 -2328
rect 1752 -2340 1758 -2334
rect 1752 -2346 1758 -2340
rect 1752 -2352 1758 -2346
rect 1752 -2358 1758 -2352
rect 1752 -2364 1758 -2358
rect 1752 -2370 1758 -2364
rect 1752 -2376 1758 -2370
rect 1752 -2382 1758 -2376
rect 1752 -2388 1758 -2382
rect 1752 -2394 1758 -2388
rect 1752 -2400 1758 -2394
rect 1752 -2406 1758 -2400
rect 1752 -2412 1758 -2406
rect 1752 -2418 1758 -2412
rect 1752 -2424 1758 -2418
rect 1752 -2430 1758 -2424
rect 1752 -2436 1758 -2430
rect 1752 -2442 1758 -2436
rect 1752 -2448 1758 -2442
rect 1752 -2454 1758 -2448
rect 1752 -2460 1758 -2454
rect 1752 -2466 1758 -2460
rect 1752 -2472 1758 -2466
rect 1752 -2478 1758 -2472
rect 1752 -2484 1758 -2478
rect 1752 -2490 1758 -2484
rect 1752 -2496 1758 -2490
rect 1752 -2502 1758 -2496
rect 1752 -2508 1758 -2502
rect 1752 -2514 1758 -2508
rect 1752 -2520 1758 -2514
rect 1752 -2526 1758 -2520
rect 1752 -2532 1758 -2526
rect 1752 -2538 1758 -2532
rect 1752 -2544 1758 -2538
rect 1752 -2550 1758 -2544
rect 1752 -2556 1758 -2550
rect 1752 -2562 1758 -2556
rect 1752 -2568 1758 -2562
rect 1752 -2574 1758 -2568
rect 1752 -2580 1758 -2574
rect 1752 -2586 1758 -2580
rect 1752 -2592 1758 -2586
rect 1752 -2598 1758 -2592
rect 1752 -2604 1758 -2598
rect 1752 -2610 1758 -2604
rect 1752 -2616 1758 -2610
rect 1752 -2622 1758 -2616
rect 1752 -2628 1758 -2622
rect 1752 -2634 1758 -2628
rect 1752 -2640 1758 -2634
rect 1752 -2646 1758 -2640
rect 1752 -2652 1758 -2646
rect 1752 -2658 1758 -2652
rect 1752 -2736 1758 -2730
rect 1752 -2742 1758 -2736
rect 1752 -2748 1758 -2742
rect 1752 -2754 1758 -2748
rect 1752 -2760 1758 -2754
rect 1752 -2766 1758 -2760
rect 1752 -2772 1758 -2766
rect 1752 -2778 1758 -2772
rect 1752 -2784 1758 -2778
rect 1752 -2790 1758 -2784
rect 1752 -2796 1758 -2790
rect 1752 -2802 1758 -2796
rect 1752 -2808 1758 -2802
rect 1752 -2814 1758 -2808
rect 1752 -2820 1758 -2814
rect 1752 -2826 1758 -2820
rect 1752 -2832 1758 -2826
rect 1752 -2838 1758 -2832
rect 1752 -2844 1758 -2838
rect 1752 -2850 1758 -2844
rect 1752 -2856 1758 -2850
rect 1752 -2862 1758 -2856
rect 1752 -2868 1758 -2862
rect 1752 -2874 1758 -2868
rect 1752 -2880 1758 -2874
rect 1752 -2886 1758 -2880
rect 1752 -2892 1758 -2886
rect 1752 -2898 1758 -2892
rect 1752 -2904 1758 -2898
rect 1752 -2910 1758 -2904
rect 1752 -2916 1758 -2910
rect 1752 -2922 1758 -2916
rect 1752 -2928 1758 -2922
rect 1752 -2934 1758 -2928
rect 1752 -2940 1758 -2934
rect 1752 -2946 1758 -2940
rect 1752 -2952 1758 -2946
rect 1752 -2958 1758 -2952
rect 1752 -2964 1758 -2958
rect 1752 -2970 1758 -2964
rect 1752 -2976 1758 -2970
rect 1752 -2982 1758 -2976
rect 1752 -2988 1758 -2982
rect 1752 -2994 1758 -2988
rect 1752 -3000 1758 -2994
rect 1752 -3006 1758 -3000
rect 1752 -3012 1758 -3006
rect 1752 -3018 1758 -3012
rect 1752 -3024 1758 -3018
rect 1752 -3030 1758 -3024
rect 1752 -3036 1758 -3030
rect 1752 -3042 1758 -3036
rect 1752 -3048 1758 -3042
rect 1752 -3054 1758 -3048
rect 1752 -3060 1758 -3054
rect 1752 -3066 1758 -3060
rect 1752 -3072 1758 -3066
rect 1752 -3078 1758 -3072
rect 1752 -3084 1758 -3078
rect 1752 -3090 1758 -3084
rect 1752 -3096 1758 -3090
rect 1752 -3102 1758 -3096
rect 1752 -3108 1758 -3102
rect 1752 -3114 1758 -3108
rect 1752 -3120 1758 -3114
rect 1752 -3126 1758 -3120
rect 1752 -3132 1758 -3126
rect 1752 -3138 1758 -3132
rect 1752 -3144 1758 -3138
rect 1752 -3150 1758 -3144
rect 1752 -3156 1758 -3150
rect 1752 -3162 1758 -3156
rect 1752 -3168 1758 -3162
rect 1752 -3174 1758 -3168
rect 1752 -3180 1758 -3174
rect 1752 -3186 1758 -3180
rect 1752 -3192 1758 -3186
rect 1752 -3198 1758 -3192
rect 1752 -3204 1758 -3198
rect 1752 -3252 1758 -3246
rect 1752 -3258 1758 -3252
rect 1752 -3264 1758 -3258
rect 1752 -3270 1758 -3264
rect 1752 -3276 1758 -3270
rect 1752 -3282 1758 -3276
rect 1752 -3288 1758 -3282
rect 1752 -3294 1758 -3288
rect 1752 -3300 1758 -3294
rect 1752 -3306 1758 -3300
rect 1752 -3312 1758 -3306
rect 1752 -3318 1758 -3312
rect 1752 -3324 1758 -3318
rect 1752 -3330 1758 -3324
rect 1752 -3336 1758 -3330
rect 1752 -3342 1758 -3336
rect 1752 -3348 1758 -3342
rect 1752 -3354 1758 -3348
rect 1752 -3360 1758 -3354
rect 1752 -3366 1758 -3360
rect 1752 -3372 1758 -3366
rect 1752 -3378 1758 -3372
rect 1752 -3384 1758 -3378
rect 1752 -3390 1758 -3384
rect 1752 -3396 1758 -3390
rect 1758 -780 1764 -774
rect 1758 -786 1764 -780
rect 1758 -792 1764 -786
rect 1758 -798 1764 -792
rect 1758 -804 1764 -798
rect 1758 -810 1764 -804
rect 1758 -816 1764 -810
rect 1758 -822 1764 -816
rect 1758 -828 1764 -822
rect 1758 -834 1764 -828
rect 1758 -840 1764 -834
rect 1758 -846 1764 -840
rect 1758 -852 1764 -846
rect 1758 -858 1764 -852
rect 1758 -864 1764 -858
rect 1758 -870 1764 -864
rect 1758 -876 1764 -870
rect 1758 -882 1764 -876
rect 1758 -888 1764 -882
rect 1758 -894 1764 -888
rect 1758 -900 1764 -894
rect 1758 -906 1764 -900
rect 1758 -912 1764 -906
rect 1758 -918 1764 -912
rect 1758 -924 1764 -918
rect 1758 -930 1764 -924
rect 1758 -936 1764 -930
rect 1758 -942 1764 -936
rect 1758 -948 1764 -942
rect 1758 -954 1764 -948
rect 1758 -960 1764 -954
rect 1758 -966 1764 -960
rect 1758 -972 1764 -966
rect 1758 -978 1764 -972
rect 1758 -984 1764 -978
rect 1758 -990 1764 -984
rect 1758 -996 1764 -990
rect 1758 -1002 1764 -996
rect 1758 -1008 1764 -1002
rect 1758 -1014 1764 -1008
rect 1758 -1020 1764 -1014
rect 1758 -1026 1764 -1020
rect 1758 -1032 1764 -1026
rect 1758 -1038 1764 -1032
rect 1758 -1044 1764 -1038
rect 1758 -1050 1764 -1044
rect 1758 -1056 1764 -1050
rect 1758 -1062 1764 -1056
rect 1758 -1068 1764 -1062
rect 1758 -1074 1764 -1068
rect 1758 -1080 1764 -1074
rect 1758 -1086 1764 -1080
rect 1758 -1092 1764 -1086
rect 1758 -1098 1764 -1092
rect 1758 -1104 1764 -1098
rect 1758 -1110 1764 -1104
rect 1758 -1116 1764 -1110
rect 1758 -1122 1764 -1116
rect 1758 -1128 1764 -1122
rect 1758 -1134 1764 -1128
rect 1758 -1140 1764 -1134
rect 1758 -1146 1764 -1140
rect 1758 -1152 1764 -1146
rect 1758 -1158 1764 -1152
rect 1758 -1164 1764 -1158
rect 1758 -1170 1764 -1164
rect 1758 -1176 1764 -1170
rect 1758 -1182 1764 -1176
rect 1758 -1188 1764 -1182
rect 1758 -1194 1764 -1188
rect 1758 -1200 1764 -1194
rect 1758 -1206 1764 -1200
rect 1758 -1212 1764 -1206
rect 1758 -1218 1764 -1212
rect 1758 -1224 1764 -1218
rect 1758 -1230 1764 -1224
rect 1758 -1236 1764 -1230
rect 1758 -1242 1764 -1236
rect 1758 -1248 1764 -1242
rect 1758 -1254 1764 -1248
rect 1758 -1260 1764 -1254
rect 1758 -1266 1764 -1260
rect 1758 -1272 1764 -1266
rect 1758 -1278 1764 -1272
rect 1758 -1284 1764 -1278
rect 1758 -1290 1764 -1284
rect 1758 -1296 1764 -1290
rect 1758 -1302 1764 -1296
rect 1758 -1308 1764 -1302
rect 1758 -1314 1764 -1308
rect 1758 -1320 1764 -1314
rect 1758 -1326 1764 -1320
rect 1758 -1332 1764 -1326
rect 1758 -1338 1764 -1332
rect 1758 -1344 1764 -1338
rect 1758 -1350 1764 -1344
rect 1758 -1356 1764 -1350
rect 1758 -1362 1764 -1356
rect 1758 -1368 1764 -1362
rect 1758 -1374 1764 -1368
rect 1758 -1380 1764 -1374
rect 1758 -1386 1764 -1380
rect 1758 -1392 1764 -1386
rect 1758 -1398 1764 -1392
rect 1758 -1404 1764 -1398
rect 1758 -1410 1764 -1404
rect 1758 -1416 1764 -1410
rect 1758 -1422 1764 -1416
rect 1758 -1428 1764 -1422
rect 1758 -1434 1764 -1428
rect 1758 -1440 1764 -1434
rect 1758 -1446 1764 -1440
rect 1758 -1452 1764 -1446
rect 1758 -1458 1764 -1452
rect 1758 -1464 1764 -1458
rect 1758 -1470 1764 -1464
rect 1758 -1476 1764 -1470
rect 1758 -1482 1764 -1476
rect 1758 -1488 1764 -1482
rect 1758 -1494 1764 -1488
rect 1758 -1500 1764 -1494
rect 1758 -1506 1764 -1500
rect 1758 -1512 1764 -1506
rect 1758 -1518 1764 -1512
rect 1758 -1524 1764 -1518
rect 1758 -1530 1764 -1524
rect 1758 -1536 1764 -1530
rect 1758 -1542 1764 -1536
rect 1758 -1548 1764 -1542
rect 1758 -1554 1764 -1548
rect 1758 -1560 1764 -1554
rect 1758 -1566 1764 -1560
rect 1758 -1572 1764 -1566
rect 1758 -1578 1764 -1572
rect 1758 -1584 1764 -1578
rect 1758 -1590 1764 -1584
rect 1758 -1596 1764 -1590
rect 1758 -1602 1764 -1596
rect 1758 -1608 1764 -1602
rect 1758 -1614 1764 -1608
rect 1758 -1620 1764 -1614
rect 1758 -1626 1764 -1620
rect 1758 -1632 1764 -1626
rect 1758 -1638 1764 -1632
rect 1758 -1644 1764 -1638
rect 1758 -1650 1764 -1644
rect 1758 -1656 1764 -1650
rect 1758 -1662 1764 -1656
rect 1758 -1668 1764 -1662
rect 1758 -1674 1764 -1668
rect 1758 -1680 1764 -1674
rect 1758 -1686 1764 -1680
rect 1758 -1692 1764 -1686
rect 1758 -1698 1764 -1692
rect 1758 -1704 1764 -1698
rect 1758 -1710 1764 -1704
rect 1758 -1716 1764 -1710
rect 1758 -1722 1764 -1716
rect 1758 -1728 1764 -1722
rect 1758 -1734 1764 -1728
rect 1758 -1740 1764 -1734
rect 1758 -1746 1764 -1740
rect 1758 -1752 1764 -1746
rect 1758 -1758 1764 -1752
rect 1758 -1764 1764 -1758
rect 1758 -1770 1764 -1764
rect 1758 -1776 1764 -1770
rect 1758 -1782 1764 -1776
rect 1758 -1788 1764 -1782
rect 1758 -1794 1764 -1788
rect 1758 -1800 1764 -1794
rect 1758 -1806 1764 -1800
rect 1758 -1812 1764 -1806
rect 1758 -1818 1764 -1812
rect 1758 -1824 1764 -1818
rect 1758 -1830 1764 -1824
rect 1758 -1836 1764 -1830
rect 1758 -1842 1764 -1836
rect 1758 -1848 1764 -1842
rect 1758 -1854 1764 -1848
rect 1758 -1860 1764 -1854
rect 1758 -1866 1764 -1860
rect 1758 -1872 1764 -1866
rect 1758 -1878 1764 -1872
rect 1758 -1884 1764 -1878
rect 1758 -1890 1764 -1884
rect 1758 -1968 1764 -1962
rect 1758 -1974 1764 -1968
rect 1758 -1980 1764 -1974
rect 1758 -1986 1764 -1980
rect 1758 -1992 1764 -1986
rect 1758 -1998 1764 -1992
rect 1758 -2004 1764 -1998
rect 1758 -2010 1764 -2004
rect 1758 -2016 1764 -2010
rect 1758 -2022 1764 -2016
rect 1758 -2028 1764 -2022
rect 1758 -2034 1764 -2028
rect 1758 -2040 1764 -2034
rect 1758 -2046 1764 -2040
rect 1758 -2052 1764 -2046
rect 1758 -2058 1764 -2052
rect 1758 -2064 1764 -2058
rect 1758 -2070 1764 -2064
rect 1758 -2076 1764 -2070
rect 1758 -2082 1764 -2076
rect 1758 -2088 1764 -2082
rect 1758 -2094 1764 -2088
rect 1758 -2100 1764 -2094
rect 1758 -2106 1764 -2100
rect 1758 -2112 1764 -2106
rect 1758 -2118 1764 -2112
rect 1758 -2124 1764 -2118
rect 1758 -2130 1764 -2124
rect 1758 -2136 1764 -2130
rect 1758 -2142 1764 -2136
rect 1758 -2148 1764 -2142
rect 1758 -2154 1764 -2148
rect 1758 -2160 1764 -2154
rect 1758 -2166 1764 -2160
rect 1758 -2172 1764 -2166
rect 1758 -2178 1764 -2172
rect 1758 -2184 1764 -2178
rect 1758 -2190 1764 -2184
rect 1758 -2196 1764 -2190
rect 1758 -2202 1764 -2196
rect 1758 -2208 1764 -2202
rect 1758 -2214 1764 -2208
rect 1758 -2220 1764 -2214
rect 1758 -2226 1764 -2220
rect 1758 -2232 1764 -2226
rect 1758 -2238 1764 -2232
rect 1758 -2244 1764 -2238
rect 1758 -2250 1764 -2244
rect 1758 -2256 1764 -2250
rect 1758 -2262 1764 -2256
rect 1758 -2268 1764 -2262
rect 1758 -2274 1764 -2268
rect 1758 -2280 1764 -2274
rect 1758 -2286 1764 -2280
rect 1758 -2292 1764 -2286
rect 1758 -2298 1764 -2292
rect 1758 -2304 1764 -2298
rect 1758 -2310 1764 -2304
rect 1758 -2316 1764 -2310
rect 1758 -2322 1764 -2316
rect 1758 -2328 1764 -2322
rect 1758 -2334 1764 -2328
rect 1758 -2340 1764 -2334
rect 1758 -2346 1764 -2340
rect 1758 -2352 1764 -2346
rect 1758 -2358 1764 -2352
rect 1758 -2364 1764 -2358
rect 1758 -2370 1764 -2364
rect 1758 -2376 1764 -2370
rect 1758 -2382 1764 -2376
rect 1758 -2388 1764 -2382
rect 1758 -2394 1764 -2388
rect 1758 -2400 1764 -2394
rect 1758 -2406 1764 -2400
rect 1758 -2412 1764 -2406
rect 1758 -2418 1764 -2412
rect 1758 -2424 1764 -2418
rect 1758 -2430 1764 -2424
rect 1758 -2436 1764 -2430
rect 1758 -2442 1764 -2436
rect 1758 -2448 1764 -2442
rect 1758 -2454 1764 -2448
rect 1758 -2460 1764 -2454
rect 1758 -2466 1764 -2460
rect 1758 -2472 1764 -2466
rect 1758 -2478 1764 -2472
rect 1758 -2484 1764 -2478
rect 1758 -2490 1764 -2484
rect 1758 -2496 1764 -2490
rect 1758 -2502 1764 -2496
rect 1758 -2508 1764 -2502
rect 1758 -2514 1764 -2508
rect 1758 -2520 1764 -2514
rect 1758 -2526 1764 -2520
rect 1758 -2532 1764 -2526
rect 1758 -2538 1764 -2532
rect 1758 -2544 1764 -2538
rect 1758 -2550 1764 -2544
rect 1758 -2556 1764 -2550
rect 1758 -2562 1764 -2556
rect 1758 -2568 1764 -2562
rect 1758 -2574 1764 -2568
rect 1758 -2580 1764 -2574
rect 1758 -2586 1764 -2580
rect 1758 -2592 1764 -2586
rect 1758 -2598 1764 -2592
rect 1758 -2604 1764 -2598
rect 1758 -2610 1764 -2604
rect 1758 -2616 1764 -2610
rect 1758 -2622 1764 -2616
rect 1758 -2628 1764 -2622
rect 1758 -2634 1764 -2628
rect 1758 -2640 1764 -2634
rect 1758 -2646 1764 -2640
rect 1758 -2652 1764 -2646
rect 1758 -2658 1764 -2652
rect 1758 -2730 1764 -2724
rect 1758 -2736 1764 -2730
rect 1758 -2742 1764 -2736
rect 1758 -2748 1764 -2742
rect 1758 -2754 1764 -2748
rect 1758 -2760 1764 -2754
rect 1758 -2766 1764 -2760
rect 1758 -2772 1764 -2766
rect 1758 -2778 1764 -2772
rect 1758 -2784 1764 -2778
rect 1758 -2790 1764 -2784
rect 1758 -2796 1764 -2790
rect 1758 -2802 1764 -2796
rect 1758 -2808 1764 -2802
rect 1758 -2814 1764 -2808
rect 1758 -2820 1764 -2814
rect 1758 -2826 1764 -2820
rect 1758 -2832 1764 -2826
rect 1758 -2838 1764 -2832
rect 1758 -2844 1764 -2838
rect 1758 -2850 1764 -2844
rect 1758 -2856 1764 -2850
rect 1758 -2862 1764 -2856
rect 1758 -2868 1764 -2862
rect 1758 -2874 1764 -2868
rect 1758 -2880 1764 -2874
rect 1758 -2886 1764 -2880
rect 1758 -2892 1764 -2886
rect 1758 -2898 1764 -2892
rect 1758 -2904 1764 -2898
rect 1758 -2910 1764 -2904
rect 1758 -2916 1764 -2910
rect 1758 -2922 1764 -2916
rect 1758 -2928 1764 -2922
rect 1758 -2934 1764 -2928
rect 1758 -2940 1764 -2934
rect 1758 -2946 1764 -2940
rect 1758 -2952 1764 -2946
rect 1758 -2958 1764 -2952
rect 1758 -2964 1764 -2958
rect 1758 -2970 1764 -2964
rect 1758 -2976 1764 -2970
rect 1758 -2982 1764 -2976
rect 1758 -2988 1764 -2982
rect 1758 -2994 1764 -2988
rect 1758 -3000 1764 -2994
rect 1758 -3006 1764 -3000
rect 1758 -3012 1764 -3006
rect 1758 -3018 1764 -3012
rect 1758 -3024 1764 -3018
rect 1758 -3030 1764 -3024
rect 1758 -3036 1764 -3030
rect 1758 -3042 1764 -3036
rect 1758 -3048 1764 -3042
rect 1758 -3054 1764 -3048
rect 1758 -3060 1764 -3054
rect 1758 -3066 1764 -3060
rect 1758 -3072 1764 -3066
rect 1758 -3078 1764 -3072
rect 1758 -3084 1764 -3078
rect 1758 -3090 1764 -3084
rect 1758 -3096 1764 -3090
rect 1758 -3102 1764 -3096
rect 1758 -3108 1764 -3102
rect 1758 -3114 1764 -3108
rect 1758 -3120 1764 -3114
rect 1758 -3126 1764 -3120
rect 1758 -3132 1764 -3126
rect 1758 -3138 1764 -3132
rect 1758 -3144 1764 -3138
rect 1758 -3150 1764 -3144
rect 1758 -3156 1764 -3150
rect 1758 -3162 1764 -3156
rect 1758 -3168 1764 -3162
rect 1758 -3174 1764 -3168
rect 1758 -3180 1764 -3174
rect 1758 -3186 1764 -3180
rect 1758 -3192 1764 -3186
rect 1758 -3198 1764 -3192
rect 1758 -3252 1764 -3246
rect 1758 -3258 1764 -3252
rect 1758 -3264 1764 -3258
rect 1758 -3270 1764 -3264
rect 1758 -3276 1764 -3270
rect 1758 -3282 1764 -3276
rect 1758 -3288 1764 -3282
rect 1758 -3294 1764 -3288
rect 1758 -3300 1764 -3294
rect 1758 -3306 1764 -3300
rect 1758 -3312 1764 -3306
rect 1758 -3318 1764 -3312
rect 1758 -3324 1764 -3318
rect 1758 -3330 1764 -3324
rect 1758 -3336 1764 -3330
rect 1758 -3342 1764 -3336
rect 1758 -3348 1764 -3342
rect 1758 -3354 1764 -3348
rect 1758 -3360 1764 -3354
rect 1758 -3366 1764 -3360
rect 1758 -3372 1764 -3366
rect 1758 -3378 1764 -3372
rect 1758 -3384 1764 -3378
rect 1758 -3390 1764 -3384
rect 1764 -768 1770 -762
rect 1764 -774 1770 -768
rect 1764 -780 1770 -774
rect 1764 -786 1770 -780
rect 1764 -792 1770 -786
rect 1764 -798 1770 -792
rect 1764 -804 1770 -798
rect 1764 -810 1770 -804
rect 1764 -816 1770 -810
rect 1764 -822 1770 -816
rect 1764 -828 1770 -822
rect 1764 -834 1770 -828
rect 1764 -840 1770 -834
rect 1764 -846 1770 -840
rect 1764 -852 1770 -846
rect 1764 -858 1770 -852
rect 1764 -864 1770 -858
rect 1764 -870 1770 -864
rect 1764 -876 1770 -870
rect 1764 -882 1770 -876
rect 1764 -888 1770 -882
rect 1764 -894 1770 -888
rect 1764 -900 1770 -894
rect 1764 -906 1770 -900
rect 1764 -912 1770 -906
rect 1764 -918 1770 -912
rect 1764 -924 1770 -918
rect 1764 -930 1770 -924
rect 1764 -936 1770 -930
rect 1764 -942 1770 -936
rect 1764 -948 1770 -942
rect 1764 -954 1770 -948
rect 1764 -960 1770 -954
rect 1764 -966 1770 -960
rect 1764 -972 1770 -966
rect 1764 -978 1770 -972
rect 1764 -984 1770 -978
rect 1764 -990 1770 -984
rect 1764 -996 1770 -990
rect 1764 -1002 1770 -996
rect 1764 -1008 1770 -1002
rect 1764 -1014 1770 -1008
rect 1764 -1020 1770 -1014
rect 1764 -1026 1770 -1020
rect 1764 -1032 1770 -1026
rect 1764 -1038 1770 -1032
rect 1764 -1044 1770 -1038
rect 1764 -1050 1770 -1044
rect 1764 -1056 1770 -1050
rect 1764 -1062 1770 -1056
rect 1764 -1068 1770 -1062
rect 1764 -1074 1770 -1068
rect 1764 -1080 1770 -1074
rect 1764 -1086 1770 -1080
rect 1764 -1092 1770 -1086
rect 1764 -1098 1770 -1092
rect 1764 -1104 1770 -1098
rect 1764 -1110 1770 -1104
rect 1764 -1116 1770 -1110
rect 1764 -1122 1770 -1116
rect 1764 -1128 1770 -1122
rect 1764 -1134 1770 -1128
rect 1764 -1140 1770 -1134
rect 1764 -1146 1770 -1140
rect 1764 -1152 1770 -1146
rect 1764 -1158 1770 -1152
rect 1764 -1164 1770 -1158
rect 1764 -1170 1770 -1164
rect 1764 -1176 1770 -1170
rect 1764 -1182 1770 -1176
rect 1764 -1188 1770 -1182
rect 1764 -1194 1770 -1188
rect 1764 -1200 1770 -1194
rect 1764 -1206 1770 -1200
rect 1764 -1212 1770 -1206
rect 1764 -1218 1770 -1212
rect 1764 -1224 1770 -1218
rect 1764 -1230 1770 -1224
rect 1764 -1236 1770 -1230
rect 1764 -1242 1770 -1236
rect 1764 -1248 1770 -1242
rect 1764 -1254 1770 -1248
rect 1764 -1260 1770 -1254
rect 1764 -1266 1770 -1260
rect 1764 -1272 1770 -1266
rect 1764 -1278 1770 -1272
rect 1764 -1284 1770 -1278
rect 1764 -1290 1770 -1284
rect 1764 -1296 1770 -1290
rect 1764 -1302 1770 -1296
rect 1764 -1308 1770 -1302
rect 1764 -1314 1770 -1308
rect 1764 -1320 1770 -1314
rect 1764 -1326 1770 -1320
rect 1764 -1332 1770 -1326
rect 1764 -1338 1770 -1332
rect 1764 -1344 1770 -1338
rect 1764 -1350 1770 -1344
rect 1764 -1356 1770 -1350
rect 1764 -1362 1770 -1356
rect 1764 -1368 1770 -1362
rect 1764 -1374 1770 -1368
rect 1764 -1380 1770 -1374
rect 1764 -1386 1770 -1380
rect 1764 -1392 1770 -1386
rect 1764 -1398 1770 -1392
rect 1764 -1404 1770 -1398
rect 1764 -1410 1770 -1404
rect 1764 -1416 1770 -1410
rect 1764 -1422 1770 -1416
rect 1764 -1428 1770 -1422
rect 1764 -1434 1770 -1428
rect 1764 -1440 1770 -1434
rect 1764 -1446 1770 -1440
rect 1764 -1452 1770 -1446
rect 1764 -1458 1770 -1452
rect 1764 -1464 1770 -1458
rect 1764 -1470 1770 -1464
rect 1764 -1476 1770 -1470
rect 1764 -1482 1770 -1476
rect 1764 -1488 1770 -1482
rect 1764 -1494 1770 -1488
rect 1764 -1500 1770 -1494
rect 1764 -1506 1770 -1500
rect 1764 -1512 1770 -1506
rect 1764 -1518 1770 -1512
rect 1764 -1524 1770 -1518
rect 1764 -1530 1770 -1524
rect 1764 -1536 1770 -1530
rect 1764 -1542 1770 -1536
rect 1764 -1548 1770 -1542
rect 1764 -1554 1770 -1548
rect 1764 -1560 1770 -1554
rect 1764 -1566 1770 -1560
rect 1764 -1572 1770 -1566
rect 1764 -1578 1770 -1572
rect 1764 -1584 1770 -1578
rect 1764 -1590 1770 -1584
rect 1764 -1596 1770 -1590
rect 1764 -1602 1770 -1596
rect 1764 -1608 1770 -1602
rect 1764 -1614 1770 -1608
rect 1764 -1620 1770 -1614
rect 1764 -1626 1770 -1620
rect 1764 -1632 1770 -1626
rect 1764 -1638 1770 -1632
rect 1764 -1644 1770 -1638
rect 1764 -1650 1770 -1644
rect 1764 -1656 1770 -1650
rect 1764 -1662 1770 -1656
rect 1764 -1668 1770 -1662
rect 1764 -1674 1770 -1668
rect 1764 -1680 1770 -1674
rect 1764 -1686 1770 -1680
rect 1764 -1692 1770 -1686
rect 1764 -1698 1770 -1692
rect 1764 -1704 1770 -1698
rect 1764 -1710 1770 -1704
rect 1764 -1716 1770 -1710
rect 1764 -1722 1770 -1716
rect 1764 -1728 1770 -1722
rect 1764 -1734 1770 -1728
rect 1764 -1740 1770 -1734
rect 1764 -1746 1770 -1740
rect 1764 -1752 1770 -1746
rect 1764 -1758 1770 -1752
rect 1764 -1764 1770 -1758
rect 1764 -1770 1770 -1764
rect 1764 -1776 1770 -1770
rect 1764 -1782 1770 -1776
rect 1764 -1788 1770 -1782
rect 1764 -1794 1770 -1788
rect 1764 -1800 1770 -1794
rect 1764 -1806 1770 -1800
rect 1764 -1812 1770 -1806
rect 1764 -1818 1770 -1812
rect 1764 -1824 1770 -1818
rect 1764 -1830 1770 -1824
rect 1764 -1836 1770 -1830
rect 1764 -1842 1770 -1836
rect 1764 -1848 1770 -1842
rect 1764 -1854 1770 -1848
rect 1764 -1860 1770 -1854
rect 1764 -1866 1770 -1860
rect 1764 -1872 1770 -1866
rect 1764 -1878 1770 -1872
rect 1764 -1884 1770 -1878
rect 1764 -1962 1770 -1956
rect 1764 -1968 1770 -1962
rect 1764 -1974 1770 -1968
rect 1764 -1980 1770 -1974
rect 1764 -1986 1770 -1980
rect 1764 -1992 1770 -1986
rect 1764 -1998 1770 -1992
rect 1764 -2004 1770 -1998
rect 1764 -2010 1770 -2004
rect 1764 -2016 1770 -2010
rect 1764 -2022 1770 -2016
rect 1764 -2028 1770 -2022
rect 1764 -2034 1770 -2028
rect 1764 -2040 1770 -2034
rect 1764 -2046 1770 -2040
rect 1764 -2052 1770 -2046
rect 1764 -2058 1770 -2052
rect 1764 -2064 1770 -2058
rect 1764 -2070 1770 -2064
rect 1764 -2076 1770 -2070
rect 1764 -2082 1770 -2076
rect 1764 -2088 1770 -2082
rect 1764 -2094 1770 -2088
rect 1764 -2100 1770 -2094
rect 1764 -2106 1770 -2100
rect 1764 -2112 1770 -2106
rect 1764 -2118 1770 -2112
rect 1764 -2124 1770 -2118
rect 1764 -2130 1770 -2124
rect 1764 -2136 1770 -2130
rect 1764 -2142 1770 -2136
rect 1764 -2148 1770 -2142
rect 1764 -2154 1770 -2148
rect 1764 -2160 1770 -2154
rect 1764 -2166 1770 -2160
rect 1764 -2172 1770 -2166
rect 1764 -2178 1770 -2172
rect 1764 -2184 1770 -2178
rect 1764 -2190 1770 -2184
rect 1764 -2196 1770 -2190
rect 1764 -2202 1770 -2196
rect 1764 -2208 1770 -2202
rect 1764 -2214 1770 -2208
rect 1764 -2220 1770 -2214
rect 1764 -2226 1770 -2220
rect 1764 -2232 1770 -2226
rect 1764 -2238 1770 -2232
rect 1764 -2244 1770 -2238
rect 1764 -2250 1770 -2244
rect 1764 -2256 1770 -2250
rect 1764 -2262 1770 -2256
rect 1764 -2268 1770 -2262
rect 1764 -2274 1770 -2268
rect 1764 -2280 1770 -2274
rect 1764 -2286 1770 -2280
rect 1764 -2292 1770 -2286
rect 1764 -2298 1770 -2292
rect 1764 -2304 1770 -2298
rect 1764 -2310 1770 -2304
rect 1764 -2316 1770 -2310
rect 1764 -2322 1770 -2316
rect 1764 -2328 1770 -2322
rect 1764 -2334 1770 -2328
rect 1764 -2340 1770 -2334
rect 1764 -2346 1770 -2340
rect 1764 -2352 1770 -2346
rect 1764 -2358 1770 -2352
rect 1764 -2364 1770 -2358
rect 1764 -2370 1770 -2364
rect 1764 -2376 1770 -2370
rect 1764 -2382 1770 -2376
rect 1764 -2388 1770 -2382
rect 1764 -2394 1770 -2388
rect 1764 -2400 1770 -2394
rect 1764 -2406 1770 -2400
rect 1764 -2412 1770 -2406
rect 1764 -2418 1770 -2412
rect 1764 -2424 1770 -2418
rect 1764 -2430 1770 -2424
rect 1764 -2436 1770 -2430
rect 1764 -2442 1770 -2436
rect 1764 -2448 1770 -2442
rect 1764 -2454 1770 -2448
rect 1764 -2460 1770 -2454
rect 1764 -2466 1770 -2460
rect 1764 -2472 1770 -2466
rect 1764 -2478 1770 -2472
rect 1764 -2484 1770 -2478
rect 1764 -2490 1770 -2484
rect 1764 -2496 1770 -2490
rect 1764 -2502 1770 -2496
rect 1764 -2508 1770 -2502
rect 1764 -2514 1770 -2508
rect 1764 -2520 1770 -2514
rect 1764 -2526 1770 -2520
rect 1764 -2532 1770 -2526
rect 1764 -2538 1770 -2532
rect 1764 -2544 1770 -2538
rect 1764 -2550 1770 -2544
rect 1764 -2556 1770 -2550
rect 1764 -2562 1770 -2556
rect 1764 -2568 1770 -2562
rect 1764 -2574 1770 -2568
rect 1764 -2580 1770 -2574
rect 1764 -2586 1770 -2580
rect 1764 -2592 1770 -2586
rect 1764 -2598 1770 -2592
rect 1764 -2604 1770 -2598
rect 1764 -2610 1770 -2604
rect 1764 -2616 1770 -2610
rect 1764 -2622 1770 -2616
rect 1764 -2628 1770 -2622
rect 1764 -2634 1770 -2628
rect 1764 -2640 1770 -2634
rect 1764 -2646 1770 -2640
rect 1764 -2652 1770 -2646
rect 1764 -2724 1770 -2718
rect 1764 -2730 1770 -2724
rect 1764 -2736 1770 -2730
rect 1764 -2742 1770 -2736
rect 1764 -2748 1770 -2742
rect 1764 -2754 1770 -2748
rect 1764 -2760 1770 -2754
rect 1764 -2766 1770 -2760
rect 1764 -2772 1770 -2766
rect 1764 -2778 1770 -2772
rect 1764 -2784 1770 -2778
rect 1764 -2790 1770 -2784
rect 1764 -2796 1770 -2790
rect 1764 -2802 1770 -2796
rect 1764 -2808 1770 -2802
rect 1764 -2814 1770 -2808
rect 1764 -2820 1770 -2814
rect 1764 -2826 1770 -2820
rect 1764 -2832 1770 -2826
rect 1764 -2838 1770 -2832
rect 1764 -2844 1770 -2838
rect 1764 -2850 1770 -2844
rect 1764 -2856 1770 -2850
rect 1764 -2862 1770 -2856
rect 1764 -2868 1770 -2862
rect 1764 -2874 1770 -2868
rect 1764 -2880 1770 -2874
rect 1764 -2886 1770 -2880
rect 1764 -2892 1770 -2886
rect 1764 -2898 1770 -2892
rect 1764 -2904 1770 -2898
rect 1764 -2910 1770 -2904
rect 1764 -2916 1770 -2910
rect 1764 -2922 1770 -2916
rect 1764 -2928 1770 -2922
rect 1764 -2934 1770 -2928
rect 1764 -2940 1770 -2934
rect 1764 -2946 1770 -2940
rect 1764 -2952 1770 -2946
rect 1764 -2958 1770 -2952
rect 1764 -2964 1770 -2958
rect 1764 -2970 1770 -2964
rect 1764 -2976 1770 -2970
rect 1764 -2982 1770 -2976
rect 1764 -2988 1770 -2982
rect 1764 -2994 1770 -2988
rect 1764 -3000 1770 -2994
rect 1764 -3006 1770 -3000
rect 1764 -3012 1770 -3006
rect 1764 -3018 1770 -3012
rect 1764 -3024 1770 -3018
rect 1764 -3030 1770 -3024
rect 1764 -3036 1770 -3030
rect 1764 -3042 1770 -3036
rect 1764 -3048 1770 -3042
rect 1764 -3054 1770 -3048
rect 1764 -3060 1770 -3054
rect 1764 -3066 1770 -3060
rect 1764 -3072 1770 -3066
rect 1764 -3078 1770 -3072
rect 1764 -3084 1770 -3078
rect 1764 -3090 1770 -3084
rect 1764 -3096 1770 -3090
rect 1764 -3102 1770 -3096
rect 1764 -3108 1770 -3102
rect 1764 -3114 1770 -3108
rect 1764 -3120 1770 -3114
rect 1764 -3126 1770 -3120
rect 1764 -3132 1770 -3126
rect 1764 -3138 1770 -3132
rect 1764 -3144 1770 -3138
rect 1764 -3150 1770 -3144
rect 1764 -3156 1770 -3150
rect 1764 -3162 1770 -3156
rect 1764 -3168 1770 -3162
rect 1764 -3174 1770 -3168
rect 1764 -3180 1770 -3174
rect 1764 -3186 1770 -3180
rect 1764 -3192 1770 -3186
rect 1764 -3198 1770 -3192
rect 1764 -3246 1770 -3240
rect 1764 -3252 1770 -3246
rect 1764 -3258 1770 -3252
rect 1764 -3264 1770 -3258
rect 1764 -3270 1770 -3264
rect 1764 -3276 1770 -3270
rect 1764 -3282 1770 -3276
rect 1764 -3288 1770 -3282
rect 1764 -3294 1770 -3288
rect 1764 -3300 1770 -3294
rect 1764 -3306 1770 -3300
rect 1764 -3312 1770 -3306
rect 1764 -3318 1770 -3312
rect 1764 -3324 1770 -3318
rect 1764 -3330 1770 -3324
rect 1764 -3336 1770 -3330
rect 1764 -3342 1770 -3336
rect 1764 -3348 1770 -3342
rect 1764 -3354 1770 -3348
rect 1764 -3360 1770 -3354
rect 1764 -3366 1770 -3360
rect 1764 -3372 1770 -3366
rect 1764 -3378 1770 -3372
rect 1764 -3384 1770 -3378
rect 1764 -3390 1770 -3384
rect 1770 -762 1776 -756
rect 1770 -768 1776 -762
rect 1770 -774 1776 -768
rect 1770 -780 1776 -774
rect 1770 -786 1776 -780
rect 1770 -792 1776 -786
rect 1770 -798 1776 -792
rect 1770 -804 1776 -798
rect 1770 -810 1776 -804
rect 1770 -816 1776 -810
rect 1770 -822 1776 -816
rect 1770 -828 1776 -822
rect 1770 -834 1776 -828
rect 1770 -840 1776 -834
rect 1770 -846 1776 -840
rect 1770 -852 1776 -846
rect 1770 -858 1776 -852
rect 1770 -864 1776 -858
rect 1770 -870 1776 -864
rect 1770 -876 1776 -870
rect 1770 -882 1776 -876
rect 1770 -888 1776 -882
rect 1770 -894 1776 -888
rect 1770 -900 1776 -894
rect 1770 -906 1776 -900
rect 1770 -912 1776 -906
rect 1770 -918 1776 -912
rect 1770 -924 1776 -918
rect 1770 -930 1776 -924
rect 1770 -936 1776 -930
rect 1770 -942 1776 -936
rect 1770 -948 1776 -942
rect 1770 -954 1776 -948
rect 1770 -960 1776 -954
rect 1770 -966 1776 -960
rect 1770 -972 1776 -966
rect 1770 -978 1776 -972
rect 1770 -984 1776 -978
rect 1770 -990 1776 -984
rect 1770 -996 1776 -990
rect 1770 -1002 1776 -996
rect 1770 -1008 1776 -1002
rect 1770 -1014 1776 -1008
rect 1770 -1020 1776 -1014
rect 1770 -1026 1776 -1020
rect 1770 -1032 1776 -1026
rect 1770 -1038 1776 -1032
rect 1770 -1044 1776 -1038
rect 1770 -1050 1776 -1044
rect 1770 -1056 1776 -1050
rect 1770 -1062 1776 -1056
rect 1770 -1068 1776 -1062
rect 1770 -1074 1776 -1068
rect 1770 -1080 1776 -1074
rect 1770 -1086 1776 -1080
rect 1770 -1092 1776 -1086
rect 1770 -1098 1776 -1092
rect 1770 -1104 1776 -1098
rect 1770 -1110 1776 -1104
rect 1770 -1116 1776 -1110
rect 1770 -1122 1776 -1116
rect 1770 -1128 1776 -1122
rect 1770 -1134 1776 -1128
rect 1770 -1140 1776 -1134
rect 1770 -1146 1776 -1140
rect 1770 -1152 1776 -1146
rect 1770 -1158 1776 -1152
rect 1770 -1164 1776 -1158
rect 1770 -1170 1776 -1164
rect 1770 -1176 1776 -1170
rect 1770 -1182 1776 -1176
rect 1770 -1188 1776 -1182
rect 1770 -1194 1776 -1188
rect 1770 -1200 1776 -1194
rect 1770 -1206 1776 -1200
rect 1770 -1212 1776 -1206
rect 1770 -1218 1776 -1212
rect 1770 -1224 1776 -1218
rect 1770 -1230 1776 -1224
rect 1770 -1236 1776 -1230
rect 1770 -1242 1776 -1236
rect 1770 -1248 1776 -1242
rect 1770 -1254 1776 -1248
rect 1770 -1260 1776 -1254
rect 1770 -1266 1776 -1260
rect 1770 -1272 1776 -1266
rect 1770 -1278 1776 -1272
rect 1770 -1284 1776 -1278
rect 1770 -1290 1776 -1284
rect 1770 -1296 1776 -1290
rect 1770 -1302 1776 -1296
rect 1770 -1308 1776 -1302
rect 1770 -1314 1776 -1308
rect 1770 -1320 1776 -1314
rect 1770 -1326 1776 -1320
rect 1770 -1332 1776 -1326
rect 1770 -1338 1776 -1332
rect 1770 -1344 1776 -1338
rect 1770 -1350 1776 -1344
rect 1770 -1356 1776 -1350
rect 1770 -1362 1776 -1356
rect 1770 -1368 1776 -1362
rect 1770 -1374 1776 -1368
rect 1770 -1380 1776 -1374
rect 1770 -1386 1776 -1380
rect 1770 -1392 1776 -1386
rect 1770 -1398 1776 -1392
rect 1770 -1404 1776 -1398
rect 1770 -1410 1776 -1404
rect 1770 -1416 1776 -1410
rect 1770 -1422 1776 -1416
rect 1770 -1428 1776 -1422
rect 1770 -1434 1776 -1428
rect 1770 -1440 1776 -1434
rect 1770 -1446 1776 -1440
rect 1770 -1452 1776 -1446
rect 1770 -1458 1776 -1452
rect 1770 -1464 1776 -1458
rect 1770 -1470 1776 -1464
rect 1770 -1476 1776 -1470
rect 1770 -1482 1776 -1476
rect 1770 -1488 1776 -1482
rect 1770 -1494 1776 -1488
rect 1770 -1500 1776 -1494
rect 1770 -1506 1776 -1500
rect 1770 -1512 1776 -1506
rect 1770 -1518 1776 -1512
rect 1770 -1524 1776 -1518
rect 1770 -1530 1776 -1524
rect 1770 -1536 1776 -1530
rect 1770 -1542 1776 -1536
rect 1770 -1548 1776 -1542
rect 1770 -1554 1776 -1548
rect 1770 -1560 1776 -1554
rect 1770 -1566 1776 -1560
rect 1770 -1572 1776 -1566
rect 1770 -1578 1776 -1572
rect 1770 -1584 1776 -1578
rect 1770 -1590 1776 -1584
rect 1770 -1596 1776 -1590
rect 1770 -1602 1776 -1596
rect 1770 -1608 1776 -1602
rect 1770 -1614 1776 -1608
rect 1770 -1620 1776 -1614
rect 1770 -1626 1776 -1620
rect 1770 -1632 1776 -1626
rect 1770 -1638 1776 -1632
rect 1770 -1644 1776 -1638
rect 1770 -1650 1776 -1644
rect 1770 -1656 1776 -1650
rect 1770 -1662 1776 -1656
rect 1770 -1668 1776 -1662
rect 1770 -1674 1776 -1668
rect 1770 -1680 1776 -1674
rect 1770 -1686 1776 -1680
rect 1770 -1692 1776 -1686
rect 1770 -1698 1776 -1692
rect 1770 -1704 1776 -1698
rect 1770 -1710 1776 -1704
rect 1770 -1716 1776 -1710
rect 1770 -1722 1776 -1716
rect 1770 -1728 1776 -1722
rect 1770 -1734 1776 -1728
rect 1770 -1740 1776 -1734
rect 1770 -1746 1776 -1740
rect 1770 -1752 1776 -1746
rect 1770 -1758 1776 -1752
rect 1770 -1764 1776 -1758
rect 1770 -1770 1776 -1764
rect 1770 -1776 1776 -1770
rect 1770 -1782 1776 -1776
rect 1770 -1788 1776 -1782
rect 1770 -1794 1776 -1788
rect 1770 -1800 1776 -1794
rect 1770 -1806 1776 -1800
rect 1770 -1812 1776 -1806
rect 1770 -1818 1776 -1812
rect 1770 -1824 1776 -1818
rect 1770 -1830 1776 -1824
rect 1770 -1836 1776 -1830
rect 1770 -1842 1776 -1836
rect 1770 -1848 1776 -1842
rect 1770 -1854 1776 -1848
rect 1770 -1860 1776 -1854
rect 1770 -1866 1776 -1860
rect 1770 -1872 1776 -1866
rect 1770 -1878 1776 -1872
rect 1770 -1956 1776 -1950
rect 1770 -1962 1776 -1956
rect 1770 -1968 1776 -1962
rect 1770 -1974 1776 -1968
rect 1770 -1980 1776 -1974
rect 1770 -1986 1776 -1980
rect 1770 -1992 1776 -1986
rect 1770 -1998 1776 -1992
rect 1770 -2004 1776 -1998
rect 1770 -2010 1776 -2004
rect 1770 -2016 1776 -2010
rect 1770 -2022 1776 -2016
rect 1770 -2028 1776 -2022
rect 1770 -2034 1776 -2028
rect 1770 -2040 1776 -2034
rect 1770 -2046 1776 -2040
rect 1770 -2052 1776 -2046
rect 1770 -2058 1776 -2052
rect 1770 -2064 1776 -2058
rect 1770 -2070 1776 -2064
rect 1770 -2076 1776 -2070
rect 1770 -2082 1776 -2076
rect 1770 -2088 1776 -2082
rect 1770 -2094 1776 -2088
rect 1770 -2100 1776 -2094
rect 1770 -2106 1776 -2100
rect 1770 -2112 1776 -2106
rect 1770 -2118 1776 -2112
rect 1770 -2124 1776 -2118
rect 1770 -2130 1776 -2124
rect 1770 -2136 1776 -2130
rect 1770 -2142 1776 -2136
rect 1770 -2148 1776 -2142
rect 1770 -2154 1776 -2148
rect 1770 -2160 1776 -2154
rect 1770 -2166 1776 -2160
rect 1770 -2172 1776 -2166
rect 1770 -2178 1776 -2172
rect 1770 -2184 1776 -2178
rect 1770 -2190 1776 -2184
rect 1770 -2196 1776 -2190
rect 1770 -2202 1776 -2196
rect 1770 -2208 1776 -2202
rect 1770 -2214 1776 -2208
rect 1770 -2220 1776 -2214
rect 1770 -2226 1776 -2220
rect 1770 -2232 1776 -2226
rect 1770 -2238 1776 -2232
rect 1770 -2244 1776 -2238
rect 1770 -2250 1776 -2244
rect 1770 -2256 1776 -2250
rect 1770 -2262 1776 -2256
rect 1770 -2268 1776 -2262
rect 1770 -2274 1776 -2268
rect 1770 -2280 1776 -2274
rect 1770 -2286 1776 -2280
rect 1770 -2292 1776 -2286
rect 1770 -2298 1776 -2292
rect 1770 -2304 1776 -2298
rect 1770 -2310 1776 -2304
rect 1770 -2316 1776 -2310
rect 1770 -2322 1776 -2316
rect 1770 -2328 1776 -2322
rect 1770 -2334 1776 -2328
rect 1770 -2340 1776 -2334
rect 1770 -2346 1776 -2340
rect 1770 -2352 1776 -2346
rect 1770 -2358 1776 -2352
rect 1770 -2364 1776 -2358
rect 1770 -2370 1776 -2364
rect 1770 -2376 1776 -2370
rect 1770 -2382 1776 -2376
rect 1770 -2388 1776 -2382
rect 1770 -2394 1776 -2388
rect 1770 -2400 1776 -2394
rect 1770 -2406 1776 -2400
rect 1770 -2412 1776 -2406
rect 1770 -2418 1776 -2412
rect 1770 -2424 1776 -2418
rect 1770 -2430 1776 -2424
rect 1770 -2436 1776 -2430
rect 1770 -2442 1776 -2436
rect 1770 -2448 1776 -2442
rect 1770 -2454 1776 -2448
rect 1770 -2460 1776 -2454
rect 1770 -2466 1776 -2460
rect 1770 -2472 1776 -2466
rect 1770 -2478 1776 -2472
rect 1770 -2484 1776 -2478
rect 1770 -2490 1776 -2484
rect 1770 -2496 1776 -2490
rect 1770 -2502 1776 -2496
rect 1770 -2508 1776 -2502
rect 1770 -2514 1776 -2508
rect 1770 -2520 1776 -2514
rect 1770 -2526 1776 -2520
rect 1770 -2532 1776 -2526
rect 1770 -2538 1776 -2532
rect 1770 -2544 1776 -2538
rect 1770 -2550 1776 -2544
rect 1770 -2556 1776 -2550
rect 1770 -2562 1776 -2556
rect 1770 -2568 1776 -2562
rect 1770 -2574 1776 -2568
rect 1770 -2580 1776 -2574
rect 1770 -2586 1776 -2580
rect 1770 -2592 1776 -2586
rect 1770 -2598 1776 -2592
rect 1770 -2604 1776 -2598
rect 1770 -2610 1776 -2604
rect 1770 -2616 1776 -2610
rect 1770 -2622 1776 -2616
rect 1770 -2628 1776 -2622
rect 1770 -2634 1776 -2628
rect 1770 -2640 1776 -2634
rect 1770 -2646 1776 -2640
rect 1770 -2724 1776 -2718
rect 1770 -2730 1776 -2724
rect 1770 -2736 1776 -2730
rect 1770 -2742 1776 -2736
rect 1770 -2748 1776 -2742
rect 1770 -2754 1776 -2748
rect 1770 -2760 1776 -2754
rect 1770 -2766 1776 -2760
rect 1770 -2772 1776 -2766
rect 1770 -2778 1776 -2772
rect 1770 -2784 1776 -2778
rect 1770 -2790 1776 -2784
rect 1770 -2796 1776 -2790
rect 1770 -2802 1776 -2796
rect 1770 -2808 1776 -2802
rect 1770 -2814 1776 -2808
rect 1770 -2820 1776 -2814
rect 1770 -2826 1776 -2820
rect 1770 -2832 1776 -2826
rect 1770 -2838 1776 -2832
rect 1770 -2844 1776 -2838
rect 1770 -2850 1776 -2844
rect 1770 -2856 1776 -2850
rect 1770 -2862 1776 -2856
rect 1770 -2868 1776 -2862
rect 1770 -2874 1776 -2868
rect 1770 -2880 1776 -2874
rect 1770 -2886 1776 -2880
rect 1770 -2892 1776 -2886
rect 1770 -2898 1776 -2892
rect 1770 -2904 1776 -2898
rect 1770 -2910 1776 -2904
rect 1770 -2916 1776 -2910
rect 1770 -2922 1776 -2916
rect 1770 -2928 1776 -2922
rect 1770 -2934 1776 -2928
rect 1770 -2940 1776 -2934
rect 1770 -2946 1776 -2940
rect 1770 -2952 1776 -2946
rect 1770 -2958 1776 -2952
rect 1770 -2964 1776 -2958
rect 1770 -2970 1776 -2964
rect 1770 -2976 1776 -2970
rect 1770 -2982 1776 -2976
rect 1770 -2988 1776 -2982
rect 1770 -2994 1776 -2988
rect 1770 -3000 1776 -2994
rect 1770 -3006 1776 -3000
rect 1770 -3012 1776 -3006
rect 1770 -3018 1776 -3012
rect 1770 -3024 1776 -3018
rect 1770 -3030 1776 -3024
rect 1770 -3036 1776 -3030
rect 1770 -3042 1776 -3036
rect 1770 -3048 1776 -3042
rect 1770 -3054 1776 -3048
rect 1770 -3060 1776 -3054
rect 1770 -3066 1776 -3060
rect 1770 -3072 1776 -3066
rect 1770 -3078 1776 -3072
rect 1770 -3084 1776 -3078
rect 1770 -3090 1776 -3084
rect 1770 -3096 1776 -3090
rect 1770 -3102 1776 -3096
rect 1770 -3108 1776 -3102
rect 1770 -3114 1776 -3108
rect 1770 -3120 1776 -3114
rect 1770 -3126 1776 -3120
rect 1770 -3132 1776 -3126
rect 1770 -3138 1776 -3132
rect 1770 -3144 1776 -3138
rect 1770 -3150 1776 -3144
rect 1770 -3156 1776 -3150
rect 1770 -3162 1776 -3156
rect 1770 -3168 1776 -3162
rect 1770 -3174 1776 -3168
rect 1770 -3180 1776 -3174
rect 1770 -3186 1776 -3180
rect 1770 -3192 1776 -3186
rect 1770 -3246 1776 -3240
rect 1770 -3252 1776 -3246
rect 1770 -3258 1776 -3252
rect 1770 -3264 1776 -3258
rect 1770 -3270 1776 -3264
rect 1770 -3276 1776 -3270
rect 1770 -3282 1776 -3276
rect 1770 -3288 1776 -3282
rect 1770 -3294 1776 -3288
rect 1770 -3300 1776 -3294
rect 1770 -3306 1776 -3300
rect 1770 -3312 1776 -3306
rect 1770 -3318 1776 -3312
rect 1770 -3324 1776 -3318
rect 1770 -3330 1776 -3324
rect 1770 -3336 1776 -3330
rect 1770 -3342 1776 -3336
rect 1770 -3348 1776 -3342
rect 1770 -3354 1776 -3348
rect 1770 -3360 1776 -3354
rect 1770 -3366 1776 -3360
rect 1770 -3372 1776 -3366
rect 1770 -3378 1776 -3372
rect 1770 -3384 1776 -3378
rect 1776 -756 1782 -750
rect 1776 -762 1782 -756
rect 1776 -768 1782 -762
rect 1776 -774 1782 -768
rect 1776 -780 1782 -774
rect 1776 -786 1782 -780
rect 1776 -792 1782 -786
rect 1776 -798 1782 -792
rect 1776 -804 1782 -798
rect 1776 -810 1782 -804
rect 1776 -816 1782 -810
rect 1776 -822 1782 -816
rect 1776 -828 1782 -822
rect 1776 -834 1782 -828
rect 1776 -840 1782 -834
rect 1776 -846 1782 -840
rect 1776 -852 1782 -846
rect 1776 -858 1782 -852
rect 1776 -864 1782 -858
rect 1776 -870 1782 -864
rect 1776 -876 1782 -870
rect 1776 -882 1782 -876
rect 1776 -888 1782 -882
rect 1776 -894 1782 -888
rect 1776 -900 1782 -894
rect 1776 -906 1782 -900
rect 1776 -912 1782 -906
rect 1776 -918 1782 -912
rect 1776 -924 1782 -918
rect 1776 -930 1782 -924
rect 1776 -936 1782 -930
rect 1776 -942 1782 -936
rect 1776 -948 1782 -942
rect 1776 -954 1782 -948
rect 1776 -960 1782 -954
rect 1776 -966 1782 -960
rect 1776 -972 1782 -966
rect 1776 -978 1782 -972
rect 1776 -984 1782 -978
rect 1776 -990 1782 -984
rect 1776 -996 1782 -990
rect 1776 -1002 1782 -996
rect 1776 -1008 1782 -1002
rect 1776 -1014 1782 -1008
rect 1776 -1020 1782 -1014
rect 1776 -1026 1782 -1020
rect 1776 -1032 1782 -1026
rect 1776 -1038 1782 -1032
rect 1776 -1044 1782 -1038
rect 1776 -1050 1782 -1044
rect 1776 -1056 1782 -1050
rect 1776 -1062 1782 -1056
rect 1776 -1068 1782 -1062
rect 1776 -1074 1782 -1068
rect 1776 -1080 1782 -1074
rect 1776 -1086 1782 -1080
rect 1776 -1092 1782 -1086
rect 1776 -1098 1782 -1092
rect 1776 -1104 1782 -1098
rect 1776 -1110 1782 -1104
rect 1776 -1116 1782 -1110
rect 1776 -1122 1782 -1116
rect 1776 -1128 1782 -1122
rect 1776 -1134 1782 -1128
rect 1776 -1140 1782 -1134
rect 1776 -1146 1782 -1140
rect 1776 -1152 1782 -1146
rect 1776 -1158 1782 -1152
rect 1776 -1164 1782 -1158
rect 1776 -1170 1782 -1164
rect 1776 -1176 1782 -1170
rect 1776 -1182 1782 -1176
rect 1776 -1188 1782 -1182
rect 1776 -1194 1782 -1188
rect 1776 -1200 1782 -1194
rect 1776 -1206 1782 -1200
rect 1776 -1212 1782 -1206
rect 1776 -1218 1782 -1212
rect 1776 -1224 1782 -1218
rect 1776 -1230 1782 -1224
rect 1776 -1236 1782 -1230
rect 1776 -1242 1782 -1236
rect 1776 -1248 1782 -1242
rect 1776 -1254 1782 -1248
rect 1776 -1260 1782 -1254
rect 1776 -1266 1782 -1260
rect 1776 -1272 1782 -1266
rect 1776 -1278 1782 -1272
rect 1776 -1284 1782 -1278
rect 1776 -1290 1782 -1284
rect 1776 -1296 1782 -1290
rect 1776 -1302 1782 -1296
rect 1776 -1308 1782 -1302
rect 1776 -1314 1782 -1308
rect 1776 -1320 1782 -1314
rect 1776 -1326 1782 -1320
rect 1776 -1332 1782 -1326
rect 1776 -1338 1782 -1332
rect 1776 -1344 1782 -1338
rect 1776 -1350 1782 -1344
rect 1776 -1356 1782 -1350
rect 1776 -1362 1782 -1356
rect 1776 -1368 1782 -1362
rect 1776 -1374 1782 -1368
rect 1776 -1380 1782 -1374
rect 1776 -1386 1782 -1380
rect 1776 -1392 1782 -1386
rect 1776 -1398 1782 -1392
rect 1776 -1404 1782 -1398
rect 1776 -1410 1782 -1404
rect 1776 -1416 1782 -1410
rect 1776 -1422 1782 -1416
rect 1776 -1428 1782 -1422
rect 1776 -1434 1782 -1428
rect 1776 -1440 1782 -1434
rect 1776 -1446 1782 -1440
rect 1776 -1452 1782 -1446
rect 1776 -1458 1782 -1452
rect 1776 -1464 1782 -1458
rect 1776 -1470 1782 -1464
rect 1776 -1476 1782 -1470
rect 1776 -1482 1782 -1476
rect 1776 -1488 1782 -1482
rect 1776 -1494 1782 -1488
rect 1776 -1500 1782 -1494
rect 1776 -1506 1782 -1500
rect 1776 -1512 1782 -1506
rect 1776 -1518 1782 -1512
rect 1776 -1524 1782 -1518
rect 1776 -1530 1782 -1524
rect 1776 -1536 1782 -1530
rect 1776 -1542 1782 -1536
rect 1776 -1548 1782 -1542
rect 1776 -1554 1782 -1548
rect 1776 -1560 1782 -1554
rect 1776 -1566 1782 -1560
rect 1776 -1572 1782 -1566
rect 1776 -1578 1782 -1572
rect 1776 -1584 1782 -1578
rect 1776 -1590 1782 -1584
rect 1776 -1596 1782 -1590
rect 1776 -1602 1782 -1596
rect 1776 -1608 1782 -1602
rect 1776 -1614 1782 -1608
rect 1776 -1620 1782 -1614
rect 1776 -1626 1782 -1620
rect 1776 -1632 1782 -1626
rect 1776 -1638 1782 -1632
rect 1776 -1644 1782 -1638
rect 1776 -1650 1782 -1644
rect 1776 -1656 1782 -1650
rect 1776 -1662 1782 -1656
rect 1776 -1668 1782 -1662
rect 1776 -1674 1782 -1668
rect 1776 -1680 1782 -1674
rect 1776 -1686 1782 -1680
rect 1776 -1692 1782 -1686
rect 1776 -1698 1782 -1692
rect 1776 -1704 1782 -1698
rect 1776 -1710 1782 -1704
rect 1776 -1716 1782 -1710
rect 1776 -1722 1782 -1716
rect 1776 -1728 1782 -1722
rect 1776 -1734 1782 -1728
rect 1776 -1740 1782 -1734
rect 1776 -1746 1782 -1740
rect 1776 -1752 1782 -1746
rect 1776 -1758 1782 -1752
rect 1776 -1764 1782 -1758
rect 1776 -1770 1782 -1764
rect 1776 -1776 1782 -1770
rect 1776 -1782 1782 -1776
rect 1776 -1788 1782 -1782
rect 1776 -1794 1782 -1788
rect 1776 -1800 1782 -1794
rect 1776 -1806 1782 -1800
rect 1776 -1812 1782 -1806
rect 1776 -1818 1782 -1812
rect 1776 -1824 1782 -1818
rect 1776 -1830 1782 -1824
rect 1776 -1836 1782 -1830
rect 1776 -1842 1782 -1836
rect 1776 -1848 1782 -1842
rect 1776 -1854 1782 -1848
rect 1776 -1860 1782 -1854
rect 1776 -1866 1782 -1860
rect 1776 -1872 1782 -1866
rect 1776 -1950 1782 -1944
rect 1776 -1956 1782 -1950
rect 1776 -1962 1782 -1956
rect 1776 -1968 1782 -1962
rect 1776 -1974 1782 -1968
rect 1776 -1980 1782 -1974
rect 1776 -1986 1782 -1980
rect 1776 -1992 1782 -1986
rect 1776 -1998 1782 -1992
rect 1776 -2004 1782 -1998
rect 1776 -2010 1782 -2004
rect 1776 -2016 1782 -2010
rect 1776 -2022 1782 -2016
rect 1776 -2028 1782 -2022
rect 1776 -2034 1782 -2028
rect 1776 -2040 1782 -2034
rect 1776 -2046 1782 -2040
rect 1776 -2052 1782 -2046
rect 1776 -2058 1782 -2052
rect 1776 -2064 1782 -2058
rect 1776 -2070 1782 -2064
rect 1776 -2076 1782 -2070
rect 1776 -2082 1782 -2076
rect 1776 -2088 1782 -2082
rect 1776 -2094 1782 -2088
rect 1776 -2100 1782 -2094
rect 1776 -2106 1782 -2100
rect 1776 -2112 1782 -2106
rect 1776 -2118 1782 -2112
rect 1776 -2124 1782 -2118
rect 1776 -2130 1782 -2124
rect 1776 -2136 1782 -2130
rect 1776 -2142 1782 -2136
rect 1776 -2148 1782 -2142
rect 1776 -2154 1782 -2148
rect 1776 -2160 1782 -2154
rect 1776 -2166 1782 -2160
rect 1776 -2172 1782 -2166
rect 1776 -2178 1782 -2172
rect 1776 -2184 1782 -2178
rect 1776 -2190 1782 -2184
rect 1776 -2196 1782 -2190
rect 1776 -2202 1782 -2196
rect 1776 -2208 1782 -2202
rect 1776 -2214 1782 -2208
rect 1776 -2220 1782 -2214
rect 1776 -2226 1782 -2220
rect 1776 -2232 1782 -2226
rect 1776 -2238 1782 -2232
rect 1776 -2244 1782 -2238
rect 1776 -2250 1782 -2244
rect 1776 -2256 1782 -2250
rect 1776 -2262 1782 -2256
rect 1776 -2268 1782 -2262
rect 1776 -2274 1782 -2268
rect 1776 -2280 1782 -2274
rect 1776 -2286 1782 -2280
rect 1776 -2292 1782 -2286
rect 1776 -2298 1782 -2292
rect 1776 -2304 1782 -2298
rect 1776 -2310 1782 -2304
rect 1776 -2316 1782 -2310
rect 1776 -2322 1782 -2316
rect 1776 -2328 1782 -2322
rect 1776 -2334 1782 -2328
rect 1776 -2340 1782 -2334
rect 1776 -2346 1782 -2340
rect 1776 -2352 1782 -2346
rect 1776 -2358 1782 -2352
rect 1776 -2364 1782 -2358
rect 1776 -2370 1782 -2364
rect 1776 -2376 1782 -2370
rect 1776 -2382 1782 -2376
rect 1776 -2388 1782 -2382
rect 1776 -2394 1782 -2388
rect 1776 -2400 1782 -2394
rect 1776 -2406 1782 -2400
rect 1776 -2412 1782 -2406
rect 1776 -2418 1782 -2412
rect 1776 -2424 1782 -2418
rect 1776 -2430 1782 -2424
rect 1776 -2436 1782 -2430
rect 1776 -2442 1782 -2436
rect 1776 -2448 1782 -2442
rect 1776 -2454 1782 -2448
rect 1776 -2460 1782 -2454
rect 1776 -2466 1782 -2460
rect 1776 -2472 1782 -2466
rect 1776 -2478 1782 -2472
rect 1776 -2484 1782 -2478
rect 1776 -2490 1782 -2484
rect 1776 -2496 1782 -2490
rect 1776 -2502 1782 -2496
rect 1776 -2508 1782 -2502
rect 1776 -2514 1782 -2508
rect 1776 -2520 1782 -2514
rect 1776 -2526 1782 -2520
rect 1776 -2532 1782 -2526
rect 1776 -2538 1782 -2532
rect 1776 -2544 1782 -2538
rect 1776 -2550 1782 -2544
rect 1776 -2556 1782 -2550
rect 1776 -2562 1782 -2556
rect 1776 -2568 1782 -2562
rect 1776 -2574 1782 -2568
rect 1776 -2580 1782 -2574
rect 1776 -2586 1782 -2580
rect 1776 -2592 1782 -2586
rect 1776 -2598 1782 -2592
rect 1776 -2604 1782 -2598
rect 1776 -2610 1782 -2604
rect 1776 -2616 1782 -2610
rect 1776 -2622 1782 -2616
rect 1776 -2628 1782 -2622
rect 1776 -2634 1782 -2628
rect 1776 -2640 1782 -2634
rect 1776 -2646 1782 -2640
rect 1776 -2718 1782 -2712
rect 1776 -2724 1782 -2718
rect 1776 -2730 1782 -2724
rect 1776 -2736 1782 -2730
rect 1776 -2742 1782 -2736
rect 1776 -2748 1782 -2742
rect 1776 -2754 1782 -2748
rect 1776 -2760 1782 -2754
rect 1776 -2766 1782 -2760
rect 1776 -2772 1782 -2766
rect 1776 -2778 1782 -2772
rect 1776 -2784 1782 -2778
rect 1776 -2790 1782 -2784
rect 1776 -2796 1782 -2790
rect 1776 -2802 1782 -2796
rect 1776 -2808 1782 -2802
rect 1776 -2814 1782 -2808
rect 1776 -2820 1782 -2814
rect 1776 -2826 1782 -2820
rect 1776 -2832 1782 -2826
rect 1776 -2838 1782 -2832
rect 1776 -2844 1782 -2838
rect 1776 -2850 1782 -2844
rect 1776 -2856 1782 -2850
rect 1776 -2862 1782 -2856
rect 1776 -2868 1782 -2862
rect 1776 -2874 1782 -2868
rect 1776 -2880 1782 -2874
rect 1776 -2886 1782 -2880
rect 1776 -2892 1782 -2886
rect 1776 -2898 1782 -2892
rect 1776 -2904 1782 -2898
rect 1776 -2910 1782 -2904
rect 1776 -2916 1782 -2910
rect 1776 -2922 1782 -2916
rect 1776 -2928 1782 -2922
rect 1776 -2934 1782 -2928
rect 1776 -2940 1782 -2934
rect 1776 -2946 1782 -2940
rect 1776 -2952 1782 -2946
rect 1776 -2958 1782 -2952
rect 1776 -2964 1782 -2958
rect 1776 -2970 1782 -2964
rect 1776 -2976 1782 -2970
rect 1776 -2982 1782 -2976
rect 1776 -2988 1782 -2982
rect 1776 -2994 1782 -2988
rect 1776 -3000 1782 -2994
rect 1776 -3006 1782 -3000
rect 1776 -3012 1782 -3006
rect 1776 -3018 1782 -3012
rect 1776 -3024 1782 -3018
rect 1776 -3030 1782 -3024
rect 1776 -3036 1782 -3030
rect 1776 -3042 1782 -3036
rect 1776 -3048 1782 -3042
rect 1776 -3054 1782 -3048
rect 1776 -3060 1782 -3054
rect 1776 -3066 1782 -3060
rect 1776 -3072 1782 -3066
rect 1776 -3078 1782 -3072
rect 1776 -3084 1782 -3078
rect 1776 -3090 1782 -3084
rect 1776 -3096 1782 -3090
rect 1776 -3102 1782 -3096
rect 1776 -3108 1782 -3102
rect 1776 -3114 1782 -3108
rect 1776 -3120 1782 -3114
rect 1776 -3126 1782 -3120
rect 1776 -3132 1782 -3126
rect 1776 -3138 1782 -3132
rect 1776 -3144 1782 -3138
rect 1776 -3150 1782 -3144
rect 1776 -3156 1782 -3150
rect 1776 -3162 1782 -3156
rect 1776 -3168 1782 -3162
rect 1776 -3174 1782 -3168
rect 1776 -3180 1782 -3174
rect 1776 -3186 1782 -3180
rect 1776 -3192 1782 -3186
rect 1776 -3240 1782 -3234
rect 1776 -3246 1782 -3240
rect 1776 -3252 1782 -3246
rect 1776 -3258 1782 -3252
rect 1776 -3264 1782 -3258
rect 1776 -3270 1782 -3264
rect 1776 -3276 1782 -3270
rect 1776 -3282 1782 -3276
rect 1776 -3288 1782 -3282
rect 1776 -3294 1782 -3288
rect 1776 -3300 1782 -3294
rect 1776 -3306 1782 -3300
rect 1776 -3312 1782 -3306
rect 1776 -3318 1782 -3312
rect 1776 -3324 1782 -3318
rect 1776 -3330 1782 -3324
rect 1776 -3336 1782 -3330
rect 1776 -3342 1782 -3336
rect 1776 -3348 1782 -3342
rect 1776 -3354 1782 -3348
rect 1776 -3360 1782 -3354
rect 1776 -3366 1782 -3360
rect 1776 -3372 1782 -3366
rect 1776 -3378 1782 -3372
rect 1776 -3384 1782 -3378
rect 1782 -744 1788 -738
rect 1782 -750 1788 -744
rect 1782 -756 1788 -750
rect 1782 -762 1788 -756
rect 1782 -768 1788 -762
rect 1782 -774 1788 -768
rect 1782 -780 1788 -774
rect 1782 -786 1788 -780
rect 1782 -792 1788 -786
rect 1782 -798 1788 -792
rect 1782 -804 1788 -798
rect 1782 -810 1788 -804
rect 1782 -816 1788 -810
rect 1782 -822 1788 -816
rect 1782 -828 1788 -822
rect 1782 -834 1788 -828
rect 1782 -840 1788 -834
rect 1782 -846 1788 -840
rect 1782 -852 1788 -846
rect 1782 -858 1788 -852
rect 1782 -864 1788 -858
rect 1782 -870 1788 -864
rect 1782 -876 1788 -870
rect 1782 -882 1788 -876
rect 1782 -888 1788 -882
rect 1782 -894 1788 -888
rect 1782 -900 1788 -894
rect 1782 -906 1788 -900
rect 1782 -912 1788 -906
rect 1782 -918 1788 -912
rect 1782 -924 1788 -918
rect 1782 -930 1788 -924
rect 1782 -936 1788 -930
rect 1782 -942 1788 -936
rect 1782 -948 1788 -942
rect 1782 -954 1788 -948
rect 1782 -960 1788 -954
rect 1782 -966 1788 -960
rect 1782 -972 1788 -966
rect 1782 -978 1788 -972
rect 1782 -984 1788 -978
rect 1782 -990 1788 -984
rect 1782 -996 1788 -990
rect 1782 -1002 1788 -996
rect 1782 -1008 1788 -1002
rect 1782 -1014 1788 -1008
rect 1782 -1020 1788 -1014
rect 1782 -1026 1788 -1020
rect 1782 -1032 1788 -1026
rect 1782 -1038 1788 -1032
rect 1782 -1044 1788 -1038
rect 1782 -1050 1788 -1044
rect 1782 -1056 1788 -1050
rect 1782 -1062 1788 -1056
rect 1782 -1068 1788 -1062
rect 1782 -1074 1788 -1068
rect 1782 -1080 1788 -1074
rect 1782 -1086 1788 -1080
rect 1782 -1092 1788 -1086
rect 1782 -1098 1788 -1092
rect 1782 -1104 1788 -1098
rect 1782 -1110 1788 -1104
rect 1782 -1116 1788 -1110
rect 1782 -1122 1788 -1116
rect 1782 -1128 1788 -1122
rect 1782 -1134 1788 -1128
rect 1782 -1140 1788 -1134
rect 1782 -1146 1788 -1140
rect 1782 -1152 1788 -1146
rect 1782 -1158 1788 -1152
rect 1782 -1164 1788 -1158
rect 1782 -1170 1788 -1164
rect 1782 -1176 1788 -1170
rect 1782 -1182 1788 -1176
rect 1782 -1188 1788 -1182
rect 1782 -1194 1788 -1188
rect 1782 -1200 1788 -1194
rect 1782 -1206 1788 -1200
rect 1782 -1212 1788 -1206
rect 1782 -1218 1788 -1212
rect 1782 -1224 1788 -1218
rect 1782 -1230 1788 -1224
rect 1782 -1236 1788 -1230
rect 1782 -1242 1788 -1236
rect 1782 -1248 1788 -1242
rect 1782 -1254 1788 -1248
rect 1782 -1260 1788 -1254
rect 1782 -1266 1788 -1260
rect 1782 -1272 1788 -1266
rect 1782 -1278 1788 -1272
rect 1782 -1284 1788 -1278
rect 1782 -1290 1788 -1284
rect 1782 -1296 1788 -1290
rect 1782 -1302 1788 -1296
rect 1782 -1308 1788 -1302
rect 1782 -1314 1788 -1308
rect 1782 -1320 1788 -1314
rect 1782 -1326 1788 -1320
rect 1782 -1332 1788 -1326
rect 1782 -1338 1788 -1332
rect 1782 -1344 1788 -1338
rect 1782 -1350 1788 -1344
rect 1782 -1356 1788 -1350
rect 1782 -1362 1788 -1356
rect 1782 -1368 1788 -1362
rect 1782 -1374 1788 -1368
rect 1782 -1380 1788 -1374
rect 1782 -1386 1788 -1380
rect 1782 -1392 1788 -1386
rect 1782 -1398 1788 -1392
rect 1782 -1404 1788 -1398
rect 1782 -1410 1788 -1404
rect 1782 -1416 1788 -1410
rect 1782 -1422 1788 -1416
rect 1782 -1428 1788 -1422
rect 1782 -1434 1788 -1428
rect 1782 -1440 1788 -1434
rect 1782 -1446 1788 -1440
rect 1782 -1452 1788 -1446
rect 1782 -1458 1788 -1452
rect 1782 -1464 1788 -1458
rect 1782 -1470 1788 -1464
rect 1782 -1476 1788 -1470
rect 1782 -1482 1788 -1476
rect 1782 -1488 1788 -1482
rect 1782 -1494 1788 -1488
rect 1782 -1500 1788 -1494
rect 1782 -1506 1788 -1500
rect 1782 -1512 1788 -1506
rect 1782 -1518 1788 -1512
rect 1782 -1524 1788 -1518
rect 1782 -1530 1788 -1524
rect 1782 -1536 1788 -1530
rect 1782 -1542 1788 -1536
rect 1782 -1548 1788 -1542
rect 1782 -1554 1788 -1548
rect 1782 -1560 1788 -1554
rect 1782 -1566 1788 -1560
rect 1782 -1572 1788 -1566
rect 1782 -1578 1788 -1572
rect 1782 -1584 1788 -1578
rect 1782 -1590 1788 -1584
rect 1782 -1596 1788 -1590
rect 1782 -1602 1788 -1596
rect 1782 -1608 1788 -1602
rect 1782 -1614 1788 -1608
rect 1782 -1620 1788 -1614
rect 1782 -1626 1788 -1620
rect 1782 -1632 1788 -1626
rect 1782 -1638 1788 -1632
rect 1782 -1644 1788 -1638
rect 1782 -1650 1788 -1644
rect 1782 -1656 1788 -1650
rect 1782 -1662 1788 -1656
rect 1782 -1668 1788 -1662
rect 1782 -1674 1788 -1668
rect 1782 -1680 1788 -1674
rect 1782 -1686 1788 -1680
rect 1782 -1692 1788 -1686
rect 1782 -1698 1788 -1692
rect 1782 -1704 1788 -1698
rect 1782 -1710 1788 -1704
rect 1782 -1716 1788 -1710
rect 1782 -1722 1788 -1716
rect 1782 -1728 1788 -1722
rect 1782 -1734 1788 -1728
rect 1782 -1740 1788 -1734
rect 1782 -1746 1788 -1740
rect 1782 -1752 1788 -1746
rect 1782 -1758 1788 -1752
rect 1782 -1764 1788 -1758
rect 1782 -1770 1788 -1764
rect 1782 -1776 1788 -1770
rect 1782 -1782 1788 -1776
rect 1782 -1788 1788 -1782
rect 1782 -1794 1788 -1788
rect 1782 -1800 1788 -1794
rect 1782 -1806 1788 -1800
rect 1782 -1812 1788 -1806
rect 1782 -1818 1788 -1812
rect 1782 -1824 1788 -1818
rect 1782 -1830 1788 -1824
rect 1782 -1836 1788 -1830
rect 1782 -1842 1788 -1836
rect 1782 -1848 1788 -1842
rect 1782 -1854 1788 -1848
rect 1782 -1860 1788 -1854
rect 1782 -1866 1788 -1860
rect 1782 -1944 1788 -1938
rect 1782 -1950 1788 -1944
rect 1782 -1956 1788 -1950
rect 1782 -1962 1788 -1956
rect 1782 -1968 1788 -1962
rect 1782 -1974 1788 -1968
rect 1782 -1980 1788 -1974
rect 1782 -1986 1788 -1980
rect 1782 -1992 1788 -1986
rect 1782 -1998 1788 -1992
rect 1782 -2004 1788 -1998
rect 1782 -2010 1788 -2004
rect 1782 -2016 1788 -2010
rect 1782 -2022 1788 -2016
rect 1782 -2028 1788 -2022
rect 1782 -2034 1788 -2028
rect 1782 -2040 1788 -2034
rect 1782 -2046 1788 -2040
rect 1782 -2052 1788 -2046
rect 1782 -2058 1788 -2052
rect 1782 -2064 1788 -2058
rect 1782 -2070 1788 -2064
rect 1782 -2076 1788 -2070
rect 1782 -2082 1788 -2076
rect 1782 -2088 1788 -2082
rect 1782 -2094 1788 -2088
rect 1782 -2100 1788 -2094
rect 1782 -2106 1788 -2100
rect 1782 -2112 1788 -2106
rect 1782 -2118 1788 -2112
rect 1782 -2124 1788 -2118
rect 1782 -2130 1788 -2124
rect 1782 -2136 1788 -2130
rect 1782 -2142 1788 -2136
rect 1782 -2148 1788 -2142
rect 1782 -2154 1788 -2148
rect 1782 -2160 1788 -2154
rect 1782 -2166 1788 -2160
rect 1782 -2172 1788 -2166
rect 1782 -2178 1788 -2172
rect 1782 -2184 1788 -2178
rect 1782 -2190 1788 -2184
rect 1782 -2196 1788 -2190
rect 1782 -2202 1788 -2196
rect 1782 -2208 1788 -2202
rect 1782 -2214 1788 -2208
rect 1782 -2220 1788 -2214
rect 1782 -2226 1788 -2220
rect 1782 -2232 1788 -2226
rect 1782 -2238 1788 -2232
rect 1782 -2244 1788 -2238
rect 1782 -2250 1788 -2244
rect 1782 -2256 1788 -2250
rect 1782 -2262 1788 -2256
rect 1782 -2268 1788 -2262
rect 1782 -2274 1788 -2268
rect 1782 -2280 1788 -2274
rect 1782 -2286 1788 -2280
rect 1782 -2292 1788 -2286
rect 1782 -2298 1788 -2292
rect 1782 -2304 1788 -2298
rect 1782 -2310 1788 -2304
rect 1782 -2316 1788 -2310
rect 1782 -2322 1788 -2316
rect 1782 -2328 1788 -2322
rect 1782 -2334 1788 -2328
rect 1782 -2340 1788 -2334
rect 1782 -2346 1788 -2340
rect 1782 -2352 1788 -2346
rect 1782 -2358 1788 -2352
rect 1782 -2364 1788 -2358
rect 1782 -2370 1788 -2364
rect 1782 -2376 1788 -2370
rect 1782 -2382 1788 -2376
rect 1782 -2388 1788 -2382
rect 1782 -2394 1788 -2388
rect 1782 -2400 1788 -2394
rect 1782 -2406 1788 -2400
rect 1782 -2412 1788 -2406
rect 1782 -2418 1788 -2412
rect 1782 -2424 1788 -2418
rect 1782 -2430 1788 -2424
rect 1782 -2436 1788 -2430
rect 1782 -2442 1788 -2436
rect 1782 -2448 1788 -2442
rect 1782 -2454 1788 -2448
rect 1782 -2460 1788 -2454
rect 1782 -2466 1788 -2460
rect 1782 -2472 1788 -2466
rect 1782 -2478 1788 -2472
rect 1782 -2484 1788 -2478
rect 1782 -2490 1788 -2484
rect 1782 -2496 1788 -2490
rect 1782 -2502 1788 -2496
rect 1782 -2508 1788 -2502
rect 1782 -2514 1788 -2508
rect 1782 -2520 1788 -2514
rect 1782 -2526 1788 -2520
rect 1782 -2532 1788 -2526
rect 1782 -2538 1788 -2532
rect 1782 -2544 1788 -2538
rect 1782 -2550 1788 -2544
rect 1782 -2556 1788 -2550
rect 1782 -2562 1788 -2556
rect 1782 -2568 1788 -2562
rect 1782 -2574 1788 -2568
rect 1782 -2580 1788 -2574
rect 1782 -2586 1788 -2580
rect 1782 -2592 1788 -2586
rect 1782 -2598 1788 -2592
rect 1782 -2604 1788 -2598
rect 1782 -2610 1788 -2604
rect 1782 -2616 1788 -2610
rect 1782 -2622 1788 -2616
rect 1782 -2628 1788 -2622
rect 1782 -2634 1788 -2628
rect 1782 -2640 1788 -2634
rect 1782 -2718 1788 -2712
rect 1782 -2724 1788 -2718
rect 1782 -2730 1788 -2724
rect 1782 -2736 1788 -2730
rect 1782 -2742 1788 -2736
rect 1782 -2748 1788 -2742
rect 1782 -2754 1788 -2748
rect 1782 -2760 1788 -2754
rect 1782 -2766 1788 -2760
rect 1782 -2772 1788 -2766
rect 1782 -2778 1788 -2772
rect 1782 -2784 1788 -2778
rect 1782 -2790 1788 -2784
rect 1782 -2796 1788 -2790
rect 1782 -2802 1788 -2796
rect 1782 -2808 1788 -2802
rect 1782 -2814 1788 -2808
rect 1782 -2820 1788 -2814
rect 1782 -2826 1788 -2820
rect 1782 -2832 1788 -2826
rect 1782 -2838 1788 -2832
rect 1782 -2844 1788 -2838
rect 1782 -2850 1788 -2844
rect 1782 -2856 1788 -2850
rect 1782 -2862 1788 -2856
rect 1782 -2868 1788 -2862
rect 1782 -2874 1788 -2868
rect 1782 -2880 1788 -2874
rect 1782 -2886 1788 -2880
rect 1782 -2892 1788 -2886
rect 1782 -2898 1788 -2892
rect 1782 -2904 1788 -2898
rect 1782 -2910 1788 -2904
rect 1782 -2916 1788 -2910
rect 1782 -2922 1788 -2916
rect 1782 -2928 1788 -2922
rect 1782 -2934 1788 -2928
rect 1782 -2940 1788 -2934
rect 1782 -2946 1788 -2940
rect 1782 -2952 1788 -2946
rect 1782 -2958 1788 -2952
rect 1782 -2964 1788 -2958
rect 1782 -2970 1788 -2964
rect 1782 -2976 1788 -2970
rect 1782 -2982 1788 -2976
rect 1782 -2988 1788 -2982
rect 1782 -2994 1788 -2988
rect 1782 -3000 1788 -2994
rect 1782 -3006 1788 -3000
rect 1782 -3012 1788 -3006
rect 1782 -3018 1788 -3012
rect 1782 -3024 1788 -3018
rect 1782 -3030 1788 -3024
rect 1782 -3036 1788 -3030
rect 1782 -3042 1788 -3036
rect 1782 -3048 1788 -3042
rect 1782 -3054 1788 -3048
rect 1782 -3060 1788 -3054
rect 1782 -3066 1788 -3060
rect 1782 -3072 1788 -3066
rect 1782 -3078 1788 -3072
rect 1782 -3084 1788 -3078
rect 1782 -3090 1788 -3084
rect 1782 -3096 1788 -3090
rect 1782 -3102 1788 -3096
rect 1782 -3108 1788 -3102
rect 1782 -3114 1788 -3108
rect 1782 -3120 1788 -3114
rect 1782 -3126 1788 -3120
rect 1782 -3132 1788 -3126
rect 1782 -3138 1788 -3132
rect 1782 -3144 1788 -3138
rect 1782 -3150 1788 -3144
rect 1782 -3156 1788 -3150
rect 1782 -3162 1788 -3156
rect 1782 -3168 1788 -3162
rect 1782 -3174 1788 -3168
rect 1782 -3180 1788 -3174
rect 1782 -3186 1788 -3180
rect 1782 -3192 1788 -3186
rect 1782 -3240 1788 -3234
rect 1782 -3246 1788 -3240
rect 1782 -3252 1788 -3246
rect 1782 -3258 1788 -3252
rect 1782 -3264 1788 -3258
rect 1782 -3270 1788 -3264
rect 1782 -3276 1788 -3270
rect 1782 -3282 1788 -3276
rect 1782 -3288 1788 -3282
rect 1782 -3294 1788 -3288
rect 1782 -3300 1788 -3294
rect 1782 -3306 1788 -3300
rect 1782 -3312 1788 -3306
rect 1782 -3318 1788 -3312
rect 1782 -3324 1788 -3318
rect 1782 -3330 1788 -3324
rect 1782 -3336 1788 -3330
rect 1782 -3342 1788 -3336
rect 1782 -3348 1788 -3342
rect 1782 -3354 1788 -3348
rect 1782 -3360 1788 -3354
rect 1782 -3366 1788 -3360
rect 1782 -3372 1788 -3366
rect 1782 -3378 1788 -3372
rect 1788 -738 1794 -732
rect 1788 -744 1794 -738
rect 1788 -750 1794 -744
rect 1788 -756 1794 -750
rect 1788 -762 1794 -756
rect 1788 -768 1794 -762
rect 1788 -774 1794 -768
rect 1788 -780 1794 -774
rect 1788 -786 1794 -780
rect 1788 -792 1794 -786
rect 1788 -798 1794 -792
rect 1788 -804 1794 -798
rect 1788 -810 1794 -804
rect 1788 -816 1794 -810
rect 1788 -822 1794 -816
rect 1788 -828 1794 -822
rect 1788 -834 1794 -828
rect 1788 -840 1794 -834
rect 1788 -846 1794 -840
rect 1788 -852 1794 -846
rect 1788 -858 1794 -852
rect 1788 -864 1794 -858
rect 1788 -870 1794 -864
rect 1788 -876 1794 -870
rect 1788 -882 1794 -876
rect 1788 -888 1794 -882
rect 1788 -894 1794 -888
rect 1788 -900 1794 -894
rect 1788 -906 1794 -900
rect 1788 -912 1794 -906
rect 1788 -918 1794 -912
rect 1788 -924 1794 -918
rect 1788 -930 1794 -924
rect 1788 -936 1794 -930
rect 1788 -942 1794 -936
rect 1788 -948 1794 -942
rect 1788 -954 1794 -948
rect 1788 -960 1794 -954
rect 1788 -966 1794 -960
rect 1788 -972 1794 -966
rect 1788 -978 1794 -972
rect 1788 -984 1794 -978
rect 1788 -990 1794 -984
rect 1788 -996 1794 -990
rect 1788 -1002 1794 -996
rect 1788 -1008 1794 -1002
rect 1788 -1014 1794 -1008
rect 1788 -1020 1794 -1014
rect 1788 -1026 1794 -1020
rect 1788 -1032 1794 -1026
rect 1788 -1038 1794 -1032
rect 1788 -1044 1794 -1038
rect 1788 -1050 1794 -1044
rect 1788 -1056 1794 -1050
rect 1788 -1062 1794 -1056
rect 1788 -1068 1794 -1062
rect 1788 -1074 1794 -1068
rect 1788 -1080 1794 -1074
rect 1788 -1086 1794 -1080
rect 1788 -1092 1794 -1086
rect 1788 -1098 1794 -1092
rect 1788 -1104 1794 -1098
rect 1788 -1110 1794 -1104
rect 1788 -1116 1794 -1110
rect 1788 -1122 1794 -1116
rect 1788 -1128 1794 -1122
rect 1788 -1134 1794 -1128
rect 1788 -1140 1794 -1134
rect 1788 -1146 1794 -1140
rect 1788 -1152 1794 -1146
rect 1788 -1158 1794 -1152
rect 1788 -1164 1794 -1158
rect 1788 -1170 1794 -1164
rect 1788 -1176 1794 -1170
rect 1788 -1182 1794 -1176
rect 1788 -1188 1794 -1182
rect 1788 -1194 1794 -1188
rect 1788 -1200 1794 -1194
rect 1788 -1206 1794 -1200
rect 1788 -1212 1794 -1206
rect 1788 -1218 1794 -1212
rect 1788 -1224 1794 -1218
rect 1788 -1230 1794 -1224
rect 1788 -1236 1794 -1230
rect 1788 -1242 1794 -1236
rect 1788 -1248 1794 -1242
rect 1788 -1254 1794 -1248
rect 1788 -1260 1794 -1254
rect 1788 -1266 1794 -1260
rect 1788 -1272 1794 -1266
rect 1788 -1278 1794 -1272
rect 1788 -1284 1794 -1278
rect 1788 -1290 1794 -1284
rect 1788 -1296 1794 -1290
rect 1788 -1302 1794 -1296
rect 1788 -1308 1794 -1302
rect 1788 -1314 1794 -1308
rect 1788 -1320 1794 -1314
rect 1788 -1326 1794 -1320
rect 1788 -1332 1794 -1326
rect 1788 -1338 1794 -1332
rect 1788 -1344 1794 -1338
rect 1788 -1350 1794 -1344
rect 1788 -1356 1794 -1350
rect 1788 -1362 1794 -1356
rect 1788 -1368 1794 -1362
rect 1788 -1374 1794 -1368
rect 1788 -1380 1794 -1374
rect 1788 -1386 1794 -1380
rect 1788 -1392 1794 -1386
rect 1788 -1398 1794 -1392
rect 1788 -1404 1794 -1398
rect 1788 -1410 1794 -1404
rect 1788 -1416 1794 -1410
rect 1788 -1422 1794 -1416
rect 1788 -1428 1794 -1422
rect 1788 -1434 1794 -1428
rect 1788 -1440 1794 -1434
rect 1788 -1446 1794 -1440
rect 1788 -1452 1794 -1446
rect 1788 -1458 1794 -1452
rect 1788 -1464 1794 -1458
rect 1788 -1470 1794 -1464
rect 1788 -1476 1794 -1470
rect 1788 -1482 1794 -1476
rect 1788 -1488 1794 -1482
rect 1788 -1494 1794 -1488
rect 1788 -1500 1794 -1494
rect 1788 -1506 1794 -1500
rect 1788 -1512 1794 -1506
rect 1788 -1518 1794 -1512
rect 1788 -1524 1794 -1518
rect 1788 -1530 1794 -1524
rect 1788 -1536 1794 -1530
rect 1788 -1542 1794 -1536
rect 1788 -1548 1794 -1542
rect 1788 -1554 1794 -1548
rect 1788 -1560 1794 -1554
rect 1788 -1566 1794 -1560
rect 1788 -1572 1794 -1566
rect 1788 -1578 1794 -1572
rect 1788 -1584 1794 -1578
rect 1788 -1590 1794 -1584
rect 1788 -1596 1794 -1590
rect 1788 -1602 1794 -1596
rect 1788 -1608 1794 -1602
rect 1788 -1614 1794 -1608
rect 1788 -1620 1794 -1614
rect 1788 -1626 1794 -1620
rect 1788 -1632 1794 -1626
rect 1788 -1638 1794 -1632
rect 1788 -1644 1794 -1638
rect 1788 -1650 1794 -1644
rect 1788 -1656 1794 -1650
rect 1788 -1662 1794 -1656
rect 1788 -1668 1794 -1662
rect 1788 -1674 1794 -1668
rect 1788 -1680 1794 -1674
rect 1788 -1686 1794 -1680
rect 1788 -1692 1794 -1686
rect 1788 -1698 1794 -1692
rect 1788 -1704 1794 -1698
rect 1788 -1710 1794 -1704
rect 1788 -1716 1794 -1710
rect 1788 -1722 1794 -1716
rect 1788 -1728 1794 -1722
rect 1788 -1734 1794 -1728
rect 1788 -1740 1794 -1734
rect 1788 -1746 1794 -1740
rect 1788 -1752 1794 -1746
rect 1788 -1758 1794 -1752
rect 1788 -1764 1794 -1758
rect 1788 -1770 1794 -1764
rect 1788 -1776 1794 -1770
rect 1788 -1782 1794 -1776
rect 1788 -1788 1794 -1782
rect 1788 -1794 1794 -1788
rect 1788 -1800 1794 -1794
rect 1788 -1806 1794 -1800
rect 1788 -1812 1794 -1806
rect 1788 -1818 1794 -1812
rect 1788 -1824 1794 -1818
rect 1788 -1830 1794 -1824
rect 1788 -1836 1794 -1830
rect 1788 -1842 1794 -1836
rect 1788 -1848 1794 -1842
rect 1788 -1854 1794 -1848
rect 1788 -1860 1794 -1854
rect 1788 -1938 1794 -1932
rect 1788 -1944 1794 -1938
rect 1788 -1950 1794 -1944
rect 1788 -1956 1794 -1950
rect 1788 -1962 1794 -1956
rect 1788 -1968 1794 -1962
rect 1788 -1974 1794 -1968
rect 1788 -1980 1794 -1974
rect 1788 -1986 1794 -1980
rect 1788 -1992 1794 -1986
rect 1788 -1998 1794 -1992
rect 1788 -2004 1794 -1998
rect 1788 -2010 1794 -2004
rect 1788 -2016 1794 -2010
rect 1788 -2022 1794 -2016
rect 1788 -2028 1794 -2022
rect 1788 -2034 1794 -2028
rect 1788 -2040 1794 -2034
rect 1788 -2046 1794 -2040
rect 1788 -2052 1794 -2046
rect 1788 -2058 1794 -2052
rect 1788 -2064 1794 -2058
rect 1788 -2070 1794 -2064
rect 1788 -2076 1794 -2070
rect 1788 -2082 1794 -2076
rect 1788 -2088 1794 -2082
rect 1788 -2094 1794 -2088
rect 1788 -2100 1794 -2094
rect 1788 -2106 1794 -2100
rect 1788 -2112 1794 -2106
rect 1788 -2118 1794 -2112
rect 1788 -2124 1794 -2118
rect 1788 -2130 1794 -2124
rect 1788 -2136 1794 -2130
rect 1788 -2142 1794 -2136
rect 1788 -2148 1794 -2142
rect 1788 -2154 1794 -2148
rect 1788 -2160 1794 -2154
rect 1788 -2166 1794 -2160
rect 1788 -2172 1794 -2166
rect 1788 -2178 1794 -2172
rect 1788 -2184 1794 -2178
rect 1788 -2190 1794 -2184
rect 1788 -2196 1794 -2190
rect 1788 -2202 1794 -2196
rect 1788 -2208 1794 -2202
rect 1788 -2214 1794 -2208
rect 1788 -2220 1794 -2214
rect 1788 -2226 1794 -2220
rect 1788 -2232 1794 -2226
rect 1788 -2238 1794 -2232
rect 1788 -2244 1794 -2238
rect 1788 -2250 1794 -2244
rect 1788 -2256 1794 -2250
rect 1788 -2262 1794 -2256
rect 1788 -2268 1794 -2262
rect 1788 -2274 1794 -2268
rect 1788 -2280 1794 -2274
rect 1788 -2286 1794 -2280
rect 1788 -2292 1794 -2286
rect 1788 -2298 1794 -2292
rect 1788 -2304 1794 -2298
rect 1788 -2310 1794 -2304
rect 1788 -2316 1794 -2310
rect 1788 -2322 1794 -2316
rect 1788 -2328 1794 -2322
rect 1788 -2334 1794 -2328
rect 1788 -2340 1794 -2334
rect 1788 -2346 1794 -2340
rect 1788 -2352 1794 -2346
rect 1788 -2358 1794 -2352
rect 1788 -2364 1794 -2358
rect 1788 -2370 1794 -2364
rect 1788 -2376 1794 -2370
rect 1788 -2382 1794 -2376
rect 1788 -2388 1794 -2382
rect 1788 -2394 1794 -2388
rect 1788 -2400 1794 -2394
rect 1788 -2406 1794 -2400
rect 1788 -2412 1794 -2406
rect 1788 -2418 1794 -2412
rect 1788 -2424 1794 -2418
rect 1788 -2430 1794 -2424
rect 1788 -2436 1794 -2430
rect 1788 -2442 1794 -2436
rect 1788 -2448 1794 -2442
rect 1788 -2454 1794 -2448
rect 1788 -2460 1794 -2454
rect 1788 -2466 1794 -2460
rect 1788 -2472 1794 -2466
rect 1788 -2478 1794 -2472
rect 1788 -2484 1794 -2478
rect 1788 -2490 1794 -2484
rect 1788 -2496 1794 -2490
rect 1788 -2502 1794 -2496
rect 1788 -2508 1794 -2502
rect 1788 -2514 1794 -2508
rect 1788 -2520 1794 -2514
rect 1788 -2526 1794 -2520
rect 1788 -2532 1794 -2526
rect 1788 -2538 1794 -2532
rect 1788 -2544 1794 -2538
rect 1788 -2550 1794 -2544
rect 1788 -2556 1794 -2550
rect 1788 -2562 1794 -2556
rect 1788 -2568 1794 -2562
rect 1788 -2574 1794 -2568
rect 1788 -2580 1794 -2574
rect 1788 -2586 1794 -2580
rect 1788 -2592 1794 -2586
rect 1788 -2598 1794 -2592
rect 1788 -2604 1794 -2598
rect 1788 -2610 1794 -2604
rect 1788 -2616 1794 -2610
rect 1788 -2622 1794 -2616
rect 1788 -2628 1794 -2622
rect 1788 -2634 1794 -2628
rect 1788 -2640 1794 -2634
rect 1788 -2712 1794 -2706
rect 1788 -2718 1794 -2712
rect 1788 -2724 1794 -2718
rect 1788 -2730 1794 -2724
rect 1788 -2736 1794 -2730
rect 1788 -2742 1794 -2736
rect 1788 -2748 1794 -2742
rect 1788 -2754 1794 -2748
rect 1788 -2760 1794 -2754
rect 1788 -2766 1794 -2760
rect 1788 -2772 1794 -2766
rect 1788 -2778 1794 -2772
rect 1788 -2784 1794 -2778
rect 1788 -2790 1794 -2784
rect 1788 -2796 1794 -2790
rect 1788 -2802 1794 -2796
rect 1788 -2808 1794 -2802
rect 1788 -2814 1794 -2808
rect 1788 -2820 1794 -2814
rect 1788 -2826 1794 -2820
rect 1788 -2832 1794 -2826
rect 1788 -2838 1794 -2832
rect 1788 -2844 1794 -2838
rect 1788 -2850 1794 -2844
rect 1788 -2856 1794 -2850
rect 1788 -2862 1794 -2856
rect 1788 -2868 1794 -2862
rect 1788 -2874 1794 -2868
rect 1788 -2880 1794 -2874
rect 1788 -2886 1794 -2880
rect 1788 -2892 1794 -2886
rect 1788 -2898 1794 -2892
rect 1788 -2904 1794 -2898
rect 1788 -2910 1794 -2904
rect 1788 -2916 1794 -2910
rect 1788 -2922 1794 -2916
rect 1788 -2928 1794 -2922
rect 1788 -2934 1794 -2928
rect 1788 -2940 1794 -2934
rect 1788 -2946 1794 -2940
rect 1788 -2952 1794 -2946
rect 1788 -2958 1794 -2952
rect 1788 -2964 1794 -2958
rect 1788 -2970 1794 -2964
rect 1788 -2976 1794 -2970
rect 1788 -2982 1794 -2976
rect 1788 -2988 1794 -2982
rect 1788 -2994 1794 -2988
rect 1788 -3000 1794 -2994
rect 1788 -3006 1794 -3000
rect 1788 -3012 1794 -3006
rect 1788 -3018 1794 -3012
rect 1788 -3024 1794 -3018
rect 1788 -3030 1794 -3024
rect 1788 -3036 1794 -3030
rect 1788 -3042 1794 -3036
rect 1788 -3048 1794 -3042
rect 1788 -3054 1794 -3048
rect 1788 -3060 1794 -3054
rect 1788 -3066 1794 -3060
rect 1788 -3072 1794 -3066
rect 1788 -3078 1794 -3072
rect 1788 -3084 1794 -3078
rect 1788 -3090 1794 -3084
rect 1788 -3096 1794 -3090
rect 1788 -3102 1794 -3096
rect 1788 -3108 1794 -3102
rect 1788 -3114 1794 -3108
rect 1788 -3120 1794 -3114
rect 1788 -3126 1794 -3120
rect 1788 -3132 1794 -3126
rect 1788 -3138 1794 -3132
rect 1788 -3144 1794 -3138
rect 1788 -3150 1794 -3144
rect 1788 -3156 1794 -3150
rect 1788 -3162 1794 -3156
rect 1788 -3168 1794 -3162
rect 1788 -3174 1794 -3168
rect 1788 -3180 1794 -3174
rect 1788 -3186 1794 -3180
rect 1788 -3240 1794 -3234
rect 1788 -3246 1794 -3240
rect 1788 -3252 1794 -3246
rect 1788 -3258 1794 -3252
rect 1788 -3264 1794 -3258
rect 1788 -3270 1794 -3264
rect 1788 -3276 1794 -3270
rect 1788 -3282 1794 -3276
rect 1788 -3288 1794 -3282
rect 1788 -3294 1794 -3288
rect 1788 -3300 1794 -3294
rect 1788 -3306 1794 -3300
rect 1788 -3312 1794 -3306
rect 1788 -3318 1794 -3312
rect 1788 -3324 1794 -3318
rect 1788 -3330 1794 -3324
rect 1788 -3336 1794 -3330
rect 1788 -3342 1794 -3336
rect 1788 -3348 1794 -3342
rect 1788 -3354 1794 -3348
rect 1788 -3360 1794 -3354
rect 1788 -3366 1794 -3360
rect 1788 -3372 1794 -3366
rect 1788 -3378 1794 -3372
rect 1794 -726 1800 -720
rect 1794 -732 1800 -726
rect 1794 -738 1800 -732
rect 1794 -744 1800 -738
rect 1794 -750 1800 -744
rect 1794 -756 1800 -750
rect 1794 -762 1800 -756
rect 1794 -768 1800 -762
rect 1794 -774 1800 -768
rect 1794 -780 1800 -774
rect 1794 -786 1800 -780
rect 1794 -792 1800 -786
rect 1794 -798 1800 -792
rect 1794 -804 1800 -798
rect 1794 -810 1800 -804
rect 1794 -816 1800 -810
rect 1794 -822 1800 -816
rect 1794 -828 1800 -822
rect 1794 -834 1800 -828
rect 1794 -840 1800 -834
rect 1794 -846 1800 -840
rect 1794 -852 1800 -846
rect 1794 -858 1800 -852
rect 1794 -864 1800 -858
rect 1794 -870 1800 -864
rect 1794 -876 1800 -870
rect 1794 -882 1800 -876
rect 1794 -888 1800 -882
rect 1794 -894 1800 -888
rect 1794 -900 1800 -894
rect 1794 -906 1800 -900
rect 1794 -912 1800 -906
rect 1794 -918 1800 -912
rect 1794 -924 1800 -918
rect 1794 -930 1800 -924
rect 1794 -936 1800 -930
rect 1794 -942 1800 -936
rect 1794 -948 1800 -942
rect 1794 -954 1800 -948
rect 1794 -960 1800 -954
rect 1794 -966 1800 -960
rect 1794 -972 1800 -966
rect 1794 -978 1800 -972
rect 1794 -984 1800 -978
rect 1794 -990 1800 -984
rect 1794 -996 1800 -990
rect 1794 -1002 1800 -996
rect 1794 -1008 1800 -1002
rect 1794 -1014 1800 -1008
rect 1794 -1020 1800 -1014
rect 1794 -1026 1800 -1020
rect 1794 -1032 1800 -1026
rect 1794 -1038 1800 -1032
rect 1794 -1044 1800 -1038
rect 1794 -1050 1800 -1044
rect 1794 -1056 1800 -1050
rect 1794 -1062 1800 -1056
rect 1794 -1068 1800 -1062
rect 1794 -1074 1800 -1068
rect 1794 -1080 1800 -1074
rect 1794 -1086 1800 -1080
rect 1794 -1092 1800 -1086
rect 1794 -1098 1800 -1092
rect 1794 -1104 1800 -1098
rect 1794 -1110 1800 -1104
rect 1794 -1116 1800 -1110
rect 1794 -1122 1800 -1116
rect 1794 -1128 1800 -1122
rect 1794 -1134 1800 -1128
rect 1794 -1140 1800 -1134
rect 1794 -1146 1800 -1140
rect 1794 -1152 1800 -1146
rect 1794 -1158 1800 -1152
rect 1794 -1164 1800 -1158
rect 1794 -1170 1800 -1164
rect 1794 -1176 1800 -1170
rect 1794 -1182 1800 -1176
rect 1794 -1188 1800 -1182
rect 1794 -1194 1800 -1188
rect 1794 -1200 1800 -1194
rect 1794 -1206 1800 -1200
rect 1794 -1212 1800 -1206
rect 1794 -1218 1800 -1212
rect 1794 -1224 1800 -1218
rect 1794 -1230 1800 -1224
rect 1794 -1236 1800 -1230
rect 1794 -1242 1800 -1236
rect 1794 -1248 1800 -1242
rect 1794 -1254 1800 -1248
rect 1794 -1260 1800 -1254
rect 1794 -1266 1800 -1260
rect 1794 -1272 1800 -1266
rect 1794 -1278 1800 -1272
rect 1794 -1284 1800 -1278
rect 1794 -1290 1800 -1284
rect 1794 -1296 1800 -1290
rect 1794 -1302 1800 -1296
rect 1794 -1308 1800 -1302
rect 1794 -1314 1800 -1308
rect 1794 -1320 1800 -1314
rect 1794 -1326 1800 -1320
rect 1794 -1332 1800 -1326
rect 1794 -1338 1800 -1332
rect 1794 -1344 1800 -1338
rect 1794 -1350 1800 -1344
rect 1794 -1356 1800 -1350
rect 1794 -1362 1800 -1356
rect 1794 -1368 1800 -1362
rect 1794 -1374 1800 -1368
rect 1794 -1380 1800 -1374
rect 1794 -1386 1800 -1380
rect 1794 -1392 1800 -1386
rect 1794 -1398 1800 -1392
rect 1794 -1404 1800 -1398
rect 1794 -1410 1800 -1404
rect 1794 -1416 1800 -1410
rect 1794 -1422 1800 -1416
rect 1794 -1428 1800 -1422
rect 1794 -1434 1800 -1428
rect 1794 -1440 1800 -1434
rect 1794 -1446 1800 -1440
rect 1794 -1452 1800 -1446
rect 1794 -1458 1800 -1452
rect 1794 -1464 1800 -1458
rect 1794 -1470 1800 -1464
rect 1794 -1476 1800 -1470
rect 1794 -1482 1800 -1476
rect 1794 -1488 1800 -1482
rect 1794 -1494 1800 -1488
rect 1794 -1500 1800 -1494
rect 1794 -1506 1800 -1500
rect 1794 -1512 1800 -1506
rect 1794 -1518 1800 -1512
rect 1794 -1524 1800 -1518
rect 1794 -1530 1800 -1524
rect 1794 -1536 1800 -1530
rect 1794 -1542 1800 -1536
rect 1794 -1548 1800 -1542
rect 1794 -1554 1800 -1548
rect 1794 -1560 1800 -1554
rect 1794 -1566 1800 -1560
rect 1794 -1572 1800 -1566
rect 1794 -1578 1800 -1572
rect 1794 -1584 1800 -1578
rect 1794 -1590 1800 -1584
rect 1794 -1596 1800 -1590
rect 1794 -1602 1800 -1596
rect 1794 -1608 1800 -1602
rect 1794 -1614 1800 -1608
rect 1794 -1620 1800 -1614
rect 1794 -1626 1800 -1620
rect 1794 -1632 1800 -1626
rect 1794 -1638 1800 -1632
rect 1794 -1644 1800 -1638
rect 1794 -1650 1800 -1644
rect 1794 -1656 1800 -1650
rect 1794 -1662 1800 -1656
rect 1794 -1668 1800 -1662
rect 1794 -1674 1800 -1668
rect 1794 -1680 1800 -1674
rect 1794 -1686 1800 -1680
rect 1794 -1692 1800 -1686
rect 1794 -1698 1800 -1692
rect 1794 -1704 1800 -1698
rect 1794 -1710 1800 -1704
rect 1794 -1716 1800 -1710
rect 1794 -1722 1800 -1716
rect 1794 -1728 1800 -1722
rect 1794 -1734 1800 -1728
rect 1794 -1740 1800 -1734
rect 1794 -1746 1800 -1740
rect 1794 -1752 1800 -1746
rect 1794 -1758 1800 -1752
rect 1794 -1764 1800 -1758
rect 1794 -1770 1800 -1764
rect 1794 -1776 1800 -1770
rect 1794 -1782 1800 -1776
rect 1794 -1788 1800 -1782
rect 1794 -1794 1800 -1788
rect 1794 -1800 1800 -1794
rect 1794 -1806 1800 -1800
rect 1794 -1812 1800 -1806
rect 1794 -1818 1800 -1812
rect 1794 -1824 1800 -1818
rect 1794 -1830 1800 -1824
rect 1794 -1836 1800 -1830
rect 1794 -1842 1800 -1836
rect 1794 -1848 1800 -1842
rect 1794 -1854 1800 -1848
rect 1794 -1932 1800 -1926
rect 1794 -1938 1800 -1932
rect 1794 -1944 1800 -1938
rect 1794 -1950 1800 -1944
rect 1794 -1956 1800 -1950
rect 1794 -1962 1800 -1956
rect 1794 -1968 1800 -1962
rect 1794 -1974 1800 -1968
rect 1794 -1980 1800 -1974
rect 1794 -1986 1800 -1980
rect 1794 -1992 1800 -1986
rect 1794 -1998 1800 -1992
rect 1794 -2004 1800 -1998
rect 1794 -2010 1800 -2004
rect 1794 -2016 1800 -2010
rect 1794 -2022 1800 -2016
rect 1794 -2028 1800 -2022
rect 1794 -2034 1800 -2028
rect 1794 -2040 1800 -2034
rect 1794 -2046 1800 -2040
rect 1794 -2052 1800 -2046
rect 1794 -2058 1800 -2052
rect 1794 -2064 1800 -2058
rect 1794 -2070 1800 -2064
rect 1794 -2076 1800 -2070
rect 1794 -2082 1800 -2076
rect 1794 -2088 1800 -2082
rect 1794 -2094 1800 -2088
rect 1794 -2100 1800 -2094
rect 1794 -2106 1800 -2100
rect 1794 -2112 1800 -2106
rect 1794 -2118 1800 -2112
rect 1794 -2124 1800 -2118
rect 1794 -2130 1800 -2124
rect 1794 -2136 1800 -2130
rect 1794 -2142 1800 -2136
rect 1794 -2148 1800 -2142
rect 1794 -2154 1800 -2148
rect 1794 -2160 1800 -2154
rect 1794 -2166 1800 -2160
rect 1794 -2172 1800 -2166
rect 1794 -2178 1800 -2172
rect 1794 -2184 1800 -2178
rect 1794 -2190 1800 -2184
rect 1794 -2196 1800 -2190
rect 1794 -2202 1800 -2196
rect 1794 -2208 1800 -2202
rect 1794 -2214 1800 -2208
rect 1794 -2220 1800 -2214
rect 1794 -2226 1800 -2220
rect 1794 -2232 1800 -2226
rect 1794 -2238 1800 -2232
rect 1794 -2244 1800 -2238
rect 1794 -2250 1800 -2244
rect 1794 -2256 1800 -2250
rect 1794 -2262 1800 -2256
rect 1794 -2268 1800 -2262
rect 1794 -2274 1800 -2268
rect 1794 -2280 1800 -2274
rect 1794 -2286 1800 -2280
rect 1794 -2292 1800 -2286
rect 1794 -2298 1800 -2292
rect 1794 -2304 1800 -2298
rect 1794 -2310 1800 -2304
rect 1794 -2316 1800 -2310
rect 1794 -2322 1800 -2316
rect 1794 -2328 1800 -2322
rect 1794 -2334 1800 -2328
rect 1794 -2340 1800 -2334
rect 1794 -2346 1800 -2340
rect 1794 -2352 1800 -2346
rect 1794 -2358 1800 -2352
rect 1794 -2364 1800 -2358
rect 1794 -2370 1800 -2364
rect 1794 -2376 1800 -2370
rect 1794 -2382 1800 -2376
rect 1794 -2388 1800 -2382
rect 1794 -2394 1800 -2388
rect 1794 -2400 1800 -2394
rect 1794 -2406 1800 -2400
rect 1794 -2412 1800 -2406
rect 1794 -2418 1800 -2412
rect 1794 -2424 1800 -2418
rect 1794 -2430 1800 -2424
rect 1794 -2436 1800 -2430
rect 1794 -2442 1800 -2436
rect 1794 -2448 1800 -2442
rect 1794 -2454 1800 -2448
rect 1794 -2460 1800 -2454
rect 1794 -2466 1800 -2460
rect 1794 -2472 1800 -2466
rect 1794 -2478 1800 -2472
rect 1794 -2484 1800 -2478
rect 1794 -2490 1800 -2484
rect 1794 -2496 1800 -2490
rect 1794 -2502 1800 -2496
rect 1794 -2508 1800 -2502
rect 1794 -2514 1800 -2508
rect 1794 -2520 1800 -2514
rect 1794 -2526 1800 -2520
rect 1794 -2532 1800 -2526
rect 1794 -2538 1800 -2532
rect 1794 -2544 1800 -2538
rect 1794 -2550 1800 -2544
rect 1794 -2556 1800 -2550
rect 1794 -2562 1800 -2556
rect 1794 -2568 1800 -2562
rect 1794 -2574 1800 -2568
rect 1794 -2580 1800 -2574
rect 1794 -2586 1800 -2580
rect 1794 -2592 1800 -2586
rect 1794 -2598 1800 -2592
rect 1794 -2604 1800 -2598
rect 1794 -2610 1800 -2604
rect 1794 -2616 1800 -2610
rect 1794 -2622 1800 -2616
rect 1794 -2628 1800 -2622
rect 1794 -2634 1800 -2628
rect 1794 -2712 1800 -2706
rect 1794 -2718 1800 -2712
rect 1794 -2724 1800 -2718
rect 1794 -2730 1800 -2724
rect 1794 -2736 1800 -2730
rect 1794 -2742 1800 -2736
rect 1794 -2748 1800 -2742
rect 1794 -2754 1800 -2748
rect 1794 -2760 1800 -2754
rect 1794 -2766 1800 -2760
rect 1794 -2772 1800 -2766
rect 1794 -2778 1800 -2772
rect 1794 -2784 1800 -2778
rect 1794 -2790 1800 -2784
rect 1794 -2796 1800 -2790
rect 1794 -2802 1800 -2796
rect 1794 -2808 1800 -2802
rect 1794 -2814 1800 -2808
rect 1794 -2820 1800 -2814
rect 1794 -2826 1800 -2820
rect 1794 -2832 1800 -2826
rect 1794 -2838 1800 -2832
rect 1794 -2844 1800 -2838
rect 1794 -2850 1800 -2844
rect 1794 -2856 1800 -2850
rect 1794 -2862 1800 -2856
rect 1794 -2868 1800 -2862
rect 1794 -2874 1800 -2868
rect 1794 -2880 1800 -2874
rect 1794 -2886 1800 -2880
rect 1794 -2892 1800 -2886
rect 1794 -2898 1800 -2892
rect 1794 -2904 1800 -2898
rect 1794 -2910 1800 -2904
rect 1794 -2916 1800 -2910
rect 1794 -2922 1800 -2916
rect 1794 -2928 1800 -2922
rect 1794 -2934 1800 -2928
rect 1794 -2940 1800 -2934
rect 1794 -2946 1800 -2940
rect 1794 -2952 1800 -2946
rect 1794 -2958 1800 -2952
rect 1794 -2964 1800 -2958
rect 1794 -2970 1800 -2964
rect 1794 -2976 1800 -2970
rect 1794 -2982 1800 -2976
rect 1794 -2988 1800 -2982
rect 1794 -2994 1800 -2988
rect 1794 -3000 1800 -2994
rect 1794 -3006 1800 -3000
rect 1794 -3012 1800 -3006
rect 1794 -3018 1800 -3012
rect 1794 -3024 1800 -3018
rect 1794 -3030 1800 -3024
rect 1794 -3036 1800 -3030
rect 1794 -3042 1800 -3036
rect 1794 -3048 1800 -3042
rect 1794 -3054 1800 -3048
rect 1794 -3060 1800 -3054
rect 1794 -3066 1800 -3060
rect 1794 -3072 1800 -3066
rect 1794 -3078 1800 -3072
rect 1794 -3084 1800 -3078
rect 1794 -3090 1800 -3084
rect 1794 -3096 1800 -3090
rect 1794 -3102 1800 -3096
rect 1794 -3108 1800 -3102
rect 1794 -3114 1800 -3108
rect 1794 -3120 1800 -3114
rect 1794 -3126 1800 -3120
rect 1794 -3132 1800 -3126
rect 1794 -3138 1800 -3132
rect 1794 -3144 1800 -3138
rect 1794 -3150 1800 -3144
rect 1794 -3156 1800 -3150
rect 1794 -3162 1800 -3156
rect 1794 -3168 1800 -3162
rect 1794 -3174 1800 -3168
rect 1794 -3180 1800 -3174
rect 1794 -3186 1800 -3180
rect 1794 -3234 1800 -3228
rect 1794 -3240 1800 -3234
rect 1794 -3246 1800 -3240
rect 1794 -3252 1800 -3246
rect 1794 -3258 1800 -3252
rect 1794 -3264 1800 -3258
rect 1794 -3270 1800 -3264
rect 1794 -3276 1800 -3270
rect 1794 -3282 1800 -3276
rect 1794 -3288 1800 -3282
rect 1794 -3294 1800 -3288
rect 1794 -3300 1800 -3294
rect 1794 -3306 1800 -3300
rect 1794 -3312 1800 -3306
rect 1794 -3318 1800 -3312
rect 1794 -3324 1800 -3318
rect 1794 -3330 1800 -3324
rect 1794 -3336 1800 -3330
rect 1794 -3342 1800 -3336
rect 1794 -3348 1800 -3342
rect 1794 -3354 1800 -3348
rect 1794 -3360 1800 -3354
rect 1794 -3366 1800 -3360
rect 1794 -3372 1800 -3366
rect 1800 -720 1806 -714
rect 1800 -726 1806 -720
rect 1800 -732 1806 -726
rect 1800 -738 1806 -732
rect 1800 -744 1806 -738
rect 1800 -750 1806 -744
rect 1800 -756 1806 -750
rect 1800 -762 1806 -756
rect 1800 -768 1806 -762
rect 1800 -774 1806 -768
rect 1800 -780 1806 -774
rect 1800 -786 1806 -780
rect 1800 -792 1806 -786
rect 1800 -798 1806 -792
rect 1800 -804 1806 -798
rect 1800 -810 1806 -804
rect 1800 -816 1806 -810
rect 1800 -822 1806 -816
rect 1800 -828 1806 -822
rect 1800 -834 1806 -828
rect 1800 -840 1806 -834
rect 1800 -846 1806 -840
rect 1800 -852 1806 -846
rect 1800 -858 1806 -852
rect 1800 -864 1806 -858
rect 1800 -870 1806 -864
rect 1800 -876 1806 -870
rect 1800 -882 1806 -876
rect 1800 -888 1806 -882
rect 1800 -894 1806 -888
rect 1800 -900 1806 -894
rect 1800 -906 1806 -900
rect 1800 -912 1806 -906
rect 1800 -918 1806 -912
rect 1800 -924 1806 -918
rect 1800 -930 1806 -924
rect 1800 -936 1806 -930
rect 1800 -942 1806 -936
rect 1800 -948 1806 -942
rect 1800 -954 1806 -948
rect 1800 -960 1806 -954
rect 1800 -966 1806 -960
rect 1800 -972 1806 -966
rect 1800 -978 1806 -972
rect 1800 -984 1806 -978
rect 1800 -990 1806 -984
rect 1800 -996 1806 -990
rect 1800 -1002 1806 -996
rect 1800 -1008 1806 -1002
rect 1800 -1014 1806 -1008
rect 1800 -1020 1806 -1014
rect 1800 -1026 1806 -1020
rect 1800 -1032 1806 -1026
rect 1800 -1038 1806 -1032
rect 1800 -1044 1806 -1038
rect 1800 -1050 1806 -1044
rect 1800 -1056 1806 -1050
rect 1800 -1062 1806 -1056
rect 1800 -1068 1806 -1062
rect 1800 -1074 1806 -1068
rect 1800 -1080 1806 -1074
rect 1800 -1086 1806 -1080
rect 1800 -1092 1806 -1086
rect 1800 -1098 1806 -1092
rect 1800 -1104 1806 -1098
rect 1800 -1110 1806 -1104
rect 1800 -1116 1806 -1110
rect 1800 -1122 1806 -1116
rect 1800 -1128 1806 -1122
rect 1800 -1134 1806 -1128
rect 1800 -1140 1806 -1134
rect 1800 -1146 1806 -1140
rect 1800 -1152 1806 -1146
rect 1800 -1158 1806 -1152
rect 1800 -1164 1806 -1158
rect 1800 -1170 1806 -1164
rect 1800 -1176 1806 -1170
rect 1800 -1182 1806 -1176
rect 1800 -1188 1806 -1182
rect 1800 -1194 1806 -1188
rect 1800 -1200 1806 -1194
rect 1800 -1206 1806 -1200
rect 1800 -1212 1806 -1206
rect 1800 -1218 1806 -1212
rect 1800 -1224 1806 -1218
rect 1800 -1230 1806 -1224
rect 1800 -1236 1806 -1230
rect 1800 -1242 1806 -1236
rect 1800 -1248 1806 -1242
rect 1800 -1254 1806 -1248
rect 1800 -1260 1806 -1254
rect 1800 -1266 1806 -1260
rect 1800 -1272 1806 -1266
rect 1800 -1278 1806 -1272
rect 1800 -1284 1806 -1278
rect 1800 -1290 1806 -1284
rect 1800 -1296 1806 -1290
rect 1800 -1302 1806 -1296
rect 1800 -1308 1806 -1302
rect 1800 -1314 1806 -1308
rect 1800 -1320 1806 -1314
rect 1800 -1326 1806 -1320
rect 1800 -1332 1806 -1326
rect 1800 -1338 1806 -1332
rect 1800 -1344 1806 -1338
rect 1800 -1350 1806 -1344
rect 1800 -1356 1806 -1350
rect 1800 -1362 1806 -1356
rect 1800 -1368 1806 -1362
rect 1800 -1374 1806 -1368
rect 1800 -1380 1806 -1374
rect 1800 -1386 1806 -1380
rect 1800 -1392 1806 -1386
rect 1800 -1398 1806 -1392
rect 1800 -1404 1806 -1398
rect 1800 -1410 1806 -1404
rect 1800 -1416 1806 -1410
rect 1800 -1422 1806 -1416
rect 1800 -1428 1806 -1422
rect 1800 -1434 1806 -1428
rect 1800 -1440 1806 -1434
rect 1800 -1446 1806 -1440
rect 1800 -1452 1806 -1446
rect 1800 -1458 1806 -1452
rect 1800 -1464 1806 -1458
rect 1800 -1470 1806 -1464
rect 1800 -1476 1806 -1470
rect 1800 -1482 1806 -1476
rect 1800 -1488 1806 -1482
rect 1800 -1494 1806 -1488
rect 1800 -1500 1806 -1494
rect 1800 -1506 1806 -1500
rect 1800 -1512 1806 -1506
rect 1800 -1518 1806 -1512
rect 1800 -1524 1806 -1518
rect 1800 -1530 1806 -1524
rect 1800 -1536 1806 -1530
rect 1800 -1542 1806 -1536
rect 1800 -1548 1806 -1542
rect 1800 -1554 1806 -1548
rect 1800 -1560 1806 -1554
rect 1800 -1566 1806 -1560
rect 1800 -1572 1806 -1566
rect 1800 -1578 1806 -1572
rect 1800 -1584 1806 -1578
rect 1800 -1590 1806 -1584
rect 1800 -1596 1806 -1590
rect 1800 -1602 1806 -1596
rect 1800 -1608 1806 -1602
rect 1800 -1614 1806 -1608
rect 1800 -1620 1806 -1614
rect 1800 -1626 1806 -1620
rect 1800 -1632 1806 -1626
rect 1800 -1638 1806 -1632
rect 1800 -1644 1806 -1638
rect 1800 -1650 1806 -1644
rect 1800 -1656 1806 -1650
rect 1800 -1662 1806 -1656
rect 1800 -1668 1806 -1662
rect 1800 -1674 1806 -1668
rect 1800 -1680 1806 -1674
rect 1800 -1686 1806 -1680
rect 1800 -1692 1806 -1686
rect 1800 -1698 1806 -1692
rect 1800 -1704 1806 -1698
rect 1800 -1710 1806 -1704
rect 1800 -1716 1806 -1710
rect 1800 -1722 1806 -1716
rect 1800 -1728 1806 -1722
rect 1800 -1734 1806 -1728
rect 1800 -1740 1806 -1734
rect 1800 -1746 1806 -1740
rect 1800 -1752 1806 -1746
rect 1800 -1758 1806 -1752
rect 1800 -1764 1806 -1758
rect 1800 -1770 1806 -1764
rect 1800 -1776 1806 -1770
rect 1800 -1782 1806 -1776
rect 1800 -1788 1806 -1782
rect 1800 -1794 1806 -1788
rect 1800 -1800 1806 -1794
rect 1800 -1806 1806 -1800
rect 1800 -1812 1806 -1806
rect 1800 -1818 1806 -1812
rect 1800 -1824 1806 -1818
rect 1800 -1830 1806 -1824
rect 1800 -1836 1806 -1830
rect 1800 -1842 1806 -1836
rect 1800 -1848 1806 -1842
rect 1800 -1926 1806 -1920
rect 1800 -1932 1806 -1926
rect 1800 -1938 1806 -1932
rect 1800 -1944 1806 -1938
rect 1800 -1950 1806 -1944
rect 1800 -1956 1806 -1950
rect 1800 -1962 1806 -1956
rect 1800 -1968 1806 -1962
rect 1800 -1974 1806 -1968
rect 1800 -1980 1806 -1974
rect 1800 -1986 1806 -1980
rect 1800 -1992 1806 -1986
rect 1800 -1998 1806 -1992
rect 1800 -2004 1806 -1998
rect 1800 -2010 1806 -2004
rect 1800 -2016 1806 -2010
rect 1800 -2022 1806 -2016
rect 1800 -2028 1806 -2022
rect 1800 -2034 1806 -2028
rect 1800 -2040 1806 -2034
rect 1800 -2046 1806 -2040
rect 1800 -2052 1806 -2046
rect 1800 -2058 1806 -2052
rect 1800 -2064 1806 -2058
rect 1800 -2070 1806 -2064
rect 1800 -2076 1806 -2070
rect 1800 -2082 1806 -2076
rect 1800 -2088 1806 -2082
rect 1800 -2094 1806 -2088
rect 1800 -2100 1806 -2094
rect 1800 -2106 1806 -2100
rect 1800 -2112 1806 -2106
rect 1800 -2118 1806 -2112
rect 1800 -2124 1806 -2118
rect 1800 -2130 1806 -2124
rect 1800 -2136 1806 -2130
rect 1800 -2142 1806 -2136
rect 1800 -2148 1806 -2142
rect 1800 -2154 1806 -2148
rect 1800 -2160 1806 -2154
rect 1800 -2166 1806 -2160
rect 1800 -2172 1806 -2166
rect 1800 -2178 1806 -2172
rect 1800 -2184 1806 -2178
rect 1800 -2190 1806 -2184
rect 1800 -2196 1806 -2190
rect 1800 -2202 1806 -2196
rect 1800 -2208 1806 -2202
rect 1800 -2214 1806 -2208
rect 1800 -2220 1806 -2214
rect 1800 -2226 1806 -2220
rect 1800 -2232 1806 -2226
rect 1800 -2238 1806 -2232
rect 1800 -2244 1806 -2238
rect 1800 -2250 1806 -2244
rect 1800 -2256 1806 -2250
rect 1800 -2262 1806 -2256
rect 1800 -2268 1806 -2262
rect 1800 -2274 1806 -2268
rect 1800 -2280 1806 -2274
rect 1800 -2286 1806 -2280
rect 1800 -2292 1806 -2286
rect 1800 -2298 1806 -2292
rect 1800 -2304 1806 -2298
rect 1800 -2310 1806 -2304
rect 1800 -2316 1806 -2310
rect 1800 -2322 1806 -2316
rect 1800 -2328 1806 -2322
rect 1800 -2334 1806 -2328
rect 1800 -2340 1806 -2334
rect 1800 -2346 1806 -2340
rect 1800 -2352 1806 -2346
rect 1800 -2358 1806 -2352
rect 1800 -2364 1806 -2358
rect 1800 -2370 1806 -2364
rect 1800 -2376 1806 -2370
rect 1800 -2382 1806 -2376
rect 1800 -2388 1806 -2382
rect 1800 -2394 1806 -2388
rect 1800 -2400 1806 -2394
rect 1800 -2406 1806 -2400
rect 1800 -2412 1806 -2406
rect 1800 -2418 1806 -2412
rect 1800 -2424 1806 -2418
rect 1800 -2430 1806 -2424
rect 1800 -2436 1806 -2430
rect 1800 -2442 1806 -2436
rect 1800 -2448 1806 -2442
rect 1800 -2454 1806 -2448
rect 1800 -2460 1806 -2454
rect 1800 -2466 1806 -2460
rect 1800 -2472 1806 -2466
rect 1800 -2478 1806 -2472
rect 1800 -2484 1806 -2478
rect 1800 -2490 1806 -2484
rect 1800 -2496 1806 -2490
rect 1800 -2502 1806 -2496
rect 1800 -2508 1806 -2502
rect 1800 -2514 1806 -2508
rect 1800 -2520 1806 -2514
rect 1800 -2526 1806 -2520
rect 1800 -2532 1806 -2526
rect 1800 -2538 1806 -2532
rect 1800 -2544 1806 -2538
rect 1800 -2550 1806 -2544
rect 1800 -2556 1806 -2550
rect 1800 -2562 1806 -2556
rect 1800 -2568 1806 -2562
rect 1800 -2574 1806 -2568
rect 1800 -2580 1806 -2574
rect 1800 -2586 1806 -2580
rect 1800 -2592 1806 -2586
rect 1800 -2598 1806 -2592
rect 1800 -2604 1806 -2598
rect 1800 -2610 1806 -2604
rect 1800 -2616 1806 -2610
rect 1800 -2622 1806 -2616
rect 1800 -2628 1806 -2622
rect 1800 -2634 1806 -2628
rect 1800 -2706 1806 -2700
rect 1800 -2712 1806 -2706
rect 1800 -2718 1806 -2712
rect 1800 -2724 1806 -2718
rect 1800 -2730 1806 -2724
rect 1800 -2736 1806 -2730
rect 1800 -2742 1806 -2736
rect 1800 -2748 1806 -2742
rect 1800 -2754 1806 -2748
rect 1800 -2760 1806 -2754
rect 1800 -2766 1806 -2760
rect 1800 -2772 1806 -2766
rect 1800 -2778 1806 -2772
rect 1800 -2784 1806 -2778
rect 1800 -2790 1806 -2784
rect 1800 -2796 1806 -2790
rect 1800 -2802 1806 -2796
rect 1800 -2808 1806 -2802
rect 1800 -2814 1806 -2808
rect 1800 -2820 1806 -2814
rect 1800 -2826 1806 -2820
rect 1800 -2832 1806 -2826
rect 1800 -2838 1806 -2832
rect 1800 -2844 1806 -2838
rect 1800 -2850 1806 -2844
rect 1800 -2856 1806 -2850
rect 1800 -2862 1806 -2856
rect 1800 -2868 1806 -2862
rect 1800 -2874 1806 -2868
rect 1800 -2880 1806 -2874
rect 1800 -2886 1806 -2880
rect 1800 -2892 1806 -2886
rect 1800 -2898 1806 -2892
rect 1800 -2904 1806 -2898
rect 1800 -2910 1806 -2904
rect 1800 -2916 1806 -2910
rect 1800 -2922 1806 -2916
rect 1800 -2928 1806 -2922
rect 1800 -2934 1806 -2928
rect 1800 -2940 1806 -2934
rect 1800 -2946 1806 -2940
rect 1800 -2952 1806 -2946
rect 1800 -2958 1806 -2952
rect 1800 -2964 1806 -2958
rect 1800 -2970 1806 -2964
rect 1800 -2976 1806 -2970
rect 1800 -2982 1806 -2976
rect 1800 -2988 1806 -2982
rect 1800 -2994 1806 -2988
rect 1800 -3000 1806 -2994
rect 1800 -3006 1806 -3000
rect 1800 -3012 1806 -3006
rect 1800 -3018 1806 -3012
rect 1800 -3024 1806 -3018
rect 1800 -3030 1806 -3024
rect 1800 -3036 1806 -3030
rect 1800 -3042 1806 -3036
rect 1800 -3048 1806 -3042
rect 1800 -3054 1806 -3048
rect 1800 -3060 1806 -3054
rect 1800 -3066 1806 -3060
rect 1800 -3072 1806 -3066
rect 1800 -3078 1806 -3072
rect 1800 -3084 1806 -3078
rect 1800 -3090 1806 -3084
rect 1800 -3096 1806 -3090
rect 1800 -3102 1806 -3096
rect 1800 -3108 1806 -3102
rect 1800 -3114 1806 -3108
rect 1800 -3120 1806 -3114
rect 1800 -3126 1806 -3120
rect 1800 -3132 1806 -3126
rect 1800 -3138 1806 -3132
rect 1800 -3144 1806 -3138
rect 1800 -3150 1806 -3144
rect 1800 -3156 1806 -3150
rect 1800 -3162 1806 -3156
rect 1800 -3168 1806 -3162
rect 1800 -3174 1806 -3168
rect 1800 -3180 1806 -3174
rect 1800 -3234 1806 -3228
rect 1800 -3240 1806 -3234
rect 1800 -3246 1806 -3240
rect 1800 -3252 1806 -3246
rect 1800 -3258 1806 -3252
rect 1800 -3264 1806 -3258
rect 1800 -3270 1806 -3264
rect 1800 -3276 1806 -3270
rect 1800 -3282 1806 -3276
rect 1800 -3288 1806 -3282
rect 1800 -3294 1806 -3288
rect 1800 -3300 1806 -3294
rect 1800 -3306 1806 -3300
rect 1800 -3312 1806 -3306
rect 1800 -3318 1806 -3312
rect 1800 -3324 1806 -3318
rect 1800 -3330 1806 -3324
rect 1800 -3336 1806 -3330
rect 1800 -3342 1806 -3336
rect 1800 -3348 1806 -3342
rect 1800 -3354 1806 -3348
rect 1800 -3360 1806 -3354
rect 1800 -3366 1806 -3360
rect 1806 -714 1812 -708
rect 1806 -720 1812 -714
rect 1806 -726 1812 -720
rect 1806 -732 1812 -726
rect 1806 -738 1812 -732
rect 1806 -744 1812 -738
rect 1806 -750 1812 -744
rect 1806 -756 1812 -750
rect 1806 -762 1812 -756
rect 1806 -768 1812 -762
rect 1806 -774 1812 -768
rect 1806 -780 1812 -774
rect 1806 -786 1812 -780
rect 1806 -792 1812 -786
rect 1806 -798 1812 -792
rect 1806 -804 1812 -798
rect 1806 -810 1812 -804
rect 1806 -816 1812 -810
rect 1806 -822 1812 -816
rect 1806 -828 1812 -822
rect 1806 -834 1812 -828
rect 1806 -840 1812 -834
rect 1806 -846 1812 -840
rect 1806 -852 1812 -846
rect 1806 -858 1812 -852
rect 1806 -864 1812 -858
rect 1806 -870 1812 -864
rect 1806 -876 1812 -870
rect 1806 -882 1812 -876
rect 1806 -888 1812 -882
rect 1806 -894 1812 -888
rect 1806 -900 1812 -894
rect 1806 -906 1812 -900
rect 1806 -912 1812 -906
rect 1806 -918 1812 -912
rect 1806 -924 1812 -918
rect 1806 -930 1812 -924
rect 1806 -936 1812 -930
rect 1806 -942 1812 -936
rect 1806 -948 1812 -942
rect 1806 -954 1812 -948
rect 1806 -960 1812 -954
rect 1806 -966 1812 -960
rect 1806 -972 1812 -966
rect 1806 -978 1812 -972
rect 1806 -984 1812 -978
rect 1806 -990 1812 -984
rect 1806 -996 1812 -990
rect 1806 -1002 1812 -996
rect 1806 -1008 1812 -1002
rect 1806 -1014 1812 -1008
rect 1806 -1020 1812 -1014
rect 1806 -1026 1812 -1020
rect 1806 -1032 1812 -1026
rect 1806 -1038 1812 -1032
rect 1806 -1044 1812 -1038
rect 1806 -1050 1812 -1044
rect 1806 -1056 1812 -1050
rect 1806 -1062 1812 -1056
rect 1806 -1068 1812 -1062
rect 1806 -1074 1812 -1068
rect 1806 -1080 1812 -1074
rect 1806 -1086 1812 -1080
rect 1806 -1092 1812 -1086
rect 1806 -1098 1812 -1092
rect 1806 -1104 1812 -1098
rect 1806 -1110 1812 -1104
rect 1806 -1116 1812 -1110
rect 1806 -1122 1812 -1116
rect 1806 -1128 1812 -1122
rect 1806 -1134 1812 -1128
rect 1806 -1140 1812 -1134
rect 1806 -1146 1812 -1140
rect 1806 -1152 1812 -1146
rect 1806 -1158 1812 -1152
rect 1806 -1164 1812 -1158
rect 1806 -1170 1812 -1164
rect 1806 -1176 1812 -1170
rect 1806 -1182 1812 -1176
rect 1806 -1188 1812 -1182
rect 1806 -1194 1812 -1188
rect 1806 -1200 1812 -1194
rect 1806 -1206 1812 -1200
rect 1806 -1212 1812 -1206
rect 1806 -1218 1812 -1212
rect 1806 -1224 1812 -1218
rect 1806 -1230 1812 -1224
rect 1806 -1236 1812 -1230
rect 1806 -1242 1812 -1236
rect 1806 -1248 1812 -1242
rect 1806 -1254 1812 -1248
rect 1806 -1260 1812 -1254
rect 1806 -1266 1812 -1260
rect 1806 -1272 1812 -1266
rect 1806 -1278 1812 -1272
rect 1806 -1284 1812 -1278
rect 1806 -1290 1812 -1284
rect 1806 -1296 1812 -1290
rect 1806 -1302 1812 -1296
rect 1806 -1308 1812 -1302
rect 1806 -1314 1812 -1308
rect 1806 -1320 1812 -1314
rect 1806 -1326 1812 -1320
rect 1806 -1332 1812 -1326
rect 1806 -1338 1812 -1332
rect 1806 -1344 1812 -1338
rect 1806 -1350 1812 -1344
rect 1806 -1356 1812 -1350
rect 1806 -1362 1812 -1356
rect 1806 -1368 1812 -1362
rect 1806 -1374 1812 -1368
rect 1806 -1380 1812 -1374
rect 1806 -1386 1812 -1380
rect 1806 -1392 1812 -1386
rect 1806 -1398 1812 -1392
rect 1806 -1404 1812 -1398
rect 1806 -1410 1812 -1404
rect 1806 -1416 1812 -1410
rect 1806 -1422 1812 -1416
rect 1806 -1428 1812 -1422
rect 1806 -1434 1812 -1428
rect 1806 -1440 1812 -1434
rect 1806 -1446 1812 -1440
rect 1806 -1452 1812 -1446
rect 1806 -1458 1812 -1452
rect 1806 -1464 1812 -1458
rect 1806 -1470 1812 -1464
rect 1806 -1476 1812 -1470
rect 1806 -1482 1812 -1476
rect 1806 -1488 1812 -1482
rect 1806 -1494 1812 -1488
rect 1806 -1500 1812 -1494
rect 1806 -1506 1812 -1500
rect 1806 -1512 1812 -1506
rect 1806 -1518 1812 -1512
rect 1806 -1524 1812 -1518
rect 1806 -1530 1812 -1524
rect 1806 -1536 1812 -1530
rect 1806 -1542 1812 -1536
rect 1806 -1548 1812 -1542
rect 1806 -1554 1812 -1548
rect 1806 -1560 1812 -1554
rect 1806 -1566 1812 -1560
rect 1806 -1572 1812 -1566
rect 1806 -1578 1812 -1572
rect 1806 -1584 1812 -1578
rect 1806 -1590 1812 -1584
rect 1806 -1596 1812 -1590
rect 1806 -1602 1812 -1596
rect 1806 -1608 1812 -1602
rect 1806 -1614 1812 -1608
rect 1806 -1620 1812 -1614
rect 1806 -1626 1812 -1620
rect 1806 -1632 1812 -1626
rect 1806 -1638 1812 -1632
rect 1806 -1644 1812 -1638
rect 1806 -1650 1812 -1644
rect 1806 -1656 1812 -1650
rect 1806 -1662 1812 -1656
rect 1806 -1668 1812 -1662
rect 1806 -1674 1812 -1668
rect 1806 -1680 1812 -1674
rect 1806 -1686 1812 -1680
rect 1806 -1692 1812 -1686
rect 1806 -1698 1812 -1692
rect 1806 -1704 1812 -1698
rect 1806 -1710 1812 -1704
rect 1806 -1716 1812 -1710
rect 1806 -1722 1812 -1716
rect 1806 -1728 1812 -1722
rect 1806 -1734 1812 -1728
rect 1806 -1740 1812 -1734
rect 1806 -1746 1812 -1740
rect 1806 -1752 1812 -1746
rect 1806 -1758 1812 -1752
rect 1806 -1764 1812 -1758
rect 1806 -1770 1812 -1764
rect 1806 -1776 1812 -1770
rect 1806 -1782 1812 -1776
rect 1806 -1788 1812 -1782
rect 1806 -1794 1812 -1788
rect 1806 -1800 1812 -1794
rect 1806 -1806 1812 -1800
rect 1806 -1812 1812 -1806
rect 1806 -1818 1812 -1812
rect 1806 -1824 1812 -1818
rect 1806 -1830 1812 -1824
rect 1806 -1836 1812 -1830
rect 1806 -1842 1812 -1836
rect 1806 -1920 1812 -1914
rect 1806 -1926 1812 -1920
rect 1806 -1932 1812 -1926
rect 1806 -1938 1812 -1932
rect 1806 -1944 1812 -1938
rect 1806 -1950 1812 -1944
rect 1806 -1956 1812 -1950
rect 1806 -1962 1812 -1956
rect 1806 -1968 1812 -1962
rect 1806 -1974 1812 -1968
rect 1806 -1980 1812 -1974
rect 1806 -1986 1812 -1980
rect 1806 -1992 1812 -1986
rect 1806 -1998 1812 -1992
rect 1806 -2004 1812 -1998
rect 1806 -2010 1812 -2004
rect 1806 -2016 1812 -2010
rect 1806 -2022 1812 -2016
rect 1806 -2028 1812 -2022
rect 1806 -2034 1812 -2028
rect 1806 -2040 1812 -2034
rect 1806 -2046 1812 -2040
rect 1806 -2052 1812 -2046
rect 1806 -2058 1812 -2052
rect 1806 -2064 1812 -2058
rect 1806 -2070 1812 -2064
rect 1806 -2076 1812 -2070
rect 1806 -2082 1812 -2076
rect 1806 -2088 1812 -2082
rect 1806 -2094 1812 -2088
rect 1806 -2100 1812 -2094
rect 1806 -2106 1812 -2100
rect 1806 -2112 1812 -2106
rect 1806 -2118 1812 -2112
rect 1806 -2124 1812 -2118
rect 1806 -2130 1812 -2124
rect 1806 -2136 1812 -2130
rect 1806 -2142 1812 -2136
rect 1806 -2148 1812 -2142
rect 1806 -2154 1812 -2148
rect 1806 -2160 1812 -2154
rect 1806 -2166 1812 -2160
rect 1806 -2172 1812 -2166
rect 1806 -2178 1812 -2172
rect 1806 -2184 1812 -2178
rect 1806 -2190 1812 -2184
rect 1806 -2196 1812 -2190
rect 1806 -2202 1812 -2196
rect 1806 -2208 1812 -2202
rect 1806 -2214 1812 -2208
rect 1806 -2220 1812 -2214
rect 1806 -2226 1812 -2220
rect 1806 -2232 1812 -2226
rect 1806 -2238 1812 -2232
rect 1806 -2244 1812 -2238
rect 1806 -2250 1812 -2244
rect 1806 -2256 1812 -2250
rect 1806 -2262 1812 -2256
rect 1806 -2268 1812 -2262
rect 1806 -2274 1812 -2268
rect 1806 -2280 1812 -2274
rect 1806 -2286 1812 -2280
rect 1806 -2292 1812 -2286
rect 1806 -2298 1812 -2292
rect 1806 -2304 1812 -2298
rect 1806 -2310 1812 -2304
rect 1806 -2316 1812 -2310
rect 1806 -2322 1812 -2316
rect 1806 -2328 1812 -2322
rect 1806 -2334 1812 -2328
rect 1806 -2340 1812 -2334
rect 1806 -2346 1812 -2340
rect 1806 -2352 1812 -2346
rect 1806 -2358 1812 -2352
rect 1806 -2364 1812 -2358
rect 1806 -2370 1812 -2364
rect 1806 -2376 1812 -2370
rect 1806 -2382 1812 -2376
rect 1806 -2388 1812 -2382
rect 1806 -2394 1812 -2388
rect 1806 -2400 1812 -2394
rect 1806 -2406 1812 -2400
rect 1806 -2412 1812 -2406
rect 1806 -2418 1812 -2412
rect 1806 -2424 1812 -2418
rect 1806 -2430 1812 -2424
rect 1806 -2436 1812 -2430
rect 1806 -2442 1812 -2436
rect 1806 -2448 1812 -2442
rect 1806 -2454 1812 -2448
rect 1806 -2460 1812 -2454
rect 1806 -2466 1812 -2460
rect 1806 -2472 1812 -2466
rect 1806 -2478 1812 -2472
rect 1806 -2484 1812 -2478
rect 1806 -2490 1812 -2484
rect 1806 -2496 1812 -2490
rect 1806 -2502 1812 -2496
rect 1806 -2508 1812 -2502
rect 1806 -2514 1812 -2508
rect 1806 -2520 1812 -2514
rect 1806 -2526 1812 -2520
rect 1806 -2532 1812 -2526
rect 1806 -2538 1812 -2532
rect 1806 -2544 1812 -2538
rect 1806 -2550 1812 -2544
rect 1806 -2556 1812 -2550
rect 1806 -2562 1812 -2556
rect 1806 -2568 1812 -2562
rect 1806 -2574 1812 -2568
rect 1806 -2580 1812 -2574
rect 1806 -2586 1812 -2580
rect 1806 -2592 1812 -2586
rect 1806 -2598 1812 -2592
rect 1806 -2604 1812 -2598
rect 1806 -2610 1812 -2604
rect 1806 -2616 1812 -2610
rect 1806 -2622 1812 -2616
rect 1806 -2628 1812 -2622
rect 1806 -2700 1812 -2694
rect 1806 -2706 1812 -2700
rect 1806 -2712 1812 -2706
rect 1806 -2718 1812 -2712
rect 1806 -2724 1812 -2718
rect 1806 -2730 1812 -2724
rect 1806 -2736 1812 -2730
rect 1806 -2742 1812 -2736
rect 1806 -2748 1812 -2742
rect 1806 -2754 1812 -2748
rect 1806 -2760 1812 -2754
rect 1806 -2766 1812 -2760
rect 1806 -2772 1812 -2766
rect 1806 -2778 1812 -2772
rect 1806 -2784 1812 -2778
rect 1806 -2790 1812 -2784
rect 1806 -2796 1812 -2790
rect 1806 -2802 1812 -2796
rect 1806 -2808 1812 -2802
rect 1806 -2814 1812 -2808
rect 1806 -2820 1812 -2814
rect 1806 -2826 1812 -2820
rect 1806 -2832 1812 -2826
rect 1806 -2838 1812 -2832
rect 1806 -2844 1812 -2838
rect 1806 -2850 1812 -2844
rect 1806 -2856 1812 -2850
rect 1806 -2862 1812 -2856
rect 1806 -2868 1812 -2862
rect 1806 -2874 1812 -2868
rect 1806 -2880 1812 -2874
rect 1806 -2886 1812 -2880
rect 1806 -2892 1812 -2886
rect 1806 -2898 1812 -2892
rect 1806 -2904 1812 -2898
rect 1806 -2910 1812 -2904
rect 1806 -2916 1812 -2910
rect 1806 -2922 1812 -2916
rect 1806 -2928 1812 -2922
rect 1806 -2934 1812 -2928
rect 1806 -2940 1812 -2934
rect 1806 -2946 1812 -2940
rect 1806 -2952 1812 -2946
rect 1806 -2958 1812 -2952
rect 1806 -2964 1812 -2958
rect 1806 -2970 1812 -2964
rect 1806 -2976 1812 -2970
rect 1806 -2982 1812 -2976
rect 1806 -2988 1812 -2982
rect 1806 -2994 1812 -2988
rect 1806 -3000 1812 -2994
rect 1806 -3006 1812 -3000
rect 1806 -3012 1812 -3006
rect 1806 -3018 1812 -3012
rect 1806 -3024 1812 -3018
rect 1806 -3030 1812 -3024
rect 1806 -3036 1812 -3030
rect 1806 -3042 1812 -3036
rect 1806 -3048 1812 -3042
rect 1806 -3054 1812 -3048
rect 1806 -3060 1812 -3054
rect 1806 -3066 1812 -3060
rect 1806 -3072 1812 -3066
rect 1806 -3078 1812 -3072
rect 1806 -3084 1812 -3078
rect 1806 -3090 1812 -3084
rect 1806 -3096 1812 -3090
rect 1806 -3102 1812 -3096
rect 1806 -3108 1812 -3102
rect 1806 -3114 1812 -3108
rect 1806 -3120 1812 -3114
rect 1806 -3126 1812 -3120
rect 1806 -3132 1812 -3126
rect 1806 -3138 1812 -3132
rect 1806 -3144 1812 -3138
rect 1806 -3150 1812 -3144
rect 1806 -3156 1812 -3150
rect 1806 -3162 1812 -3156
rect 1806 -3168 1812 -3162
rect 1806 -3174 1812 -3168
rect 1806 -3180 1812 -3174
rect 1806 -3234 1812 -3228
rect 1806 -3240 1812 -3234
rect 1806 -3246 1812 -3240
rect 1806 -3252 1812 -3246
rect 1806 -3258 1812 -3252
rect 1806 -3264 1812 -3258
rect 1806 -3270 1812 -3264
rect 1806 -3276 1812 -3270
rect 1806 -3282 1812 -3276
rect 1806 -3288 1812 -3282
rect 1806 -3294 1812 -3288
rect 1806 -3300 1812 -3294
rect 1806 -3306 1812 -3300
rect 1806 -3312 1812 -3306
rect 1806 -3318 1812 -3312
rect 1806 -3324 1812 -3318
rect 1806 -3330 1812 -3324
rect 1806 -3336 1812 -3330
rect 1806 -3342 1812 -3336
rect 1806 -3348 1812 -3342
rect 1806 -3354 1812 -3348
rect 1806 -3360 1812 -3354
rect 1806 -3366 1812 -3360
rect 1812 -702 1818 -696
rect 1812 -708 1818 -702
rect 1812 -714 1818 -708
rect 1812 -720 1818 -714
rect 1812 -726 1818 -720
rect 1812 -732 1818 -726
rect 1812 -738 1818 -732
rect 1812 -744 1818 -738
rect 1812 -750 1818 -744
rect 1812 -756 1818 -750
rect 1812 -762 1818 -756
rect 1812 -768 1818 -762
rect 1812 -774 1818 -768
rect 1812 -780 1818 -774
rect 1812 -786 1818 -780
rect 1812 -792 1818 -786
rect 1812 -798 1818 -792
rect 1812 -804 1818 -798
rect 1812 -810 1818 -804
rect 1812 -816 1818 -810
rect 1812 -822 1818 -816
rect 1812 -828 1818 -822
rect 1812 -834 1818 -828
rect 1812 -840 1818 -834
rect 1812 -846 1818 -840
rect 1812 -852 1818 -846
rect 1812 -858 1818 -852
rect 1812 -864 1818 -858
rect 1812 -870 1818 -864
rect 1812 -876 1818 -870
rect 1812 -882 1818 -876
rect 1812 -888 1818 -882
rect 1812 -894 1818 -888
rect 1812 -900 1818 -894
rect 1812 -906 1818 -900
rect 1812 -912 1818 -906
rect 1812 -918 1818 -912
rect 1812 -924 1818 -918
rect 1812 -930 1818 -924
rect 1812 -936 1818 -930
rect 1812 -942 1818 -936
rect 1812 -948 1818 -942
rect 1812 -954 1818 -948
rect 1812 -960 1818 -954
rect 1812 -966 1818 -960
rect 1812 -972 1818 -966
rect 1812 -978 1818 -972
rect 1812 -984 1818 -978
rect 1812 -990 1818 -984
rect 1812 -996 1818 -990
rect 1812 -1002 1818 -996
rect 1812 -1008 1818 -1002
rect 1812 -1014 1818 -1008
rect 1812 -1020 1818 -1014
rect 1812 -1026 1818 -1020
rect 1812 -1032 1818 -1026
rect 1812 -1038 1818 -1032
rect 1812 -1044 1818 -1038
rect 1812 -1050 1818 -1044
rect 1812 -1056 1818 -1050
rect 1812 -1062 1818 -1056
rect 1812 -1068 1818 -1062
rect 1812 -1074 1818 -1068
rect 1812 -1080 1818 -1074
rect 1812 -1086 1818 -1080
rect 1812 -1092 1818 -1086
rect 1812 -1098 1818 -1092
rect 1812 -1104 1818 -1098
rect 1812 -1110 1818 -1104
rect 1812 -1116 1818 -1110
rect 1812 -1122 1818 -1116
rect 1812 -1128 1818 -1122
rect 1812 -1134 1818 -1128
rect 1812 -1140 1818 -1134
rect 1812 -1146 1818 -1140
rect 1812 -1152 1818 -1146
rect 1812 -1158 1818 -1152
rect 1812 -1164 1818 -1158
rect 1812 -1170 1818 -1164
rect 1812 -1176 1818 -1170
rect 1812 -1182 1818 -1176
rect 1812 -1188 1818 -1182
rect 1812 -1194 1818 -1188
rect 1812 -1200 1818 -1194
rect 1812 -1206 1818 -1200
rect 1812 -1212 1818 -1206
rect 1812 -1218 1818 -1212
rect 1812 -1224 1818 -1218
rect 1812 -1230 1818 -1224
rect 1812 -1236 1818 -1230
rect 1812 -1242 1818 -1236
rect 1812 -1248 1818 -1242
rect 1812 -1254 1818 -1248
rect 1812 -1260 1818 -1254
rect 1812 -1266 1818 -1260
rect 1812 -1272 1818 -1266
rect 1812 -1278 1818 -1272
rect 1812 -1284 1818 -1278
rect 1812 -1290 1818 -1284
rect 1812 -1296 1818 -1290
rect 1812 -1302 1818 -1296
rect 1812 -1308 1818 -1302
rect 1812 -1314 1818 -1308
rect 1812 -1320 1818 -1314
rect 1812 -1326 1818 -1320
rect 1812 -1332 1818 -1326
rect 1812 -1338 1818 -1332
rect 1812 -1344 1818 -1338
rect 1812 -1350 1818 -1344
rect 1812 -1356 1818 -1350
rect 1812 -1362 1818 -1356
rect 1812 -1368 1818 -1362
rect 1812 -1374 1818 -1368
rect 1812 -1380 1818 -1374
rect 1812 -1386 1818 -1380
rect 1812 -1392 1818 -1386
rect 1812 -1398 1818 -1392
rect 1812 -1404 1818 -1398
rect 1812 -1410 1818 -1404
rect 1812 -1416 1818 -1410
rect 1812 -1422 1818 -1416
rect 1812 -1428 1818 -1422
rect 1812 -1434 1818 -1428
rect 1812 -1440 1818 -1434
rect 1812 -1446 1818 -1440
rect 1812 -1452 1818 -1446
rect 1812 -1458 1818 -1452
rect 1812 -1464 1818 -1458
rect 1812 -1470 1818 -1464
rect 1812 -1476 1818 -1470
rect 1812 -1482 1818 -1476
rect 1812 -1488 1818 -1482
rect 1812 -1494 1818 -1488
rect 1812 -1500 1818 -1494
rect 1812 -1506 1818 -1500
rect 1812 -1512 1818 -1506
rect 1812 -1518 1818 -1512
rect 1812 -1524 1818 -1518
rect 1812 -1530 1818 -1524
rect 1812 -1536 1818 -1530
rect 1812 -1542 1818 -1536
rect 1812 -1548 1818 -1542
rect 1812 -1554 1818 -1548
rect 1812 -1560 1818 -1554
rect 1812 -1566 1818 -1560
rect 1812 -1572 1818 -1566
rect 1812 -1578 1818 -1572
rect 1812 -1584 1818 -1578
rect 1812 -1590 1818 -1584
rect 1812 -1596 1818 -1590
rect 1812 -1602 1818 -1596
rect 1812 -1608 1818 -1602
rect 1812 -1614 1818 -1608
rect 1812 -1620 1818 -1614
rect 1812 -1626 1818 -1620
rect 1812 -1632 1818 -1626
rect 1812 -1638 1818 -1632
rect 1812 -1644 1818 -1638
rect 1812 -1650 1818 -1644
rect 1812 -1656 1818 -1650
rect 1812 -1662 1818 -1656
rect 1812 -1668 1818 -1662
rect 1812 -1674 1818 -1668
rect 1812 -1680 1818 -1674
rect 1812 -1686 1818 -1680
rect 1812 -1692 1818 -1686
rect 1812 -1698 1818 -1692
rect 1812 -1704 1818 -1698
rect 1812 -1710 1818 -1704
rect 1812 -1716 1818 -1710
rect 1812 -1722 1818 -1716
rect 1812 -1728 1818 -1722
rect 1812 -1734 1818 -1728
rect 1812 -1740 1818 -1734
rect 1812 -1746 1818 -1740
rect 1812 -1752 1818 -1746
rect 1812 -1758 1818 -1752
rect 1812 -1764 1818 -1758
rect 1812 -1770 1818 -1764
rect 1812 -1776 1818 -1770
rect 1812 -1782 1818 -1776
rect 1812 -1788 1818 -1782
rect 1812 -1794 1818 -1788
rect 1812 -1800 1818 -1794
rect 1812 -1806 1818 -1800
rect 1812 -1812 1818 -1806
rect 1812 -1818 1818 -1812
rect 1812 -1824 1818 -1818
rect 1812 -1830 1818 -1824
rect 1812 -1836 1818 -1830
rect 1812 -1914 1818 -1908
rect 1812 -1920 1818 -1914
rect 1812 -1926 1818 -1920
rect 1812 -1932 1818 -1926
rect 1812 -1938 1818 -1932
rect 1812 -1944 1818 -1938
rect 1812 -1950 1818 -1944
rect 1812 -1956 1818 -1950
rect 1812 -1962 1818 -1956
rect 1812 -1968 1818 -1962
rect 1812 -1974 1818 -1968
rect 1812 -1980 1818 -1974
rect 1812 -1986 1818 -1980
rect 1812 -1992 1818 -1986
rect 1812 -1998 1818 -1992
rect 1812 -2004 1818 -1998
rect 1812 -2010 1818 -2004
rect 1812 -2016 1818 -2010
rect 1812 -2022 1818 -2016
rect 1812 -2028 1818 -2022
rect 1812 -2034 1818 -2028
rect 1812 -2040 1818 -2034
rect 1812 -2046 1818 -2040
rect 1812 -2052 1818 -2046
rect 1812 -2058 1818 -2052
rect 1812 -2064 1818 -2058
rect 1812 -2070 1818 -2064
rect 1812 -2076 1818 -2070
rect 1812 -2082 1818 -2076
rect 1812 -2088 1818 -2082
rect 1812 -2094 1818 -2088
rect 1812 -2100 1818 -2094
rect 1812 -2106 1818 -2100
rect 1812 -2112 1818 -2106
rect 1812 -2118 1818 -2112
rect 1812 -2124 1818 -2118
rect 1812 -2130 1818 -2124
rect 1812 -2136 1818 -2130
rect 1812 -2142 1818 -2136
rect 1812 -2148 1818 -2142
rect 1812 -2154 1818 -2148
rect 1812 -2160 1818 -2154
rect 1812 -2166 1818 -2160
rect 1812 -2172 1818 -2166
rect 1812 -2178 1818 -2172
rect 1812 -2184 1818 -2178
rect 1812 -2190 1818 -2184
rect 1812 -2196 1818 -2190
rect 1812 -2202 1818 -2196
rect 1812 -2208 1818 -2202
rect 1812 -2214 1818 -2208
rect 1812 -2220 1818 -2214
rect 1812 -2226 1818 -2220
rect 1812 -2232 1818 -2226
rect 1812 -2238 1818 -2232
rect 1812 -2244 1818 -2238
rect 1812 -2250 1818 -2244
rect 1812 -2256 1818 -2250
rect 1812 -2262 1818 -2256
rect 1812 -2268 1818 -2262
rect 1812 -2274 1818 -2268
rect 1812 -2280 1818 -2274
rect 1812 -2286 1818 -2280
rect 1812 -2292 1818 -2286
rect 1812 -2298 1818 -2292
rect 1812 -2304 1818 -2298
rect 1812 -2310 1818 -2304
rect 1812 -2316 1818 -2310
rect 1812 -2322 1818 -2316
rect 1812 -2328 1818 -2322
rect 1812 -2334 1818 -2328
rect 1812 -2340 1818 -2334
rect 1812 -2346 1818 -2340
rect 1812 -2352 1818 -2346
rect 1812 -2358 1818 -2352
rect 1812 -2364 1818 -2358
rect 1812 -2370 1818 -2364
rect 1812 -2376 1818 -2370
rect 1812 -2382 1818 -2376
rect 1812 -2388 1818 -2382
rect 1812 -2394 1818 -2388
rect 1812 -2400 1818 -2394
rect 1812 -2406 1818 -2400
rect 1812 -2412 1818 -2406
rect 1812 -2418 1818 -2412
rect 1812 -2424 1818 -2418
rect 1812 -2430 1818 -2424
rect 1812 -2436 1818 -2430
rect 1812 -2442 1818 -2436
rect 1812 -2448 1818 -2442
rect 1812 -2454 1818 -2448
rect 1812 -2460 1818 -2454
rect 1812 -2466 1818 -2460
rect 1812 -2472 1818 -2466
rect 1812 -2478 1818 -2472
rect 1812 -2484 1818 -2478
rect 1812 -2490 1818 -2484
rect 1812 -2496 1818 -2490
rect 1812 -2502 1818 -2496
rect 1812 -2508 1818 -2502
rect 1812 -2514 1818 -2508
rect 1812 -2520 1818 -2514
rect 1812 -2526 1818 -2520
rect 1812 -2532 1818 -2526
rect 1812 -2538 1818 -2532
rect 1812 -2544 1818 -2538
rect 1812 -2550 1818 -2544
rect 1812 -2556 1818 -2550
rect 1812 -2562 1818 -2556
rect 1812 -2568 1818 -2562
rect 1812 -2574 1818 -2568
rect 1812 -2580 1818 -2574
rect 1812 -2586 1818 -2580
rect 1812 -2592 1818 -2586
rect 1812 -2598 1818 -2592
rect 1812 -2604 1818 -2598
rect 1812 -2610 1818 -2604
rect 1812 -2616 1818 -2610
rect 1812 -2622 1818 -2616
rect 1812 -2628 1818 -2622
rect 1812 -2700 1818 -2694
rect 1812 -2706 1818 -2700
rect 1812 -2712 1818 -2706
rect 1812 -2718 1818 -2712
rect 1812 -2724 1818 -2718
rect 1812 -2730 1818 -2724
rect 1812 -2736 1818 -2730
rect 1812 -2742 1818 -2736
rect 1812 -2748 1818 -2742
rect 1812 -2754 1818 -2748
rect 1812 -2760 1818 -2754
rect 1812 -2766 1818 -2760
rect 1812 -2772 1818 -2766
rect 1812 -2778 1818 -2772
rect 1812 -2784 1818 -2778
rect 1812 -2790 1818 -2784
rect 1812 -2796 1818 -2790
rect 1812 -2802 1818 -2796
rect 1812 -2808 1818 -2802
rect 1812 -2814 1818 -2808
rect 1812 -2820 1818 -2814
rect 1812 -2826 1818 -2820
rect 1812 -2832 1818 -2826
rect 1812 -2838 1818 -2832
rect 1812 -2844 1818 -2838
rect 1812 -2850 1818 -2844
rect 1812 -2856 1818 -2850
rect 1812 -2862 1818 -2856
rect 1812 -2868 1818 -2862
rect 1812 -2874 1818 -2868
rect 1812 -2880 1818 -2874
rect 1812 -2886 1818 -2880
rect 1812 -2892 1818 -2886
rect 1812 -2898 1818 -2892
rect 1812 -2904 1818 -2898
rect 1812 -2910 1818 -2904
rect 1812 -2916 1818 -2910
rect 1812 -2922 1818 -2916
rect 1812 -2928 1818 -2922
rect 1812 -2934 1818 -2928
rect 1812 -2940 1818 -2934
rect 1812 -2946 1818 -2940
rect 1812 -2952 1818 -2946
rect 1812 -2958 1818 -2952
rect 1812 -2964 1818 -2958
rect 1812 -2970 1818 -2964
rect 1812 -2976 1818 -2970
rect 1812 -2982 1818 -2976
rect 1812 -2988 1818 -2982
rect 1812 -2994 1818 -2988
rect 1812 -3000 1818 -2994
rect 1812 -3006 1818 -3000
rect 1812 -3012 1818 -3006
rect 1812 -3018 1818 -3012
rect 1812 -3024 1818 -3018
rect 1812 -3030 1818 -3024
rect 1812 -3036 1818 -3030
rect 1812 -3042 1818 -3036
rect 1812 -3048 1818 -3042
rect 1812 -3054 1818 -3048
rect 1812 -3060 1818 -3054
rect 1812 -3066 1818 -3060
rect 1812 -3072 1818 -3066
rect 1812 -3078 1818 -3072
rect 1812 -3084 1818 -3078
rect 1812 -3090 1818 -3084
rect 1812 -3096 1818 -3090
rect 1812 -3102 1818 -3096
rect 1812 -3108 1818 -3102
rect 1812 -3114 1818 -3108
rect 1812 -3120 1818 -3114
rect 1812 -3126 1818 -3120
rect 1812 -3132 1818 -3126
rect 1812 -3138 1818 -3132
rect 1812 -3144 1818 -3138
rect 1812 -3150 1818 -3144
rect 1812 -3156 1818 -3150
rect 1812 -3162 1818 -3156
rect 1812 -3168 1818 -3162
rect 1812 -3174 1818 -3168
rect 1812 -3180 1818 -3174
rect 1812 -3228 1818 -3222
rect 1812 -3234 1818 -3228
rect 1812 -3240 1818 -3234
rect 1812 -3246 1818 -3240
rect 1812 -3252 1818 -3246
rect 1812 -3258 1818 -3252
rect 1812 -3264 1818 -3258
rect 1812 -3270 1818 -3264
rect 1812 -3276 1818 -3270
rect 1812 -3282 1818 -3276
rect 1812 -3288 1818 -3282
rect 1812 -3294 1818 -3288
rect 1812 -3300 1818 -3294
rect 1812 -3306 1818 -3300
rect 1812 -3312 1818 -3306
rect 1812 -3318 1818 -3312
rect 1812 -3324 1818 -3318
rect 1812 -3330 1818 -3324
rect 1812 -3336 1818 -3330
rect 1812 -3342 1818 -3336
rect 1812 -3348 1818 -3342
rect 1812 -3354 1818 -3348
rect 1812 -3360 1818 -3354
rect 1818 -696 1824 -690
rect 1818 -702 1824 -696
rect 1818 -708 1824 -702
rect 1818 -714 1824 -708
rect 1818 -720 1824 -714
rect 1818 -726 1824 -720
rect 1818 -732 1824 -726
rect 1818 -738 1824 -732
rect 1818 -744 1824 -738
rect 1818 -750 1824 -744
rect 1818 -756 1824 -750
rect 1818 -762 1824 -756
rect 1818 -768 1824 -762
rect 1818 -774 1824 -768
rect 1818 -780 1824 -774
rect 1818 -786 1824 -780
rect 1818 -792 1824 -786
rect 1818 -798 1824 -792
rect 1818 -804 1824 -798
rect 1818 -810 1824 -804
rect 1818 -816 1824 -810
rect 1818 -822 1824 -816
rect 1818 -828 1824 -822
rect 1818 -834 1824 -828
rect 1818 -840 1824 -834
rect 1818 -846 1824 -840
rect 1818 -852 1824 -846
rect 1818 -858 1824 -852
rect 1818 -864 1824 -858
rect 1818 -870 1824 -864
rect 1818 -876 1824 -870
rect 1818 -882 1824 -876
rect 1818 -888 1824 -882
rect 1818 -894 1824 -888
rect 1818 -900 1824 -894
rect 1818 -906 1824 -900
rect 1818 -912 1824 -906
rect 1818 -918 1824 -912
rect 1818 -924 1824 -918
rect 1818 -930 1824 -924
rect 1818 -936 1824 -930
rect 1818 -942 1824 -936
rect 1818 -948 1824 -942
rect 1818 -954 1824 -948
rect 1818 -960 1824 -954
rect 1818 -966 1824 -960
rect 1818 -972 1824 -966
rect 1818 -978 1824 -972
rect 1818 -984 1824 -978
rect 1818 -990 1824 -984
rect 1818 -996 1824 -990
rect 1818 -1002 1824 -996
rect 1818 -1008 1824 -1002
rect 1818 -1014 1824 -1008
rect 1818 -1020 1824 -1014
rect 1818 -1026 1824 -1020
rect 1818 -1032 1824 -1026
rect 1818 -1038 1824 -1032
rect 1818 -1044 1824 -1038
rect 1818 -1050 1824 -1044
rect 1818 -1056 1824 -1050
rect 1818 -1062 1824 -1056
rect 1818 -1068 1824 -1062
rect 1818 -1074 1824 -1068
rect 1818 -1080 1824 -1074
rect 1818 -1086 1824 -1080
rect 1818 -1092 1824 -1086
rect 1818 -1098 1824 -1092
rect 1818 -1104 1824 -1098
rect 1818 -1110 1824 -1104
rect 1818 -1116 1824 -1110
rect 1818 -1122 1824 -1116
rect 1818 -1128 1824 -1122
rect 1818 -1134 1824 -1128
rect 1818 -1140 1824 -1134
rect 1818 -1146 1824 -1140
rect 1818 -1152 1824 -1146
rect 1818 -1158 1824 -1152
rect 1818 -1164 1824 -1158
rect 1818 -1170 1824 -1164
rect 1818 -1176 1824 -1170
rect 1818 -1182 1824 -1176
rect 1818 -1188 1824 -1182
rect 1818 -1194 1824 -1188
rect 1818 -1200 1824 -1194
rect 1818 -1206 1824 -1200
rect 1818 -1212 1824 -1206
rect 1818 -1218 1824 -1212
rect 1818 -1224 1824 -1218
rect 1818 -1230 1824 -1224
rect 1818 -1236 1824 -1230
rect 1818 -1242 1824 -1236
rect 1818 -1248 1824 -1242
rect 1818 -1254 1824 -1248
rect 1818 -1260 1824 -1254
rect 1818 -1266 1824 -1260
rect 1818 -1272 1824 -1266
rect 1818 -1278 1824 -1272
rect 1818 -1284 1824 -1278
rect 1818 -1290 1824 -1284
rect 1818 -1296 1824 -1290
rect 1818 -1302 1824 -1296
rect 1818 -1308 1824 -1302
rect 1818 -1314 1824 -1308
rect 1818 -1320 1824 -1314
rect 1818 -1326 1824 -1320
rect 1818 -1332 1824 -1326
rect 1818 -1338 1824 -1332
rect 1818 -1344 1824 -1338
rect 1818 -1350 1824 -1344
rect 1818 -1356 1824 -1350
rect 1818 -1362 1824 -1356
rect 1818 -1368 1824 -1362
rect 1818 -1374 1824 -1368
rect 1818 -1380 1824 -1374
rect 1818 -1386 1824 -1380
rect 1818 -1392 1824 -1386
rect 1818 -1398 1824 -1392
rect 1818 -1404 1824 -1398
rect 1818 -1410 1824 -1404
rect 1818 -1416 1824 -1410
rect 1818 -1422 1824 -1416
rect 1818 -1428 1824 -1422
rect 1818 -1434 1824 -1428
rect 1818 -1440 1824 -1434
rect 1818 -1446 1824 -1440
rect 1818 -1452 1824 -1446
rect 1818 -1458 1824 -1452
rect 1818 -1464 1824 -1458
rect 1818 -1470 1824 -1464
rect 1818 -1476 1824 -1470
rect 1818 -1482 1824 -1476
rect 1818 -1488 1824 -1482
rect 1818 -1494 1824 -1488
rect 1818 -1500 1824 -1494
rect 1818 -1506 1824 -1500
rect 1818 -1512 1824 -1506
rect 1818 -1518 1824 -1512
rect 1818 -1524 1824 -1518
rect 1818 -1530 1824 -1524
rect 1818 -1536 1824 -1530
rect 1818 -1542 1824 -1536
rect 1818 -1548 1824 -1542
rect 1818 -1554 1824 -1548
rect 1818 -1560 1824 -1554
rect 1818 -1566 1824 -1560
rect 1818 -1572 1824 -1566
rect 1818 -1578 1824 -1572
rect 1818 -1584 1824 -1578
rect 1818 -1590 1824 -1584
rect 1818 -1596 1824 -1590
rect 1818 -1602 1824 -1596
rect 1818 -1608 1824 -1602
rect 1818 -1614 1824 -1608
rect 1818 -1620 1824 -1614
rect 1818 -1626 1824 -1620
rect 1818 -1632 1824 -1626
rect 1818 -1638 1824 -1632
rect 1818 -1644 1824 -1638
rect 1818 -1650 1824 -1644
rect 1818 -1656 1824 -1650
rect 1818 -1662 1824 -1656
rect 1818 -1668 1824 -1662
rect 1818 -1674 1824 -1668
rect 1818 -1680 1824 -1674
rect 1818 -1686 1824 -1680
rect 1818 -1692 1824 -1686
rect 1818 -1698 1824 -1692
rect 1818 -1704 1824 -1698
rect 1818 -1710 1824 -1704
rect 1818 -1716 1824 -1710
rect 1818 -1722 1824 -1716
rect 1818 -1728 1824 -1722
rect 1818 -1734 1824 -1728
rect 1818 -1740 1824 -1734
rect 1818 -1746 1824 -1740
rect 1818 -1752 1824 -1746
rect 1818 -1758 1824 -1752
rect 1818 -1764 1824 -1758
rect 1818 -1770 1824 -1764
rect 1818 -1776 1824 -1770
rect 1818 -1782 1824 -1776
rect 1818 -1788 1824 -1782
rect 1818 -1794 1824 -1788
rect 1818 -1800 1824 -1794
rect 1818 -1806 1824 -1800
rect 1818 -1812 1824 -1806
rect 1818 -1818 1824 -1812
rect 1818 -1824 1824 -1818
rect 1818 -1830 1824 -1824
rect 1818 -1908 1824 -1902
rect 1818 -1914 1824 -1908
rect 1818 -1920 1824 -1914
rect 1818 -1926 1824 -1920
rect 1818 -1932 1824 -1926
rect 1818 -1938 1824 -1932
rect 1818 -1944 1824 -1938
rect 1818 -1950 1824 -1944
rect 1818 -1956 1824 -1950
rect 1818 -1962 1824 -1956
rect 1818 -1968 1824 -1962
rect 1818 -1974 1824 -1968
rect 1818 -1980 1824 -1974
rect 1818 -1986 1824 -1980
rect 1818 -1992 1824 -1986
rect 1818 -1998 1824 -1992
rect 1818 -2004 1824 -1998
rect 1818 -2010 1824 -2004
rect 1818 -2016 1824 -2010
rect 1818 -2022 1824 -2016
rect 1818 -2028 1824 -2022
rect 1818 -2034 1824 -2028
rect 1818 -2040 1824 -2034
rect 1818 -2046 1824 -2040
rect 1818 -2052 1824 -2046
rect 1818 -2058 1824 -2052
rect 1818 -2064 1824 -2058
rect 1818 -2070 1824 -2064
rect 1818 -2076 1824 -2070
rect 1818 -2082 1824 -2076
rect 1818 -2088 1824 -2082
rect 1818 -2094 1824 -2088
rect 1818 -2100 1824 -2094
rect 1818 -2106 1824 -2100
rect 1818 -2112 1824 -2106
rect 1818 -2118 1824 -2112
rect 1818 -2124 1824 -2118
rect 1818 -2130 1824 -2124
rect 1818 -2136 1824 -2130
rect 1818 -2142 1824 -2136
rect 1818 -2148 1824 -2142
rect 1818 -2154 1824 -2148
rect 1818 -2160 1824 -2154
rect 1818 -2166 1824 -2160
rect 1818 -2172 1824 -2166
rect 1818 -2178 1824 -2172
rect 1818 -2184 1824 -2178
rect 1818 -2190 1824 -2184
rect 1818 -2196 1824 -2190
rect 1818 -2202 1824 -2196
rect 1818 -2208 1824 -2202
rect 1818 -2214 1824 -2208
rect 1818 -2220 1824 -2214
rect 1818 -2226 1824 -2220
rect 1818 -2232 1824 -2226
rect 1818 -2238 1824 -2232
rect 1818 -2244 1824 -2238
rect 1818 -2250 1824 -2244
rect 1818 -2256 1824 -2250
rect 1818 -2262 1824 -2256
rect 1818 -2268 1824 -2262
rect 1818 -2274 1824 -2268
rect 1818 -2280 1824 -2274
rect 1818 -2286 1824 -2280
rect 1818 -2292 1824 -2286
rect 1818 -2298 1824 -2292
rect 1818 -2304 1824 -2298
rect 1818 -2310 1824 -2304
rect 1818 -2316 1824 -2310
rect 1818 -2322 1824 -2316
rect 1818 -2328 1824 -2322
rect 1818 -2334 1824 -2328
rect 1818 -2340 1824 -2334
rect 1818 -2346 1824 -2340
rect 1818 -2352 1824 -2346
rect 1818 -2358 1824 -2352
rect 1818 -2364 1824 -2358
rect 1818 -2370 1824 -2364
rect 1818 -2376 1824 -2370
rect 1818 -2382 1824 -2376
rect 1818 -2388 1824 -2382
rect 1818 -2394 1824 -2388
rect 1818 -2400 1824 -2394
rect 1818 -2406 1824 -2400
rect 1818 -2412 1824 -2406
rect 1818 -2418 1824 -2412
rect 1818 -2424 1824 -2418
rect 1818 -2430 1824 -2424
rect 1818 -2436 1824 -2430
rect 1818 -2442 1824 -2436
rect 1818 -2448 1824 -2442
rect 1818 -2454 1824 -2448
rect 1818 -2460 1824 -2454
rect 1818 -2466 1824 -2460
rect 1818 -2472 1824 -2466
rect 1818 -2478 1824 -2472
rect 1818 -2484 1824 -2478
rect 1818 -2490 1824 -2484
rect 1818 -2496 1824 -2490
rect 1818 -2502 1824 -2496
rect 1818 -2508 1824 -2502
rect 1818 -2514 1824 -2508
rect 1818 -2520 1824 -2514
rect 1818 -2526 1824 -2520
rect 1818 -2532 1824 -2526
rect 1818 -2538 1824 -2532
rect 1818 -2544 1824 -2538
rect 1818 -2550 1824 -2544
rect 1818 -2556 1824 -2550
rect 1818 -2562 1824 -2556
rect 1818 -2568 1824 -2562
rect 1818 -2574 1824 -2568
rect 1818 -2580 1824 -2574
rect 1818 -2586 1824 -2580
rect 1818 -2592 1824 -2586
rect 1818 -2598 1824 -2592
rect 1818 -2604 1824 -2598
rect 1818 -2610 1824 -2604
rect 1818 -2616 1824 -2610
rect 1818 -2622 1824 -2616
rect 1818 -2694 1824 -2688
rect 1818 -2700 1824 -2694
rect 1818 -2706 1824 -2700
rect 1818 -2712 1824 -2706
rect 1818 -2718 1824 -2712
rect 1818 -2724 1824 -2718
rect 1818 -2730 1824 -2724
rect 1818 -2736 1824 -2730
rect 1818 -2742 1824 -2736
rect 1818 -2748 1824 -2742
rect 1818 -2754 1824 -2748
rect 1818 -2760 1824 -2754
rect 1818 -2766 1824 -2760
rect 1818 -2772 1824 -2766
rect 1818 -2778 1824 -2772
rect 1818 -2784 1824 -2778
rect 1818 -2790 1824 -2784
rect 1818 -2796 1824 -2790
rect 1818 -2802 1824 -2796
rect 1818 -2808 1824 -2802
rect 1818 -2814 1824 -2808
rect 1818 -2820 1824 -2814
rect 1818 -2826 1824 -2820
rect 1818 -2832 1824 -2826
rect 1818 -2838 1824 -2832
rect 1818 -2844 1824 -2838
rect 1818 -2850 1824 -2844
rect 1818 -2856 1824 -2850
rect 1818 -2862 1824 -2856
rect 1818 -2868 1824 -2862
rect 1818 -2874 1824 -2868
rect 1818 -2880 1824 -2874
rect 1818 -2886 1824 -2880
rect 1818 -2892 1824 -2886
rect 1818 -2898 1824 -2892
rect 1818 -2904 1824 -2898
rect 1818 -2910 1824 -2904
rect 1818 -2916 1824 -2910
rect 1818 -2922 1824 -2916
rect 1818 -2928 1824 -2922
rect 1818 -2934 1824 -2928
rect 1818 -2940 1824 -2934
rect 1818 -2946 1824 -2940
rect 1818 -2952 1824 -2946
rect 1818 -2958 1824 -2952
rect 1818 -2964 1824 -2958
rect 1818 -2970 1824 -2964
rect 1818 -2976 1824 -2970
rect 1818 -2982 1824 -2976
rect 1818 -2988 1824 -2982
rect 1818 -2994 1824 -2988
rect 1818 -3000 1824 -2994
rect 1818 -3006 1824 -3000
rect 1818 -3012 1824 -3006
rect 1818 -3018 1824 -3012
rect 1818 -3024 1824 -3018
rect 1818 -3030 1824 -3024
rect 1818 -3036 1824 -3030
rect 1818 -3042 1824 -3036
rect 1818 -3048 1824 -3042
rect 1818 -3054 1824 -3048
rect 1818 -3060 1824 -3054
rect 1818 -3066 1824 -3060
rect 1818 -3072 1824 -3066
rect 1818 -3078 1824 -3072
rect 1818 -3084 1824 -3078
rect 1818 -3090 1824 -3084
rect 1818 -3096 1824 -3090
rect 1818 -3102 1824 -3096
rect 1818 -3108 1824 -3102
rect 1818 -3114 1824 -3108
rect 1818 -3120 1824 -3114
rect 1818 -3126 1824 -3120
rect 1818 -3132 1824 -3126
rect 1818 -3138 1824 -3132
rect 1818 -3144 1824 -3138
rect 1818 -3150 1824 -3144
rect 1818 -3156 1824 -3150
rect 1818 -3162 1824 -3156
rect 1818 -3168 1824 -3162
rect 1818 -3174 1824 -3168
rect 1818 -3228 1824 -3222
rect 1818 -3234 1824 -3228
rect 1818 -3240 1824 -3234
rect 1818 -3246 1824 -3240
rect 1818 -3252 1824 -3246
rect 1818 -3258 1824 -3252
rect 1818 -3264 1824 -3258
rect 1818 -3270 1824 -3264
rect 1818 -3276 1824 -3270
rect 1818 -3282 1824 -3276
rect 1818 -3288 1824 -3282
rect 1818 -3294 1824 -3288
rect 1818 -3300 1824 -3294
rect 1818 -3306 1824 -3300
rect 1818 -3312 1824 -3306
rect 1818 -3318 1824 -3312
rect 1818 -3324 1824 -3318
rect 1818 -3330 1824 -3324
rect 1818 -3336 1824 -3330
rect 1818 -3342 1824 -3336
rect 1818 -3348 1824 -3342
rect 1818 -3354 1824 -3348
rect 1818 -3360 1824 -3354
rect 1824 -684 1830 -678
rect 1824 -690 1830 -684
rect 1824 -696 1830 -690
rect 1824 -702 1830 -696
rect 1824 -708 1830 -702
rect 1824 -714 1830 -708
rect 1824 -720 1830 -714
rect 1824 -726 1830 -720
rect 1824 -732 1830 -726
rect 1824 -738 1830 -732
rect 1824 -744 1830 -738
rect 1824 -750 1830 -744
rect 1824 -756 1830 -750
rect 1824 -762 1830 -756
rect 1824 -768 1830 -762
rect 1824 -774 1830 -768
rect 1824 -780 1830 -774
rect 1824 -786 1830 -780
rect 1824 -792 1830 -786
rect 1824 -798 1830 -792
rect 1824 -804 1830 -798
rect 1824 -810 1830 -804
rect 1824 -816 1830 -810
rect 1824 -822 1830 -816
rect 1824 -828 1830 -822
rect 1824 -834 1830 -828
rect 1824 -840 1830 -834
rect 1824 -846 1830 -840
rect 1824 -852 1830 -846
rect 1824 -858 1830 -852
rect 1824 -864 1830 -858
rect 1824 -870 1830 -864
rect 1824 -876 1830 -870
rect 1824 -882 1830 -876
rect 1824 -888 1830 -882
rect 1824 -894 1830 -888
rect 1824 -900 1830 -894
rect 1824 -906 1830 -900
rect 1824 -912 1830 -906
rect 1824 -918 1830 -912
rect 1824 -924 1830 -918
rect 1824 -930 1830 -924
rect 1824 -936 1830 -930
rect 1824 -942 1830 -936
rect 1824 -948 1830 -942
rect 1824 -954 1830 -948
rect 1824 -960 1830 -954
rect 1824 -966 1830 -960
rect 1824 -972 1830 -966
rect 1824 -978 1830 -972
rect 1824 -984 1830 -978
rect 1824 -990 1830 -984
rect 1824 -996 1830 -990
rect 1824 -1002 1830 -996
rect 1824 -1008 1830 -1002
rect 1824 -1014 1830 -1008
rect 1824 -1020 1830 -1014
rect 1824 -1026 1830 -1020
rect 1824 -1032 1830 -1026
rect 1824 -1038 1830 -1032
rect 1824 -1044 1830 -1038
rect 1824 -1050 1830 -1044
rect 1824 -1056 1830 -1050
rect 1824 -1062 1830 -1056
rect 1824 -1068 1830 -1062
rect 1824 -1074 1830 -1068
rect 1824 -1080 1830 -1074
rect 1824 -1086 1830 -1080
rect 1824 -1092 1830 -1086
rect 1824 -1098 1830 -1092
rect 1824 -1104 1830 -1098
rect 1824 -1110 1830 -1104
rect 1824 -1116 1830 -1110
rect 1824 -1122 1830 -1116
rect 1824 -1128 1830 -1122
rect 1824 -1134 1830 -1128
rect 1824 -1140 1830 -1134
rect 1824 -1146 1830 -1140
rect 1824 -1152 1830 -1146
rect 1824 -1158 1830 -1152
rect 1824 -1164 1830 -1158
rect 1824 -1170 1830 -1164
rect 1824 -1176 1830 -1170
rect 1824 -1182 1830 -1176
rect 1824 -1188 1830 -1182
rect 1824 -1194 1830 -1188
rect 1824 -1200 1830 -1194
rect 1824 -1206 1830 -1200
rect 1824 -1212 1830 -1206
rect 1824 -1218 1830 -1212
rect 1824 -1224 1830 -1218
rect 1824 -1230 1830 -1224
rect 1824 -1236 1830 -1230
rect 1824 -1242 1830 -1236
rect 1824 -1248 1830 -1242
rect 1824 -1254 1830 -1248
rect 1824 -1260 1830 -1254
rect 1824 -1266 1830 -1260
rect 1824 -1272 1830 -1266
rect 1824 -1278 1830 -1272
rect 1824 -1284 1830 -1278
rect 1824 -1290 1830 -1284
rect 1824 -1296 1830 -1290
rect 1824 -1302 1830 -1296
rect 1824 -1308 1830 -1302
rect 1824 -1314 1830 -1308
rect 1824 -1320 1830 -1314
rect 1824 -1326 1830 -1320
rect 1824 -1332 1830 -1326
rect 1824 -1338 1830 -1332
rect 1824 -1344 1830 -1338
rect 1824 -1350 1830 -1344
rect 1824 -1356 1830 -1350
rect 1824 -1362 1830 -1356
rect 1824 -1368 1830 -1362
rect 1824 -1374 1830 -1368
rect 1824 -1380 1830 -1374
rect 1824 -1386 1830 -1380
rect 1824 -1392 1830 -1386
rect 1824 -1398 1830 -1392
rect 1824 -1404 1830 -1398
rect 1824 -1410 1830 -1404
rect 1824 -1416 1830 -1410
rect 1824 -1422 1830 -1416
rect 1824 -1428 1830 -1422
rect 1824 -1434 1830 -1428
rect 1824 -1440 1830 -1434
rect 1824 -1446 1830 -1440
rect 1824 -1452 1830 -1446
rect 1824 -1458 1830 -1452
rect 1824 -1464 1830 -1458
rect 1824 -1470 1830 -1464
rect 1824 -1476 1830 -1470
rect 1824 -1482 1830 -1476
rect 1824 -1488 1830 -1482
rect 1824 -1494 1830 -1488
rect 1824 -1500 1830 -1494
rect 1824 -1506 1830 -1500
rect 1824 -1512 1830 -1506
rect 1824 -1518 1830 -1512
rect 1824 -1524 1830 -1518
rect 1824 -1530 1830 -1524
rect 1824 -1536 1830 -1530
rect 1824 -1542 1830 -1536
rect 1824 -1548 1830 -1542
rect 1824 -1554 1830 -1548
rect 1824 -1560 1830 -1554
rect 1824 -1566 1830 -1560
rect 1824 -1572 1830 -1566
rect 1824 -1578 1830 -1572
rect 1824 -1584 1830 -1578
rect 1824 -1590 1830 -1584
rect 1824 -1596 1830 -1590
rect 1824 -1602 1830 -1596
rect 1824 -1608 1830 -1602
rect 1824 -1614 1830 -1608
rect 1824 -1620 1830 -1614
rect 1824 -1626 1830 -1620
rect 1824 -1632 1830 -1626
rect 1824 -1638 1830 -1632
rect 1824 -1644 1830 -1638
rect 1824 -1650 1830 -1644
rect 1824 -1656 1830 -1650
rect 1824 -1662 1830 -1656
rect 1824 -1668 1830 -1662
rect 1824 -1674 1830 -1668
rect 1824 -1680 1830 -1674
rect 1824 -1686 1830 -1680
rect 1824 -1692 1830 -1686
rect 1824 -1698 1830 -1692
rect 1824 -1704 1830 -1698
rect 1824 -1710 1830 -1704
rect 1824 -1716 1830 -1710
rect 1824 -1722 1830 -1716
rect 1824 -1728 1830 -1722
rect 1824 -1734 1830 -1728
rect 1824 -1740 1830 -1734
rect 1824 -1746 1830 -1740
rect 1824 -1752 1830 -1746
rect 1824 -1758 1830 -1752
rect 1824 -1764 1830 -1758
rect 1824 -1770 1830 -1764
rect 1824 -1776 1830 -1770
rect 1824 -1782 1830 -1776
rect 1824 -1788 1830 -1782
rect 1824 -1794 1830 -1788
rect 1824 -1800 1830 -1794
rect 1824 -1806 1830 -1800
rect 1824 -1812 1830 -1806
rect 1824 -1818 1830 -1812
rect 1824 -1824 1830 -1818
rect 1824 -1902 1830 -1896
rect 1824 -1908 1830 -1902
rect 1824 -1914 1830 -1908
rect 1824 -1920 1830 -1914
rect 1824 -1926 1830 -1920
rect 1824 -1932 1830 -1926
rect 1824 -1938 1830 -1932
rect 1824 -1944 1830 -1938
rect 1824 -1950 1830 -1944
rect 1824 -1956 1830 -1950
rect 1824 -1962 1830 -1956
rect 1824 -1968 1830 -1962
rect 1824 -1974 1830 -1968
rect 1824 -1980 1830 -1974
rect 1824 -1986 1830 -1980
rect 1824 -1992 1830 -1986
rect 1824 -1998 1830 -1992
rect 1824 -2004 1830 -1998
rect 1824 -2010 1830 -2004
rect 1824 -2016 1830 -2010
rect 1824 -2022 1830 -2016
rect 1824 -2028 1830 -2022
rect 1824 -2034 1830 -2028
rect 1824 -2040 1830 -2034
rect 1824 -2046 1830 -2040
rect 1824 -2052 1830 -2046
rect 1824 -2058 1830 -2052
rect 1824 -2064 1830 -2058
rect 1824 -2070 1830 -2064
rect 1824 -2076 1830 -2070
rect 1824 -2082 1830 -2076
rect 1824 -2088 1830 -2082
rect 1824 -2094 1830 -2088
rect 1824 -2100 1830 -2094
rect 1824 -2106 1830 -2100
rect 1824 -2112 1830 -2106
rect 1824 -2118 1830 -2112
rect 1824 -2124 1830 -2118
rect 1824 -2130 1830 -2124
rect 1824 -2136 1830 -2130
rect 1824 -2142 1830 -2136
rect 1824 -2148 1830 -2142
rect 1824 -2154 1830 -2148
rect 1824 -2160 1830 -2154
rect 1824 -2166 1830 -2160
rect 1824 -2172 1830 -2166
rect 1824 -2178 1830 -2172
rect 1824 -2184 1830 -2178
rect 1824 -2190 1830 -2184
rect 1824 -2196 1830 -2190
rect 1824 -2202 1830 -2196
rect 1824 -2208 1830 -2202
rect 1824 -2214 1830 -2208
rect 1824 -2220 1830 -2214
rect 1824 -2226 1830 -2220
rect 1824 -2232 1830 -2226
rect 1824 -2238 1830 -2232
rect 1824 -2244 1830 -2238
rect 1824 -2250 1830 -2244
rect 1824 -2256 1830 -2250
rect 1824 -2262 1830 -2256
rect 1824 -2268 1830 -2262
rect 1824 -2274 1830 -2268
rect 1824 -2280 1830 -2274
rect 1824 -2286 1830 -2280
rect 1824 -2292 1830 -2286
rect 1824 -2298 1830 -2292
rect 1824 -2304 1830 -2298
rect 1824 -2310 1830 -2304
rect 1824 -2316 1830 -2310
rect 1824 -2322 1830 -2316
rect 1824 -2328 1830 -2322
rect 1824 -2334 1830 -2328
rect 1824 -2340 1830 -2334
rect 1824 -2346 1830 -2340
rect 1824 -2352 1830 -2346
rect 1824 -2358 1830 -2352
rect 1824 -2364 1830 -2358
rect 1824 -2370 1830 -2364
rect 1824 -2376 1830 -2370
rect 1824 -2382 1830 -2376
rect 1824 -2388 1830 -2382
rect 1824 -2394 1830 -2388
rect 1824 -2400 1830 -2394
rect 1824 -2406 1830 -2400
rect 1824 -2412 1830 -2406
rect 1824 -2418 1830 -2412
rect 1824 -2424 1830 -2418
rect 1824 -2430 1830 -2424
rect 1824 -2436 1830 -2430
rect 1824 -2442 1830 -2436
rect 1824 -2448 1830 -2442
rect 1824 -2454 1830 -2448
rect 1824 -2460 1830 -2454
rect 1824 -2466 1830 -2460
rect 1824 -2472 1830 -2466
rect 1824 -2478 1830 -2472
rect 1824 -2484 1830 -2478
rect 1824 -2490 1830 -2484
rect 1824 -2496 1830 -2490
rect 1824 -2502 1830 -2496
rect 1824 -2508 1830 -2502
rect 1824 -2514 1830 -2508
rect 1824 -2520 1830 -2514
rect 1824 -2526 1830 -2520
rect 1824 -2532 1830 -2526
rect 1824 -2538 1830 -2532
rect 1824 -2544 1830 -2538
rect 1824 -2550 1830 -2544
rect 1824 -2556 1830 -2550
rect 1824 -2562 1830 -2556
rect 1824 -2568 1830 -2562
rect 1824 -2574 1830 -2568
rect 1824 -2580 1830 -2574
rect 1824 -2586 1830 -2580
rect 1824 -2592 1830 -2586
rect 1824 -2598 1830 -2592
rect 1824 -2604 1830 -2598
rect 1824 -2610 1830 -2604
rect 1824 -2616 1830 -2610
rect 1824 -2622 1830 -2616
rect 1824 -2694 1830 -2688
rect 1824 -2700 1830 -2694
rect 1824 -2706 1830 -2700
rect 1824 -2712 1830 -2706
rect 1824 -2718 1830 -2712
rect 1824 -2724 1830 -2718
rect 1824 -2730 1830 -2724
rect 1824 -2736 1830 -2730
rect 1824 -2742 1830 -2736
rect 1824 -2748 1830 -2742
rect 1824 -2754 1830 -2748
rect 1824 -2760 1830 -2754
rect 1824 -2766 1830 -2760
rect 1824 -2772 1830 -2766
rect 1824 -2778 1830 -2772
rect 1824 -2784 1830 -2778
rect 1824 -2790 1830 -2784
rect 1824 -2796 1830 -2790
rect 1824 -2802 1830 -2796
rect 1824 -2808 1830 -2802
rect 1824 -2814 1830 -2808
rect 1824 -2820 1830 -2814
rect 1824 -2826 1830 -2820
rect 1824 -2832 1830 -2826
rect 1824 -2838 1830 -2832
rect 1824 -2844 1830 -2838
rect 1824 -2850 1830 -2844
rect 1824 -2856 1830 -2850
rect 1824 -2862 1830 -2856
rect 1824 -2868 1830 -2862
rect 1824 -2874 1830 -2868
rect 1824 -2880 1830 -2874
rect 1824 -2886 1830 -2880
rect 1824 -2892 1830 -2886
rect 1824 -2898 1830 -2892
rect 1824 -2904 1830 -2898
rect 1824 -2910 1830 -2904
rect 1824 -2916 1830 -2910
rect 1824 -2922 1830 -2916
rect 1824 -2928 1830 -2922
rect 1824 -2934 1830 -2928
rect 1824 -2940 1830 -2934
rect 1824 -2946 1830 -2940
rect 1824 -2952 1830 -2946
rect 1824 -2958 1830 -2952
rect 1824 -2964 1830 -2958
rect 1824 -2970 1830 -2964
rect 1824 -2976 1830 -2970
rect 1824 -2982 1830 -2976
rect 1824 -2988 1830 -2982
rect 1824 -2994 1830 -2988
rect 1824 -3000 1830 -2994
rect 1824 -3006 1830 -3000
rect 1824 -3012 1830 -3006
rect 1824 -3018 1830 -3012
rect 1824 -3024 1830 -3018
rect 1824 -3030 1830 -3024
rect 1824 -3036 1830 -3030
rect 1824 -3042 1830 -3036
rect 1824 -3048 1830 -3042
rect 1824 -3054 1830 -3048
rect 1824 -3060 1830 -3054
rect 1824 -3066 1830 -3060
rect 1824 -3072 1830 -3066
rect 1824 -3078 1830 -3072
rect 1824 -3084 1830 -3078
rect 1824 -3090 1830 -3084
rect 1824 -3096 1830 -3090
rect 1824 -3102 1830 -3096
rect 1824 -3108 1830 -3102
rect 1824 -3114 1830 -3108
rect 1824 -3120 1830 -3114
rect 1824 -3126 1830 -3120
rect 1824 -3132 1830 -3126
rect 1824 -3138 1830 -3132
rect 1824 -3144 1830 -3138
rect 1824 -3150 1830 -3144
rect 1824 -3156 1830 -3150
rect 1824 -3162 1830 -3156
rect 1824 -3168 1830 -3162
rect 1824 -3174 1830 -3168
rect 1824 -3222 1830 -3216
rect 1824 -3228 1830 -3222
rect 1824 -3234 1830 -3228
rect 1824 -3240 1830 -3234
rect 1824 -3246 1830 -3240
rect 1824 -3252 1830 -3246
rect 1824 -3258 1830 -3252
rect 1824 -3264 1830 -3258
rect 1824 -3270 1830 -3264
rect 1824 -3276 1830 -3270
rect 1824 -3282 1830 -3276
rect 1824 -3288 1830 -3282
rect 1824 -3294 1830 -3288
rect 1824 -3300 1830 -3294
rect 1824 -3306 1830 -3300
rect 1824 -3312 1830 -3306
rect 1824 -3318 1830 -3312
rect 1824 -3324 1830 -3318
rect 1824 -3330 1830 -3324
rect 1824 -3336 1830 -3330
rect 1824 -3342 1830 -3336
rect 1824 -3348 1830 -3342
rect 1824 -3354 1830 -3348
rect 1830 -678 1836 -672
rect 1830 -684 1836 -678
rect 1830 -690 1836 -684
rect 1830 -696 1836 -690
rect 1830 -702 1836 -696
rect 1830 -708 1836 -702
rect 1830 -714 1836 -708
rect 1830 -720 1836 -714
rect 1830 -726 1836 -720
rect 1830 -732 1836 -726
rect 1830 -738 1836 -732
rect 1830 -744 1836 -738
rect 1830 -750 1836 -744
rect 1830 -756 1836 -750
rect 1830 -762 1836 -756
rect 1830 -768 1836 -762
rect 1830 -774 1836 -768
rect 1830 -780 1836 -774
rect 1830 -786 1836 -780
rect 1830 -792 1836 -786
rect 1830 -798 1836 -792
rect 1830 -804 1836 -798
rect 1830 -810 1836 -804
rect 1830 -816 1836 -810
rect 1830 -822 1836 -816
rect 1830 -828 1836 -822
rect 1830 -834 1836 -828
rect 1830 -840 1836 -834
rect 1830 -846 1836 -840
rect 1830 -852 1836 -846
rect 1830 -858 1836 -852
rect 1830 -864 1836 -858
rect 1830 -870 1836 -864
rect 1830 -876 1836 -870
rect 1830 -882 1836 -876
rect 1830 -888 1836 -882
rect 1830 -894 1836 -888
rect 1830 -900 1836 -894
rect 1830 -906 1836 -900
rect 1830 -912 1836 -906
rect 1830 -918 1836 -912
rect 1830 -924 1836 -918
rect 1830 -930 1836 -924
rect 1830 -936 1836 -930
rect 1830 -942 1836 -936
rect 1830 -948 1836 -942
rect 1830 -954 1836 -948
rect 1830 -960 1836 -954
rect 1830 -966 1836 -960
rect 1830 -972 1836 -966
rect 1830 -978 1836 -972
rect 1830 -984 1836 -978
rect 1830 -990 1836 -984
rect 1830 -996 1836 -990
rect 1830 -1002 1836 -996
rect 1830 -1008 1836 -1002
rect 1830 -1014 1836 -1008
rect 1830 -1020 1836 -1014
rect 1830 -1026 1836 -1020
rect 1830 -1032 1836 -1026
rect 1830 -1038 1836 -1032
rect 1830 -1044 1836 -1038
rect 1830 -1050 1836 -1044
rect 1830 -1056 1836 -1050
rect 1830 -1062 1836 -1056
rect 1830 -1068 1836 -1062
rect 1830 -1074 1836 -1068
rect 1830 -1080 1836 -1074
rect 1830 -1086 1836 -1080
rect 1830 -1092 1836 -1086
rect 1830 -1098 1836 -1092
rect 1830 -1104 1836 -1098
rect 1830 -1110 1836 -1104
rect 1830 -1116 1836 -1110
rect 1830 -1122 1836 -1116
rect 1830 -1128 1836 -1122
rect 1830 -1134 1836 -1128
rect 1830 -1140 1836 -1134
rect 1830 -1146 1836 -1140
rect 1830 -1152 1836 -1146
rect 1830 -1158 1836 -1152
rect 1830 -1164 1836 -1158
rect 1830 -1170 1836 -1164
rect 1830 -1176 1836 -1170
rect 1830 -1182 1836 -1176
rect 1830 -1188 1836 -1182
rect 1830 -1194 1836 -1188
rect 1830 -1200 1836 -1194
rect 1830 -1206 1836 -1200
rect 1830 -1212 1836 -1206
rect 1830 -1218 1836 -1212
rect 1830 -1224 1836 -1218
rect 1830 -1230 1836 -1224
rect 1830 -1236 1836 -1230
rect 1830 -1242 1836 -1236
rect 1830 -1248 1836 -1242
rect 1830 -1254 1836 -1248
rect 1830 -1260 1836 -1254
rect 1830 -1266 1836 -1260
rect 1830 -1272 1836 -1266
rect 1830 -1278 1836 -1272
rect 1830 -1284 1836 -1278
rect 1830 -1290 1836 -1284
rect 1830 -1296 1836 -1290
rect 1830 -1302 1836 -1296
rect 1830 -1308 1836 -1302
rect 1830 -1314 1836 -1308
rect 1830 -1320 1836 -1314
rect 1830 -1326 1836 -1320
rect 1830 -1332 1836 -1326
rect 1830 -1338 1836 -1332
rect 1830 -1344 1836 -1338
rect 1830 -1350 1836 -1344
rect 1830 -1356 1836 -1350
rect 1830 -1362 1836 -1356
rect 1830 -1368 1836 -1362
rect 1830 -1374 1836 -1368
rect 1830 -1380 1836 -1374
rect 1830 -1386 1836 -1380
rect 1830 -1392 1836 -1386
rect 1830 -1398 1836 -1392
rect 1830 -1404 1836 -1398
rect 1830 -1410 1836 -1404
rect 1830 -1416 1836 -1410
rect 1830 -1422 1836 -1416
rect 1830 -1428 1836 -1422
rect 1830 -1434 1836 -1428
rect 1830 -1440 1836 -1434
rect 1830 -1446 1836 -1440
rect 1830 -1452 1836 -1446
rect 1830 -1458 1836 -1452
rect 1830 -1464 1836 -1458
rect 1830 -1470 1836 -1464
rect 1830 -1476 1836 -1470
rect 1830 -1482 1836 -1476
rect 1830 -1488 1836 -1482
rect 1830 -1494 1836 -1488
rect 1830 -1500 1836 -1494
rect 1830 -1506 1836 -1500
rect 1830 -1512 1836 -1506
rect 1830 -1518 1836 -1512
rect 1830 -1524 1836 -1518
rect 1830 -1530 1836 -1524
rect 1830 -1536 1836 -1530
rect 1830 -1542 1836 -1536
rect 1830 -1548 1836 -1542
rect 1830 -1554 1836 -1548
rect 1830 -1560 1836 -1554
rect 1830 -1566 1836 -1560
rect 1830 -1572 1836 -1566
rect 1830 -1578 1836 -1572
rect 1830 -1584 1836 -1578
rect 1830 -1590 1836 -1584
rect 1830 -1596 1836 -1590
rect 1830 -1602 1836 -1596
rect 1830 -1608 1836 -1602
rect 1830 -1614 1836 -1608
rect 1830 -1620 1836 -1614
rect 1830 -1626 1836 -1620
rect 1830 -1632 1836 -1626
rect 1830 -1638 1836 -1632
rect 1830 -1644 1836 -1638
rect 1830 -1650 1836 -1644
rect 1830 -1656 1836 -1650
rect 1830 -1662 1836 -1656
rect 1830 -1668 1836 -1662
rect 1830 -1674 1836 -1668
rect 1830 -1680 1836 -1674
rect 1830 -1686 1836 -1680
rect 1830 -1692 1836 -1686
rect 1830 -1698 1836 -1692
rect 1830 -1704 1836 -1698
rect 1830 -1710 1836 -1704
rect 1830 -1716 1836 -1710
rect 1830 -1722 1836 -1716
rect 1830 -1728 1836 -1722
rect 1830 -1734 1836 -1728
rect 1830 -1740 1836 -1734
rect 1830 -1746 1836 -1740
rect 1830 -1752 1836 -1746
rect 1830 -1758 1836 -1752
rect 1830 -1764 1836 -1758
rect 1830 -1770 1836 -1764
rect 1830 -1776 1836 -1770
rect 1830 -1782 1836 -1776
rect 1830 -1788 1836 -1782
rect 1830 -1794 1836 -1788
rect 1830 -1800 1836 -1794
rect 1830 -1806 1836 -1800
rect 1830 -1812 1836 -1806
rect 1830 -1818 1836 -1812
rect 1830 -1896 1836 -1890
rect 1830 -1902 1836 -1896
rect 1830 -1908 1836 -1902
rect 1830 -1914 1836 -1908
rect 1830 -1920 1836 -1914
rect 1830 -1926 1836 -1920
rect 1830 -1932 1836 -1926
rect 1830 -1938 1836 -1932
rect 1830 -1944 1836 -1938
rect 1830 -1950 1836 -1944
rect 1830 -1956 1836 -1950
rect 1830 -1962 1836 -1956
rect 1830 -1968 1836 -1962
rect 1830 -1974 1836 -1968
rect 1830 -1980 1836 -1974
rect 1830 -1986 1836 -1980
rect 1830 -1992 1836 -1986
rect 1830 -1998 1836 -1992
rect 1830 -2004 1836 -1998
rect 1830 -2010 1836 -2004
rect 1830 -2016 1836 -2010
rect 1830 -2022 1836 -2016
rect 1830 -2028 1836 -2022
rect 1830 -2034 1836 -2028
rect 1830 -2040 1836 -2034
rect 1830 -2046 1836 -2040
rect 1830 -2052 1836 -2046
rect 1830 -2058 1836 -2052
rect 1830 -2064 1836 -2058
rect 1830 -2070 1836 -2064
rect 1830 -2076 1836 -2070
rect 1830 -2082 1836 -2076
rect 1830 -2088 1836 -2082
rect 1830 -2094 1836 -2088
rect 1830 -2100 1836 -2094
rect 1830 -2106 1836 -2100
rect 1830 -2112 1836 -2106
rect 1830 -2118 1836 -2112
rect 1830 -2124 1836 -2118
rect 1830 -2130 1836 -2124
rect 1830 -2136 1836 -2130
rect 1830 -2142 1836 -2136
rect 1830 -2148 1836 -2142
rect 1830 -2154 1836 -2148
rect 1830 -2160 1836 -2154
rect 1830 -2166 1836 -2160
rect 1830 -2172 1836 -2166
rect 1830 -2178 1836 -2172
rect 1830 -2184 1836 -2178
rect 1830 -2190 1836 -2184
rect 1830 -2196 1836 -2190
rect 1830 -2202 1836 -2196
rect 1830 -2208 1836 -2202
rect 1830 -2214 1836 -2208
rect 1830 -2220 1836 -2214
rect 1830 -2226 1836 -2220
rect 1830 -2232 1836 -2226
rect 1830 -2238 1836 -2232
rect 1830 -2244 1836 -2238
rect 1830 -2250 1836 -2244
rect 1830 -2256 1836 -2250
rect 1830 -2262 1836 -2256
rect 1830 -2268 1836 -2262
rect 1830 -2274 1836 -2268
rect 1830 -2280 1836 -2274
rect 1830 -2286 1836 -2280
rect 1830 -2292 1836 -2286
rect 1830 -2298 1836 -2292
rect 1830 -2304 1836 -2298
rect 1830 -2310 1836 -2304
rect 1830 -2316 1836 -2310
rect 1830 -2322 1836 -2316
rect 1830 -2328 1836 -2322
rect 1830 -2334 1836 -2328
rect 1830 -2340 1836 -2334
rect 1830 -2346 1836 -2340
rect 1830 -2352 1836 -2346
rect 1830 -2358 1836 -2352
rect 1830 -2364 1836 -2358
rect 1830 -2370 1836 -2364
rect 1830 -2376 1836 -2370
rect 1830 -2382 1836 -2376
rect 1830 -2388 1836 -2382
rect 1830 -2394 1836 -2388
rect 1830 -2400 1836 -2394
rect 1830 -2406 1836 -2400
rect 1830 -2412 1836 -2406
rect 1830 -2418 1836 -2412
rect 1830 -2424 1836 -2418
rect 1830 -2430 1836 -2424
rect 1830 -2436 1836 -2430
rect 1830 -2442 1836 -2436
rect 1830 -2448 1836 -2442
rect 1830 -2454 1836 -2448
rect 1830 -2460 1836 -2454
rect 1830 -2466 1836 -2460
rect 1830 -2472 1836 -2466
rect 1830 -2478 1836 -2472
rect 1830 -2484 1836 -2478
rect 1830 -2490 1836 -2484
rect 1830 -2496 1836 -2490
rect 1830 -2502 1836 -2496
rect 1830 -2508 1836 -2502
rect 1830 -2514 1836 -2508
rect 1830 -2520 1836 -2514
rect 1830 -2526 1836 -2520
rect 1830 -2532 1836 -2526
rect 1830 -2538 1836 -2532
rect 1830 -2544 1836 -2538
rect 1830 -2550 1836 -2544
rect 1830 -2556 1836 -2550
rect 1830 -2562 1836 -2556
rect 1830 -2568 1836 -2562
rect 1830 -2574 1836 -2568
rect 1830 -2580 1836 -2574
rect 1830 -2586 1836 -2580
rect 1830 -2592 1836 -2586
rect 1830 -2598 1836 -2592
rect 1830 -2604 1836 -2598
rect 1830 -2610 1836 -2604
rect 1830 -2616 1836 -2610
rect 1830 -2688 1836 -2682
rect 1830 -2694 1836 -2688
rect 1830 -2700 1836 -2694
rect 1830 -2706 1836 -2700
rect 1830 -2712 1836 -2706
rect 1830 -2718 1836 -2712
rect 1830 -2724 1836 -2718
rect 1830 -2730 1836 -2724
rect 1830 -2736 1836 -2730
rect 1830 -2742 1836 -2736
rect 1830 -2748 1836 -2742
rect 1830 -2754 1836 -2748
rect 1830 -2760 1836 -2754
rect 1830 -2766 1836 -2760
rect 1830 -2772 1836 -2766
rect 1830 -2778 1836 -2772
rect 1830 -2784 1836 -2778
rect 1830 -2790 1836 -2784
rect 1830 -2796 1836 -2790
rect 1830 -2802 1836 -2796
rect 1830 -2808 1836 -2802
rect 1830 -2814 1836 -2808
rect 1830 -2820 1836 -2814
rect 1830 -2826 1836 -2820
rect 1830 -2832 1836 -2826
rect 1830 -2838 1836 -2832
rect 1830 -2844 1836 -2838
rect 1830 -2850 1836 -2844
rect 1830 -2856 1836 -2850
rect 1830 -2862 1836 -2856
rect 1830 -2868 1836 -2862
rect 1830 -2874 1836 -2868
rect 1830 -2880 1836 -2874
rect 1830 -2886 1836 -2880
rect 1830 -2892 1836 -2886
rect 1830 -2898 1836 -2892
rect 1830 -2904 1836 -2898
rect 1830 -2910 1836 -2904
rect 1830 -2916 1836 -2910
rect 1830 -2922 1836 -2916
rect 1830 -2928 1836 -2922
rect 1830 -2934 1836 -2928
rect 1830 -2940 1836 -2934
rect 1830 -2946 1836 -2940
rect 1830 -2952 1836 -2946
rect 1830 -2958 1836 -2952
rect 1830 -2964 1836 -2958
rect 1830 -2970 1836 -2964
rect 1830 -2976 1836 -2970
rect 1830 -2982 1836 -2976
rect 1830 -2988 1836 -2982
rect 1830 -2994 1836 -2988
rect 1830 -3000 1836 -2994
rect 1830 -3006 1836 -3000
rect 1830 -3012 1836 -3006
rect 1830 -3018 1836 -3012
rect 1830 -3024 1836 -3018
rect 1830 -3030 1836 -3024
rect 1830 -3036 1836 -3030
rect 1830 -3042 1836 -3036
rect 1830 -3048 1836 -3042
rect 1830 -3054 1836 -3048
rect 1830 -3060 1836 -3054
rect 1830 -3066 1836 -3060
rect 1830 -3072 1836 -3066
rect 1830 -3078 1836 -3072
rect 1830 -3084 1836 -3078
rect 1830 -3090 1836 -3084
rect 1830 -3096 1836 -3090
rect 1830 -3102 1836 -3096
rect 1830 -3108 1836 -3102
rect 1830 -3114 1836 -3108
rect 1830 -3120 1836 -3114
rect 1830 -3126 1836 -3120
rect 1830 -3132 1836 -3126
rect 1830 -3138 1836 -3132
rect 1830 -3144 1836 -3138
rect 1830 -3150 1836 -3144
rect 1830 -3156 1836 -3150
rect 1830 -3162 1836 -3156
rect 1830 -3168 1836 -3162
rect 1830 -3174 1836 -3168
rect 1830 -3222 1836 -3216
rect 1830 -3228 1836 -3222
rect 1830 -3234 1836 -3228
rect 1830 -3240 1836 -3234
rect 1830 -3246 1836 -3240
rect 1830 -3252 1836 -3246
rect 1830 -3258 1836 -3252
rect 1830 -3264 1836 -3258
rect 1830 -3270 1836 -3264
rect 1830 -3276 1836 -3270
rect 1830 -3282 1836 -3276
rect 1830 -3288 1836 -3282
rect 1830 -3294 1836 -3288
rect 1830 -3300 1836 -3294
rect 1830 -3306 1836 -3300
rect 1830 -3312 1836 -3306
rect 1830 -3318 1836 -3312
rect 1830 -3324 1836 -3318
rect 1830 -3330 1836 -3324
rect 1830 -3336 1836 -3330
rect 1830 -3342 1836 -3336
rect 1830 -3348 1836 -3342
rect 1836 -672 1842 -666
rect 1836 -678 1842 -672
rect 1836 -684 1842 -678
rect 1836 -690 1842 -684
rect 1836 -696 1842 -690
rect 1836 -702 1842 -696
rect 1836 -708 1842 -702
rect 1836 -714 1842 -708
rect 1836 -720 1842 -714
rect 1836 -726 1842 -720
rect 1836 -732 1842 -726
rect 1836 -738 1842 -732
rect 1836 -744 1842 -738
rect 1836 -750 1842 -744
rect 1836 -756 1842 -750
rect 1836 -762 1842 -756
rect 1836 -768 1842 -762
rect 1836 -774 1842 -768
rect 1836 -780 1842 -774
rect 1836 -786 1842 -780
rect 1836 -792 1842 -786
rect 1836 -798 1842 -792
rect 1836 -804 1842 -798
rect 1836 -810 1842 -804
rect 1836 -816 1842 -810
rect 1836 -822 1842 -816
rect 1836 -828 1842 -822
rect 1836 -834 1842 -828
rect 1836 -840 1842 -834
rect 1836 -846 1842 -840
rect 1836 -852 1842 -846
rect 1836 -858 1842 -852
rect 1836 -864 1842 -858
rect 1836 -870 1842 -864
rect 1836 -876 1842 -870
rect 1836 -882 1842 -876
rect 1836 -888 1842 -882
rect 1836 -894 1842 -888
rect 1836 -900 1842 -894
rect 1836 -906 1842 -900
rect 1836 -912 1842 -906
rect 1836 -918 1842 -912
rect 1836 -924 1842 -918
rect 1836 -930 1842 -924
rect 1836 -936 1842 -930
rect 1836 -942 1842 -936
rect 1836 -948 1842 -942
rect 1836 -954 1842 -948
rect 1836 -960 1842 -954
rect 1836 -966 1842 -960
rect 1836 -972 1842 -966
rect 1836 -978 1842 -972
rect 1836 -984 1842 -978
rect 1836 -990 1842 -984
rect 1836 -996 1842 -990
rect 1836 -1002 1842 -996
rect 1836 -1008 1842 -1002
rect 1836 -1014 1842 -1008
rect 1836 -1020 1842 -1014
rect 1836 -1026 1842 -1020
rect 1836 -1032 1842 -1026
rect 1836 -1038 1842 -1032
rect 1836 -1044 1842 -1038
rect 1836 -1050 1842 -1044
rect 1836 -1056 1842 -1050
rect 1836 -1062 1842 -1056
rect 1836 -1068 1842 -1062
rect 1836 -1074 1842 -1068
rect 1836 -1080 1842 -1074
rect 1836 -1086 1842 -1080
rect 1836 -1092 1842 -1086
rect 1836 -1098 1842 -1092
rect 1836 -1104 1842 -1098
rect 1836 -1110 1842 -1104
rect 1836 -1116 1842 -1110
rect 1836 -1122 1842 -1116
rect 1836 -1128 1842 -1122
rect 1836 -1134 1842 -1128
rect 1836 -1140 1842 -1134
rect 1836 -1146 1842 -1140
rect 1836 -1152 1842 -1146
rect 1836 -1158 1842 -1152
rect 1836 -1164 1842 -1158
rect 1836 -1170 1842 -1164
rect 1836 -1176 1842 -1170
rect 1836 -1182 1842 -1176
rect 1836 -1188 1842 -1182
rect 1836 -1194 1842 -1188
rect 1836 -1200 1842 -1194
rect 1836 -1206 1842 -1200
rect 1836 -1212 1842 -1206
rect 1836 -1218 1842 -1212
rect 1836 -1224 1842 -1218
rect 1836 -1230 1842 -1224
rect 1836 -1236 1842 -1230
rect 1836 -1242 1842 -1236
rect 1836 -1248 1842 -1242
rect 1836 -1254 1842 -1248
rect 1836 -1260 1842 -1254
rect 1836 -1266 1842 -1260
rect 1836 -1272 1842 -1266
rect 1836 -1278 1842 -1272
rect 1836 -1284 1842 -1278
rect 1836 -1290 1842 -1284
rect 1836 -1296 1842 -1290
rect 1836 -1302 1842 -1296
rect 1836 -1308 1842 -1302
rect 1836 -1314 1842 -1308
rect 1836 -1320 1842 -1314
rect 1836 -1326 1842 -1320
rect 1836 -1332 1842 -1326
rect 1836 -1338 1842 -1332
rect 1836 -1344 1842 -1338
rect 1836 -1350 1842 -1344
rect 1836 -1356 1842 -1350
rect 1836 -1362 1842 -1356
rect 1836 -1368 1842 -1362
rect 1836 -1374 1842 -1368
rect 1836 -1380 1842 -1374
rect 1836 -1386 1842 -1380
rect 1836 -1392 1842 -1386
rect 1836 -1398 1842 -1392
rect 1836 -1404 1842 -1398
rect 1836 -1410 1842 -1404
rect 1836 -1416 1842 -1410
rect 1836 -1422 1842 -1416
rect 1836 -1428 1842 -1422
rect 1836 -1434 1842 -1428
rect 1836 -1440 1842 -1434
rect 1836 -1446 1842 -1440
rect 1836 -1452 1842 -1446
rect 1836 -1458 1842 -1452
rect 1836 -1464 1842 -1458
rect 1836 -1470 1842 -1464
rect 1836 -1476 1842 -1470
rect 1836 -1482 1842 -1476
rect 1836 -1488 1842 -1482
rect 1836 -1494 1842 -1488
rect 1836 -1500 1842 -1494
rect 1836 -1506 1842 -1500
rect 1836 -1512 1842 -1506
rect 1836 -1518 1842 -1512
rect 1836 -1524 1842 -1518
rect 1836 -1530 1842 -1524
rect 1836 -1536 1842 -1530
rect 1836 -1542 1842 -1536
rect 1836 -1548 1842 -1542
rect 1836 -1554 1842 -1548
rect 1836 -1560 1842 -1554
rect 1836 -1566 1842 -1560
rect 1836 -1572 1842 -1566
rect 1836 -1578 1842 -1572
rect 1836 -1584 1842 -1578
rect 1836 -1590 1842 -1584
rect 1836 -1596 1842 -1590
rect 1836 -1602 1842 -1596
rect 1836 -1608 1842 -1602
rect 1836 -1614 1842 -1608
rect 1836 -1620 1842 -1614
rect 1836 -1626 1842 -1620
rect 1836 -1632 1842 -1626
rect 1836 -1638 1842 -1632
rect 1836 -1644 1842 -1638
rect 1836 -1650 1842 -1644
rect 1836 -1656 1842 -1650
rect 1836 -1662 1842 -1656
rect 1836 -1668 1842 -1662
rect 1836 -1674 1842 -1668
rect 1836 -1680 1842 -1674
rect 1836 -1686 1842 -1680
rect 1836 -1692 1842 -1686
rect 1836 -1698 1842 -1692
rect 1836 -1704 1842 -1698
rect 1836 -1710 1842 -1704
rect 1836 -1716 1842 -1710
rect 1836 -1722 1842 -1716
rect 1836 -1728 1842 -1722
rect 1836 -1734 1842 -1728
rect 1836 -1740 1842 -1734
rect 1836 -1746 1842 -1740
rect 1836 -1752 1842 -1746
rect 1836 -1758 1842 -1752
rect 1836 -1764 1842 -1758
rect 1836 -1770 1842 -1764
rect 1836 -1776 1842 -1770
rect 1836 -1782 1842 -1776
rect 1836 -1788 1842 -1782
rect 1836 -1794 1842 -1788
rect 1836 -1800 1842 -1794
rect 1836 -1806 1842 -1800
rect 1836 -1812 1842 -1806
rect 1836 -1890 1842 -1884
rect 1836 -1896 1842 -1890
rect 1836 -1902 1842 -1896
rect 1836 -1908 1842 -1902
rect 1836 -1914 1842 -1908
rect 1836 -1920 1842 -1914
rect 1836 -1926 1842 -1920
rect 1836 -1932 1842 -1926
rect 1836 -1938 1842 -1932
rect 1836 -1944 1842 -1938
rect 1836 -1950 1842 -1944
rect 1836 -1956 1842 -1950
rect 1836 -1962 1842 -1956
rect 1836 -1968 1842 -1962
rect 1836 -1974 1842 -1968
rect 1836 -1980 1842 -1974
rect 1836 -1986 1842 -1980
rect 1836 -1992 1842 -1986
rect 1836 -1998 1842 -1992
rect 1836 -2004 1842 -1998
rect 1836 -2010 1842 -2004
rect 1836 -2016 1842 -2010
rect 1836 -2022 1842 -2016
rect 1836 -2028 1842 -2022
rect 1836 -2034 1842 -2028
rect 1836 -2040 1842 -2034
rect 1836 -2046 1842 -2040
rect 1836 -2052 1842 -2046
rect 1836 -2058 1842 -2052
rect 1836 -2064 1842 -2058
rect 1836 -2070 1842 -2064
rect 1836 -2076 1842 -2070
rect 1836 -2082 1842 -2076
rect 1836 -2088 1842 -2082
rect 1836 -2094 1842 -2088
rect 1836 -2100 1842 -2094
rect 1836 -2106 1842 -2100
rect 1836 -2112 1842 -2106
rect 1836 -2118 1842 -2112
rect 1836 -2124 1842 -2118
rect 1836 -2130 1842 -2124
rect 1836 -2136 1842 -2130
rect 1836 -2142 1842 -2136
rect 1836 -2148 1842 -2142
rect 1836 -2154 1842 -2148
rect 1836 -2160 1842 -2154
rect 1836 -2166 1842 -2160
rect 1836 -2172 1842 -2166
rect 1836 -2178 1842 -2172
rect 1836 -2184 1842 -2178
rect 1836 -2190 1842 -2184
rect 1836 -2196 1842 -2190
rect 1836 -2202 1842 -2196
rect 1836 -2208 1842 -2202
rect 1836 -2214 1842 -2208
rect 1836 -2220 1842 -2214
rect 1836 -2226 1842 -2220
rect 1836 -2232 1842 -2226
rect 1836 -2238 1842 -2232
rect 1836 -2244 1842 -2238
rect 1836 -2250 1842 -2244
rect 1836 -2256 1842 -2250
rect 1836 -2262 1842 -2256
rect 1836 -2268 1842 -2262
rect 1836 -2274 1842 -2268
rect 1836 -2280 1842 -2274
rect 1836 -2286 1842 -2280
rect 1836 -2292 1842 -2286
rect 1836 -2298 1842 -2292
rect 1836 -2304 1842 -2298
rect 1836 -2310 1842 -2304
rect 1836 -2316 1842 -2310
rect 1836 -2322 1842 -2316
rect 1836 -2328 1842 -2322
rect 1836 -2334 1842 -2328
rect 1836 -2340 1842 -2334
rect 1836 -2346 1842 -2340
rect 1836 -2352 1842 -2346
rect 1836 -2358 1842 -2352
rect 1836 -2364 1842 -2358
rect 1836 -2370 1842 -2364
rect 1836 -2376 1842 -2370
rect 1836 -2382 1842 -2376
rect 1836 -2388 1842 -2382
rect 1836 -2394 1842 -2388
rect 1836 -2400 1842 -2394
rect 1836 -2406 1842 -2400
rect 1836 -2412 1842 -2406
rect 1836 -2418 1842 -2412
rect 1836 -2424 1842 -2418
rect 1836 -2430 1842 -2424
rect 1836 -2436 1842 -2430
rect 1836 -2442 1842 -2436
rect 1836 -2448 1842 -2442
rect 1836 -2454 1842 -2448
rect 1836 -2460 1842 -2454
rect 1836 -2466 1842 -2460
rect 1836 -2472 1842 -2466
rect 1836 -2478 1842 -2472
rect 1836 -2484 1842 -2478
rect 1836 -2490 1842 -2484
rect 1836 -2496 1842 -2490
rect 1836 -2502 1842 -2496
rect 1836 -2508 1842 -2502
rect 1836 -2514 1842 -2508
rect 1836 -2520 1842 -2514
rect 1836 -2526 1842 -2520
rect 1836 -2532 1842 -2526
rect 1836 -2538 1842 -2532
rect 1836 -2544 1842 -2538
rect 1836 -2550 1842 -2544
rect 1836 -2556 1842 -2550
rect 1836 -2562 1842 -2556
rect 1836 -2568 1842 -2562
rect 1836 -2574 1842 -2568
rect 1836 -2580 1842 -2574
rect 1836 -2586 1842 -2580
rect 1836 -2592 1842 -2586
rect 1836 -2598 1842 -2592
rect 1836 -2604 1842 -2598
rect 1836 -2610 1842 -2604
rect 1836 -2688 1842 -2682
rect 1836 -2694 1842 -2688
rect 1836 -2700 1842 -2694
rect 1836 -2706 1842 -2700
rect 1836 -2712 1842 -2706
rect 1836 -2718 1842 -2712
rect 1836 -2724 1842 -2718
rect 1836 -2730 1842 -2724
rect 1836 -2736 1842 -2730
rect 1836 -2742 1842 -2736
rect 1836 -2748 1842 -2742
rect 1836 -2754 1842 -2748
rect 1836 -2760 1842 -2754
rect 1836 -2766 1842 -2760
rect 1836 -2772 1842 -2766
rect 1836 -2778 1842 -2772
rect 1836 -2784 1842 -2778
rect 1836 -2790 1842 -2784
rect 1836 -2796 1842 -2790
rect 1836 -2802 1842 -2796
rect 1836 -2808 1842 -2802
rect 1836 -2814 1842 -2808
rect 1836 -2820 1842 -2814
rect 1836 -2826 1842 -2820
rect 1836 -2832 1842 -2826
rect 1836 -2838 1842 -2832
rect 1836 -2844 1842 -2838
rect 1836 -2850 1842 -2844
rect 1836 -2856 1842 -2850
rect 1836 -2862 1842 -2856
rect 1836 -2868 1842 -2862
rect 1836 -2874 1842 -2868
rect 1836 -2880 1842 -2874
rect 1836 -2886 1842 -2880
rect 1836 -2892 1842 -2886
rect 1836 -2898 1842 -2892
rect 1836 -2904 1842 -2898
rect 1836 -2910 1842 -2904
rect 1836 -2916 1842 -2910
rect 1836 -2922 1842 -2916
rect 1836 -2928 1842 -2922
rect 1836 -2934 1842 -2928
rect 1836 -2940 1842 -2934
rect 1836 -2946 1842 -2940
rect 1836 -2952 1842 -2946
rect 1836 -2958 1842 -2952
rect 1836 -2964 1842 -2958
rect 1836 -2970 1842 -2964
rect 1836 -2976 1842 -2970
rect 1836 -2982 1842 -2976
rect 1836 -2988 1842 -2982
rect 1836 -2994 1842 -2988
rect 1836 -3000 1842 -2994
rect 1836 -3006 1842 -3000
rect 1836 -3012 1842 -3006
rect 1836 -3018 1842 -3012
rect 1836 -3024 1842 -3018
rect 1836 -3030 1842 -3024
rect 1836 -3036 1842 -3030
rect 1836 -3042 1842 -3036
rect 1836 -3048 1842 -3042
rect 1836 -3054 1842 -3048
rect 1836 -3060 1842 -3054
rect 1836 -3066 1842 -3060
rect 1836 -3072 1842 -3066
rect 1836 -3078 1842 -3072
rect 1836 -3084 1842 -3078
rect 1836 -3090 1842 -3084
rect 1836 -3096 1842 -3090
rect 1836 -3102 1842 -3096
rect 1836 -3108 1842 -3102
rect 1836 -3114 1842 -3108
rect 1836 -3120 1842 -3114
rect 1836 -3126 1842 -3120
rect 1836 -3132 1842 -3126
rect 1836 -3138 1842 -3132
rect 1836 -3144 1842 -3138
rect 1836 -3150 1842 -3144
rect 1836 -3156 1842 -3150
rect 1836 -3162 1842 -3156
rect 1836 -3168 1842 -3162
rect 1836 -3222 1842 -3216
rect 1836 -3228 1842 -3222
rect 1836 -3234 1842 -3228
rect 1836 -3240 1842 -3234
rect 1836 -3246 1842 -3240
rect 1836 -3252 1842 -3246
rect 1836 -3258 1842 -3252
rect 1836 -3264 1842 -3258
rect 1836 -3270 1842 -3264
rect 1836 -3276 1842 -3270
rect 1836 -3282 1842 -3276
rect 1836 -3288 1842 -3282
rect 1836 -3294 1842 -3288
rect 1836 -3300 1842 -3294
rect 1836 -3306 1842 -3300
rect 1836 -3312 1842 -3306
rect 1836 -3318 1842 -3312
rect 1836 -3324 1842 -3318
rect 1836 -3330 1842 -3324
rect 1836 -3336 1842 -3330
rect 1836 -3342 1842 -3336
rect 1836 -3348 1842 -3342
rect 1842 -660 1848 -654
rect 1842 -666 1848 -660
rect 1842 -672 1848 -666
rect 1842 -678 1848 -672
rect 1842 -684 1848 -678
rect 1842 -690 1848 -684
rect 1842 -696 1848 -690
rect 1842 -702 1848 -696
rect 1842 -708 1848 -702
rect 1842 -714 1848 -708
rect 1842 -720 1848 -714
rect 1842 -726 1848 -720
rect 1842 -732 1848 -726
rect 1842 -738 1848 -732
rect 1842 -744 1848 -738
rect 1842 -750 1848 -744
rect 1842 -756 1848 -750
rect 1842 -762 1848 -756
rect 1842 -768 1848 -762
rect 1842 -774 1848 -768
rect 1842 -780 1848 -774
rect 1842 -786 1848 -780
rect 1842 -792 1848 -786
rect 1842 -798 1848 -792
rect 1842 -804 1848 -798
rect 1842 -810 1848 -804
rect 1842 -816 1848 -810
rect 1842 -822 1848 -816
rect 1842 -828 1848 -822
rect 1842 -834 1848 -828
rect 1842 -840 1848 -834
rect 1842 -846 1848 -840
rect 1842 -852 1848 -846
rect 1842 -858 1848 -852
rect 1842 -864 1848 -858
rect 1842 -870 1848 -864
rect 1842 -876 1848 -870
rect 1842 -882 1848 -876
rect 1842 -888 1848 -882
rect 1842 -894 1848 -888
rect 1842 -900 1848 -894
rect 1842 -906 1848 -900
rect 1842 -912 1848 -906
rect 1842 -918 1848 -912
rect 1842 -924 1848 -918
rect 1842 -930 1848 -924
rect 1842 -936 1848 -930
rect 1842 -942 1848 -936
rect 1842 -948 1848 -942
rect 1842 -954 1848 -948
rect 1842 -960 1848 -954
rect 1842 -966 1848 -960
rect 1842 -972 1848 -966
rect 1842 -978 1848 -972
rect 1842 -984 1848 -978
rect 1842 -990 1848 -984
rect 1842 -996 1848 -990
rect 1842 -1002 1848 -996
rect 1842 -1008 1848 -1002
rect 1842 -1014 1848 -1008
rect 1842 -1020 1848 -1014
rect 1842 -1026 1848 -1020
rect 1842 -1032 1848 -1026
rect 1842 -1038 1848 -1032
rect 1842 -1044 1848 -1038
rect 1842 -1050 1848 -1044
rect 1842 -1056 1848 -1050
rect 1842 -1062 1848 -1056
rect 1842 -1068 1848 -1062
rect 1842 -1074 1848 -1068
rect 1842 -1080 1848 -1074
rect 1842 -1086 1848 -1080
rect 1842 -1092 1848 -1086
rect 1842 -1098 1848 -1092
rect 1842 -1104 1848 -1098
rect 1842 -1110 1848 -1104
rect 1842 -1116 1848 -1110
rect 1842 -1122 1848 -1116
rect 1842 -1128 1848 -1122
rect 1842 -1134 1848 -1128
rect 1842 -1140 1848 -1134
rect 1842 -1146 1848 -1140
rect 1842 -1152 1848 -1146
rect 1842 -1158 1848 -1152
rect 1842 -1164 1848 -1158
rect 1842 -1170 1848 -1164
rect 1842 -1176 1848 -1170
rect 1842 -1182 1848 -1176
rect 1842 -1188 1848 -1182
rect 1842 -1194 1848 -1188
rect 1842 -1200 1848 -1194
rect 1842 -1206 1848 -1200
rect 1842 -1212 1848 -1206
rect 1842 -1218 1848 -1212
rect 1842 -1224 1848 -1218
rect 1842 -1230 1848 -1224
rect 1842 -1236 1848 -1230
rect 1842 -1242 1848 -1236
rect 1842 -1248 1848 -1242
rect 1842 -1254 1848 -1248
rect 1842 -1260 1848 -1254
rect 1842 -1266 1848 -1260
rect 1842 -1272 1848 -1266
rect 1842 -1278 1848 -1272
rect 1842 -1284 1848 -1278
rect 1842 -1290 1848 -1284
rect 1842 -1296 1848 -1290
rect 1842 -1302 1848 -1296
rect 1842 -1308 1848 -1302
rect 1842 -1314 1848 -1308
rect 1842 -1320 1848 -1314
rect 1842 -1326 1848 -1320
rect 1842 -1332 1848 -1326
rect 1842 -1338 1848 -1332
rect 1842 -1344 1848 -1338
rect 1842 -1350 1848 -1344
rect 1842 -1356 1848 -1350
rect 1842 -1362 1848 -1356
rect 1842 -1368 1848 -1362
rect 1842 -1374 1848 -1368
rect 1842 -1380 1848 -1374
rect 1842 -1386 1848 -1380
rect 1842 -1392 1848 -1386
rect 1842 -1398 1848 -1392
rect 1842 -1404 1848 -1398
rect 1842 -1410 1848 -1404
rect 1842 -1416 1848 -1410
rect 1842 -1422 1848 -1416
rect 1842 -1428 1848 -1422
rect 1842 -1434 1848 -1428
rect 1842 -1440 1848 -1434
rect 1842 -1446 1848 -1440
rect 1842 -1452 1848 -1446
rect 1842 -1458 1848 -1452
rect 1842 -1464 1848 -1458
rect 1842 -1470 1848 -1464
rect 1842 -1476 1848 -1470
rect 1842 -1482 1848 -1476
rect 1842 -1488 1848 -1482
rect 1842 -1494 1848 -1488
rect 1842 -1500 1848 -1494
rect 1842 -1506 1848 -1500
rect 1842 -1512 1848 -1506
rect 1842 -1518 1848 -1512
rect 1842 -1524 1848 -1518
rect 1842 -1530 1848 -1524
rect 1842 -1536 1848 -1530
rect 1842 -1542 1848 -1536
rect 1842 -1548 1848 -1542
rect 1842 -1554 1848 -1548
rect 1842 -1560 1848 -1554
rect 1842 -1566 1848 -1560
rect 1842 -1572 1848 -1566
rect 1842 -1578 1848 -1572
rect 1842 -1584 1848 -1578
rect 1842 -1590 1848 -1584
rect 1842 -1596 1848 -1590
rect 1842 -1602 1848 -1596
rect 1842 -1608 1848 -1602
rect 1842 -1614 1848 -1608
rect 1842 -1620 1848 -1614
rect 1842 -1626 1848 -1620
rect 1842 -1632 1848 -1626
rect 1842 -1638 1848 -1632
rect 1842 -1644 1848 -1638
rect 1842 -1650 1848 -1644
rect 1842 -1656 1848 -1650
rect 1842 -1662 1848 -1656
rect 1842 -1668 1848 -1662
rect 1842 -1674 1848 -1668
rect 1842 -1680 1848 -1674
rect 1842 -1686 1848 -1680
rect 1842 -1692 1848 -1686
rect 1842 -1698 1848 -1692
rect 1842 -1704 1848 -1698
rect 1842 -1710 1848 -1704
rect 1842 -1716 1848 -1710
rect 1842 -1722 1848 -1716
rect 1842 -1728 1848 -1722
rect 1842 -1734 1848 -1728
rect 1842 -1740 1848 -1734
rect 1842 -1746 1848 -1740
rect 1842 -1752 1848 -1746
rect 1842 -1758 1848 -1752
rect 1842 -1764 1848 -1758
rect 1842 -1770 1848 -1764
rect 1842 -1776 1848 -1770
rect 1842 -1782 1848 -1776
rect 1842 -1788 1848 -1782
rect 1842 -1794 1848 -1788
rect 1842 -1800 1848 -1794
rect 1842 -1806 1848 -1800
rect 1842 -1884 1848 -1878
rect 1842 -1890 1848 -1884
rect 1842 -1896 1848 -1890
rect 1842 -1902 1848 -1896
rect 1842 -1908 1848 -1902
rect 1842 -1914 1848 -1908
rect 1842 -1920 1848 -1914
rect 1842 -1926 1848 -1920
rect 1842 -1932 1848 -1926
rect 1842 -1938 1848 -1932
rect 1842 -1944 1848 -1938
rect 1842 -1950 1848 -1944
rect 1842 -1956 1848 -1950
rect 1842 -1962 1848 -1956
rect 1842 -1968 1848 -1962
rect 1842 -1974 1848 -1968
rect 1842 -1980 1848 -1974
rect 1842 -1986 1848 -1980
rect 1842 -1992 1848 -1986
rect 1842 -1998 1848 -1992
rect 1842 -2004 1848 -1998
rect 1842 -2010 1848 -2004
rect 1842 -2016 1848 -2010
rect 1842 -2022 1848 -2016
rect 1842 -2028 1848 -2022
rect 1842 -2034 1848 -2028
rect 1842 -2040 1848 -2034
rect 1842 -2046 1848 -2040
rect 1842 -2052 1848 -2046
rect 1842 -2058 1848 -2052
rect 1842 -2064 1848 -2058
rect 1842 -2070 1848 -2064
rect 1842 -2076 1848 -2070
rect 1842 -2082 1848 -2076
rect 1842 -2088 1848 -2082
rect 1842 -2094 1848 -2088
rect 1842 -2100 1848 -2094
rect 1842 -2106 1848 -2100
rect 1842 -2112 1848 -2106
rect 1842 -2118 1848 -2112
rect 1842 -2124 1848 -2118
rect 1842 -2130 1848 -2124
rect 1842 -2136 1848 -2130
rect 1842 -2142 1848 -2136
rect 1842 -2148 1848 -2142
rect 1842 -2154 1848 -2148
rect 1842 -2160 1848 -2154
rect 1842 -2166 1848 -2160
rect 1842 -2172 1848 -2166
rect 1842 -2178 1848 -2172
rect 1842 -2184 1848 -2178
rect 1842 -2190 1848 -2184
rect 1842 -2196 1848 -2190
rect 1842 -2202 1848 -2196
rect 1842 -2208 1848 -2202
rect 1842 -2214 1848 -2208
rect 1842 -2220 1848 -2214
rect 1842 -2226 1848 -2220
rect 1842 -2232 1848 -2226
rect 1842 -2238 1848 -2232
rect 1842 -2244 1848 -2238
rect 1842 -2250 1848 -2244
rect 1842 -2256 1848 -2250
rect 1842 -2262 1848 -2256
rect 1842 -2268 1848 -2262
rect 1842 -2274 1848 -2268
rect 1842 -2280 1848 -2274
rect 1842 -2286 1848 -2280
rect 1842 -2292 1848 -2286
rect 1842 -2298 1848 -2292
rect 1842 -2304 1848 -2298
rect 1842 -2310 1848 -2304
rect 1842 -2316 1848 -2310
rect 1842 -2322 1848 -2316
rect 1842 -2328 1848 -2322
rect 1842 -2334 1848 -2328
rect 1842 -2340 1848 -2334
rect 1842 -2346 1848 -2340
rect 1842 -2352 1848 -2346
rect 1842 -2358 1848 -2352
rect 1842 -2364 1848 -2358
rect 1842 -2370 1848 -2364
rect 1842 -2376 1848 -2370
rect 1842 -2382 1848 -2376
rect 1842 -2388 1848 -2382
rect 1842 -2394 1848 -2388
rect 1842 -2400 1848 -2394
rect 1842 -2406 1848 -2400
rect 1842 -2412 1848 -2406
rect 1842 -2418 1848 -2412
rect 1842 -2424 1848 -2418
rect 1842 -2430 1848 -2424
rect 1842 -2436 1848 -2430
rect 1842 -2442 1848 -2436
rect 1842 -2448 1848 -2442
rect 1842 -2454 1848 -2448
rect 1842 -2460 1848 -2454
rect 1842 -2466 1848 -2460
rect 1842 -2472 1848 -2466
rect 1842 -2478 1848 -2472
rect 1842 -2484 1848 -2478
rect 1842 -2490 1848 -2484
rect 1842 -2496 1848 -2490
rect 1842 -2502 1848 -2496
rect 1842 -2508 1848 -2502
rect 1842 -2514 1848 -2508
rect 1842 -2520 1848 -2514
rect 1842 -2526 1848 -2520
rect 1842 -2532 1848 -2526
rect 1842 -2538 1848 -2532
rect 1842 -2544 1848 -2538
rect 1842 -2550 1848 -2544
rect 1842 -2556 1848 -2550
rect 1842 -2562 1848 -2556
rect 1842 -2568 1848 -2562
rect 1842 -2574 1848 -2568
rect 1842 -2580 1848 -2574
rect 1842 -2586 1848 -2580
rect 1842 -2592 1848 -2586
rect 1842 -2598 1848 -2592
rect 1842 -2604 1848 -2598
rect 1842 -2610 1848 -2604
rect 1842 -2682 1848 -2676
rect 1842 -2688 1848 -2682
rect 1842 -2694 1848 -2688
rect 1842 -2700 1848 -2694
rect 1842 -2706 1848 -2700
rect 1842 -2712 1848 -2706
rect 1842 -2718 1848 -2712
rect 1842 -2724 1848 -2718
rect 1842 -2730 1848 -2724
rect 1842 -2736 1848 -2730
rect 1842 -2742 1848 -2736
rect 1842 -2748 1848 -2742
rect 1842 -2754 1848 -2748
rect 1842 -2760 1848 -2754
rect 1842 -2766 1848 -2760
rect 1842 -2772 1848 -2766
rect 1842 -2778 1848 -2772
rect 1842 -2784 1848 -2778
rect 1842 -2790 1848 -2784
rect 1842 -2796 1848 -2790
rect 1842 -2802 1848 -2796
rect 1842 -2808 1848 -2802
rect 1842 -2814 1848 -2808
rect 1842 -2820 1848 -2814
rect 1842 -2826 1848 -2820
rect 1842 -2832 1848 -2826
rect 1842 -2838 1848 -2832
rect 1842 -2844 1848 -2838
rect 1842 -2850 1848 -2844
rect 1842 -2856 1848 -2850
rect 1842 -2862 1848 -2856
rect 1842 -2868 1848 -2862
rect 1842 -2874 1848 -2868
rect 1842 -2880 1848 -2874
rect 1842 -2886 1848 -2880
rect 1842 -2892 1848 -2886
rect 1842 -2898 1848 -2892
rect 1842 -2904 1848 -2898
rect 1842 -2910 1848 -2904
rect 1842 -2916 1848 -2910
rect 1842 -2922 1848 -2916
rect 1842 -2928 1848 -2922
rect 1842 -2934 1848 -2928
rect 1842 -2940 1848 -2934
rect 1842 -2946 1848 -2940
rect 1842 -2952 1848 -2946
rect 1842 -2958 1848 -2952
rect 1842 -2964 1848 -2958
rect 1842 -2970 1848 -2964
rect 1842 -2976 1848 -2970
rect 1842 -2982 1848 -2976
rect 1842 -2988 1848 -2982
rect 1842 -2994 1848 -2988
rect 1842 -3000 1848 -2994
rect 1842 -3006 1848 -3000
rect 1842 -3012 1848 -3006
rect 1842 -3018 1848 -3012
rect 1842 -3024 1848 -3018
rect 1842 -3030 1848 -3024
rect 1842 -3036 1848 -3030
rect 1842 -3042 1848 -3036
rect 1842 -3048 1848 -3042
rect 1842 -3054 1848 -3048
rect 1842 -3060 1848 -3054
rect 1842 -3066 1848 -3060
rect 1842 -3072 1848 -3066
rect 1842 -3078 1848 -3072
rect 1842 -3084 1848 -3078
rect 1842 -3090 1848 -3084
rect 1842 -3096 1848 -3090
rect 1842 -3102 1848 -3096
rect 1842 -3108 1848 -3102
rect 1842 -3114 1848 -3108
rect 1842 -3120 1848 -3114
rect 1842 -3126 1848 -3120
rect 1842 -3132 1848 -3126
rect 1842 -3138 1848 -3132
rect 1842 -3144 1848 -3138
rect 1842 -3150 1848 -3144
rect 1842 -3156 1848 -3150
rect 1842 -3162 1848 -3156
rect 1842 -3168 1848 -3162
rect 1842 -3216 1848 -3210
rect 1842 -3222 1848 -3216
rect 1842 -3228 1848 -3222
rect 1842 -3234 1848 -3228
rect 1842 -3240 1848 -3234
rect 1842 -3246 1848 -3240
rect 1842 -3252 1848 -3246
rect 1842 -3258 1848 -3252
rect 1842 -3264 1848 -3258
rect 1842 -3270 1848 -3264
rect 1842 -3276 1848 -3270
rect 1842 -3282 1848 -3276
rect 1842 -3288 1848 -3282
rect 1842 -3294 1848 -3288
rect 1842 -3300 1848 -3294
rect 1842 -3306 1848 -3300
rect 1842 -3312 1848 -3306
rect 1842 -3318 1848 -3312
rect 1842 -3324 1848 -3318
rect 1842 -3330 1848 -3324
rect 1842 -3336 1848 -3330
rect 1842 -3342 1848 -3336
rect 1848 -654 1854 -648
rect 1848 -660 1854 -654
rect 1848 -666 1854 -660
rect 1848 -672 1854 -666
rect 1848 -678 1854 -672
rect 1848 -684 1854 -678
rect 1848 -690 1854 -684
rect 1848 -696 1854 -690
rect 1848 -702 1854 -696
rect 1848 -708 1854 -702
rect 1848 -714 1854 -708
rect 1848 -720 1854 -714
rect 1848 -726 1854 -720
rect 1848 -732 1854 -726
rect 1848 -738 1854 -732
rect 1848 -744 1854 -738
rect 1848 -750 1854 -744
rect 1848 -756 1854 -750
rect 1848 -762 1854 -756
rect 1848 -768 1854 -762
rect 1848 -774 1854 -768
rect 1848 -780 1854 -774
rect 1848 -786 1854 -780
rect 1848 -792 1854 -786
rect 1848 -798 1854 -792
rect 1848 -804 1854 -798
rect 1848 -810 1854 -804
rect 1848 -816 1854 -810
rect 1848 -822 1854 -816
rect 1848 -828 1854 -822
rect 1848 -834 1854 -828
rect 1848 -840 1854 -834
rect 1848 -846 1854 -840
rect 1848 -852 1854 -846
rect 1848 -858 1854 -852
rect 1848 -864 1854 -858
rect 1848 -870 1854 -864
rect 1848 -876 1854 -870
rect 1848 -882 1854 -876
rect 1848 -888 1854 -882
rect 1848 -894 1854 -888
rect 1848 -900 1854 -894
rect 1848 -906 1854 -900
rect 1848 -912 1854 -906
rect 1848 -918 1854 -912
rect 1848 -924 1854 -918
rect 1848 -930 1854 -924
rect 1848 -936 1854 -930
rect 1848 -942 1854 -936
rect 1848 -948 1854 -942
rect 1848 -954 1854 -948
rect 1848 -960 1854 -954
rect 1848 -966 1854 -960
rect 1848 -972 1854 -966
rect 1848 -978 1854 -972
rect 1848 -984 1854 -978
rect 1848 -990 1854 -984
rect 1848 -996 1854 -990
rect 1848 -1002 1854 -996
rect 1848 -1008 1854 -1002
rect 1848 -1014 1854 -1008
rect 1848 -1020 1854 -1014
rect 1848 -1026 1854 -1020
rect 1848 -1032 1854 -1026
rect 1848 -1038 1854 -1032
rect 1848 -1044 1854 -1038
rect 1848 -1050 1854 -1044
rect 1848 -1056 1854 -1050
rect 1848 -1062 1854 -1056
rect 1848 -1068 1854 -1062
rect 1848 -1074 1854 -1068
rect 1848 -1080 1854 -1074
rect 1848 -1086 1854 -1080
rect 1848 -1092 1854 -1086
rect 1848 -1098 1854 -1092
rect 1848 -1104 1854 -1098
rect 1848 -1110 1854 -1104
rect 1848 -1116 1854 -1110
rect 1848 -1122 1854 -1116
rect 1848 -1128 1854 -1122
rect 1848 -1134 1854 -1128
rect 1848 -1140 1854 -1134
rect 1848 -1146 1854 -1140
rect 1848 -1152 1854 -1146
rect 1848 -1158 1854 -1152
rect 1848 -1164 1854 -1158
rect 1848 -1170 1854 -1164
rect 1848 -1176 1854 -1170
rect 1848 -1182 1854 -1176
rect 1848 -1188 1854 -1182
rect 1848 -1194 1854 -1188
rect 1848 -1200 1854 -1194
rect 1848 -1206 1854 -1200
rect 1848 -1212 1854 -1206
rect 1848 -1218 1854 -1212
rect 1848 -1224 1854 -1218
rect 1848 -1230 1854 -1224
rect 1848 -1236 1854 -1230
rect 1848 -1242 1854 -1236
rect 1848 -1248 1854 -1242
rect 1848 -1254 1854 -1248
rect 1848 -1260 1854 -1254
rect 1848 -1266 1854 -1260
rect 1848 -1272 1854 -1266
rect 1848 -1278 1854 -1272
rect 1848 -1284 1854 -1278
rect 1848 -1290 1854 -1284
rect 1848 -1296 1854 -1290
rect 1848 -1302 1854 -1296
rect 1848 -1308 1854 -1302
rect 1848 -1314 1854 -1308
rect 1848 -1320 1854 -1314
rect 1848 -1326 1854 -1320
rect 1848 -1332 1854 -1326
rect 1848 -1338 1854 -1332
rect 1848 -1344 1854 -1338
rect 1848 -1350 1854 -1344
rect 1848 -1356 1854 -1350
rect 1848 -1362 1854 -1356
rect 1848 -1368 1854 -1362
rect 1848 -1374 1854 -1368
rect 1848 -1380 1854 -1374
rect 1848 -1386 1854 -1380
rect 1848 -1392 1854 -1386
rect 1848 -1398 1854 -1392
rect 1848 -1404 1854 -1398
rect 1848 -1410 1854 -1404
rect 1848 -1416 1854 -1410
rect 1848 -1422 1854 -1416
rect 1848 -1428 1854 -1422
rect 1848 -1434 1854 -1428
rect 1848 -1440 1854 -1434
rect 1848 -1446 1854 -1440
rect 1848 -1452 1854 -1446
rect 1848 -1458 1854 -1452
rect 1848 -1464 1854 -1458
rect 1848 -1470 1854 -1464
rect 1848 -1476 1854 -1470
rect 1848 -1482 1854 -1476
rect 1848 -1488 1854 -1482
rect 1848 -1494 1854 -1488
rect 1848 -1500 1854 -1494
rect 1848 -1506 1854 -1500
rect 1848 -1512 1854 -1506
rect 1848 -1518 1854 -1512
rect 1848 -1524 1854 -1518
rect 1848 -1530 1854 -1524
rect 1848 -1536 1854 -1530
rect 1848 -1542 1854 -1536
rect 1848 -1548 1854 -1542
rect 1848 -1554 1854 -1548
rect 1848 -1560 1854 -1554
rect 1848 -1566 1854 -1560
rect 1848 -1572 1854 -1566
rect 1848 -1578 1854 -1572
rect 1848 -1584 1854 -1578
rect 1848 -1590 1854 -1584
rect 1848 -1596 1854 -1590
rect 1848 -1602 1854 -1596
rect 1848 -1608 1854 -1602
rect 1848 -1614 1854 -1608
rect 1848 -1620 1854 -1614
rect 1848 -1626 1854 -1620
rect 1848 -1632 1854 -1626
rect 1848 -1638 1854 -1632
rect 1848 -1644 1854 -1638
rect 1848 -1650 1854 -1644
rect 1848 -1656 1854 -1650
rect 1848 -1662 1854 -1656
rect 1848 -1668 1854 -1662
rect 1848 -1674 1854 -1668
rect 1848 -1680 1854 -1674
rect 1848 -1686 1854 -1680
rect 1848 -1692 1854 -1686
rect 1848 -1698 1854 -1692
rect 1848 -1704 1854 -1698
rect 1848 -1710 1854 -1704
rect 1848 -1716 1854 -1710
rect 1848 -1722 1854 -1716
rect 1848 -1728 1854 -1722
rect 1848 -1734 1854 -1728
rect 1848 -1740 1854 -1734
rect 1848 -1746 1854 -1740
rect 1848 -1752 1854 -1746
rect 1848 -1758 1854 -1752
rect 1848 -1764 1854 -1758
rect 1848 -1770 1854 -1764
rect 1848 -1776 1854 -1770
rect 1848 -1782 1854 -1776
rect 1848 -1788 1854 -1782
rect 1848 -1794 1854 -1788
rect 1848 -1800 1854 -1794
rect 1848 -1878 1854 -1872
rect 1848 -1884 1854 -1878
rect 1848 -1890 1854 -1884
rect 1848 -1896 1854 -1890
rect 1848 -1902 1854 -1896
rect 1848 -1908 1854 -1902
rect 1848 -1914 1854 -1908
rect 1848 -1920 1854 -1914
rect 1848 -1926 1854 -1920
rect 1848 -1932 1854 -1926
rect 1848 -1938 1854 -1932
rect 1848 -1944 1854 -1938
rect 1848 -1950 1854 -1944
rect 1848 -1956 1854 -1950
rect 1848 -1962 1854 -1956
rect 1848 -1968 1854 -1962
rect 1848 -1974 1854 -1968
rect 1848 -1980 1854 -1974
rect 1848 -1986 1854 -1980
rect 1848 -1992 1854 -1986
rect 1848 -1998 1854 -1992
rect 1848 -2004 1854 -1998
rect 1848 -2010 1854 -2004
rect 1848 -2016 1854 -2010
rect 1848 -2022 1854 -2016
rect 1848 -2028 1854 -2022
rect 1848 -2034 1854 -2028
rect 1848 -2040 1854 -2034
rect 1848 -2046 1854 -2040
rect 1848 -2052 1854 -2046
rect 1848 -2058 1854 -2052
rect 1848 -2064 1854 -2058
rect 1848 -2070 1854 -2064
rect 1848 -2076 1854 -2070
rect 1848 -2082 1854 -2076
rect 1848 -2088 1854 -2082
rect 1848 -2094 1854 -2088
rect 1848 -2100 1854 -2094
rect 1848 -2106 1854 -2100
rect 1848 -2112 1854 -2106
rect 1848 -2118 1854 -2112
rect 1848 -2124 1854 -2118
rect 1848 -2130 1854 -2124
rect 1848 -2136 1854 -2130
rect 1848 -2142 1854 -2136
rect 1848 -2148 1854 -2142
rect 1848 -2154 1854 -2148
rect 1848 -2160 1854 -2154
rect 1848 -2166 1854 -2160
rect 1848 -2172 1854 -2166
rect 1848 -2178 1854 -2172
rect 1848 -2184 1854 -2178
rect 1848 -2190 1854 -2184
rect 1848 -2196 1854 -2190
rect 1848 -2202 1854 -2196
rect 1848 -2208 1854 -2202
rect 1848 -2214 1854 -2208
rect 1848 -2220 1854 -2214
rect 1848 -2226 1854 -2220
rect 1848 -2232 1854 -2226
rect 1848 -2238 1854 -2232
rect 1848 -2244 1854 -2238
rect 1848 -2250 1854 -2244
rect 1848 -2256 1854 -2250
rect 1848 -2262 1854 -2256
rect 1848 -2268 1854 -2262
rect 1848 -2274 1854 -2268
rect 1848 -2280 1854 -2274
rect 1848 -2286 1854 -2280
rect 1848 -2292 1854 -2286
rect 1848 -2298 1854 -2292
rect 1848 -2304 1854 -2298
rect 1848 -2310 1854 -2304
rect 1848 -2316 1854 -2310
rect 1848 -2322 1854 -2316
rect 1848 -2328 1854 -2322
rect 1848 -2334 1854 -2328
rect 1848 -2340 1854 -2334
rect 1848 -2346 1854 -2340
rect 1848 -2352 1854 -2346
rect 1848 -2358 1854 -2352
rect 1848 -2364 1854 -2358
rect 1848 -2370 1854 -2364
rect 1848 -2376 1854 -2370
rect 1848 -2382 1854 -2376
rect 1848 -2388 1854 -2382
rect 1848 -2394 1854 -2388
rect 1848 -2400 1854 -2394
rect 1848 -2406 1854 -2400
rect 1848 -2412 1854 -2406
rect 1848 -2418 1854 -2412
rect 1848 -2424 1854 -2418
rect 1848 -2430 1854 -2424
rect 1848 -2436 1854 -2430
rect 1848 -2442 1854 -2436
rect 1848 -2448 1854 -2442
rect 1848 -2454 1854 -2448
rect 1848 -2460 1854 -2454
rect 1848 -2466 1854 -2460
rect 1848 -2472 1854 -2466
rect 1848 -2478 1854 -2472
rect 1848 -2484 1854 -2478
rect 1848 -2490 1854 -2484
rect 1848 -2496 1854 -2490
rect 1848 -2502 1854 -2496
rect 1848 -2508 1854 -2502
rect 1848 -2514 1854 -2508
rect 1848 -2520 1854 -2514
rect 1848 -2526 1854 -2520
rect 1848 -2532 1854 -2526
rect 1848 -2538 1854 -2532
rect 1848 -2544 1854 -2538
rect 1848 -2550 1854 -2544
rect 1848 -2556 1854 -2550
rect 1848 -2562 1854 -2556
rect 1848 -2568 1854 -2562
rect 1848 -2574 1854 -2568
rect 1848 -2580 1854 -2574
rect 1848 -2586 1854 -2580
rect 1848 -2592 1854 -2586
rect 1848 -2598 1854 -2592
rect 1848 -2604 1854 -2598
rect 1848 -2682 1854 -2676
rect 1848 -2688 1854 -2682
rect 1848 -2694 1854 -2688
rect 1848 -2700 1854 -2694
rect 1848 -2706 1854 -2700
rect 1848 -2712 1854 -2706
rect 1848 -2718 1854 -2712
rect 1848 -2724 1854 -2718
rect 1848 -2730 1854 -2724
rect 1848 -2736 1854 -2730
rect 1848 -2742 1854 -2736
rect 1848 -2748 1854 -2742
rect 1848 -2754 1854 -2748
rect 1848 -2760 1854 -2754
rect 1848 -2766 1854 -2760
rect 1848 -2772 1854 -2766
rect 1848 -2778 1854 -2772
rect 1848 -2784 1854 -2778
rect 1848 -2790 1854 -2784
rect 1848 -2796 1854 -2790
rect 1848 -2802 1854 -2796
rect 1848 -2808 1854 -2802
rect 1848 -2814 1854 -2808
rect 1848 -2820 1854 -2814
rect 1848 -2826 1854 -2820
rect 1848 -2832 1854 -2826
rect 1848 -2838 1854 -2832
rect 1848 -2844 1854 -2838
rect 1848 -2850 1854 -2844
rect 1848 -2856 1854 -2850
rect 1848 -2862 1854 -2856
rect 1848 -2868 1854 -2862
rect 1848 -2874 1854 -2868
rect 1848 -2880 1854 -2874
rect 1848 -2886 1854 -2880
rect 1848 -2892 1854 -2886
rect 1848 -2898 1854 -2892
rect 1848 -2904 1854 -2898
rect 1848 -2910 1854 -2904
rect 1848 -2916 1854 -2910
rect 1848 -2922 1854 -2916
rect 1848 -2928 1854 -2922
rect 1848 -2934 1854 -2928
rect 1848 -2940 1854 -2934
rect 1848 -2946 1854 -2940
rect 1848 -2952 1854 -2946
rect 1848 -2958 1854 -2952
rect 1848 -2964 1854 -2958
rect 1848 -2970 1854 -2964
rect 1848 -2976 1854 -2970
rect 1848 -2982 1854 -2976
rect 1848 -2988 1854 -2982
rect 1848 -2994 1854 -2988
rect 1848 -3000 1854 -2994
rect 1848 -3006 1854 -3000
rect 1848 -3012 1854 -3006
rect 1848 -3018 1854 -3012
rect 1848 -3024 1854 -3018
rect 1848 -3030 1854 -3024
rect 1848 -3036 1854 -3030
rect 1848 -3042 1854 -3036
rect 1848 -3048 1854 -3042
rect 1848 -3054 1854 -3048
rect 1848 -3060 1854 -3054
rect 1848 -3066 1854 -3060
rect 1848 -3072 1854 -3066
rect 1848 -3078 1854 -3072
rect 1848 -3084 1854 -3078
rect 1848 -3090 1854 -3084
rect 1848 -3096 1854 -3090
rect 1848 -3102 1854 -3096
rect 1848 -3108 1854 -3102
rect 1848 -3114 1854 -3108
rect 1848 -3120 1854 -3114
rect 1848 -3126 1854 -3120
rect 1848 -3132 1854 -3126
rect 1848 -3138 1854 -3132
rect 1848 -3144 1854 -3138
rect 1848 -3150 1854 -3144
rect 1848 -3156 1854 -3150
rect 1848 -3162 1854 -3156
rect 1848 -3216 1854 -3210
rect 1848 -3222 1854 -3216
rect 1848 -3228 1854 -3222
rect 1848 -3234 1854 -3228
rect 1848 -3240 1854 -3234
rect 1848 -3246 1854 -3240
rect 1848 -3252 1854 -3246
rect 1848 -3258 1854 -3252
rect 1848 -3264 1854 -3258
rect 1848 -3270 1854 -3264
rect 1848 -3276 1854 -3270
rect 1848 -3282 1854 -3276
rect 1848 -3288 1854 -3282
rect 1848 -3294 1854 -3288
rect 1848 -3300 1854 -3294
rect 1848 -3306 1854 -3300
rect 1848 -3312 1854 -3306
rect 1848 -3318 1854 -3312
rect 1848 -3324 1854 -3318
rect 1848 -3330 1854 -3324
rect 1848 -3336 1854 -3330
rect 1854 -648 1860 -642
rect 1854 -654 1860 -648
rect 1854 -660 1860 -654
rect 1854 -666 1860 -660
rect 1854 -672 1860 -666
rect 1854 -678 1860 -672
rect 1854 -684 1860 -678
rect 1854 -690 1860 -684
rect 1854 -696 1860 -690
rect 1854 -702 1860 -696
rect 1854 -708 1860 -702
rect 1854 -714 1860 -708
rect 1854 -720 1860 -714
rect 1854 -726 1860 -720
rect 1854 -732 1860 -726
rect 1854 -738 1860 -732
rect 1854 -744 1860 -738
rect 1854 -750 1860 -744
rect 1854 -756 1860 -750
rect 1854 -762 1860 -756
rect 1854 -768 1860 -762
rect 1854 -774 1860 -768
rect 1854 -780 1860 -774
rect 1854 -786 1860 -780
rect 1854 -792 1860 -786
rect 1854 -798 1860 -792
rect 1854 -804 1860 -798
rect 1854 -810 1860 -804
rect 1854 -816 1860 -810
rect 1854 -822 1860 -816
rect 1854 -828 1860 -822
rect 1854 -834 1860 -828
rect 1854 -840 1860 -834
rect 1854 -846 1860 -840
rect 1854 -852 1860 -846
rect 1854 -858 1860 -852
rect 1854 -864 1860 -858
rect 1854 -870 1860 -864
rect 1854 -876 1860 -870
rect 1854 -882 1860 -876
rect 1854 -888 1860 -882
rect 1854 -894 1860 -888
rect 1854 -900 1860 -894
rect 1854 -906 1860 -900
rect 1854 -912 1860 -906
rect 1854 -918 1860 -912
rect 1854 -924 1860 -918
rect 1854 -930 1860 -924
rect 1854 -936 1860 -930
rect 1854 -942 1860 -936
rect 1854 -948 1860 -942
rect 1854 -954 1860 -948
rect 1854 -960 1860 -954
rect 1854 -966 1860 -960
rect 1854 -972 1860 -966
rect 1854 -978 1860 -972
rect 1854 -984 1860 -978
rect 1854 -990 1860 -984
rect 1854 -996 1860 -990
rect 1854 -1002 1860 -996
rect 1854 -1008 1860 -1002
rect 1854 -1014 1860 -1008
rect 1854 -1020 1860 -1014
rect 1854 -1026 1860 -1020
rect 1854 -1032 1860 -1026
rect 1854 -1038 1860 -1032
rect 1854 -1044 1860 -1038
rect 1854 -1050 1860 -1044
rect 1854 -1056 1860 -1050
rect 1854 -1062 1860 -1056
rect 1854 -1068 1860 -1062
rect 1854 -1074 1860 -1068
rect 1854 -1080 1860 -1074
rect 1854 -1086 1860 -1080
rect 1854 -1092 1860 -1086
rect 1854 -1098 1860 -1092
rect 1854 -1104 1860 -1098
rect 1854 -1110 1860 -1104
rect 1854 -1116 1860 -1110
rect 1854 -1122 1860 -1116
rect 1854 -1128 1860 -1122
rect 1854 -1134 1860 -1128
rect 1854 -1140 1860 -1134
rect 1854 -1146 1860 -1140
rect 1854 -1152 1860 -1146
rect 1854 -1158 1860 -1152
rect 1854 -1164 1860 -1158
rect 1854 -1170 1860 -1164
rect 1854 -1176 1860 -1170
rect 1854 -1182 1860 -1176
rect 1854 -1188 1860 -1182
rect 1854 -1194 1860 -1188
rect 1854 -1200 1860 -1194
rect 1854 -1206 1860 -1200
rect 1854 -1212 1860 -1206
rect 1854 -1218 1860 -1212
rect 1854 -1224 1860 -1218
rect 1854 -1230 1860 -1224
rect 1854 -1236 1860 -1230
rect 1854 -1242 1860 -1236
rect 1854 -1248 1860 -1242
rect 1854 -1254 1860 -1248
rect 1854 -1260 1860 -1254
rect 1854 -1266 1860 -1260
rect 1854 -1272 1860 -1266
rect 1854 -1278 1860 -1272
rect 1854 -1284 1860 -1278
rect 1854 -1290 1860 -1284
rect 1854 -1296 1860 -1290
rect 1854 -1302 1860 -1296
rect 1854 -1308 1860 -1302
rect 1854 -1314 1860 -1308
rect 1854 -1320 1860 -1314
rect 1854 -1326 1860 -1320
rect 1854 -1332 1860 -1326
rect 1854 -1338 1860 -1332
rect 1854 -1344 1860 -1338
rect 1854 -1350 1860 -1344
rect 1854 -1356 1860 -1350
rect 1854 -1362 1860 -1356
rect 1854 -1368 1860 -1362
rect 1854 -1374 1860 -1368
rect 1854 -1380 1860 -1374
rect 1854 -1386 1860 -1380
rect 1854 -1392 1860 -1386
rect 1854 -1398 1860 -1392
rect 1854 -1404 1860 -1398
rect 1854 -1410 1860 -1404
rect 1854 -1416 1860 -1410
rect 1854 -1422 1860 -1416
rect 1854 -1428 1860 -1422
rect 1854 -1434 1860 -1428
rect 1854 -1440 1860 -1434
rect 1854 -1446 1860 -1440
rect 1854 -1452 1860 -1446
rect 1854 -1458 1860 -1452
rect 1854 -1464 1860 -1458
rect 1854 -1470 1860 -1464
rect 1854 -1476 1860 -1470
rect 1854 -1482 1860 -1476
rect 1854 -1488 1860 -1482
rect 1854 -1494 1860 -1488
rect 1854 -1500 1860 -1494
rect 1854 -1506 1860 -1500
rect 1854 -1512 1860 -1506
rect 1854 -1518 1860 -1512
rect 1854 -1524 1860 -1518
rect 1854 -1530 1860 -1524
rect 1854 -1536 1860 -1530
rect 1854 -1542 1860 -1536
rect 1854 -1548 1860 -1542
rect 1854 -1554 1860 -1548
rect 1854 -1560 1860 -1554
rect 1854 -1566 1860 -1560
rect 1854 -1572 1860 -1566
rect 1854 -1578 1860 -1572
rect 1854 -1584 1860 -1578
rect 1854 -1590 1860 -1584
rect 1854 -1596 1860 -1590
rect 1854 -1602 1860 -1596
rect 1854 -1608 1860 -1602
rect 1854 -1614 1860 -1608
rect 1854 -1620 1860 -1614
rect 1854 -1626 1860 -1620
rect 1854 -1632 1860 -1626
rect 1854 -1638 1860 -1632
rect 1854 -1644 1860 -1638
rect 1854 -1650 1860 -1644
rect 1854 -1656 1860 -1650
rect 1854 -1662 1860 -1656
rect 1854 -1668 1860 -1662
rect 1854 -1674 1860 -1668
rect 1854 -1680 1860 -1674
rect 1854 -1686 1860 -1680
rect 1854 -1692 1860 -1686
rect 1854 -1698 1860 -1692
rect 1854 -1704 1860 -1698
rect 1854 -1710 1860 -1704
rect 1854 -1716 1860 -1710
rect 1854 -1722 1860 -1716
rect 1854 -1728 1860 -1722
rect 1854 -1734 1860 -1728
rect 1854 -1740 1860 -1734
rect 1854 -1746 1860 -1740
rect 1854 -1752 1860 -1746
rect 1854 -1758 1860 -1752
rect 1854 -1764 1860 -1758
rect 1854 -1770 1860 -1764
rect 1854 -1776 1860 -1770
rect 1854 -1782 1860 -1776
rect 1854 -1788 1860 -1782
rect 1854 -1794 1860 -1788
rect 1854 -1872 1860 -1866
rect 1854 -1878 1860 -1872
rect 1854 -1884 1860 -1878
rect 1854 -1890 1860 -1884
rect 1854 -1896 1860 -1890
rect 1854 -1902 1860 -1896
rect 1854 -1908 1860 -1902
rect 1854 -1914 1860 -1908
rect 1854 -1920 1860 -1914
rect 1854 -1926 1860 -1920
rect 1854 -1932 1860 -1926
rect 1854 -1938 1860 -1932
rect 1854 -1944 1860 -1938
rect 1854 -1950 1860 -1944
rect 1854 -1956 1860 -1950
rect 1854 -1962 1860 -1956
rect 1854 -1968 1860 -1962
rect 1854 -1974 1860 -1968
rect 1854 -1980 1860 -1974
rect 1854 -1986 1860 -1980
rect 1854 -1992 1860 -1986
rect 1854 -1998 1860 -1992
rect 1854 -2004 1860 -1998
rect 1854 -2010 1860 -2004
rect 1854 -2016 1860 -2010
rect 1854 -2022 1860 -2016
rect 1854 -2028 1860 -2022
rect 1854 -2034 1860 -2028
rect 1854 -2040 1860 -2034
rect 1854 -2046 1860 -2040
rect 1854 -2052 1860 -2046
rect 1854 -2058 1860 -2052
rect 1854 -2064 1860 -2058
rect 1854 -2070 1860 -2064
rect 1854 -2076 1860 -2070
rect 1854 -2082 1860 -2076
rect 1854 -2088 1860 -2082
rect 1854 -2094 1860 -2088
rect 1854 -2100 1860 -2094
rect 1854 -2106 1860 -2100
rect 1854 -2112 1860 -2106
rect 1854 -2118 1860 -2112
rect 1854 -2124 1860 -2118
rect 1854 -2130 1860 -2124
rect 1854 -2136 1860 -2130
rect 1854 -2142 1860 -2136
rect 1854 -2148 1860 -2142
rect 1854 -2154 1860 -2148
rect 1854 -2160 1860 -2154
rect 1854 -2166 1860 -2160
rect 1854 -2172 1860 -2166
rect 1854 -2178 1860 -2172
rect 1854 -2184 1860 -2178
rect 1854 -2190 1860 -2184
rect 1854 -2196 1860 -2190
rect 1854 -2202 1860 -2196
rect 1854 -2208 1860 -2202
rect 1854 -2214 1860 -2208
rect 1854 -2220 1860 -2214
rect 1854 -2226 1860 -2220
rect 1854 -2232 1860 -2226
rect 1854 -2238 1860 -2232
rect 1854 -2244 1860 -2238
rect 1854 -2250 1860 -2244
rect 1854 -2256 1860 -2250
rect 1854 -2262 1860 -2256
rect 1854 -2268 1860 -2262
rect 1854 -2274 1860 -2268
rect 1854 -2280 1860 -2274
rect 1854 -2286 1860 -2280
rect 1854 -2292 1860 -2286
rect 1854 -2298 1860 -2292
rect 1854 -2304 1860 -2298
rect 1854 -2310 1860 -2304
rect 1854 -2316 1860 -2310
rect 1854 -2322 1860 -2316
rect 1854 -2328 1860 -2322
rect 1854 -2334 1860 -2328
rect 1854 -2340 1860 -2334
rect 1854 -2346 1860 -2340
rect 1854 -2352 1860 -2346
rect 1854 -2358 1860 -2352
rect 1854 -2364 1860 -2358
rect 1854 -2370 1860 -2364
rect 1854 -2376 1860 -2370
rect 1854 -2382 1860 -2376
rect 1854 -2388 1860 -2382
rect 1854 -2394 1860 -2388
rect 1854 -2400 1860 -2394
rect 1854 -2406 1860 -2400
rect 1854 -2412 1860 -2406
rect 1854 -2418 1860 -2412
rect 1854 -2424 1860 -2418
rect 1854 -2430 1860 -2424
rect 1854 -2436 1860 -2430
rect 1854 -2442 1860 -2436
rect 1854 -2448 1860 -2442
rect 1854 -2454 1860 -2448
rect 1854 -2460 1860 -2454
rect 1854 -2466 1860 -2460
rect 1854 -2472 1860 -2466
rect 1854 -2478 1860 -2472
rect 1854 -2484 1860 -2478
rect 1854 -2490 1860 -2484
rect 1854 -2496 1860 -2490
rect 1854 -2502 1860 -2496
rect 1854 -2508 1860 -2502
rect 1854 -2514 1860 -2508
rect 1854 -2520 1860 -2514
rect 1854 -2526 1860 -2520
rect 1854 -2532 1860 -2526
rect 1854 -2538 1860 -2532
rect 1854 -2544 1860 -2538
rect 1854 -2550 1860 -2544
rect 1854 -2556 1860 -2550
rect 1854 -2562 1860 -2556
rect 1854 -2568 1860 -2562
rect 1854 -2574 1860 -2568
rect 1854 -2580 1860 -2574
rect 1854 -2586 1860 -2580
rect 1854 -2592 1860 -2586
rect 1854 -2598 1860 -2592
rect 1854 -2604 1860 -2598
rect 1854 -2676 1860 -2670
rect 1854 -2682 1860 -2676
rect 1854 -2688 1860 -2682
rect 1854 -2694 1860 -2688
rect 1854 -2700 1860 -2694
rect 1854 -2706 1860 -2700
rect 1854 -2712 1860 -2706
rect 1854 -2718 1860 -2712
rect 1854 -2724 1860 -2718
rect 1854 -2730 1860 -2724
rect 1854 -2736 1860 -2730
rect 1854 -2742 1860 -2736
rect 1854 -2748 1860 -2742
rect 1854 -2754 1860 -2748
rect 1854 -2760 1860 -2754
rect 1854 -2766 1860 -2760
rect 1854 -2772 1860 -2766
rect 1854 -2778 1860 -2772
rect 1854 -2784 1860 -2778
rect 1854 -2790 1860 -2784
rect 1854 -2796 1860 -2790
rect 1854 -2802 1860 -2796
rect 1854 -2808 1860 -2802
rect 1854 -2814 1860 -2808
rect 1854 -2820 1860 -2814
rect 1854 -2826 1860 -2820
rect 1854 -2832 1860 -2826
rect 1854 -2838 1860 -2832
rect 1854 -2844 1860 -2838
rect 1854 -2850 1860 -2844
rect 1854 -2856 1860 -2850
rect 1854 -2862 1860 -2856
rect 1854 -2868 1860 -2862
rect 1854 -2874 1860 -2868
rect 1854 -2880 1860 -2874
rect 1854 -2886 1860 -2880
rect 1854 -2892 1860 -2886
rect 1854 -2898 1860 -2892
rect 1854 -2904 1860 -2898
rect 1854 -2910 1860 -2904
rect 1854 -2916 1860 -2910
rect 1854 -2922 1860 -2916
rect 1854 -2928 1860 -2922
rect 1854 -2934 1860 -2928
rect 1854 -2940 1860 -2934
rect 1854 -2946 1860 -2940
rect 1854 -2952 1860 -2946
rect 1854 -2958 1860 -2952
rect 1854 -2964 1860 -2958
rect 1854 -2970 1860 -2964
rect 1854 -2976 1860 -2970
rect 1854 -2982 1860 -2976
rect 1854 -2988 1860 -2982
rect 1854 -2994 1860 -2988
rect 1854 -3000 1860 -2994
rect 1854 -3006 1860 -3000
rect 1854 -3012 1860 -3006
rect 1854 -3018 1860 -3012
rect 1854 -3024 1860 -3018
rect 1854 -3030 1860 -3024
rect 1854 -3036 1860 -3030
rect 1854 -3042 1860 -3036
rect 1854 -3048 1860 -3042
rect 1854 -3054 1860 -3048
rect 1854 -3060 1860 -3054
rect 1854 -3066 1860 -3060
rect 1854 -3072 1860 -3066
rect 1854 -3078 1860 -3072
rect 1854 -3084 1860 -3078
rect 1854 -3090 1860 -3084
rect 1854 -3096 1860 -3090
rect 1854 -3102 1860 -3096
rect 1854 -3108 1860 -3102
rect 1854 -3114 1860 -3108
rect 1854 -3120 1860 -3114
rect 1854 -3126 1860 -3120
rect 1854 -3132 1860 -3126
rect 1854 -3138 1860 -3132
rect 1854 -3144 1860 -3138
rect 1854 -3150 1860 -3144
rect 1854 -3156 1860 -3150
rect 1854 -3162 1860 -3156
rect 1854 -3216 1860 -3210
rect 1854 -3222 1860 -3216
rect 1854 -3228 1860 -3222
rect 1854 -3234 1860 -3228
rect 1854 -3240 1860 -3234
rect 1854 -3246 1860 -3240
rect 1854 -3252 1860 -3246
rect 1854 -3258 1860 -3252
rect 1854 -3264 1860 -3258
rect 1854 -3270 1860 -3264
rect 1854 -3276 1860 -3270
rect 1854 -3282 1860 -3276
rect 1854 -3288 1860 -3282
rect 1854 -3294 1860 -3288
rect 1854 -3300 1860 -3294
rect 1854 -3306 1860 -3300
rect 1854 -3312 1860 -3306
rect 1854 -3318 1860 -3312
rect 1854 -3324 1860 -3318
rect 1854 -3330 1860 -3324
rect 1854 -3336 1860 -3330
rect 1860 -636 1866 -630
rect 1860 -642 1866 -636
rect 1860 -648 1866 -642
rect 1860 -654 1866 -648
rect 1860 -660 1866 -654
rect 1860 -666 1866 -660
rect 1860 -672 1866 -666
rect 1860 -678 1866 -672
rect 1860 -684 1866 -678
rect 1860 -690 1866 -684
rect 1860 -696 1866 -690
rect 1860 -702 1866 -696
rect 1860 -708 1866 -702
rect 1860 -714 1866 -708
rect 1860 -720 1866 -714
rect 1860 -726 1866 -720
rect 1860 -732 1866 -726
rect 1860 -738 1866 -732
rect 1860 -744 1866 -738
rect 1860 -750 1866 -744
rect 1860 -756 1866 -750
rect 1860 -762 1866 -756
rect 1860 -768 1866 -762
rect 1860 -774 1866 -768
rect 1860 -780 1866 -774
rect 1860 -786 1866 -780
rect 1860 -792 1866 -786
rect 1860 -798 1866 -792
rect 1860 -804 1866 -798
rect 1860 -810 1866 -804
rect 1860 -816 1866 -810
rect 1860 -822 1866 -816
rect 1860 -828 1866 -822
rect 1860 -834 1866 -828
rect 1860 -840 1866 -834
rect 1860 -846 1866 -840
rect 1860 -852 1866 -846
rect 1860 -858 1866 -852
rect 1860 -864 1866 -858
rect 1860 -870 1866 -864
rect 1860 -876 1866 -870
rect 1860 -882 1866 -876
rect 1860 -888 1866 -882
rect 1860 -894 1866 -888
rect 1860 -900 1866 -894
rect 1860 -906 1866 -900
rect 1860 -912 1866 -906
rect 1860 -918 1866 -912
rect 1860 -924 1866 -918
rect 1860 -930 1866 -924
rect 1860 -936 1866 -930
rect 1860 -942 1866 -936
rect 1860 -948 1866 -942
rect 1860 -954 1866 -948
rect 1860 -960 1866 -954
rect 1860 -966 1866 -960
rect 1860 -972 1866 -966
rect 1860 -978 1866 -972
rect 1860 -984 1866 -978
rect 1860 -990 1866 -984
rect 1860 -996 1866 -990
rect 1860 -1002 1866 -996
rect 1860 -1008 1866 -1002
rect 1860 -1014 1866 -1008
rect 1860 -1020 1866 -1014
rect 1860 -1026 1866 -1020
rect 1860 -1032 1866 -1026
rect 1860 -1038 1866 -1032
rect 1860 -1044 1866 -1038
rect 1860 -1050 1866 -1044
rect 1860 -1056 1866 -1050
rect 1860 -1062 1866 -1056
rect 1860 -1068 1866 -1062
rect 1860 -1074 1866 -1068
rect 1860 -1080 1866 -1074
rect 1860 -1086 1866 -1080
rect 1860 -1092 1866 -1086
rect 1860 -1098 1866 -1092
rect 1860 -1104 1866 -1098
rect 1860 -1110 1866 -1104
rect 1860 -1116 1866 -1110
rect 1860 -1122 1866 -1116
rect 1860 -1128 1866 -1122
rect 1860 -1134 1866 -1128
rect 1860 -1140 1866 -1134
rect 1860 -1146 1866 -1140
rect 1860 -1152 1866 -1146
rect 1860 -1158 1866 -1152
rect 1860 -1164 1866 -1158
rect 1860 -1170 1866 -1164
rect 1860 -1176 1866 -1170
rect 1860 -1182 1866 -1176
rect 1860 -1188 1866 -1182
rect 1860 -1194 1866 -1188
rect 1860 -1200 1866 -1194
rect 1860 -1206 1866 -1200
rect 1860 -1212 1866 -1206
rect 1860 -1218 1866 -1212
rect 1860 -1224 1866 -1218
rect 1860 -1230 1866 -1224
rect 1860 -1236 1866 -1230
rect 1860 -1242 1866 -1236
rect 1860 -1248 1866 -1242
rect 1860 -1254 1866 -1248
rect 1860 -1260 1866 -1254
rect 1860 -1266 1866 -1260
rect 1860 -1272 1866 -1266
rect 1860 -1278 1866 -1272
rect 1860 -1284 1866 -1278
rect 1860 -1290 1866 -1284
rect 1860 -1296 1866 -1290
rect 1860 -1302 1866 -1296
rect 1860 -1308 1866 -1302
rect 1860 -1314 1866 -1308
rect 1860 -1320 1866 -1314
rect 1860 -1326 1866 -1320
rect 1860 -1332 1866 -1326
rect 1860 -1338 1866 -1332
rect 1860 -1344 1866 -1338
rect 1860 -1350 1866 -1344
rect 1860 -1356 1866 -1350
rect 1860 -1362 1866 -1356
rect 1860 -1368 1866 -1362
rect 1860 -1374 1866 -1368
rect 1860 -1380 1866 -1374
rect 1860 -1386 1866 -1380
rect 1860 -1392 1866 -1386
rect 1860 -1398 1866 -1392
rect 1860 -1404 1866 -1398
rect 1860 -1410 1866 -1404
rect 1860 -1416 1866 -1410
rect 1860 -1422 1866 -1416
rect 1860 -1428 1866 -1422
rect 1860 -1434 1866 -1428
rect 1860 -1440 1866 -1434
rect 1860 -1446 1866 -1440
rect 1860 -1452 1866 -1446
rect 1860 -1458 1866 -1452
rect 1860 -1464 1866 -1458
rect 1860 -1470 1866 -1464
rect 1860 -1476 1866 -1470
rect 1860 -1482 1866 -1476
rect 1860 -1488 1866 -1482
rect 1860 -1494 1866 -1488
rect 1860 -1500 1866 -1494
rect 1860 -1506 1866 -1500
rect 1860 -1512 1866 -1506
rect 1860 -1518 1866 -1512
rect 1860 -1524 1866 -1518
rect 1860 -1530 1866 -1524
rect 1860 -1536 1866 -1530
rect 1860 -1542 1866 -1536
rect 1860 -1548 1866 -1542
rect 1860 -1554 1866 -1548
rect 1860 -1560 1866 -1554
rect 1860 -1566 1866 -1560
rect 1860 -1572 1866 -1566
rect 1860 -1578 1866 -1572
rect 1860 -1584 1866 -1578
rect 1860 -1590 1866 -1584
rect 1860 -1596 1866 -1590
rect 1860 -1602 1866 -1596
rect 1860 -1608 1866 -1602
rect 1860 -1614 1866 -1608
rect 1860 -1620 1866 -1614
rect 1860 -1626 1866 -1620
rect 1860 -1632 1866 -1626
rect 1860 -1638 1866 -1632
rect 1860 -1644 1866 -1638
rect 1860 -1650 1866 -1644
rect 1860 -1656 1866 -1650
rect 1860 -1662 1866 -1656
rect 1860 -1668 1866 -1662
rect 1860 -1674 1866 -1668
rect 1860 -1680 1866 -1674
rect 1860 -1686 1866 -1680
rect 1860 -1692 1866 -1686
rect 1860 -1698 1866 -1692
rect 1860 -1704 1866 -1698
rect 1860 -1710 1866 -1704
rect 1860 -1716 1866 -1710
rect 1860 -1722 1866 -1716
rect 1860 -1728 1866 -1722
rect 1860 -1734 1866 -1728
rect 1860 -1740 1866 -1734
rect 1860 -1746 1866 -1740
rect 1860 -1752 1866 -1746
rect 1860 -1758 1866 -1752
rect 1860 -1764 1866 -1758
rect 1860 -1770 1866 -1764
rect 1860 -1776 1866 -1770
rect 1860 -1782 1866 -1776
rect 1860 -1788 1866 -1782
rect 1860 -1866 1866 -1860
rect 1860 -1872 1866 -1866
rect 1860 -1878 1866 -1872
rect 1860 -1884 1866 -1878
rect 1860 -1890 1866 -1884
rect 1860 -1896 1866 -1890
rect 1860 -1902 1866 -1896
rect 1860 -1908 1866 -1902
rect 1860 -1914 1866 -1908
rect 1860 -1920 1866 -1914
rect 1860 -1926 1866 -1920
rect 1860 -1932 1866 -1926
rect 1860 -1938 1866 -1932
rect 1860 -1944 1866 -1938
rect 1860 -1950 1866 -1944
rect 1860 -1956 1866 -1950
rect 1860 -1962 1866 -1956
rect 1860 -1968 1866 -1962
rect 1860 -1974 1866 -1968
rect 1860 -1980 1866 -1974
rect 1860 -1986 1866 -1980
rect 1860 -1992 1866 -1986
rect 1860 -1998 1866 -1992
rect 1860 -2004 1866 -1998
rect 1860 -2010 1866 -2004
rect 1860 -2016 1866 -2010
rect 1860 -2022 1866 -2016
rect 1860 -2028 1866 -2022
rect 1860 -2034 1866 -2028
rect 1860 -2040 1866 -2034
rect 1860 -2046 1866 -2040
rect 1860 -2052 1866 -2046
rect 1860 -2058 1866 -2052
rect 1860 -2064 1866 -2058
rect 1860 -2070 1866 -2064
rect 1860 -2076 1866 -2070
rect 1860 -2082 1866 -2076
rect 1860 -2088 1866 -2082
rect 1860 -2094 1866 -2088
rect 1860 -2100 1866 -2094
rect 1860 -2106 1866 -2100
rect 1860 -2112 1866 -2106
rect 1860 -2118 1866 -2112
rect 1860 -2124 1866 -2118
rect 1860 -2130 1866 -2124
rect 1860 -2136 1866 -2130
rect 1860 -2142 1866 -2136
rect 1860 -2148 1866 -2142
rect 1860 -2154 1866 -2148
rect 1860 -2160 1866 -2154
rect 1860 -2166 1866 -2160
rect 1860 -2172 1866 -2166
rect 1860 -2178 1866 -2172
rect 1860 -2184 1866 -2178
rect 1860 -2190 1866 -2184
rect 1860 -2196 1866 -2190
rect 1860 -2202 1866 -2196
rect 1860 -2208 1866 -2202
rect 1860 -2214 1866 -2208
rect 1860 -2220 1866 -2214
rect 1860 -2226 1866 -2220
rect 1860 -2232 1866 -2226
rect 1860 -2238 1866 -2232
rect 1860 -2244 1866 -2238
rect 1860 -2250 1866 -2244
rect 1860 -2256 1866 -2250
rect 1860 -2262 1866 -2256
rect 1860 -2268 1866 -2262
rect 1860 -2274 1866 -2268
rect 1860 -2280 1866 -2274
rect 1860 -2286 1866 -2280
rect 1860 -2292 1866 -2286
rect 1860 -2298 1866 -2292
rect 1860 -2304 1866 -2298
rect 1860 -2310 1866 -2304
rect 1860 -2316 1866 -2310
rect 1860 -2322 1866 -2316
rect 1860 -2328 1866 -2322
rect 1860 -2334 1866 -2328
rect 1860 -2340 1866 -2334
rect 1860 -2346 1866 -2340
rect 1860 -2352 1866 -2346
rect 1860 -2358 1866 -2352
rect 1860 -2364 1866 -2358
rect 1860 -2370 1866 -2364
rect 1860 -2376 1866 -2370
rect 1860 -2382 1866 -2376
rect 1860 -2388 1866 -2382
rect 1860 -2394 1866 -2388
rect 1860 -2400 1866 -2394
rect 1860 -2406 1866 -2400
rect 1860 -2412 1866 -2406
rect 1860 -2418 1866 -2412
rect 1860 -2424 1866 -2418
rect 1860 -2430 1866 -2424
rect 1860 -2436 1866 -2430
rect 1860 -2442 1866 -2436
rect 1860 -2448 1866 -2442
rect 1860 -2454 1866 -2448
rect 1860 -2460 1866 -2454
rect 1860 -2466 1866 -2460
rect 1860 -2472 1866 -2466
rect 1860 -2478 1866 -2472
rect 1860 -2484 1866 -2478
rect 1860 -2490 1866 -2484
rect 1860 -2496 1866 -2490
rect 1860 -2502 1866 -2496
rect 1860 -2508 1866 -2502
rect 1860 -2514 1866 -2508
rect 1860 -2520 1866 -2514
rect 1860 -2526 1866 -2520
rect 1860 -2532 1866 -2526
rect 1860 -2538 1866 -2532
rect 1860 -2544 1866 -2538
rect 1860 -2550 1866 -2544
rect 1860 -2556 1866 -2550
rect 1860 -2562 1866 -2556
rect 1860 -2568 1866 -2562
rect 1860 -2574 1866 -2568
rect 1860 -2580 1866 -2574
rect 1860 -2586 1866 -2580
rect 1860 -2592 1866 -2586
rect 1860 -2598 1866 -2592
rect 1860 -2676 1866 -2670
rect 1860 -2682 1866 -2676
rect 1860 -2688 1866 -2682
rect 1860 -2694 1866 -2688
rect 1860 -2700 1866 -2694
rect 1860 -2706 1866 -2700
rect 1860 -2712 1866 -2706
rect 1860 -2718 1866 -2712
rect 1860 -2724 1866 -2718
rect 1860 -2730 1866 -2724
rect 1860 -2736 1866 -2730
rect 1860 -2742 1866 -2736
rect 1860 -2748 1866 -2742
rect 1860 -2754 1866 -2748
rect 1860 -2760 1866 -2754
rect 1860 -2766 1866 -2760
rect 1860 -2772 1866 -2766
rect 1860 -2778 1866 -2772
rect 1860 -2784 1866 -2778
rect 1860 -2790 1866 -2784
rect 1860 -2796 1866 -2790
rect 1860 -2802 1866 -2796
rect 1860 -2808 1866 -2802
rect 1860 -2814 1866 -2808
rect 1860 -2820 1866 -2814
rect 1860 -2826 1866 -2820
rect 1860 -2832 1866 -2826
rect 1860 -2838 1866 -2832
rect 1860 -2844 1866 -2838
rect 1860 -2850 1866 -2844
rect 1860 -2856 1866 -2850
rect 1860 -2862 1866 -2856
rect 1860 -2868 1866 -2862
rect 1860 -2874 1866 -2868
rect 1860 -2880 1866 -2874
rect 1860 -2886 1866 -2880
rect 1860 -2892 1866 -2886
rect 1860 -2898 1866 -2892
rect 1860 -2904 1866 -2898
rect 1860 -2910 1866 -2904
rect 1860 -2916 1866 -2910
rect 1860 -2922 1866 -2916
rect 1860 -2928 1866 -2922
rect 1860 -2934 1866 -2928
rect 1860 -2940 1866 -2934
rect 1860 -2946 1866 -2940
rect 1860 -2952 1866 -2946
rect 1860 -2958 1866 -2952
rect 1860 -2964 1866 -2958
rect 1860 -2970 1866 -2964
rect 1860 -2976 1866 -2970
rect 1860 -2982 1866 -2976
rect 1860 -2988 1866 -2982
rect 1860 -2994 1866 -2988
rect 1860 -3000 1866 -2994
rect 1860 -3006 1866 -3000
rect 1860 -3012 1866 -3006
rect 1860 -3018 1866 -3012
rect 1860 -3024 1866 -3018
rect 1860 -3030 1866 -3024
rect 1860 -3036 1866 -3030
rect 1860 -3042 1866 -3036
rect 1860 -3048 1866 -3042
rect 1860 -3054 1866 -3048
rect 1860 -3060 1866 -3054
rect 1860 -3066 1866 -3060
rect 1860 -3072 1866 -3066
rect 1860 -3078 1866 -3072
rect 1860 -3084 1866 -3078
rect 1860 -3090 1866 -3084
rect 1860 -3096 1866 -3090
rect 1860 -3102 1866 -3096
rect 1860 -3108 1866 -3102
rect 1860 -3114 1866 -3108
rect 1860 -3120 1866 -3114
rect 1860 -3126 1866 -3120
rect 1860 -3132 1866 -3126
rect 1860 -3138 1866 -3132
rect 1860 -3144 1866 -3138
rect 1860 -3150 1866 -3144
rect 1860 -3156 1866 -3150
rect 1860 -3162 1866 -3156
rect 1860 -3210 1866 -3204
rect 1860 -3216 1866 -3210
rect 1860 -3222 1866 -3216
rect 1860 -3228 1866 -3222
rect 1860 -3234 1866 -3228
rect 1860 -3240 1866 -3234
rect 1860 -3246 1866 -3240
rect 1860 -3252 1866 -3246
rect 1860 -3258 1866 -3252
rect 1860 -3264 1866 -3258
rect 1860 -3270 1866 -3264
rect 1860 -3276 1866 -3270
rect 1860 -3282 1866 -3276
rect 1860 -3288 1866 -3282
rect 1860 -3294 1866 -3288
rect 1860 -3300 1866 -3294
rect 1860 -3306 1866 -3300
rect 1860 -3312 1866 -3306
rect 1860 -3318 1866 -3312
rect 1860 -3324 1866 -3318
rect 1860 -3330 1866 -3324
rect 1866 -630 1872 -624
rect 1866 -636 1872 -630
rect 1866 -642 1872 -636
rect 1866 -648 1872 -642
rect 1866 -654 1872 -648
rect 1866 -660 1872 -654
rect 1866 -666 1872 -660
rect 1866 -672 1872 -666
rect 1866 -678 1872 -672
rect 1866 -684 1872 -678
rect 1866 -690 1872 -684
rect 1866 -696 1872 -690
rect 1866 -702 1872 -696
rect 1866 -708 1872 -702
rect 1866 -714 1872 -708
rect 1866 -720 1872 -714
rect 1866 -726 1872 -720
rect 1866 -732 1872 -726
rect 1866 -738 1872 -732
rect 1866 -744 1872 -738
rect 1866 -750 1872 -744
rect 1866 -756 1872 -750
rect 1866 -762 1872 -756
rect 1866 -768 1872 -762
rect 1866 -774 1872 -768
rect 1866 -780 1872 -774
rect 1866 -786 1872 -780
rect 1866 -792 1872 -786
rect 1866 -798 1872 -792
rect 1866 -804 1872 -798
rect 1866 -810 1872 -804
rect 1866 -816 1872 -810
rect 1866 -822 1872 -816
rect 1866 -828 1872 -822
rect 1866 -834 1872 -828
rect 1866 -840 1872 -834
rect 1866 -846 1872 -840
rect 1866 -852 1872 -846
rect 1866 -858 1872 -852
rect 1866 -864 1872 -858
rect 1866 -870 1872 -864
rect 1866 -876 1872 -870
rect 1866 -882 1872 -876
rect 1866 -888 1872 -882
rect 1866 -894 1872 -888
rect 1866 -900 1872 -894
rect 1866 -906 1872 -900
rect 1866 -912 1872 -906
rect 1866 -918 1872 -912
rect 1866 -924 1872 -918
rect 1866 -930 1872 -924
rect 1866 -936 1872 -930
rect 1866 -942 1872 -936
rect 1866 -948 1872 -942
rect 1866 -954 1872 -948
rect 1866 -960 1872 -954
rect 1866 -966 1872 -960
rect 1866 -972 1872 -966
rect 1866 -978 1872 -972
rect 1866 -984 1872 -978
rect 1866 -990 1872 -984
rect 1866 -996 1872 -990
rect 1866 -1002 1872 -996
rect 1866 -1008 1872 -1002
rect 1866 -1014 1872 -1008
rect 1866 -1020 1872 -1014
rect 1866 -1026 1872 -1020
rect 1866 -1032 1872 -1026
rect 1866 -1038 1872 -1032
rect 1866 -1044 1872 -1038
rect 1866 -1050 1872 -1044
rect 1866 -1056 1872 -1050
rect 1866 -1062 1872 -1056
rect 1866 -1068 1872 -1062
rect 1866 -1074 1872 -1068
rect 1866 -1080 1872 -1074
rect 1866 -1086 1872 -1080
rect 1866 -1092 1872 -1086
rect 1866 -1098 1872 -1092
rect 1866 -1104 1872 -1098
rect 1866 -1110 1872 -1104
rect 1866 -1116 1872 -1110
rect 1866 -1122 1872 -1116
rect 1866 -1128 1872 -1122
rect 1866 -1134 1872 -1128
rect 1866 -1140 1872 -1134
rect 1866 -1146 1872 -1140
rect 1866 -1152 1872 -1146
rect 1866 -1158 1872 -1152
rect 1866 -1164 1872 -1158
rect 1866 -1170 1872 -1164
rect 1866 -1176 1872 -1170
rect 1866 -1182 1872 -1176
rect 1866 -1188 1872 -1182
rect 1866 -1194 1872 -1188
rect 1866 -1200 1872 -1194
rect 1866 -1206 1872 -1200
rect 1866 -1212 1872 -1206
rect 1866 -1218 1872 -1212
rect 1866 -1224 1872 -1218
rect 1866 -1230 1872 -1224
rect 1866 -1236 1872 -1230
rect 1866 -1242 1872 -1236
rect 1866 -1248 1872 -1242
rect 1866 -1254 1872 -1248
rect 1866 -1260 1872 -1254
rect 1866 -1266 1872 -1260
rect 1866 -1272 1872 -1266
rect 1866 -1278 1872 -1272
rect 1866 -1284 1872 -1278
rect 1866 -1290 1872 -1284
rect 1866 -1296 1872 -1290
rect 1866 -1302 1872 -1296
rect 1866 -1308 1872 -1302
rect 1866 -1314 1872 -1308
rect 1866 -1320 1872 -1314
rect 1866 -1326 1872 -1320
rect 1866 -1332 1872 -1326
rect 1866 -1338 1872 -1332
rect 1866 -1344 1872 -1338
rect 1866 -1350 1872 -1344
rect 1866 -1356 1872 -1350
rect 1866 -1362 1872 -1356
rect 1866 -1368 1872 -1362
rect 1866 -1374 1872 -1368
rect 1866 -1380 1872 -1374
rect 1866 -1386 1872 -1380
rect 1866 -1392 1872 -1386
rect 1866 -1398 1872 -1392
rect 1866 -1404 1872 -1398
rect 1866 -1410 1872 -1404
rect 1866 -1416 1872 -1410
rect 1866 -1422 1872 -1416
rect 1866 -1428 1872 -1422
rect 1866 -1434 1872 -1428
rect 1866 -1440 1872 -1434
rect 1866 -1446 1872 -1440
rect 1866 -1452 1872 -1446
rect 1866 -1458 1872 -1452
rect 1866 -1464 1872 -1458
rect 1866 -1470 1872 -1464
rect 1866 -1476 1872 -1470
rect 1866 -1482 1872 -1476
rect 1866 -1488 1872 -1482
rect 1866 -1494 1872 -1488
rect 1866 -1500 1872 -1494
rect 1866 -1506 1872 -1500
rect 1866 -1512 1872 -1506
rect 1866 -1518 1872 -1512
rect 1866 -1524 1872 -1518
rect 1866 -1530 1872 -1524
rect 1866 -1536 1872 -1530
rect 1866 -1542 1872 -1536
rect 1866 -1548 1872 -1542
rect 1866 -1554 1872 -1548
rect 1866 -1560 1872 -1554
rect 1866 -1566 1872 -1560
rect 1866 -1572 1872 -1566
rect 1866 -1578 1872 -1572
rect 1866 -1584 1872 -1578
rect 1866 -1590 1872 -1584
rect 1866 -1596 1872 -1590
rect 1866 -1602 1872 -1596
rect 1866 -1608 1872 -1602
rect 1866 -1614 1872 -1608
rect 1866 -1620 1872 -1614
rect 1866 -1626 1872 -1620
rect 1866 -1632 1872 -1626
rect 1866 -1638 1872 -1632
rect 1866 -1644 1872 -1638
rect 1866 -1650 1872 -1644
rect 1866 -1656 1872 -1650
rect 1866 -1662 1872 -1656
rect 1866 -1668 1872 -1662
rect 1866 -1674 1872 -1668
rect 1866 -1680 1872 -1674
rect 1866 -1686 1872 -1680
rect 1866 -1692 1872 -1686
rect 1866 -1698 1872 -1692
rect 1866 -1704 1872 -1698
rect 1866 -1710 1872 -1704
rect 1866 -1716 1872 -1710
rect 1866 -1722 1872 -1716
rect 1866 -1728 1872 -1722
rect 1866 -1734 1872 -1728
rect 1866 -1740 1872 -1734
rect 1866 -1746 1872 -1740
rect 1866 -1752 1872 -1746
rect 1866 -1758 1872 -1752
rect 1866 -1764 1872 -1758
rect 1866 -1770 1872 -1764
rect 1866 -1776 1872 -1770
rect 1866 -1782 1872 -1776
rect 1866 -1860 1872 -1854
rect 1866 -1866 1872 -1860
rect 1866 -1872 1872 -1866
rect 1866 -1878 1872 -1872
rect 1866 -1884 1872 -1878
rect 1866 -1890 1872 -1884
rect 1866 -1896 1872 -1890
rect 1866 -1902 1872 -1896
rect 1866 -1908 1872 -1902
rect 1866 -1914 1872 -1908
rect 1866 -1920 1872 -1914
rect 1866 -1926 1872 -1920
rect 1866 -1932 1872 -1926
rect 1866 -1938 1872 -1932
rect 1866 -1944 1872 -1938
rect 1866 -1950 1872 -1944
rect 1866 -1956 1872 -1950
rect 1866 -1962 1872 -1956
rect 1866 -1968 1872 -1962
rect 1866 -1974 1872 -1968
rect 1866 -1980 1872 -1974
rect 1866 -1986 1872 -1980
rect 1866 -1992 1872 -1986
rect 1866 -1998 1872 -1992
rect 1866 -2004 1872 -1998
rect 1866 -2010 1872 -2004
rect 1866 -2016 1872 -2010
rect 1866 -2022 1872 -2016
rect 1866 -2028 1872 -2022
rect 1866 -2034 1872 -2028
rect 1866 -2040 1872 -2034
rect 1866 -2046 1872 -2040
rect 1866 -2052 1872 -2046
rect 1866 -2058 1872 -2052
rect 1866 -2064 1872 -2058
rect 1866 -2070 1872 -2064
rect 1866 -2076 1872 -2070
rect 1866 -2082 1872 -2076
rect 1866 -2088 1872 -2082
rect 1866 -2094 1872 -2088
rect 1866 -2100 1872 -2094
rect 1866 -2106 1872 -2100
rect 1866 -2112 1872 -2106
rect 1866 -2118 1872 -2112
rect 1866 -2124 1872 -2118
rect 1866 -2130 1872 -2124
rect 1866 -2136 1872 -2130
rect 1866 -2142 1872 -2136
rect 1866 -2148 1872 -2142
rect 1866 -2154 1872 -2148
rect 1866 -2160 1872 -2154
rect 1866 -2166 1872 -2160
rect 1866 -2172 1872 -2166
rect 1866 -2178 1872 -2172
rect 1866 -2184 1872 -2178
rect 1866 -2190 1872 -2184
rect 1866 -2196 1872 -2190
rect 1866 -2202 1872 -2196
rect 1866 -2208 1872 -2202
rect 1866 -2214 1872 -2208
rect 1866 -2220 1872 -2214
rect 1866 -2226 1872 -2220
rect 1866 -2232 1872 -2226
rect 1866 -2238 1872 -2232
rect 1866 -2244 1872 -2238
rect 1866 -2250 1872 -2244
rect 1866 -2256 1872 -2250
rect 1866 -2262 1872 -2256
rect 1866 -2268 1872 -2262
rect 1866 -2274 1872 -2268
rect 1866 -2280 1872 -2274
rect 1866 -2286 1872 -2280
rect 1866 -2292 1872 -2286
rect 1866 -2298 1872 -2292
rect 1866 -2304 1872 -2298
rect 1866 -2310 1872 -2304
rect 1866 -2316 1872 -2310
rect 1866 -2322 1872 -2316
rect 1866 -2328 1872 -2322
rect 1866 -2334 1872 -2328
rect 1866 -2340 1872 -2334
rect 1866 -2346 1872 -2340
rect 1866 -2352 1872 -2346
rect 1866 -2358 1872 -2352
rect 1866 -2364 1872 -2358
rect 1866 -2370 1872 -2364
rect 1866 -2376 1872 -2370
rect 1866 -2382 1872 -2376
rect 1866 -2388 1872 -2382
rect 1866 -2394 1872 -2388
rect 1866 -2400 1872 -2394
rect 1866 -2406 1872 -2400
rect 1866 -2412 1872 -2406
rect 1866 -2418 1872 -2412
rect 1866 -2424 1872 -2418
rect 1866 -2430 1872 -2424
rect 1866 -2436 1872 -2430
rect 1866 -2442 1872 -2436
rect 1866 -2448 1872 -2442
rect 1866 -2454 1872 -2448
rect 1866 -2460 1872 -2454
rect 1866 -2466 1872 -2460
rect 1866 -2472 1872 -2466
rect 1866 -2478 1872 -2472
rect 1866 -2484 1872 -2478
rect 1866 -2490 1872 -2484
rect 1866 -2496 1872 -2490
rect 1866 -2502 1872 -2496
rect 1866 -2508 1872 -2502
rect 1866 -2514 1872 -2508
rect 1866 -2520 1872 -2514
rect 1866 -2526 1872 -2520
rect 1866 -2532 1872 -2526
rect 1866 -2538 1872 -2532
rect 1866 -2544 1872 -2538
rect 1866 -2550 1872 -2544
rect 1866 -2556 1872 -2550
rect 1866 -2562 1872 -2556
rect 1866 -2568 1872 -2562
rect 1866 -2574 1872 -2568
rect 1866 -2580 1872 -2574
rect 1866 -2586 1872 -2580
rect 1866 -2592 1872 -2586
rect 1866 -2598 1872 -2592
rect 1866 -2670 1872 -2664
rect 1866 -2676 1872 -2670
rect 1866 -2682 1872 -2676
rect 1866 -2688 1872 -2682
rect 1866 -2694 1872 -2688
rect 1866 -2700 1872 -2694
rect 1866 -2706 1872 -2700
rect 1866 -2712 1872 -2706
rect 1866 -2718 1872 -2712
rect 1866 -2724 1872 -2718
rect 1866 -2730 1872 -2724
rect 1866 -2736 1872 -2730
rect 1866 -2742 1872 -2736
rect 1866 -2748 1872 -2742
rect 1866 -2754 1872 -2748
rect 1866 -2760 1872 -2754
rect 1866 -2766 1872 -2760
rect 1866 -2772 1872 -2766
rect 1866 -2778 1872 -2772
rect 1866 -2784 1872 -2778
rect 1866 -2790 1872 -2784
rect 1866 -2796 1872 -2790
rect 1866 -2802 1872 -2796
rect 1866 -2808 1872 -2802
rect 1866 -2814 1872 -2808
rect 1866 -2820 1872 -2814
rect 1866 -2826 1872 -2820
rect 1866 -2832 1872 -2826
rect 1866 -2838 1872 -2832
rect 1866 -2844 1872 -2838
rect 1866 -2850 1872 -2844
rect 1866 -2856 1872 -2850
rect 1866 -2862 1872 -2856
rect 1866 -2868 1872 -2862
rect 1866 -2874 1872 -2868
rect 1866 -2880 1872 -2874
rect 1866 -2886 1872 -2880
rect 1866 -2892 1872 -2886
rect 1866 -2898 1872 -2892
rect 1866 -2904 1872 -2898
rect 1866 -2910 1872 -2904
rect 1866 -2916 1872 -2910
rect 1866 -2922 1872 -2916
rect 1866 -2928 1872 -2922
rect 1866 -2934 1872 -2928
rect 1866 -2940 1872 -2934
rect 1866 -2946 1872 -2940
rect 1866 -2952 1872 -2946
rect 1866 -2958 1872 -2952
rect 1866 -2964 1872 -2958
rect 1866 -2970 1872 -2964
rect 1866 -2976 1872 -2970
rect 1866 -2982 1872 -2976
rect 1866 -2988 1872 -2982
rect 1866 -2994 1872 -2988
rect 1866 -3000 1872 -2994
rect 1866 -3006 1872 -3000
rect 1866 -3012 1872 -3006
rect 1866 -3018 1872 -3012
rect 1866 -3024 1872 -3018
rect 1866 -3030 1872 -3024
rect 1866 -3036 1872 -3030
rect 1866 -3042 1872 -3036
rect 1866 -3048 1872 -3042
rect 1866 -3054 1872 -3048
rect 1866 -3060 1872 -3054
rect 1866 -3066 1872 -3060
rect 1866 -3072 1872 -3066
rect 1866 -3078 1872 -3072
rect 1866 -3084 1872 -3078
rect 1866 -3090 1872 -3084
rect 1866 -3096 1872 -3090
rect 1866 -3102 1872 -3096
rect 1866 -3108 1872 -3102
rect 1866 -3114 1872 -3108
rect 1866 -3120 1872 -3114
rect 1866 -3126 1872 -3120
rect 1866 -3132 1872 -3126
rect 1866 -3138 1872 -3132
rect 1866 -3144 1872 -3138
rect 1866 -3150 1872 -3144
rect 1866 -3156 1872 -3150
rect 1866 -3210 1872 -3204
rect 1866 -3216 1872 -3210
rect 1866 -3222 1872 -3216
rect 1866 -3228 1872 -3222
rect 1866 -3234 1872 -3228
rect 1866 -3240 1872 -3234
rect 1866 -3246 1872 -3240
rect 1866 -3252 1872 -3246
rect 1866 -3258 1872 -3252
rect 1866 -3264 1872 -3258
rect 1866 -3270 1872 -3264
rect 1866 -3276 1872 -3270
rect 1866 -3282 1872 -3276
rect 1866 -3288 1872 -3282
rect 1866 -3294 1872 -3288
rect 1866 -3300 1872 -3294
rect 1866 -3306 1872 -3300
rect 1866 -3312 1872 -3306
rect 1866 -3318 1872 -3312
rect 1866 -3324 1872 -3318
rect 1872 -618 1878 -612
rect 1872 -624 1878 -618
rect 1872 -630 1878 -624
rect 1872 -636 1878 -630
rect 1872 -642 1878 -636
rect 1872 -648 1878 -642
rect 1872 -654 1878 -648
rect 1872 -660 1878 -654
rect 1872 -666 1878 -660
rect 1872 -672 1878 -666
rect 1872 -678 1878 -672
rect 1872 -684 1878 -678
rect 1872 -690 1878 -684
rect 1872 -696 1878 -690
rect 1872 -702 1878 -696
rect 1872 -708 1878 -702
rect 1872 -714 1878 -708
rect 1872 -720 1878 -714
rect 1872 -726 1878 -720
rect 1872 -732 1878 -726
rect 1872 -738 1878 -732
rect 1872 -744 1878 -738
rect 1872 -750 1878 -744
rect 1872 -756 1878 -750
rect 1872 -762 1878 -756
rect 1872 -768 1878 -762
rect 1872 -774 1878 -768
rect 1872 -780 1878 -774
rect 1872 -786 1878 -780
rect 1872 -792 1878 -786
rect 1872 -798 1878 -792
rect 1872 -804 1878 -798
rect 1872 -810 1878 -804
rect 1872 -816 1878 -810
rect 1872 -822 1878 -816
rect 1872 -828 1878 -822
rect 1872 -834 1878 -828
rect 1872 -840 1878 -834
rect 1872 -846 1878 -840
rect 1872 -852 1878 -846
rect 1872 -858 1878 -852
rect 1872 -864 1878 -858
rect 1872 -870 1878 -864
rect 1872 -876 1878 -870
rect 1872 -882 1878 -876
rect 1872 -888 1878 -882
rect 1872 -894 1878 -888
rect 1872 -900 1878 -894
rect 1872 -906 1878 -900
rect 1872 -912 1878 -906
rect 1872 -918 1878 -912
rect 1872 -924 1878 -918
rect 1872 -930 1878 -924
rect 1872 -936 1878 -930
rect 1872 -942 1878 -936
rect 1872 -948 1878 -942
rect 1872 -954 1878 -948
rect 1872 -960 1878 -954
rect 1872 -966 1878 -960
rect 1872 -972 1878 -966
rect 1872 -978 1878 -972
rect 1872 -984 1878 -978
rect 1872 -990 1878 -984
rect 1872 -996 1878 -990
rect 1872 -1002 1878 -996
rect 1872 -1008 1878 -1002
rect 1872 -1014 1878 -1008
rect 1872 -1020 1878 -1014
rect 1872 -1026 1878 -1020
rect 1872 -1032 1878 -1026
rect 1872 -1038 1878 -1032
rect 1872 -1044 1878 -1038
rect 1872 -1050 1878 -1044
rect 1872 -1056 1878 -1050
rect 1872 -1062 1878 -1056
rect 1872 -1068 1878 -1062
rect 1872 -1074 1878 -1068
rect 1872 -1080 1878 -1074
rect 1872 -1086 1878 -1080
rect 1872 -1092 1878 -1086
rect 1872 -1098 1878 -1092
rect 1872 -1104 1878 -1098
rect 1872 -1110 1878 -1104
rect 1872 -1116 1878 -1110
rect 1872 -1122 1878 -1116
rect 1872 -1128 1878 -1122
rect 1872 -1134 1878 -1128
rect 1872 -1140 1878 -1134
rect 1872 -1146 1878 -1140
rect 1872 -1152 1878 -1146
rect 1872 -1158 1878 -1152
rect 1872 -1164 1878 -1158
rect 1872 -1170 1878 -1164
rect 1872 -1176 1878 -1170
rect 1872 -1182 1878 -1176
rect 1872 -1188 1878 -1182
rect 1872 -1194 1878 -1188
rect 1872 -1200 1878 -1194
rect 1872 -1206 1878 -1200
rect 1872 -1212 1878 -1206
rect 1872 -1218 1878 -1212
rect 1872 -1224 1878 -1218
rect 1872 -1230 1878 -1224
rect 1872 -1236 1878 -1230
rect 1872 -1242 1878 -1236
rect 1872 -1248 1878 -1242
rect 1872 -1254 1878 -1248
rect 1872 -1260 1878 -1254
rect 1872 -1266 1878 -1260
rect 1872 -1272 1878 -1266
rect 1872 -1278 1878 -1272
rect 1872 -1284 1878 -1278
rect 1872 -1290 1878 -1284
rect 1872 -1296 1878 -1290
rect 1872 -1302 1878 -1296
rect 1872 -1308 1878 -1302
rect 1872 -1314 1878 -1308
rect 1872 -1320 1878 -1314
rect 1872 -1326 1878 -1320
rect 1872 -1332 1878 -1326
rect 1872 -1338 1878 -1332
rect 1872 -1344 1878 -1338
rect 1872 -1350 1878 -1344
rect 1872 -1356 1878 -1350
rect 1872 -1362 1878 -1356
rect 1872 -1368 1878 -1362
rect 1872 -1374 1878 -1368
rect 1872 -1380 1878 -1374
rect 1872 -1386 1878 -1380
rect 1872 -1392 1878 -1386
rect 1872 -1398 1878 -1392
rect 1872 -1404 1878 -1398
rect 1872 -1410 1878 -1404
rect 1872 -1416 1878 -1410
rect 1872 -1422 1878 -1416
rect 1872 -1428 1878 -1422
rect 1872 -1434 1878 -1428
rect 1872 -1440 1878 -1434
rect 1872 -1446 1878 -1440
rect 1872 -1452 1878 -1446
rect 1872 -1458 1878 -1452
rect 1872 -1464 1878 -1458
rect 1872 -1470 1878 -1464
rect 1872 -1476 1878 -1470
rect 1872 -1482 1878 -1476
rect 1872 -1488 1878 -1482
rect 1872 -1494 1878 -1488
rect 1872 -1500 1878 -1494
rect 1872 -1506 1878 -1500
rect 1872 -1512 1878 -1506
rect 1872 -1518 1878 -1512
rect 1872 -1524 1878 -1518
rect 1872 -1530 1878 -1524
rect 1872 -1536 1878 -1530
rect 1872 -1542 1878 -1536
rect 1872 -1548 1878 -1542
rect 1872 -1554 1878 -1548
rect 1872 -1560 1878 -1554
rect 1872 -1566 1878 -1560
rect 1872 -1572 1878 -1566
rect 1872 -1578 1878 -1572
rect 1872 -1584 1878 -1578
rect 1872 -1590 1878 -1584
rect 1872 -1596 1878 -1590
rect 1872 -1602 1878 -1596
rect 1872 -1608 1878 -1602
rect 1872 -1614 1878 -1608
rect 1872 -1620 1878 -1614
rect 1872 -1626 1878 -1620
rect 1872 -1632 1878 -1626
rect 1872 -1638 1878 -1632
rect 1872 -1644 1878 -1638
rect 1872 -1650 1878 -1644
rect 1872 -1656 1878 -1650
rect 1872 -1662 1878 -1656
rect 1872 -1668 1878 -1662
rect 1872 -1674 1878 -1668
rect 1872 -1680 1878 -1674
rect 1872 -1686 1878 -1680
rect 1872 -1692 1878 -1686
rect 1872 -1698 1878 -1692
rect 1872 -1704 1878 -1698
rect 1872 -1710 1878 -1704
rect 1872 -1716 1878 -1710
rect 1872 -1722 1878 -1716
rect 1872 -1728 1878 -1722
rect 1872 -1734 1878 -1728
rect 1872 -1740 1878 -1734
rect 1872 -1746 1878 -1740
rect 1872 -1752 1878 -1746
rect 1872 -1758 1878 -1752
rect 1872 -1764 1878 -1758
rect 1872 -1770 1878 -1764
rect 1872 -1776 1878 -1770
rect 1872 -1854 1878 -1848
rect 1872 -1860 1878 -1854
rect 1872 -1866 1878 -1860
rect 1872 -1872 1878 -1866
rect 1872 -1878 1878 -1872
rect 1872 -1884 1878 -1878
rect 1872 -1890 1878 -1884
rect 1872 -1896 1878 -1890
rect 1872 -1902 1878 -1896
rect 1872 -1908 1878 -1902
rect 1872 -1914 1878 -1908
rect 1872 -1920 1878 -1914
rect 1872 -1926 1878 -1920
rect 1872 -1932 1878 -1926
rect 1872 -1938 1878 -1932
rect 1872 -1944 1878 -1938
rect 1872 -1950 1878 -1944
rect 1872 -1956 1878 -1950
rect 1872 -1962 1878 -1956
rect 1872 -1968 1878 -1962
rect 1872 -1974 1878 -1968
rect 1872 -1980 1878 -1974
rect 1872 -1986 1878 -1980
rect 1872 -1992 1878 -1986
rect 1872 -1998 1878 -1992
rect 1872 -2004 1878 -1998
rect 1872 -2010 1878 -2004
rect 1872 -2016 1878 -2010
rect 1872 -2022 1878 -2016
rect 1872 -2028 1878 -2022
rect 1872 -2034 1878 -2028
rect 1872 -2040 1878 -2034
rect 1872 -2046 1878 -2040
rect 1872 -2052 1878 -2046
rect 1872 -2058 1878 -2052
rect 1872 -2064 1878 -2058
rect 1872 -2070 1878 -2064
rect 1872 -2076 1878 -2070
rect 1872 -2082 1878 -2076
rect 1872 -2088 1878 -2082
rect 1872 -2094 1878 -2088
rect 1872 -2100 1878 -2094
rect 1872 -2106 1878 -2100
rect 1872 -2112 1878 -2106
rect 1872 -2118 1878 -2112
rect 1872 -2124 1878 -2118
rect 1872 -2130 1878 -2124
rect 1872 -2136 1878 -2130
rect 1872 -2142 1878 -2136
rect 1872 -2148 1878 -2142
rect 1872 -2154 1878 -2148
rect 1872 -2160 1878 -2154
rect 1872 -2166 1878 -2160
rect 1872 -2172 1878 -2166
rect 1872 -2178 1878 -2172
rect 1872 -2184 1878 -2178
rect 1872 -2190 1878 -2184
rect 1872 -2196 1878 -2190
rect 1872 -2202 1878 -2196
rect 1872 -2208 1878 -2202
rect 1872 -2214 1878 -2208
rect 1872 -2220 1878 -2214
rect 1872 -2226 1878 -2220
rect 1872 -2232 1878 -2226
rect 1872 -2238 1878 -2232
rect 1872 -2244 1878 -2238
rect 1872 -2250 1878 -2244
rect 1872 -2256 1878 -2250
rect 1872 -2262 1878 -2256
rect 1872 -2268 1878 -2262
rect 1872 -2274 1878 -2268
rect 1872 -2280 1878 -2274
rect 1872 -2286 1878 -2280
rect 1872 -2292 1878 -2286
rect 1872 -2298 1878 -2292
rect 1872 -2304 1878 -2298
rect 1872 -2310 1878 -2304
rect 1872 -2316 1878 -2310
rect 1872 -2322 1878 -2316
rect 1872 -2328 1878 -2322
rect 1872 -2334 1878 -2328
rect 1872 -2340 1878 -2334
rect 1872 -2346 1878 -2340
rect 1872 -2352 1878 -2346
rect 1872 -2358 1878 -2352
rect 1872 -2364 1878 -2358
rect 1872 -2370 1878 -2364
rect 1872 -2376 1878 -2370
rect 1872 -2382 1878 -2376
rect 1872 -2388 1878 -2382
rect 1872 -2394 1878 -2388
rect 1872 -2400 1878 -2394
rect 1872 -2406 1878 -2400
rect 1872 -2412 1878 -2406
rect 1872 -2418 1878 -2412
rect 1872 -2424 1878 -2418
rect 1872 -2430 1878 -2424
rect 1872 -2436 1878 -2430
rect 1872 -2442 1878 -2436
rect 1872 -2448 1878 -2442
rect 1872 -2454 1878 -2448
rect 1872 -2460 1878 -2454
rect 1872 -2466 1878 -2460
rect 1872 -2472 1878 -2466
rect 1872 -2478 1878 -2472
rect 1872 -2484 1878 -2478
rect 1872 -2490 1878 -2484
rect 1872 -2496 1878 -2490
rect 1872 -2502 1878 -2496
rect 1872 -2508 1878 -2502
rect 1872 -2514 1878 -2508
rect 1872 -2520 1878 -2514
rect 1872 -2526 1878 -2520
rect 1872 -2532 1878 -2526
rect 1872 -2538 1878 -2532
rect 1872 -2544 1878 -2538
rect 1872 -2550 1878 -2544
rect 1872 -2556 1878 -2550
rect 1872 -2562 1878 -2556
rect 1872 -2568 1878 -2562
rect 1872 -2574 1878 -2568
rect 1872 -2580 1878 -2574
rect 1872 -2586 1878 -2580
rect 1872 -2592 1878 -2586
rect 1872 -2670 1878 -2664
rect 1872 -2676 1878 -2670
rect 1872 -2682 1878 -2676
rect 1872 -2688 1878 -2682
rect 1872 -2694 1878 -2688
rect 1872 -2700 1878 -2694
rect 1872 -2706 1878 -2700
rect 1872 -2712 1878 -2706
rect 1872 -2718 1878 -2712
rect 1872 -2724 1878 -2718
rect 1872 -2730 1878 -2724
rect 1872 -2736 1878 -2730
rect 1872 -2742 1878 -2736
rect 1872 -2748 1878 -2742
rect 1872 -2754 1878 -2748
rect 1872 -2760 1878 -2754
rect 1872 -2766 1878 -2760
rect 1872 -2772 1878 -2766
rect 1872 -2778 1878 -2772
rect 1872 -2784 1878 -2778
rect 1872 -2790 1878 -2784
rect 1872 -2796 1878 -2790
rect 1872 -2802 1878 -2796
rect 1872 -2808 1878 -2802
rect 1872 -2814 1878 -2808
rect 1872 -2820 1878 -2814
rect 1872 -2826 1878 -2820
rect 1872 -2832 1878 -2826
rect 1872 -2838 1878 -2832
rect 1872 -2844 1878 -2838
rect 1872 -2850 1878 -2844
rect 1872 -2856 1878 -2850
rect 1872 -2862 1878 -2856
rect 1872 -2868 1878 -2862
rect 1872 -2874 1878 -2868
rect 1872 -2880 1878 -2874
rect 1872 -2886 1878 -2880
rect 1872 -2892 1878 -2886
rect 1872 -2898 1878 -2892
rect 1872 -2904 1878 -2898
rect 1872 -2910 1878 -2904
rect 1872 -2916 1878 -2910
rect 1872 -2922 1878 -2916
rect 1872 -2928 1878 -2922
rect 1872 -2934 1878 -2928
rect 1872 -2940 1878 -2934
rect 1872 -2946 1878 -2940
rect 1872 -2952 1878 -2946
rect 1872 -2958 1878 -2952
rect 1872 -2964 1878 -2958
rect 1872 -2970 1878 -2964
rect 1872 -2976 1878 -2970
rect 1872 -2982 1878 -2976
rect 1872 -2988 1878 -2982
rect 1872 -2994 1878 -2988
rect 1872 -3000 1878 -2994
rect 1872 -3006 1878 -3000
rect 1872 -3012 1878 -3006
rect 1872 -3018 1878 -3012
rect 1872 -3024 1878 -3018
rect 1872 -3030 1878 -3024
rect 1872 -3036 1878 -3030
rect 1872 -3042 1878 -3036
rect 1872 -3048 1878 -3042
rect 1872 -3054 1878 -3048
rect 1872 -3060 1878 -3054
rect 1872 -3066 1878 -3060
rect 1872 -3072 1878 -3066
rect 1872 -3078 1878 -3072
rect 1872 -3084 1878 -3078
rect 1872 -3090 1878 -3084
rect 1872 -3096 1878 -3090
rect 1872 -3102 1878 -3096
rect 1872 -3108 1878 -3102
rect 1872 -3114 1878 -3108
rect 1872 -3120 1878 -3114
rect 1872 -3126 1878 -3120
rect 1872 -3132 1878 -3126
rect 1872 -3138 1878 -3132
rect 1872 -3144 1878 -3138
rect 1872 -3150 1878 -3144
rect 1872 -3156 1878 -3150
rect 1872 -3204 1878 -3198
rect 1872 -3210 1878 -3204
rect 1872 -3216 1878 -3210
rect 1872 -3222 1878 -3216
rect 1872 -3228 1878 -3222
rect 1872 -3234 1878 -3228
rect 1872 -3240 1878 -3234
rect 1872 -3246 1878 -3240
rect 1872 -3252 1878 -3246
rect 1872 -3258 1878 -3252
rect 1872 -3264 1878 -3258
rect 1872 -3270 1878 -3264
rect 1872 -3276 1878 -3270
rect 1872 -3282 1878 -3276
rect 1872 -3288 1878 -3282
rect 1872 -3294 1878 -3288
rect 1872 -3300 1878 -3294
rect 1872 -3306 1878 -3300
rect 1872 -3312 1878 -3306
rect 1872 -3318 1878 -3312
rect 1872 -3324 1878 -3318
rect 1878 -612 1884 -606
rect 1878 -618 1884 -612
rect 1878 -624 1884 -618
rect 1878 -630 1884 -624
rect 1878 -636 1884 -630
rect 1878 -642 1884 -636
rect 1878 -648 1884 -642
rect 1878 -654 1884 -648
rect 1878 -660 1884 -654
rect 1878 -666 1884 -660
rect 1878 -672 1884 -666
rect 1878 -678 1884 -672
rect 1878 -684 1884 -678
rect 1878 -690 1884 -684
rect 1878 -696 1884 -690
rect 1878 -702 1884 -696
rect 1878 -708 1884 -702
rect 1878 -714 1884 -708
rect 1878 -720 1884 -714
rect 1878 -726 1884 -720
rect 1878 -732 1884 -726
rect 1878 -738 1884 -732
rect 1878 -744 1884 -738
rect 1878 -750 1884 -744
rect 1878 -756 1884 -750
rect 1878 -762 1884 -756
rect 1878 -768 1884 -762
rect 1878 -774 1884 -768
rect 1878 -780 1884 -774
rect 1878 -786 1884 -780
rect 1878 -792 1884 -786
rect 1878 -798 1884 -792
rect 1878 -804 1884 -798
rect 1878 -810 1884 -804
rect 1878 -816 1884 -810
rect 1878 -822 1884 -816
rect 1878 -828 1884 -822
rect 1878 -834 1884 -828
rect 1878 -840 1884 -834
rect 1878 -846 1884 -840
rect 1878 -852 1884 -846
rect 1878 -858 1884 -852
rect 1878 -864 1884 -858
rect 1878 -870 1884 -864
rect 1878 -876 1884 -870
rect 1878 -882 1884 -876
rect 1878 -888 1884 -882
rect 1878 -894 1884 -888
rect 1878 -900 1884 -894
rect 1878 -906 1884 -900
rect 1878 -912 1884 -906
rect 1878 -918 1884 -912
rect 1878 -924 1884 -918
rect 1878 -930 1884 -924
rect 1878 -936 1884 -930
rect 1878 -942 1884 -936
rect 1878 -948 1884 -942
rect 1878 -954 1884 -948
rect 1878 -960 1884 -954
rect 1878 -966 1884 -960
rect 1878 -972 1884 -966
rect 1878 -978 1884 -972
rect 1878 -984 1884 -978
rect 1878 -990 1884 -984
rect 1878 -996 1884 -990
rect 1878 -1002 1884 -996
rect 1878 -1008 1884 -1002
rect 1878 -1014 1884 -1008
rect 1878 -1020 1884 -1014
rect 1878 -1026 1884 -1020
rect 1878 -1032 1884 -1026
rect 1878 -1038 1884 -1032
rect 1878 -1044 1884 -1038
rect 1878 -1050 1884 -1044
rect 1878 -1056 1884 -1050
rect 1878 -1062 1884 -1056
rect 1878 -1068 1884 -1062
rect 1878 -1074 1884 -1068
rect 1878 -1080 1884 -1074
rect 1878 -1086 1884 -1080
rect 1878 -1092 1884 -1086
rect 1878 -1098 1884 -1092
rect 1878 -1104 1884 -1098
rect 1878 -1110 1884 -1104
rect 1878 -1116 1884 -1110
rect 1878 -1122 1884 -1116
rect 1878 -1128 1884 -1122
rect 1878 -1134 1884 -1128
rect 1878 -1140 1884 -1134
rect 1878 -1146 1884 -1140
rect 1878 -1152 1884 -1146
rect 1878 -1158 1884 -1152
rect 1878 -1164 1884 -1158
rect 1878 -1170 1884 -1164
rect 1878 -1176 1884 -1170
rect 1878 -1182 1884 -1176
rect 1878 -1188 1884 -1182
rect 1878 -1194 1884 -1188
rect 1878 -1200 1884 -1194
rect 1878 -1206 1884 -1200
rect 1878 -1212 1884 -1206
rect 1878 -1218 1884 -1212
rect 1878 -1224 1884 -1218
rect 1878 -1230 1884 -1224
rect 1878 -1236 1884 -1230
rect 1878 -1242 1884 -1236
rect 1878 -1248 1884 -1242
rect 1878 -1254 1884 -1248
rect 1878 -1260 1884 -1254
rect 1878 -1266 1884 -1260
rect 1878 -1272 1884 -1266
rect 1878 -1278 1884 -1272
rect 1878 -1284 1884 -1278
rect 1878 -1290 1884 -1284
rect 1878 -1296 1884 -1290
rect 1878 -1302 1884 -1296
rect 1878 -1308 1884 -1302
rect 1878 -1314 1884 -1308
rect 1878 -1320 1884 -1314
rect 1878 -1326 1884 -1320
rect 1878 -1332 1884 -1326
rect 1878 -1338 1884 -1332
rect 1878 -1344 1884 -1338
rect 1878 -1350 1884 -1344
rect 1878 -1356 1884 -1350
rect 1878 -1362 1884 -1356
rect 1878 -1368 1884 -1362
rect 1878 -1374 1884 -1368
rect 1878 -1380 1884 -1374
rect 1878 -1386 1884 -1380
rect 1878 -1392 1884 -1386
rect 1878 -1398 1884 -1392
rect 1878 -1404 1884 -1398
rect 1878 -1410 1884 -1404
rect 1878 -1416 1884 -1410
rect 1878 -1422 1884 -1416
rect 1878 -1428 1884 -1422
rect 1878 -1434 1884 -1428
rect 1878 -1440 1884 -1434
rect 1878 -1446 1884 -1440
rect 1878 -1452 1884 -1446
rect 1878 -1458 1884 -1452
rect 1878 -1464 1884 -1458
rect 1878 -1470 1884 -1464
rect 1878 -1476 1884 -1470
rect 1878 -1482 1884 -1476
rect 1878 -1488 1884 -1482
rect 1878 -1494 1884 -1488
rect 1878 -1500 1884 -1494
rect 1878 -1506 1884 -1500
rect 1878 -1512 1884 -1506
rect 1878 -1518 1884 -1512
rect 1878 -1524 1884 -1518
rect 1878 -1530 1884 -1524
rect 1878 -1536 1884 -1530
rect 1878 -1542 1884 -1536
rect 1878 -1548 1884 -1542
rect 1878 -1554 1884 -1548
rect 1878 -1560 1884 -1554
rect 1878 -1566 1884 -1560
rect 1878 -1572 1884 -1566
rect 1878 -1578 1884 -1572
rect 1878 -1584 1884 -1578
rect 1878 -1590 1884 -1584
rect 1878 -1596 1884 -1590
rect 1878 -1602 1884 -1596
rect 1878 -1608 1884 -1602
rect 1878 -1614 1884 -1608
rect 1878 -1620 1884 -1614
rect 1878 -1626 1884 -1620
rect 1878 -1632 1884 -1626
rect 1878 -1638 1884 -1632
rect 1878 -1644 1884 -1638
rect 1878 -1650 1884 -1644
rect 1878 -1656 1884 -1650
rect 1878 -1662 1884 -1656
rect 1878 -1668 1884 -1662
rect 1878 -1674 1884 -1668
rect 1878 -1680 1884 -1674
rect 1878 -1686 1884 -1680
rect 1878 -1692 1884 -1686
rect 1878 -1698 1884 -1692
rect 1878 -1704 1884 -1698
rect 1878 -1710 1884 -1704
rect 1878 -1716 1884 -1710
rect 1878 -1722 1884 -1716
rect 1878 -1728 1884 -1722
rect 1878 -1734 1884 -1728
rect 1878 -1740 1884 -1734
rect 1878 -1746 1884 -1740
rect 1878 -1752 1884 -1746
rect 1878 -1758 1884 -1752
rect 1878 -1764 1884 -1758
rect 1878 -1770 1884 -1764
rect 1878 -1848 1884 -1842
rect 1878 -1854 1884 -1848
rect 1878 -1860 1884 -1854
rect 1878 -1866 1884 -1860
rect 1878 -1872 1884 -1866
rect 1878 -1878 1884 -1872
rect 1878 -1884 1884 -1878
rect 1878 -1890 1884 -1884
rect 1878 -1896 1884 -1890
rect 1878 -1902 1884 -1896
rect 1878 -1908 1884 -1902
rect 1878 -1914 1884 -1908
rect 1878 -1920 1884 -1914
rect 1878 -1926 1884 -1920
rect 1878 -1932 1884 -1926
rect 1878 -1938 1884 -1932
rect 1878 -1944 1884 -1938
rect 1878 -1950 1884 -1944
rect 1878 -1956 1884 -1950
rect 1878 -1962 1884 -1956
rect 1878 -1968 1884 -1962
rect 1878 -1974 1884 -1968
rect 1878 -1980 1884 -1974
rect 1878 -1986 1884 -1980
rect 1878 -1992 1884 -1986
rect 1878 -1998 1884 -1992
rect 1878 -2004 1884 -1998
rect 1878 -2010 1884 -2004
rect 1878 -2016 1884 -2010
rect 1878 -2022 1884 -2016
rect 1878 -2028 1884 -2022
rect 1878 -2034 1884 -2028
rect 1878 -2040 1884 -2034
rect 1878 -2046 1884 -2040
rect 1878 -2052 1884 -2046
rect 1878 -2058 1884 -2052
rect 1878 -2064 1884 -2058
rect 1878 -2070 1884 -2064
rect 1878 -2076 1884 -2070
rect 1878 -2082 1884 -2076
rect 1878 -2088 1884 -2082
rect 1878 -2094 1884 -2088
rect 1878 -2100 1884 -2094
rect 1878 -2106 1884 -2100
rect 1878 -2112 1884 -2106
rect 1878 -2118 1884 -2112
rect 1878 -2124 1884 -2118
rect 1878 -2130 1884 -2124
rect 1878 -2136 1884 -2130
rect 1878 -2142 1884 -2136
rect 1878 -2148 1884 -2142
rect 1878 -2154 1884 -2148
rect 1878 -2160 1884 -2154
rect 1878 -2166 1884 -2160
rect 1878 -2172 1884 -2166
rect 1878 -2178 1884 -2172
rect 1878 -2184 1884 -2178
rect 1878 -2190 1884 -2184
rect 1878 -2196 1884 -2190
rect 1878 -2202 1884 -2196
rect 1878 -2208 1884 -2202
rect 1878 -2214 1884 -2208
rect 1878 -2220 1884 -2214
rect 1878 -2226 1884 -2220
rect 1878 -2232 1884 -2226
rect 1878 -2238 1884 -2232
rect 1878 -2244 1884 -2238
rect 1878 -2250 1884 -2244
rect 1878 -2256 1884 -2250
rect 1878 -2262 1884 -2256
rect 1878 -2268 1884 -2262
rect 1878 -2274 1884 -2268
rect 1878 -2280 1884 -2274
rect 1878 -2286 1884 -2280
rect 1878 -2292 1884 -2286
rect 1878 -2298 1884 -2292
rect 1878 -2304 1884 -2298
rect 1878 -2310 1884 -2304
rect 1878 -2316 1884 -2310
rect 1878 -2322 1884 -2316
rect 1878 -2328 1884 -2322
rect 1878 -2334 1884 -2328
rect 1878 -2340 1884 -2334
rect 1878 -2346 1884 -2340
rect 1878 -2352 1884 -2346
rect 1878 -2358 1884 -2352
rect 1878 -2364 1884 -2358
rect 1878 -2370 1884 -2364
rect 1878 -2376 1884 -2370
rect 1878 -2382 1884 -2376
rect 1878 -2388 1884 -2382
rect 1878 -2394 1884 -2388
rect 1878 -2400 1884 -2394
rect 1878 -2406 1884 -2400
rect 1878 -2412 1884 -2406
rect 1878 -2418 1884 -2412
rect 1878 -2424 1884 -2418
rect 1878 -2430 1884 -2424
rect 1878 -2436 1884 -2430
rect 1878 -2442 1884 -2436
rect 1878 -2448 1884 -2442
rect 1878 -2454 1884 -2448
rect 1878 -2460 1884 -2454
rect 1878 -2466 1884 -2460
rect 1878 -2472 1884 -2466
rect 1878 -2478 1884 -2472
rect 1878 -2484 1884 -2478
rect 1878 -2490 1884 -2484
rect 1878 -2496 1884 -2490
rect 1878 -2502 1884 -2496
rect 1878 -2508 1884 -2502
rect 1878 -2514 1884 -2508
rect 1878 -2520 1884 -2514
rect 1878 -2526 1884 -2520
rect 1878 -2532 1884 -2526
rect 1878 -2538 1884 -2532
rect 1878 -2544 1884 -2538
rect 1878 -2550 1884 -2544
rect 1878 -2556 1884 -2550
rect 1878 -2562 1884 -2556
rect 1878 -2568 1884 -2562
rect 1878 -2574 1884 -2568
rect 1878 -2580 1884 -2574
rect 1878 -2586 1884 -2580
rect 1878 -2592 1884 -2586
rect 1878 -2664 1884 -2658
rect 1878 -2670 1884 -2664
rect 1878 -2676 1884 -2670
rect 1878 -2682 1884 -2676
rect 1878 -2688 1884 -2682
rect 1878 -2694 1884 -2688
rect 1878 -2700 1884 -2694
rect 1878 -2706 1884 -2700
rect 1878 -2712 1884 -2706
rect 1878 -2718 1884 -2712
rect 1878 -2724 1884 -2718
rect 1878 -2730 1884 -2724
rect 1878 -2736 1884 -2730
rect 1878 -2742 1884 -2736
rect 1878 -2748 1884 -2742
rect 1878 -2754 1884 -2748
rect 1878 -2760 1884 -2754
rect 1878 -2766 1884 -2760
rect 1878 -2772 1884 -2766
rect 1878 -2778 1884 -2772
rect 1878 -2784 1884 -2778
rect 1878 -2790 1884 -2784
rect 1878 -2796 1884 -2790
rect 1878 -2802 1884 -2796
rect 1878 -2808 1884 -2802
rect 1878 -2814 1884 -2808
rect 1878 -2820 1884 -2814
rect 1878 -2826 1884 -2820
rect 1878 -2832 1884 -2826
rect 1878 -2838 1884 -2832
rect 1878 -2844 1884 -2838
rect 1878 -2850 1884 -2844
rect 1878 -2856 1884 -2850
rect 1878 -2862 1884 -2856
rect 1878 -2868 1884 -2862
rect 1878 -2874 1884 -2868
rect 1878 -2880 1884 -2874
rect 1878 -2886 1884 -2880
rect 1878 -2892 1884 -2886
rect 1878 -2898 1884 -2892
rect 1878 -2904 1884 -2898
rect 1878 -2910 1884 -2904
rect 1878 -2916 1884 -2910
rect 1878 -2922 1884 -2916
rect 1878 -2928 1884 -2922
rect 1878 -2934 1884 -2928
rect 1878 -2940 1884 -2934
rect 1878 -2946 1884 -2940
rect 1878 -2952 1884 -2946
rect 1878 -2958 1884 -2952
rect 1878 -2964 1884 -2958
rect 1878 -2970 1884 -2964
rect 1878 -2976 1884 -2970
rect 1878 -2982 1884 -2976
rect 1878 -2988 1884 -2982
rect 1878 -2994 1884 -2988
rect 1878 -3000 1884 -2994
rect 1878 -3006 1884 -3000
rect 1878 -3012 1884 -3006
rect 1878 -3018 1884 -3012
rect 1878 -3024 1884 -3018
rect 1878 -3030 1884 -3024
rect 1878 -3036 1884 -3030
rect 1878 -3042 1884 -3036
rect 1878 -3048 1884 -3042
rect 1878 -3054 1884 -3048
rect 1878 -3060 1884 -3054
rect 1878 -3066 1884 -3060
rect 1878 -3072 1884 -3066
rect 1878 -3078 1884 -3072
rect 1878 -3084 1884 -3078
rect 1878 -3090 1884 -3084
rect 1878 -3096 1884 -3090
rect 1878 -3102 1884 -3096
rect 1878 -3108 1884 -3102
rect 1878 -3114 1884 -3108
rect 1878 -3120 1884 -3114
rect 1878 -3126 1884 -3120
rect 1878 -3132 1884 -3126
rect 1878 -3138 1884 -3132
rect 1878 -3144 1884 -3138
rect 1878 -3150 1884 -3144
rect 1878 -3204 1884 -3198
rect 1878 -3210 1884 -3204
rect 1878 -3216 1884 -3210
rect 1878 -3222 1884 -3216
rect 1878 -3228 1884 -3222
rect 1878 -3234 1884 -3228
rect 1878 -3240 1884 -3234
rect 1878 -3246 1884 -3240
rect 1878 -3252 1884 -3246
rect 1878 -3258 1884 -3252
rect 1878 -3264 1884 -3258
rect 1878 -3270 1884 -3264
rect 1878 -3276 1884 -3270
rect 1878 -3282 1884 -3276
rect 1878 -3288 1884 -3282
rect 1878 -3294 1884 -3288
rect 1878 -3300 1884 -3294
rect 1878 -3306 1884 -3300
rect 1878 -3312 1884 -3306
rect 1878 -3318 1884 -3312
rect 1884 -606 1890 -600
rect 1884 -612 1890 -606
rect 1884 -618 1890 -612
rect 1884 -624 1890 -618
rect 1884 -630 1890 -624
rect 1884 -636 1890 -630
rect 1884 -642 1890 -636
rect 1884 -648 1890 -642
rect 1884 -654 1890 -648
rect 1884 -660 1890 -654
rect 1884 -666 1890 -660
rect 1884 -672 1890 -666
rect 1884 -678 1890 -672
rect 1884 -684 1890 -678
rect 1884 -690 1890 -684
rect 1884 -696 1890 -690
rect 1884 -702 1890 -696
rect 1884 -708 1890 -702
rect 1884 -714 1890 -708
rect 1884 -720 1890 -714
rect 1884 -726 1890 -720
rect 1884 -732 1890 -726
rect 1884 -738 1890 -732
rect 1884 -744 1890 -738
rect 1884 -750 1890 -744
rect 1884 -756 1890 -750
rect 1884 -762 1890 -756
rect 1884 -768 1890 -762
rect 1884 -774 1890 -768
rect 1884 -780 1890 -774
rect 1884 -786 1890 -780
rect 1884 -792 1890 -786
rect 1884 -798 1890 -792
rect 1884 -804 1890 -798
rect 1884 -810 1890 -804
rect 1884 -816 1890 -810
rect 1884 -822 1890 -816
rect 1884 -828 1890 -822
rect 1884 -834 1890 -828
rect 1884 -840 1890 -834
rect 1884 -846 1890 -840
rect 1884 -852 1890 -846
rect 1884 -858 1890 -852
rect 1884 -864 1890 -858
rect 1884 -870 1890 -864
rect 1884 -876 1890 -870
rect 1884 -882 1890 -876
rect 1884 -888 1890 -882
rect 1884 -894 1890 -888
rect 1884 -900 1890 -894
rect 1884 -906 1890 -900
rect 1884 -912 1890 -906
rect 1884 -918 1890 -912
rect 1884 -924 1890 -918
rect 1884 -930 1890 -924
rect 1884 -936 1890 -930
rect 1884 -942 1890 -936
rect 1884 -948 1890 -942
rect 1884 -954 1890 -948
rect 1884 -960 1890 -954
rect 1884 -966 1890 -960
rect 1884 -972 1890 -966
rect 1884 -978 1890 -972
rect 1884 -984 1890 -978
rect 1884 -990 1890 -984
rect 1884 -996 1890 -990
rect 1884 -1002 1890 -996
rect 1884 -1008 1890 -1002
rect 1884 -1014 1890 -1008
rect 1884 -1020 1890 -1014
rect 1884 -1026 1890 -1020
rect 1884 -1032 1890 -1026
rect 1884 -1038 1890 -1032
rect 1884 -1044 1890 -1038
rect 1884 -1050 1890 -1044
rect 1884 -1056 1890 -1050
rect 1884 -1062 1890 -1056
rect 1884 -1068 1890 -1062
rect 1884 -1074 1890 -1068
rect 1884 -1080 1890 -1074
rect 1884 -1086 1890 -1080
rect 1884 -1092 1890 -1086
rect 1884 -1098 1890 -1092
rect 1884 -1104 1890 -1098
rect 1884 -1110 1890 -1104
rect 1884 -1116 1890 -1110
rect 1884 -1122 1890 -1116
rect 1884 -1128 1890 -1122
rect 1884 -1134 1890 -1128
rect 1884 -1140 1890 -1134
rect 1884 -1146 1890 -1140
rect 1884 -1152 1890 -1146
rect 1884 -1158 1890 -1152
rect 1884 -1164 1890 -1158
rect 1884 -1170 1890 -1164
rect 1884 -1176 1890 -1170
rect 1884 -1182 1890 -1176
rect 1884 -1188 1890 -1182
rect 1884 -1194 1890 -1188
rect 1884 -1200 1890 -1194
rect 1884 -1206 1890 -1200
rect 1884 -1212 1890 -1206
rect 1884 -1218 1890 -1212
rect 1884 -1224 1890 -1218
rect 1884 -1230 1890 -1224
rect 1884 -1236 1890 -1230
rect 1884 -1242 1890 -1236
rect 1884 -1248 1890 -1242
rect 1884 -1254 1890 -1248
rect 1884 -1260 1890 -1254
rect 1884 -1266 1890 -1260
rect 1884 -1272 1890 -1266
rect 1884 -1278 1890 -1272
rect 1884 -1284 1890 -1278
rect 1884 -1290 1890 -1284
rect 1884 -1296 1890 -1290
rect 1884 -1302 1890 -1296
rect 1884 -1308 1890 -1302
rect 1884 -1314 1890 -1308
rect 1884 -1320 1890 -1314
rect 1884 -1326 1890 -1320
rect 1884 -1332 1890 -1326
rect 1884 -1338 1890 -1332
rect 1884 -1344 1890 -1338
rect 1884 -1350 1890 -1344
rect 1884 -1356 1890 -1350
rect 1884 -1362 1890 -1356
rect 1884 -1368 1890 -1362
rect 1884 -1374 1890 -1368
rect 1884 -1380 1890 -1374
rect 1884 -1386 1890 -1380
rect 1884 -1392 1890 -1386
rect 1884 -1398 1890 -1392
rect 1884 -1404 1890 -1398
rect 1884 -1410 1890 -1404
rect 1884 -1416 1890 -1410
rect 1884 -1422 1890 -1416
rect 1884 -1428 1890 -1422
rect 1884 -1434 1890 -1428
rect 1884 -1440 1890 -1434
rect 1884 -1446 1890 -1440
rect 1884 -1452 1890 -1446
rect 1884 -1458 1890 -1452
rect 1884 -1464 1890 -1458
rect 1884 -1470 1890 -1464
rect 1884 -1476 1890 -1470
rect 1884 -1482 1890 -1476
rect 1884 -1488 1890 -1482
rect 1884 -1494 1890 -1488
rect 1884 -1500 1890 -1494
rect 1884 -1506 1890 -1500
rect 1884 -1512 1890 -1506
rect 1884 -1518 1890 -1512
rect 1884 -1524 1890 -1518
rect 1884 -1530 1890 -1524
rect 1884 -1536 1890 -1530
rect 1884 -1542 1890 -1536
rect 1884 -1548 1890 -1542
rect 1884 -1554 1890 -1548
rect 1884 -1560 1890 -1554
rect 1884 -1566 1890 -1560
rect 1884 -1572 1890 -1566
rect 1884 -1578 1890 -1572
rect 1884 -1584 1890 -1578
rect 1884 -1590 1890 -1584
rect 1884 -1596 1890 -1590
rect 1884 -1602 1890 -1596
rect 1884 -1608 1890 -1602
rect 1884 -1614 1890 -1608
rect 1884 -1620 1890 -1614
rect 1884 -1626 1890 -1620
rect 1884 -1632 1890 -1626
rect 1884 -1638 1890 -1632
rect 1884 -1644 1890 -1638
rect 1884 -1650 1890 -1644
rect 1884 -1656 1890 -1650
rect 1884 -1662 1890 -1656
rect 1884 -1668 1890 -1662
rect 1884 -1674 1890 -1668
rect 1884 -1680 1890 -1674
rect 1884 -1686 1890 -1680
rect 1884 -1692 1890 -1686
rect 1884 -1698 1890 -1692
rect 1884 -1704 1890 -1698
rect 1884 -1710 1890 -1704
rect 1884 -1716 1890 -1710
rect 1884 -1722 1890 -1716
rect 1884 -1728 1890 -1722
rect 1884 -1734 1890 -1728
rect 1884 -1740 1890 -1734
rect 1884 -1746 1890 -1740
rect 1884 -1752 1890 -1746
rect 1884 -1758 1890 -1752
rect 1884 -1764 1890 -1758
rect 1884 -1842 1890 -1836
rect 1884 -1848 1890 -1842
rect 1884 -1854 1890 -1848
rect 1884 -1860 1890 -1854
rect 1884 -1866 1890 -1860
rect 1884 -1872 1890 -1866
rect 1884 -1878 1890 -1872
rect 1884 -1884 1890 -1878
rect 1884 -1890 1890 -1884
rect 1884 -1896 1890 -1890
rect 1884 -1902 1890 -1896
rect 1884 -1908 1890 -1902
rect 1884 -1914 1890 -1908
rect 1884 -1920 1890 -1914
rect 1884 -1926 1890 -1920
rect 1884 -1932 1890 -1926
rect 1884 -1938 1890 -1932
rect 1884 -1944 1890 -1938
rect 1884 -1950 1890 -1944
rect 1884 -1956 1890 -1950
rect 1884 -1962 1890 -1956
rect 1884 -1968 1890 -1962
rect 1884 -1974 1890 -1968
rect 1884 -1980 1890 -1974
rect 1884 -1986 1890 -1980
rect 1884 -1992 1890 -1986
rect 1884 -1998 1890 -1992
rect 1884 -2004 1890 -1998
rect 1884 -2010 1890 -2004
rect 1884 -2016 1890 -2010
rect 1884 -2022 1890 -2016
rect 1884 -2028 1890 -2022
rect 1884 -2034 1890 -2028
rect 1884 -2040 1890 -2034
rect 1884 -2046 1890 -2040
rect 1884 -2052 1890 -2046
rect 1884 -2058 1890 -2052
rect 1884 -2064 1890 -2058
rect 1884 -2070 1890 -2064
rect 1884 -2076 1890 -2070
rect 1884 -2082 1890 -2076
rect 1884 -2088 1890 -2082
rect 1884 -2094 1890 -2088
rect 1884 -2100 1890 -2094
rect 1884 -2106 1890 -2100
rect 1884 -2112 1890 -2106
rect 1884 -2118 1890 -2112
rect 1884 -2124 1890 -2118
rect 1884 -2130 1890 -2124
rect 1884 -2136 1890 -2130
rect 1884 -2142 1890 -2136
rect 1884 -2148 1890 -2142
rect 1884 -2154 1890 -2148
rect 1884 -2160 1890 -2154
rect 1884 -2166 1890 -2160
rect 1884 -2172 1890 -2166
rect 1884 -2178 1890 -2172
rect 1884 -2184 1890 -2178
rect 1884 -2190 1890 -2184
rect 1884 -2196 1890 -2190
rect 1884 -2202 1890 -2196
rect 1884 -2208 1890 -2202
rect 1884 -2214 1890 -2208
rect 1884 -2220 1890 -2214
rect 1884 -2226 1890 -2220
rect 1884 -2232 1890 -2226
rect 1884 -2238 1890 -2232
rect 1884 -2244 1890 -2238
rect 1884 -2250 1890 -2244
rect 1884 -2256 1890 -2250
rect 1884 -2262 1890 -2256
rect 1884 -2268 1890 -2262
rect 1884 -2274 1890 -2268
rect 1884 -2280 1890 -2274
rect 1884 -2286 1890 -2280
rect 1884 -2292 1890 -2286
rect 1884 -2298 1890 -2292
rect 1884 -2304 1890 -2298
rect 1884 -2310 1890 -2304
rect 1884 -2316 1890 -2310
rect 1884 -2322 1890 -2316
rect 1884 -2328 1890 -2322
rect 1884 -2334 1890 -2328
rect 1884 -2340 1890 -2334
rect 1884 -2346 1890 -2340
rect 1884 -2352 1890 -2346
rect 1884 -2358 1890 -2352
rect 1884 -2364 1890 -2358
rect 1884 -2370 1890 -2364
rect 1884 -2376 1890 -2370
rect 1884 -2382 1890 -2376
rect 1884 -2388 1890 -2382
rect 1884 -2394 1890 -2388
rect 1884 -2400 1890 -2394
rect 1884 -2406 1890 -2400
rect 1884 -2412 1890 -2406
rect 1884 -2418 1890 -2412
rect 1884 -2424 1890 -2418
rect 1884 -2430 1890 -2424
rect 1884 -2436 1890 -2430
rect 1884 -2442 1890 -2436
rect 1884 -2448 1890 -2442
rect 1884 -2454 1890 -2448
rect 1884 -2460 1890 -2454
rect 1884 -2466 1890 -2460
rect 1884 -2472 1890 -2466
rect 1884 -2478 1890 -2472
rect 1884 -2484 1890 -2478
rect 1884 -2490 1890 -2484
rect 1884 -2496 1890 -2490
rect 1884 -2502 1890 -2496
rect 1884 -2508 1890 -2502
rect 1884 -2514 1890 -2508
rect 1884 -2520 1890 -2514
rect 1884 -2526 1890 -2520
rect 1884 -2532 1890 -2526
rect 1884 -2538 1890 -2532
rect 1884 -2544 1890 -2538
rect 1884 -2550 1890 -2544
rect 1884 -2556 1890 -2550
rect 1884 -2562 1890 -2556
rect 1884 -2568 1890 -2562
rect 1884 -2574 1890 -2568
rect 1884 -2580 1890 -2574
rect 1884 -2586 1890 -2580
rect 1884 -2664 1890 -2658
rect 1884 -2670 1890 -2664
rect 1884 -2676 1890 -2670
rect 1884 -2682 1890 -2676
rect 1884 -2688 1890 -2682
rect 1884 -2694 1890 -2688
rect 1884 -2700 1890 -2694
rect 1884 -2706 1890 -2700
rect 1884 -2712 1890 -2706
rect 1884 -2718 1890 -2712
rect 1884 -2724 1890 -2718
rect 1884 -2730 1890 -2724
rect 1884 -2736 1890 -2730
rect 1884 -2742 1890 -2736
rect 1884 -2748 1890 -2742
rect 1884 -2754 1890 -2748
rect 1884 -2760 1890 -2754
rect 1884 -2766 1890 -2760
rect 1884 -2772 1890 -2766
rect 1884 -2778 1890 -2772
rect 1884 -2784 1890 -2778
rect 1884 -2790 1890 -2784
rect 1884 -2796 1890 -2790
rect 1884 -2802 1890 -2796
rect 1884 -2808 1890 -2802
rect 1884 -2814 1890 -2808
rect 1884 -2820 1890 -2814
rect 1884 -2826 1890 -2820
rect 1884 -2832 1890 -2826
rect 1884 -2838 1890 -2832
rect 1884 -2844 1890 -2838
rect 1884 -2850 1890 -2844
rect 1884 -2856 1890 -2850
rect 1884 -2862 1890 -2856
rect 1884 -2868 1890 -2862
rect 1884 -2874 1890 -2868
rect 1884 -2880 1890 -2874
rect 1884 -2886 1890 -2880
rect 1884 -2892 1890 -2886
rect 1884 -2898 1890 -2892
rect 1884 -2904 1890 -2898
rect 1884 -2910 1890 -2904
rect 1884 -2916 1890 -2910
rect 1884 -2922 1890 -2916
rect 1884 -2928 1890 -2922
rect 1884 -2934 1890 -2928
rect 1884 -2940 1890 -2934
rect 1884 -2946 1890 -2940
rect 1884 -2952 1890 -2946
rect 1884 -2958 1890 -2952
rect 1884 -2964 1890 -2958
rect 1884 -2970 1890 -2964
rect 1884 -2976 1890 -2970
rect 1884 -2982 1890 -2976
rect 1884 -2988 1890 -2982
rect 1884 -2994 1890 -2988
rect 1884 -3000 1890 -2994
rect 1884 -3006 1890 -3000
rect 1884 -3012 1890 -3006
rect 1884 -3018 1890 -3012
rect 1884 -3024 1890 -3018
rect 1884 -3030 1890 -3024
rect 1884 -3036 1890 -3030
rect 1884 -3042 1890 -3036
rect 1884 -3048 1890 -3042
rect 1884 -3054 1890 -3048
rect 1884 -3060 1890 -3054
rect 1884 -3066 1890 -3060
rect 1884 -3072 1890 -3066
rect 1884 -3078 1890 -3072
rect 1884 -3084 1890 -3078
rect 1884 -3090 1890 -3084
rect 1884 -3096 1890 -3090
rect 1884 -3102 1890 -3096
rect 1884 -3108 1890 -3102
rect 1884 -3114 1890 -3108
rect 1884 -3120 1890 -3114
rect 1884 -3126 1890 -3120
rect 1884 -3132 1890 -3126
rect 1884 -3138 1890 -3132
rect 1884 -3144 1890 -3138
rect 1884 -3150 1890 -3144
rect 1884 -3204 1890 -3198
rect 1884 -3210 1890 -3204
rect 1884 -3216 1890 -3210
rect 1884 -3222 1890 -3216
rect 1884 -3228 1890 -3222
rect 1884 -3234 1890 -3228
rect 1884 -3240 1890 -3234
rect 1884 -3246 1890 -3240
rect 1884 -3252 1890 -3246
rect 1884 -3258 1890 -3252
rect 1884 -3264 1890 -3258
rect 1884 -3270 1890 -3264
rect 1884 -3276 1890 -3270
rect 1884 -3282 1890 -3276
rect 1884 -3288 1890 -3282
rect 1884 -3294 1890 -3288
rect 1884 -3300 1890 -3294
rect 1884 -3306 1890 -3300
rect 1884 -3312 1890 -3306
rect 1890 -594 1896 -588
rect 1890 -600 1896 -594
rect 1890 -606 1896 -600
rect 1890 -612 1896 -606
rect 1890 -618 1896 -612
rect 1890 -624 1896 -618
rect 1890 -630 1896 -624
rect 1890 -636 1896 -630
rect 1890 -642 1896 -636
rect 1890 -648 1896 -642
rect 1890 -654 1896 -648
rect 1890 -660 1896 -654
rect 1890 -666 1896 -660
rect 1890 -672 1896 -666
rect 1890 -678 1896 -672
rect 1890 -684 1896 -678
rect 1890 -690 1896 -684
rect 1890 -696 1896 -690
rect 1890 -702 1896 -696
rect 1890 -708 1896 -702
rect 1890 -714 1896 -708
rect 1890 -720 1896 -714
rect 1890 -726 1896 -720
rect 1890 -732 1896 -726
rect 1890 -738 1896 -732
rect 1890 -744 1896 -738
rect 1890 -750 1896 -744
rect 1890 -756 1896 -750
rect 1890 -762 1896 -756
rect 1890 -768 1896 -762
rect 1890 -774 1896 -768
rect 1890 -780 1896 -774
rect 1890 -786 1896 -780
rect 1890 -792 1896 -786
rect 1890 -798 1896 -792
rect 1890 -804 1896 -798
rect 1890 -810 1896 -804
rect 1890 -816 1896 -810
rect 1890 -822 1896 -816
rect 1890 -828 1896 -822
rect 1890 -834 1896 -828
rect 1890 -840 1896 -834
rect 1890 -846 1896 -840
rect 1890 -852 1896 -846
rect 1890 -858 1896 -852
rect 1890 -864 1896 -858
rect 1890 -870 1896 -864
rect 1890 -876 1896 -870
rect 1890 -882 1896 -876
rect 1890 -888 1896 -882
rect 1890 -894 1896 -888
rect 1890 -900 1896 -894
rect 1890 -906 1896 -900
rect 1890 -912 1896 -906
rect 1890 -918 1896 -912
rect 1890 -924 1896 -918
rect 1890 -930 1896 -924
rect 1890 -936 1896 -930
rect 1890 -942 1896 -936
rect 1890 -948 1896 -942
rect 1890 -954 1896 -948
rect 1890 -960 1896 -954
rect 1890 -966 1896 -960
rect 1890 -972 1896 -966
rect 1890 -978 1896 -972
rect 1890 -984 1896 -978
rect 1890 -990 1896 -984
rect 1890 -996 1896 -990
rect 1890 -1002 1896 -996
rect 1890 -1008 1896 -1002
rect 1890 -1014 1896 -1008
rect 1890 -1020 1896 -1014
rect 1890 -1026 1896 -1020
rect 1890 -1032 1896 -1026
rect 1890 -1038 1896 -1032
rect 1890 -1044 1896 -1038
rect 1890 -1050 1896 -1044
rect 1890 -1056 1896 -1050
rect 1890 -1062 1896 -1056
rect 1890 -1068 1896 -1062
rect 1890 -1074 1896 -1068
rect 1890 -1080 1896 -1074
rect 1890 -1086 1896 -1080
rect 1890 -1092 1896 -1086
rect 1890 -1098 1896 -1092
rect 1890 -1104 1896 -1098
rect 1890 -1110 1896 -1104
rect 1890 -1116 1896 -1110
rect 1890 -1122 1896 -1116
rect 1890 -1128 1896 -1122
rect 1890 -1134 1896 -1128
rect 1890 -1140 1896 -1134
rect 1890 -1146 1896 -1140
rect 1890 -1152 1896 -1146
rect 1890 -1158 1896 -1152
rect 1890 -1164 1896 -1158
rect 1890 -1170 1896 -1164
rect 1890 -1176 1896 -1170
rect 1890 -1182 1896 -1176
rect 1890 -1188 1896 -1182
rect 1890 -1194 1896 -1188
rect 1890 -1200 1896 -1194
rect 1890 -1206 1896 -1200
rect 1890 -1212 1896 -1206
rect 1890 -1218 1896 -1212
rect 1890 -1224 1896 -1218
rect 1890 -1230 1896 -1224
rect 1890 -1236 1896 -1230
rect 1890 -1242 1896 -1236
rect 1890 -1248 1896 -1242
rect 1890 -1254 1896 -1248
rect 1890 -1260 1896 -1254
rect 1890 -1266 1896 -1260
rect 1890 -1272 1896 -1266
rect 1890 -1278 1896 -1272
rect 1890 -1284 1896 -1278
rect 1890 -1290 1896 -1284
rect 1890 -1296 1896 -1290
rect 1890 -1302 1896 -1296
rect 1890 -1308 1896 -1302
rect 1890 -1314 1896 -1308
rect 1890 -1320 1896 -1314
rect 1890 -1326 1896 -1320
rect 1890 -1332 1896 -1326
rect 1890 -1338 1896 -1332
rect 1890 -1344 1896 -1338
rect 1890 -1350 1896 -1344
rect 1890 -1356 1896 -1350
rect 1890 -1362 1896 -1356
rect 1890 -1368 1896 -1362
rect 1890 -1374 1896 -1368
rect 1890 -1380 1896 -1374
rect 1890 -1386 1896 -1380
rect 1890 -1392 1896 -1386
rect 1890 -1398 1896 -1392
rect 1890 -1404 1896 -1398
rect 1890 -1410 1896 -1404
rect 1890 -1416 1896 -1410
rect 1890 -1422 1896 -1416
rect 1890 -1428 1896 -1422
rect 1890 -1434 1896 -1428
rect 1890 -1440 1896 -1434
rect 1890 -1446 1896 -1440
rect 1890 -1452 1896 -1446
rect 1890 -1458 1896 -1452
rect 1890 -1464 1896 -1458
rect 1890 -1470 1896 -1464
rect 1890 -1476 1896 -1470
rect 1890 -1482 1896 -1476
rect 1890 -1488 1896 -1482
rect 1890 -1494 1896 -1488
rect 1890 -1500 1896 -1494
rect 1890 -1506 1896 -1500
rect 1890 -1512 1896 -1506
rect 1890 -1518 1896 -1512
rect 1890 -1524 1896 -1518
rect 1890 -1530 1896 -1524
rect 1890 -1536 1896 -1530
rect 1890 -1542 1896 -1536
rect 1890 -1548 1896 -1542
rect 1890 -1554 1896 -1548
rect 1890 -1560 1896 -1554
rect 1890 -1566 1896 -1560
rect 1890 -1572 1896 -1566
rect 1890 -1578 1896 -1572
rect 1890 -1584 1896 -1578
rect 1890 -1590 1896 -1584
rect 1890 -1596 1896 -1590
rect 1890 -1602 1896 -1596
rect 1890 -1608 1896 -1602
rect 1890 -1614 1896 -1608
rect 1890 -1620 1896 -1614
rect 1890 -1626 1896 -1620
rect 1890 -1632 1896 -1626
rect 1890 -1638 1896 -1632
rect 1890 -1644 1896 -1638
rect 1890 -1650 1896 -1644
rect 1890 -1656 1896 -1650
rect 1890 -1662 1896 -1656
rect 1890 -1668 1896 -1662
rect 1890 -1674 1896 -1668
rect 1890 -1680 1896 -1674
rect 1890 -1686 1896 -1680
rect 1890 -1692 1896 -1686
rect 1890 -1698 1896 -1692
rect 1890 -1704 1896 -1698
rect 1890 -1710 1896 -1704
rect 1890 -1716 1896 -1710
rect 1890 -1722 1896 -1716
rect 1890 -1728 1896 -1722
rect 1890 -1734 1896 -1728
rect 1890 -1740 1896 -1734
rect 1890 -1746 1896 -1740
rect 1890 -1752 1896 -1746
rect 1890 -1758 1896 -1752
rect 1890 -1836 1896 -1830
rect 1890 -1842 1896 -1836
rect 1890 -1848 1896 -1842
rect 1890 -1854 1896 -1848
rect 1890 -1860 1896 -1854
rect 1890 -1866 1896 -1860
rect 1890 -1872 1896 -1866
rect 1890 -1878 1896 -1872
rect 1890 -1884 1896 -1878
rect 1890 -1890 1896 -1884
rect 1890 -1896 1896 -1890
rect 1890 -1902 1896 -1896
rect 1890 -1908 1896 -1902
rect 1890 -1914 1896 -1908
rect 1890 -1920 1896 -1914
rect 1890 -1926 1896 -1920
rect 1890 -1932 1896 -1926
rect 1890 -1938 1896 -1932
rect 1890 -1944 1896 -1938
rect 1890 -1950 1896 -1944
rect 1890 -1956 1896 -1950
rect 1890 -1962 1896 -1956
rect 1890 -1968 1896 -1962
rect 1890 -1974 1896 -1968
rect 1890 -1980 1896 -1974
rect 1890 -1986 1896 -1980
rect 1890 -1992 1896 -1986
rect 1890 -1998 1896 -1992
rect 1890 -2004 1896 -1998
rect 1890 -2010 1896 -2004
rect 1890 -2016 1896 -2010
rect 1890 -2022 1896 -2016
rect 1890 -2028 1896 -2022
rect 1890 -2034 1896 -2028
rect 1890 -2040 1896 -2034
rect 1890 -2046 1896 -2040
rect 1890 -2052 1896 -2046
rect 1890 -2058 1896 -2052
rect 1890 -2064 1896 -2058
rect 1890 -2070 1896 -2064
rect 1890 -2076 1896 -2070
rect 1890 -2082 1896 -2076
rect 1890 -2088 1896 -2082
rect 1890 -2094 1896 -2088
rect 1890 -2100 1896 -2094
rect 1890 -2106 1896 -2100
rect 1890 -2112 1896 -2106
rect 1890 -2118 1896 -2112
rect 1890 -2124 1896 -2118
rect 1890 -2130 1896 -2124
rect 1890 -2136 1896 -2130
rect 1890 -2142 1896 -2136
rect 1890 -2148 1896 -2142
rect 1890 -2154 1896 -2148
rect 1890 -2160 1896 -2154
rect 1890 -2166 1896 -2160
rect 1890 -2172 1896 -2166
rect 1890 -2178 1896 -2172
rect 1890 -2184 1896 -2178
rect 1890 -2190 1896 -2184
rect 1890 -2196 1896 -2190
rect 1890 -2202 1896 -2196
rect 1890 -2208 1896 -2202
rect 1890 -2214 1896 -2208
rect 1890 -2220 1896 -2214
rect 1890 -2226 1896 -2220
rect 1890 -2232 1896 -2226
rect 1890 -2238 1896 -2232
rect 1890 -2244 1896 -2238
rect 1890 -2250 1896 -2244
rect 1890 -2256 1896 -2250
rect 1890 -2262 1896 -2256
rect 1890 -2268 1896 -2262
rect 1890 -2274 1896 -2268
rect 1890 -2280 1896 -2274
rect 1890 -2286 1896 -2280
rect 1890 -2292 1896 -2286
rect 1890 -2298 1896 -2292
rect 1890 -2304 1896 -2298
rect 1890 -2310 1896 -2304
rect 1890 -2316 1896 -2310
rect 1890 -2322 1896 -2316
rect 1890 -2328 1896 -2322
rect 1890 -2334 1896 -2328
rect 1890 -2340 1896 -2334
rect 1890 -2346 1896 -2340
rect 1890 -2352 1896 -2346
rect 1890 -2358 1896 -2352
rect 1890 -2364 1896 -2358
rect 1890 -2370 1896 -2364
rect 1890 -2376 1896 -2370
rect 1890 -2382 1896 -2376
rect 1890 -2388 1896 -2382
rect 1890 -2394 1896 -2388
rect 1890 -2400 1896 -2394
rect 1890 -2406 1896 -2400
rect 1890 -2412 1896 -2406
rect 1890 -2418 1896 -2412
rect 1890 -2424 1896 -2418
rect 1890 -2430 1896 -2424
rect 1890 -2436 1896 -2430
rect 1890 -2442 1896 -2436
rect 1890 -2448 1896 -2442
rect 1890 -2454 1896 -2448
rect 1890 -2460 1896 -2454
rect 1890 -2466 1896 -2460
rect 1890 -2472 1896 -2466
rect 1890 -2478 1896 -2472
rect 1890 -2484 1896 -2478
rect 1890 -2490 1896 -2484
rect 1890 -2496 1896 -2490
rect 1890 -2502 1896 -2496
rect 1890 -2508 1896 -2502
rect 1890 -2514 1896 -2508
rect 1890 -2520 1896 -2514
rect 1890 -2526 1896 -2520
rect 1890 -2532 1896 -2526
rect 1890 -2538 1896 -2532
rect 1890 -2544 1896 -2538
rect 1890 -2550 1896 -2544
rect 1890 -2556 1896 -2550
rect 1890 -2562 1896 -2556
rect 1890 -2568 1896 -2562
rect 1890 -2574 1896 -2568
rect 1890 -2580 1896 -2574
rect 1890 -2586 1896 -2580
rect 1890 -2658 1896 -2652
rect 1890 -2664 1896 -2658
rect 1890 -2670 1896 -2664
rect 1890 -2676 1896 -2670
rect 1890 -2682 1896 -2676
rect 1890 -2688 1896 -2682
rect 1890 -2694 1896 -2688
rect 1890 -2700 1896 -2694
rect 1890 -2706 1896 -2700
rect 1890 -2712 1896 -2706
rect 1890 -2718 1896 -2712
rect 1890 -2724 1896 -2718
rect 1890 -2730 1896 -2724
rect 1890 -2736 1896 -2730
rect 1890 -2742 1896 -2736
rect 1890 -2748 1896 -2742
rect 1890 -2754 1896 -2748
rect 1890 -2760 1896 -2754
rect 1890 -2766 1896 -2760
rect 1890 -2772 1896 -2766
rect 1890 -2778 1896 -2772
rect 1890 -2784 1896 -2778
rect 1890 -2790 1896 -2784
rect 1890 -2796 1896 -2790
rect 1890 -2802 1896 -2796
rect 1890 -2808 1896 -2802
rect 1890 -2814 1896 -2808
rect 1890 -2820 1896 -2814
rect 1890 -2826 1896 -2820
rect 1890 -2832 1896 -2826
rect 1890 -2838 1896 -2832
rect 1890 -2844 1896 -2838
rect 1890 -2850 1896 -2844
rect 1890 -2856 1896 -2850
rect 1890 -2862 1896 -2856
rect 1890 -2868 1896 -2862
rect 1890 -2874 1896 -2868
rect 1890 -2880 1896 -2874
rect 1890 -2886 1896 -2880
rect 1890 -2892 1896 -2886
rect 1890 -2898 1896 -2892
rect 1890 -2904 1896 -2898
rect 1890 -2910 1896 -2904
rect 1890 -2916 1896 -2910
rect 1890 -2922 1896 -2916
rect 1890 -2928 1896 -2922
rect 1890 -2934 1896 -2928
rect 1890 -2940 1896 -2934
rect 1890 -2946 1896 -2940
rect 1890 -2952 1896 -2946
rect 1890 -2958 1896 -2952
rect 1890 -2964 1896 -2958
rect 1890 -2970 1896 -2964
rect 1890 -2976 1896 -2970
rect 1890 -2982 1896 -2976
rect 1890 -2988 1896 -2982
rect 1890 -2994 1896 -2988
rect 1890 -3000 1896 -2994
rect 1890 -3006 1896 -3000
rect 1890 -3012 1896 -3006
rect 1890 -3018 1896 -3012
rect 1890 -3024 1896 -3018
rect 1890 -3030 1896 -3024
rect 1890 -3036 1896 -3030
rect 1890 -3042 1896 -3036
rect 1890 -3048 1896 -3042
rect 1890 -3054 1896 -3048
rect 1890 -3060 1896 -3054
rect 1890 -3066 1896 -3060
rect 1890 -3072 1896 -3066
rect 1890 -3078 1896 -3072
rect 1890 -3084 1896 -3078
rect 1890 -3090 1896 -3084
rect 1890 -3096 1896 -3090
rect 1890 -3102 1896 -3096
rect 1890 -3108 1896 -3102
rect 1890 -3114 1896 -3108
rect 1890 -3120 1896 -3114
rect 1890 -3126 1896 -3120
rect 1890 -3132 1896 -3126
rect 1890 -3138 1896 -3132
rect 1890 -3144 1896 -3138
rect 1890 -3150 1896 -3144
rect 1890 -3198 1896 -3192
rect 1890 -3204 1896 -3198
rect 1890 -3210 1896 -3204
rect 1890 -3216 1896 -3210
rect 1890 -3222 1896 -3216
rect 1890 -3228 1896 -3222
rect 1890 -3234 1896 -3228
rect 1890 -3240 1896 -3234
rect 1890 -3246 1896 -3240
rect 1890 -3252 1896 -3246
rect 1890 -3258 1896 -3252
rect 1890 -3264 1896 -3258
rect 1890 -3270 1896 -3264
rect 1890 -3276 1896 -3270
rect 1890 -3282 1896 -3276
rect 1890 -3288 1896 -3282
rect 1890 -3294 1896 -3288
rect 1890 -3300 1896 -3294
rect 1890 -3306 1896 -3300
rect 1890 -3312 1896 -3306
rect 1896 -588 1902 -582
rect 1896 -594 1902 -588
rect 1896 -600 1902 -594
rect 1896 -606 1902 -600
rect 1896 -612 1902 -606
rect 1896 -618 1902 -612
rect 1896 -624 1902 -618
rect 1896 -630 1902 -624
rect 1896 -636 1902 -630
rect 1896 -642 1902 -636
rect 1896 -648 1902 -642
rect 1896 -654 1902 -648
rect 1896 -660 1902 -654
rect 1896 -666 1902 -660
rect 1896 -672 1902 -666
rect 1896 -678 1902 -672
rect 1896 -684 1902 -678
rect 1896 -690 1902 -684
rect 1896 -696 1902 -690
rect 1896 -702 1902 -696
rect 1896 -708 1902 -702
rect 1896 -714 1902 -708
rect 1896 -720 1902 -714
rect 1896 -726 1902 -720
rect 1896 -732 1902 -726
rect 1896 -738 1902 -732
rect 1896 -744 1902 -738
rect 1896 -750 1902 -744
rect 1896 -756 1902 -750
rect 1896 -762 1902 -756
rect 1896 -768 1902 -762
rect 1896 -774 1902 -768
rect 1896 -780 1902 -774
rect 1896 -786 1902 -780
rect 1896 -792 1902 -786
rect 1896 -798 1902 -792
rect 1896 -804 1902 -798
rect 1896 -810 1902 -804
rect 1896 -816 1902 -810
rect 1896 -822 1902 -816
rect 1896 -828 1902 -822
rect 1896 -834 1902 -828
rect 1896 -840 1902 -834
rect 1896 -846 1902 -840
rect 1896 -852 1902 -846
rect 1896 -858 1902 -852
rect 1896 -864 1902 -858
rect 1896 -870 1902 -864
rect 1896 -876 1902 -870
rect 1896 -882 1902 -876
rect 1896 -888 1902 -882
rect 1896 -894 1902 -888
rect 1896 -900 1902 -894
rect 1896 -906 1902 -900
rect 1896 -912 1902 -906
rect 1896 -918 1902 -912
rect 1896 -924 1902 -918
rect 1896 -930 1902 -924
rect 1896 -936 1902 -930
rect 1896 -942 1902 -936
rect 1896 -948 1902 -942
rect 1896 -954 1902 -948
rect 1896 -960 1902 -954
rect 1896 -966 1902 -960
rect 1896 -972 1902 -966
rect 1896 -978 1902 -972
rect 1896 -984 1902 -978
rect 1896 -990 1902 -984
rect 1896 -996 1902 -990
rect 1896 -1002 1902 -996
rect 1896 -1008 1902 -1002
rect 1896 -1014 1902 -1008
rect 1896 -1020 1902 -1014
rect 1896 -1026 1902 -1020
rect 1896 -1032 1902 -1026
rect 1896 -1038 1902 -1032
rect 1896 -1044 1902 -1038
rect 1896 -1050 1902 -1044
rect 1896 -1056 1902 -1050
rect 1896 -1062 1902 -1056
rect 1896 -1068 1902 -1062
rect 1896 -1074 1902 -1068
rect 1896 -1080 1902 -1074
rect 1896 -1086 1902 -1080
rect 1896 -1092 1902 -1086
rect 1896 -1098 1902 -1092
rect 1896 -1104 1902 -1098
rect 1896 -1110 1902 -1104
rect 1896 -1116 1902 -1110
rect 1896 -1122 1902 -1116
rect 1896 -1128 1902 -1122
rect 1896 -1134 1902 -1128
rect 1896 -1140 1902 -1134
rect 1896 -1146 1902 -1140
rect 1896 -1152 1902 -1146
rect 1896 -1158 1902 -1152
rect 1896 -1164 1902 -1158
rect 1896 -1170 1902 -1164
rect 1896 -1176 1902 -1170
rect 1896 -1182 1902 -1176
rect 1896 -1188 1902 -1182
rect 1896 -1194 1902 -1188
rect 1896 -1200 1902 -1194
rect 1896 -1206 1902 -1200
rect 1896 -1212 1902 -1206
rect 1896 -1218 1902 -1212
rect 1896 -1224 1902 -1218
rect 1896 -1230 1902 -1224
rect 1896 -1236 1902 -1230
rect 1896 -1242 1902 -1236
rect 1896 -1248 1902 -1242
rect 1896 -1254 1902 -1248
rect 1896 -1260 1902 -1254
rect 1896 -1266 1902 -1260
rect 1896 -1272 1902 -1266
rect 1896 -1278 1902 -1272
rect 1896 -1284 1902 -1278
rect 1896 -1290 1902 -1284
rect 1896 -1296 1902 -1290
rect 1896 -1302 1902 -1296
rect 1896 -1308 1902 -1302
rect 1896 -1314 1902 -1308
rect 1896 -1320 1902 -1314
rect 1896 -1326 1902 -1320
rect 1896 -1332 1902 -1326
rect 1896 -1338 1902 -1332
rect 1896 -1344 1902 -1338
rect 1896 -1350 1902 -1344
rect 1896 -1356 1902 -1350
rect 1896 -1362 1902 -1356
rect 1896 -1368 1902 -1362
rect 1896 -1374 1902 -1368
rect 1896 -1380 1902 -1374
rect 1896 -1386 1902 -1380
rect 1896 -1392 1902 -1386
rect 1896 -1398 1902 -1392
rect 1896 -1404 1902 -1398
rect 1896 -1410 1902 -1404
rect 1896 -1416 1902 -1410
rect 1896 -1422 1902 -1416
rect 1896 -1428 1902 -1422
rect 1896 -1434 1902 -1428
rect 1896 -1440 1902 -1434
rect 1896 -1446 1902 -1440
rect 1896 -1452 1902 -1446
rect 1896 -1458 1902 -1452
rect 1896 -1464 1902 -1458
rect 1896 -1470 1902 -1464
rect 1896 -1476 1902 -1470
rect 1896 -1482 1902 -1476
rect 1896 -1488 1902 -1482
rect 1896 -1494 1902 -1488
rect 1896 -1500 1902 -1494
rect 1896 -1506 1902 -1500
rect 1896 -1512 1902 -1506
rect 1896 -1518 1902 -1512
rect 1896 -1524 1902 -1518
rect 1896 -1530 1902 -1524
rect 1896 -1536 1902 -1530
rect 1896 -1542 1902 -1536
rect 1896 -1548 1902 -1542
rect 1896 -1554 1902 -1548
rect 1896 -1560 1902 -1554
rect 1896 -1566 1902 -1560
rect 1896 -1572 1902 -1566
rect 1896 -1578 1902 -1572
rect 1896 -1584 1902 -1578
rect 1896 -1590 1902 -1584
rect 1896 -1596 1902 -1590
rect 1896 -1602 1902 -1596
rect 1896 -1608 1902 -1602
rect 1896 -1614 1902 -1608
rect 1896 -1620 1902 -1614
rect 1896 -1626 1902 -1620
rect 1896 -1632 1902 -1626
rect 1896 -1638 1902 -1632
rect 1896 -1644 1902 -1638
rect 1896 -1650 1902 -1644
rect 1896 -1656 1902 -1650
rect 1896 -1662 1902 -1656
rect 1896 -1668 1902 -1662
rect 1896 -1674 1902 -1668
rect 1896 -1680 1902 -1674
rect 1896 -1686 1902 -1680
rect 1896 -1692 1902 -1686
rect 1896 -1698 1902 -1692
rect 1896 -1704 1902 -1698
rect 1896 -1710 1902 -1704
rect 1896 -1716 1902 -1710
rect 1896 -1722 1902 -1716
rect 1896 -1728 1902 -1722
rect 1896 -1734 1902 -1728
rect 1896 -1740 1902 -1734
rect 1896 -1746 1902 -1740
rect 1896 -1752 1902 -1746
rect 1896 -1830 1902 -1824
rect 1896 -1836 1902 -1830
rect 1896 -1842 1902 -1836
rect 1896 -1848 1902 -1842
rect 1896 -1854 1902 -1848
rect 1896 -1860 1902 -1854
rect 1896 -1866 1902 -1860
rect 1896 -1872 1902 -1866
rect 1896 -1878 1902 -1872
rect 1896 -1884 1902 -1878
rect 1896 -1890 1902 -1884
rect 1896 -1896 1902 -1890
rect 1896 -1902 1902 -1896
rect 1896 -1908 1902 -1902
rect 1896 -1914 1902 -1908
rect 1896 -1920 1902 -1914
rect 1896 -1926 1902 -1920
rect 1896 -1932 1902 -1926
rect 1896 -1938 1902 -1932
rect 1896 -1944 1902 -1938
rect 1896 -1950 1902 -1944
rect 1896 -1956 1902 -1950
rect 1896 -1962 1902 -1956
rect 1896 -1968 1902 -1962
rect 1896 -1974 1902 -1968
rect 1896 -1980 1902 -1974
rect 1896 -1986 1902 -1980
rect 1896 -1992 1902 -1986
rect 1896 -1998 1902 -1992
rect 1896 -2004 1902 -1998
rect 1896 -2010 1902 -2004
rect 1896 -2016 1902 -2010
rect 1896 -2022 1902 -2016
rect 1896 -2028 1902 -2022
rect 1896 -2034 1902 -2028
rect 1896 -2040 1902 -2034
rect 1896 -2046 1902 -2040
rect 1896 -2052 1902 -2046
rect 1896 -2058 1902 -2052
rect 1896 -2064 1902 -2058
rect 1896 -2070 1902 -2064
rect 1896 -2076 1902 -2070
rect 1896 -2082 1902 -2076
rect 1896 -2088 1902 -2082
rect 1896 -2094 1902 -2088
rect 1896 -2100 1902 -2094
rect 1896 -2106 1902 -2100
rect 1896 -2112 1902 -2106
rect 1896 -2118 1902 -2112
rect 1896 -2124 1902 -2118
rect 1896 -2130 1902 -2124
rect 1896 -2136 1902 -2130
rect 1896 -2142 1902 -2136
rect 1896 -2148 1902 -2142
rect 1896 -2154 1902 -2148
rect 1896 -2160 1902 -2154
rect 1896 -2166 1902 -2160
rect 1896 -2172 1902 -2166
rect 1896 -2178 1902 -2172
rect 1896 -2184 1902 -2178
rect 1896 -2190 1902 -2184
rect 1896 -2196 1902 -2190
rect 1896 -2202 1902 -2196
rect 1896 -2208 1902 -2202
rect 1896 -2214 1902 -2208
rect 1896 -2220 1902 -2214
rect 1896 -2226 1902 -2220
rect 1896 -2232 1902 -2226
rect 1896 -2238 1902 -2232
rect 1896 -2244 1902 -2238
rect 1896 -2250 1902 -2244
rect 1896 -2256 1902 -2250
rect 1896 -2262 1902 -2256
rect 1896 -2268 1902 -2262
rect 1896 -2274 1902 -2268
rect 1896 -2280 1902 -2274
rect 1896 -2286 1902 -2280
rect 1896 -2292 1902 -2286
rect 1896 -2298 1902 -2292
rect 1896 -2304 1902 -2298
rect 1896 -2310 1902 -2304
rect 1896 -2316 1902 -2310
rect 1896 -2322 1902 -2316
rect 1896 -2328 1902 -2322
rect 1896 -2334 1902 -2328
rect 1896 -2340 1902 -2334
rect 1896 -2346 1902 -2340
rect 1896 -2352 1902 -2346
rect 1896 -2358 1902 -2352
rect 1896 -2364 1902 -2358
rect 1896 -2370 1902 -2364
rect 1896 -2376 1902 -2370
rect 1896 -2382 1902 -2376
rect 1896 -2388 1902 -2382
rect 1896 -2394 1902 -2388
rect 1896 -2400 1902 -2394
rect 1896 -2406 1902 -2400
rect 1896 -2412 1902 -2406
rect 1896 -2418 1902 -2412
rect 1896 -2424 1902 -2418
rect 1896 -2430 1902 -2424
rect 1896 -2436 1902 -2430
rect 1896 -2442 1902 -2436
rect 1896 -2448 1902 -2442
rect 1896 -2454 1902 -2448
rect 1896 -2460 1902 -2454
rect 1896 -2466 1902 -2460
rect 1896 -2472 1902 -2466
rect 1896 -2478 1902 -2472
rect 1896 -2484 1902 -2478
rect 1896 -2490 1902 -2484
rect 1896 -2496 1902 -2490
rect 1896 -2502 1902 -2496
rect 1896 -2508 1902 -2502
rect 1896 -2514 1902 -2508
rect 1896 -2520 1902 -2514
rect 1896 -2526 1902 -2520
rect 1896 -2532 1902 -2526
rect 1896 -2538 1902 -2532
rect 1896 -2544 1902 -2538
rect 1896 -2550 1902 -2544
rect 1896 -2556 1902 -2550
rect 1896 -2562 1902 -2556
rect 1896 -2568 1902 -2562
rect 1896 -2574 1902 -2568
rect 1896 -2580 1902 -2574
rect 1896 -2658 1902 -2652
rect 1896 -2664 1902 -2658
rect 1896 -2670 1902 -2664
rect 1896 -2676 1902 -2670
rect 1896 -2682 1902 -2676
rect 1896 -2688 1902 -2682
rect 1896 -2694 1902 -2688
rect 1896 -2700 1902 -2694
rect 1896 -2706 1902 -2700
rect 1896 -2712 1902 -2706
rect 1896 -2718 1902 -2712
rect 1896 -2724 1902 -2718
rect 1896 -2730 1902 -2724
rect 1896 -2736 1902 -2730
rect 1896 -2742 1902 -2736
rect 1896 -2748 1902 -2742
rect 1896 -2754 1902 -2748
rect 1896 -2760 1902 -2754
rect 1896 -2766 1902 -2760
rect 1896 -2772 1902 -2766
rect 1896 -2778 1902 -2772
rect 1896 -2784 1902 -2778
rect 1896 -2790 1902 -2784
rect 1896 -2796 1902 -2790
rect 1896 -2802 1902 -2796
rect 1896 -2808 1902 -2802
rect 1896 -2814 1902 -2808
rect 1896 -2820 1902 -2814
rect 1896 -2826 1902 -2820
rect 1896 -2832 1902 -2826
rect 1896 -2838 1902 -2832
rect 1896 -2844 1902 -2838
rect 1896 -2850 1902 -2844
rect 1896 -2856 1902 -2850
rect 1896 -2862 1902 -2856
rect 1896 -2868 1902 -2862
rect 1896 -2874 1902 -2868
rect 1896 -2880 1902 -2874
rect 1896 -2886 1902 -2880
rect 1896 -2892 1902 -2886
rect 1896 -2898 1902 -2892
rect 1896 -2904 1902 -2898
rect 1896 -2910 1902 -2904
rect 1896 -2916 1902 -2910
rect 1896 -2922 1902 -2916
rect 1896 -2928 1902 -2922
rect 1896 -2934 1902 -2928
rect 1896 -2940 1902 -2934
rect 1896 -2946 1902 -2940
rect 1896 -2952 1902 -2946
rect 1896 -2958 1902 -2952
rect 1896 -2964 1902 -2958
rect 1896 -2970 1902 -2964
rect 1896 -2976 1902 -2970
rect 1896 -2982 1902 -2976
rect 1896 -2988 1902 -2982
rect 1896 -2994 1902 -2988
rect 1896 -3000 1902 -2994
rect 1896 -3006 1902 -3000
rect 1896 -3012 1902 -3006
rect 1896 -3018 1902 -3012
rect 1896 -3024 1902 -3018
rect 1896 -3030 1902 -3024
rect 1896 -3036 1902 -3030
rect 1896 -3042 1902 -3036
rect 1896 -3048 1902 -3042
rect 1896 -3054 1902 -3048
rect 1896 -3060 1902 -3054
rect 1896 -3066 1902 -3060
rect 1896 -3072 1902 -3066
rect 1896 -3078 1902 -3072
rect 1896 -3084 1902 -3078
rect 1896 -3090 1902 -3084
rect 1896 -3096 1902 -3090
rect 1896 -3102 1902 -3096
rect 1896 -3108 1902 -3102
rect 1896 -3114 1902 -3108
rect 1896 -3120 1902 -3114
rect 1896 -3126 1902 -3120
rect 1896 -3132 1902 -3126
rect 1896 -3138 1902 -3132
rect 1896 -3144 1902 -3138
rect 1896 -3198 1902 -3192
rect 1896 -3204 1902 -3198
rect 1896 -3210 1902 -3204
rect 1896 -3216 1902 -3210
rect 1896 -3222 1902 -3216
rect 1896 -3228 1902 -3222
rect 1896 -3234 1902 -3228
rect 1896 -3240 1902 -3234
rect 1896 -3246 1902 -3240
rect 1896 -3252 1902 -3246
rect 1896 -3258 1902 -3252
rect 1896 -3264 1902 -3258
rect 1896 -3270 1902 -3264
rect 1896 -3276 1902 -3270
rect 1896 -3282 1902 -3276
rect 1896 -3288 1902 -3282
rect 1896 -3294 1902 -3288
rect 1896 -3300 1902 -3294
rect 1896 -3306 1902 -3300
rect 1902 -582 1908 -576
rect 1902 -588 1908 -582
rect 1902 -594 1908 -588
rect 1902 -600 1908 -594
rect 1902 -606 1908 -600
rect 1902 -612 1908 -606
rect 1902 -618 1908 -612
rect 1902 -624 1908 -618
rect 1902 -630 1908 -624
rect 1902 -636 1908 -630
rect 1902 -642 1908 -636
rect 1902 -648 1908 -642
rect 1902 -654 1908 -648
rect 1902 -660 1908 -654
rect 1902 -666 1908 -660
rect 1902 -672 1908 -666
rect 1902 -678 1908 -672
rect 1902 -684 1908 -678
rect 1902 -690 1908 -684
rect 1902 -696 1908 -690
rect 1902 -702 1908 -696
rect 1902 -708 1908 -702
rect 1902 -714 1908 -708
rect 1902 -720 1908 -714
rect 1902 -726 1908 -720
rect 1902 -732 1908 -726
rect 1902 -738 1908 -732
rect 1902 -744 1908 -738
rect 1902 -750 1908 -744
rect 1902 -756 1908 -750
rect 1902 -762 1908 -756
rect 1902 -768 1908 -762
rect 1902 -774 1908 -768
rect 1902 -780 1908 -774
rect 1902 -786 1908 -780
rect 1902 -792 1908 -786
rect 1902 -798 1908 -792
rect 1902 -804 1908 -798
rect 1902 -810 1908 -804
rect 1902 -816 1908 -810
rect 1902 -822 1908 -816
rect 1902 -828 1908 -822
rect 1902 -834 1908 -828
rect 1902 -840 1908 -834
rect 1902 -846 1908 -840
rect 1902 -852 1908 -846
rect 1902 -858 1908 -852
rect 1902 -864 1908 -858
rect 1902 -870 1908 -864
rect 1902 -876 1908 -870
rect 1902 -882 1908 -876
rect 1902 -888 1908 -882
rect 1902 -894 1908 -888
rect 1902 -900 1908 -894
rect 1902 -906 1908 -900
rect 1902 -912 1908 -906
rect 1902 -918 1908 -912
rect 1902 -924 1908 -918
rect 1902 -930 1908 -924
rect 1902 -936 1908 -930
rect 1902 -942 1908 -936
rect 1902 -948 1908 -942
rect 1902 -954 1908 -948
rect 1902 -960 1908 -954
rect 1902 -966 1908 -960
rect 1902 -972 1908 -966
rect 1902 -978 1908 -972
rect 1902 -984 1908 -978
rect 1902 -990 1908 -984
rect 1902 -996 1908 -990
rect 1902 -1002 1908 -996
rect 1902 -1008 1908 -1002
rect 1902 -1014 1908 -1008
rect 1902 -1020 1908 -1014
rect 1902 -1026 1908 -1020
rect 1902 -1032 1908 -1026
rect 1902 -1038 1908 -1032
rect 1902 -1044 1908 -1038
rect 1902 -1050 1908 -1044
rect 1902 -1056 1908 -1050
rect 1902 -1062 1908 -1056
rect 1902 -1068 1908 -1062
rect 1902 -1074 1908 -1068
rect 1902 -1080 1908 -1074
rect 1902 -1086 1908 -1080
rect 1902 -1092 1908 -1086
rect 1902 -1098 1908 -1092
rect 1902 -1104 1908 -1098
rect 1902 -1110 1908 -1104
rect 1902 -1116 1908 -1110
rect 1902 -1122 1908 -1116
rect 1902 -1128 1908 -1122
rect 1902 -1134 1908 -1128
rect 1902 -1140 1908 -1134
rect 1902 -1146 1908 -1140
rect 1902 -1152 1908 -1146
rect 1902 -1158 1908 -1152
rect 1902 -1164 1908 -1158
rect 1902 -1170 1908 -1164
rect 1902 -1176 1908 -1170
rect 1902 -1182 1908 -1176
rect 1902 -1188 1908 -1182
rect 1902 -1194 1908 -1188
rect 1902 -1200 1908 -1194
rect 1902 -1206 1908 -1200
rect 1902 -1212 1908 -1206
rect 1902 -1218 1908 -1212
rect 1902 -1224 1908 -1218
rect 1902 -1230 1908 -1224
rect 1902 -1236 1908 -1230
rect 1902 -1242 1908 -1236
rect 1902 -1248 1908 -1242
rect 1902 -1254 1908 -1248
rect 1902 -1260 1908 -1254
rect 1902 -1266 1908 -1260
rect 1902 -1272 1908 -1266
rect 1902 -1278 1908 -1272
rect 1902 -1284 1908 -1278
rect 1902 -1290 1908 -1284
rect 1902 -1296 1908 -1290
rect 1902 -1302 1908 -1296
rect 1902 -1308 1908 -1302
rect 1902 -1314 1908 -1308
rect 1902 -1320 1908 -1314
rect 1902 -1326 1908 -1320
rect 1902 -1332 1908 -1326
rect 1902 -1338 1908 -1332
rect 1902 -1344 1908 -1338
rect 1902 -1350 1908 -1344
rect 1902 -1356 1908 -1350
rect 1902 -1362 1908 -1356
rect 1902 -1368 1908 -1362
rect 1902 -1374 1908 -1368
rect 1902 -1380 1908 -1374
rect 1902 -1386 1908 -1380
rect 1902 -1392 1908 -1386
rect 1902 -1398 1908 -1392
rect 1902 -1404 1908 -1398
rect 1902 -1410 1908 -1404
rect 1902 -1416 1908 -1410
rect 1902 -1422 1908 -1416
rect 1902 -1428 1908 -1422
rect 1902 -1434 1908 -1428
rect 1902 -1440 1908 -1434
rect 1902 -1446 1908 -1440
rect 1902 -1452 1908 -1446
rect 1902 -1458 1908 -1452
rect 1902 -1464 1908 -1458
rect 1902 -1470 1908 -1464
rect 1902 -1476 1908 -1470
rect 1902 -1482 1908 -1476
rect 1902 -1488 1908 -1482
rect 1902 -1494 1908 -1488
rect 1902 -1500 1908 -1494
rect 1902 -1506 1908 -1500
rect 1902 -1512 1908 -1506
rect 1902 -1518 1908 -1512
rect 1902 -1524 1908 -1518
rect 1902 -1530 1908 -1524
rect 1902 -1536 1908 -1530
rect 1902 -1542 1908 -1536
rect 1902 -1548 1908 -1542
rect 1902 -1554 1908 -1548
rect 1902 -1560 1908 -1554
rect 1902 -1566 1908 -1560
rect 1902 -1572 1908 -1566
rect 1902 -1578 1908 -1572
rect 1902 -1584 1908 -1578
rect 1902 -1590 1908 -1584
rect 1902 -1596 1908 -1590
rect 1902 -1602 1908 -1596
rect 1902 -1608 1908 -1602
rect 1902 -1614 1908 -1608
rect 1902 -1620 1908 -1614
rect 1902 -1626 1908 -1620
rect 1902 -1632 1908 -1626
rect 1902 -1638 1908 -1632
rect 1902 -1644 1908 -1638
rect 1902 -1650 1908 -1644
rect 1902 -1656 1908 -1650
rect 1902 -1662 1908 -1656
rect 1902 -1668 1908 -1662
rect 1902 -1674 1908 -1668
rect 1902 -1680 1908 -1674
rect 1902 -1686 1908 -1680
rect 1902 -1692 1908 -1686
rect 1902 -1698 1908 -1692
rect 1902 -1704 1908 -1698
rect 1902 -1710 1908 -1704
rect 1902 -1716 1908 -1710
rect 1902 -1722 1908 -1716
rect 1902 -1728 1908 -1722
rect 1902 -1734 1908 -1728
rect 1902 -1740 1908 -1734
rect 1902 -1746 1908 -1740
rect 1902 -1824 1908 -1818
rect 1902 -1830 1908 -1824
rect 1902 -1836 1908 -1830
rect 1902 -1842 1908 -1836
rect 1902 -1848 1908 -1842
rect 1902 -1854 1908 -1848
rect 1902 -1860 1908 -1854
rect 1902 -1866 1908 -1860
rect 1902 -1872 1908 -1866
rect 1902 -1878 1908 -1872
rect 1902 -1884 1908 -1878
rect 1902 -1890 1908 -1884
rect 1902 -1896 1908 -1890
rect 1902 -1902 1908 -1896
rect 1902 -1908 1908 -1902
rect 1902 -1914 1908 -1908
rect 1902 -1920 1908 -1914
rect 1902 -1926 1908 -1920
rect 1902 -1932 1908 -1926
rect 1902 -1938 1908 -1932
rect 1902 -1944 1908 -1938
rect 1902 -1950 1908 -1944
rect 1902 -1956 1908 -1950
rect 1902 -1962 1908 -1956
rect 1902 -1968 1908 -1962
rect 1902 -1974 1908 -1968
rect 1902 -1980 1908 -1974
rect 1902 -1986 1908 -1980
rect 1902 -1992 1908 -1986
rect 1902 -1998 1908 -1992
rect 1902 -2004 1908 -1998
rect 1902 -2010 1908 -2004
rect 1902 -2016 1908 -2010
rect 1902 -2022 1908 -2016
rect 1902 -2028 1908 -2022
rect 1902 -2034 1908 -2028
rect 1902 -2040 1908 -2034
rect 1902 -2046 1908 -2040
rect 1902 -2052 1908 -2046
rect 1902 -2058 1908 -2052
rect 1902 -2064 1908 -2058
rect 1902 -2070 1908 -2064
rect 1902 -2076 1908 -2070
rect 1902 -2082 1908 -2076
rect 1902 -2088 1908 -2082
rect 1902 -2094 1908 -2088
rect 1902 -2100 1908 -2094
rect 1902 -2106 1908 -2100
rect 1902 -2112 1908 -2106
rect 1902 -2118 1908 -2112
rect 1902 -2124 1908 -2118
rect 1902 -2130 1908 -2124
rect 1902 -2136 1908 -2130
rect 1902 -2142 1908 -2136
rect 1902 -2148 1908 -2142
rect 1902 -2154 1908 -2148
rect 1902 -2160 1908 -2154
rect 1902 -2166 1908 -2160
rect 1902 -2172 1908 -2166
rect 1902 -2178 1908 -2172
rect 1902 -2184 1908 -2178
rect 1902 -2190 1908 -2184
rect 1902 -2196 1908 -2190
rect 1902 -2202 1908 -2196
rect 1902 -2208 1908 -2202
rect 1902 -2214 1908 -2208
rect 1902 -2220 1908 -2214
rect 1902 -2226 1908 -2220
rect 1902 -2232 1908 -2226
rect 1902 -2238 1908 -2232
rect 1902 -2244 1908 -2238
rect 1902 -2250 1908 -2244
rect 1902 -2256 1908 -2250
rect 1902 -2262 1908 -2256
rect 1902 -2268 1908 -2262
rect 1902 -2274 1908 -2268
rect 1902 -2280 1908 -2274
rect 1902 -2286 1908 -2280
rect 1902 -2292 1908 -2286
rect 1902 -2298 1908 -2292
rect 1902 -2304 1908 -2298
rect 1902 -2310 1908 -2304
rect 1902 -2316 1908 -2310
rect 1902 -2322 1908 -2316
rect 1902 -2328 1908 -2322
rect 1902 -2334 1908 -2328
rect 1902 -2340 1908 -2334
rect 1902 -2346 1908 -2340
rect 1902 -2352 1908 -2346
rect 1902 -2358 1908 -2352
rect 1902 -2364 1908 -2358
rect 1902 -2370 1908 -2364
rect 1902 -2376 1908 -2370
rect 1902 -2382 1908 -2376
rect 1902 -2388 1908 -2382
rect 1902 -2394 1908 -2388
rect 1902 -2400 1908 -2394
rect 1902 -2406 1908 -2400
rect 1902 -2412 1908 -2406
rect 1902 -2418 1908 -2412
rect 1902 -2424 1908 -2418
rect 1902 -2430 1908 -2424
rect 1902 -2436 1908 -2430
rect 1902 -2442 1908 -2436
rect 1902 -2448 1908 -2442
rect 1902 -2454 1908 -2448
rect 1902 -2460 1908 -2454
rect 1902 -2466 1908 -2460
rect 1902 -2472 1908 -2466
rect 1902 -2478 1908 -2472
rect 1902 -2484 1908 -2478
rect 1902 -2490 1908 -2484
rect 1902 -2496 1908 -2490
rect 1902 -2502 1908 -2496
rect 1902 -2508 1908 -2502
rect 1902 -2514 1908 -2508
rect 1902 -2520 1908 -2514
rect 1902 -2526 1908 -2520
rect 1902 -2532 1908 -2526
rect 1902 -2538 1908 -2532
rect 1902 -2544 1908 -2538
rect 1902 -2550 1908 -2544
rect 1902 -2556 1908 -2550
rect 1902 -2562 1908 -2556
rect 1902 -2568 1908 -2562
rect 1902 -2574 1908 -2568
rect 1902 -2580 1908 -2574
rect 1902 -2652 1908 -2646
rect 1902 -2658 1908 -2652
rect 1902 -2664 1908 -2658
rect 1902 -2670 1908 -2664
rect 1902 -2676 1908 -2670
rect 1902 -2682 1908 -2676
rect 1902 -2688 1908 -2682
rect 1902 -2694 1908 -2688
rect 1902 -2700 1908 -2694
rect 1902 -2706 1908 -2700
rect 1902 -2712 1908 -2706
rect 1902 -2718 1908 -2712
rect 1902 -2724 1908 -2718
rect 1902 -2730 1908 -2724
rect 1902 -2736 1908 -2730
rect 1902 -2742 1908 -2736
rect 1902 -2748 1908 -2742
rect 1902 -2754 1908 -2748
rect 1902 -2760 1908 -2754
rect 1902 -2766 1908 -2760
rect 1902 -2772 1908 -2766
rect 1902 -2778 1908 -2772
rect 1902 -2784 1908 -2778
rect 1902 -2790 1908 -2784
rect 1902 -2796 1908 -2790
rect 1902 -2802 1908 -2796
rect 1902 -2808 1908 -2802
rect 1902 -2814 1908 -2808
rect 1902 -2820 1908 -2814
rect 1902 -2826 1908 -2820
rect 1902 -2832 1908 -2826
rect 1902 -2838 1908 -2832
rect 1902 -2844 1908 -2838
rect 1902 -2850 1908 -2844
rect 1902 -2856 1908 -2850
rect 1902 -2862 1908 -2856
rect 1902 -2868 1908 -2862
rect 1902 -2874 1908 -2868
rect 1902 -2880 1908 -2874
rect 1902 -2886 1908 -2880
rect 1902 -2892 1908 -2886
rect 1902 -2898 1908 -2892
rect 1902 -2904 1908 -2898
rect 1902 -2910 1908 -2904
rect 1902 -2916 1908 -2910
rect 1902 -2922 1908 -2916
rect 1902 -2928 1908 -2922
rect 1902 -2934 1908 -2928
rect 1902 -2940 1908 -2934
rect 1902 -2946 1908 -2940
rect 1902 -2952 1908 -2946
rect 1902 -2958 1908 -2952
rect 1902 -2964 1908 -2958
rect 1902 -2970 1908 -2964
rect 1902 -2976 1908 -2970
rect 1902 -2982 1908 -2976
rect 1902 -2988 1908 -2982
rect 1902 -2994 1908 -2988
rect 1902 -3000 1908 -2994
rect 1902 -3006 1908 -3000
rect 1902 -3012 1908 -3006
rect 1902 -3018 1908 -3012
rect 1902 -3024 1908 -3018
rect 1902 -3030 1908 -3024
rect 1902 -3036 1908 -3030
rect 1902 -3042 1908 -3036
rect 1902 -3048 1908 -3042
rect 1902 -3054 1908 -3048
rect 1902 -3060 1908 -3054
rect 1902 -3066 1908 -3060
rect 1902 -3072 1908 -3066
rect 1902 -3078 1908 -3072
rect 1902 -3084 1908 -3078
rect 1902 -3090 1908 -3084
rect 1902 -3096 1908 -3090
rect 1902 -3102 1908 -3096
rect 1902 -3108 1908 -3102
rect 1902 -3114 1908 -3108
rect 1902 -3120 1908 -3114
rect 1902 -3126 1908 -3120
rect 1902 -3132 1908 -3126
rect 1902 -3138 1908 -3132
rect 1902 -3144 1908 -3138
rect 1902 -3198 1908 -3192
rect 1902 -3204 1908 -3198
rect 1902 -3210 1908 -3204
rect 1902 -3216 1908 -3210
rect 1902 -3222 1908 -3216
rect 1902 -3228 1908 -3222
rect 1902 -3234 1908 -3228
rect 1902 -3240 1908 -3234
rect 1902 -3246 1908 -3240
rect 1902 -3252 1908 -3246
rect 1902 -3258 1908 -3252
rect 1902 -3264 1908 -3258
rect 1902 -3270 1908 -3264
rect 1902 -3276 1908 -3270
rect 1902 -3282 1908 -3276
rect 1902 -3288 1908 -3282
rect 1902 -3294 1908 -3288
rect 1902 -3300 1908 -3294
rect 1908 -570 1914 -564
rect 1908 -576 1914 -570
rect 1908 -582 1914 -576
rect 1908 -588 1914 -582
rect 1908 -594 1914 -588
rect 1908 -600 1914 -594
rect 1908 -606 1914 -600
rect 1908 -612 1914 -606
rect 1908 -618 1914 -612
rect 1908 -624 1914 -618
rect 1908 -630 1914 -624
rect 1908 -636 1914 -630
rect 1908 -642 1914 -636
rect 1908 -648 1914 -642
rect 1908 -654 1914 -648
rect 1908 -660 1914 -654
rect 1908 -666 1914 -660
rect 1908 -672 1914 -666
rect 1908 -678 1914 -672
rect 1908 -684 1914 -678
rect 1908 -690 1914 -684
rect 1908 -696 1914 -690
rect 1908 -702 1914 -696
rect 1908 -708 1914 -702
rect 1908 -714 1914 -708
rect 1908 -720 1914 -714
rect 1908 -726 1914 -720
rect 1908 -732 1914 -726
rect 1908 -738 1914 -732
rect 1908 -744 1914 -738
rect 1908 -750 1914 -744
rect 1908 -756 1914 -750
rect 1908 -762 1914 -756
rect 1908 -768 1914 -762
rect 1908 -774 1914 -768
rect 1908 -780 1914 -774
rect 1908 -786 1914 -780
rect 1908 -792 1914 -786
rect 1908 -798 1914 -792
rect 1908 -804 1914 -798
rect 1908 -810 1914 -804
rect 1908 -816 1914 -810
rect 1908 -822 1914 -816
rect 1908 -828 1914 -822
rect 1908 -834 1914 -828
rect 1908 -840 1914 -834
rect 1908 -846 1914 -840
rect 1908 -852 1914 -846
rect 1908 -858 1914 -852
rect 1908 -864 1914 -858
rect 1908 -870 1914 -864
rect 1908 -876 1914 -870
rect 1908 -882 1914 -876
rect 1908 -888 1914 -882
rect 1908 -894 1914 -888
rect 1908 -900 1914 -894
rect 1908 -906 1914 -900
rect 1908 -912 1914 -906
rect 1908 -918 1914 -912
rect 1908 -924 1914 -918
rect 1908 -930 1914 -924
rect 1908 -936 1914 -930
rect 1908 -942 1914 -936
rect 1908 -948 1914 -942
rect 1908 -954 1914 -948
rect 1908 -960 1914 -954
rect 1908 -966 1914 -960
rect 1908 -972 1914 -966
rect 1908 -978 1914 -972
rect 1908 -984 1914 -978
rect 1908 -990 1914 -984
rect 1908 -996 1914 -990
rect 1908 -1002 1914 -996
rect 1908 -1008 1914 -1002
rect 1908 -1014 1914 -1008
rect 1908 -1020 1914 -1014
rect 1908 -1026 1914 -1020
rect 1908 -1032 1914 -1026
rect 1908 -1038 1914 -1032
rect 1908 -1044 1914 -1038
rect 1908 -1050 1914 -1044
rect 1908 -1056 1914 -1050
rect 1908 -1062 1914 -1056
rect 1908 -1068 1914 -1062
rect 1908 -1074 1914 -1068
rect 1908 -1080 1914 -1074
rect 1908 -1086 1914 -1080
rect 1908 -1092 1914 -1086
rect 1908 -1098 1914 -1092
rect 1908 -1104 1914 -1098
rect 1908 -1110 1914 -1104
rect 1908 -1116 1914 -1110
rect 1908 -1122 1914 -1116
rect 1908 -1128 1914 -1122
rect 1908 -1134 1914 -1128
rect 1908 -1140 1914 -1134
rect 1908 -1146 1914 -1140
rect 1908 -1152 1914 -1146
rect 1908 -1158 1914 -1152
rect 1908 -1164 1914 -1158
rect 1908 -1170 1914 -1164
rect 1908 -1176 1914 -1170
rect 1908 -1182 1914 -1176
rect 1908 -1188 1914 -1182
rect 1908 -1194 1914 -1188
rect 1908 -1200 1914 -1194
rect 1908 -1206 1914 -1200
rect 1908 -1212 1914 -1206
rect 1908 -1218 1914 -1212
rect 1908 -1224 1914 -1218
rect 1908 -1230 1914 -1224
rect 1908 -1236 1914 -1230
rect 1908 -1242 1914 -1236
rect 1908 -1248 1914 -1242
rect 1908 -1254 1914 -1248
rect 1908 -1260 1914 -1254
rect 1908 -1266 1914 -1260
rect 1908 -1272 1914 -1266
rect 1908 -1278 1914 -1272
rect 1908 -1284 1914 -1278
rect 1908 -1290 1914 -1284
rect 1908 -1296 1914 -1290
rect 1908 -1302 1914 -1296
rect 1908 -1308 1914 -1302
rect 1908 -1314 1914 -1308
rect 1908 -1320 1914 -1314
rect 1908 -1326 1914 -1320
rect 1908 -1332 1914 -1326
rect 1908 -1338 1914 -1332
rect 1908 -1344 1914 -1338
rect 1908 -1350 1914 -1344
rect 1908 -1356 1914 -1350
rect 1908 -1362 1914 -1356
rect 1908 -1368 1914 -1362
rect 1908 -1374 1914 -1368
rect 1908 -1380 1914 -1374
rect 1908 -1386 1914 -1380
rect 1908 -1392 1914 -1386
rect 1908 -1398 1914 -1392
rect 1908 -1404 1914 -1398
rect 1908 -1410 1914 -1404
rect 1908 -1416 1914 -1410
rect 1908 -1422 1914 -1416
rect 1908 -1428 1914 -1422
rect 1908 -1434 1914 -1428
rect 1908 -1440 1914 -1434
rect 1908 -1446 1914 -1440
rect 1908 -1452 1914 -1446
rect 1908 -1458 1914 -1452
rect 1908 -1464 1914 -1458
rect 1908 -1470 1914 -1464
rect 1908 -1476 1914 -1470
rect 1908 -1482 1914 -1476
rect 1908 -1488 1914 -1482
rect 1908 -1494 1914 -1488
rect 1908 -1500 1914 -1494
rect 1908 -1506 1914 -1500
rect 1908 -1512 1914 -1506
rect 1908 -1518 1914 -1512
rect 1908 -1524 1914 -1518
rect 1908 -1530 1914 -1524
rect 1908 -1536 1914 -1530
rect 1908 -1542 1914 -1536
rect 1908 -1548 1914 -1542
rect 1908 -1554 1914 -1548
rect 1908 -1560 1914 -1554
rect 1908 -1566 1914 -1560
rect 1908 -1572 1914 -1566
rect 1908 -1578 1914 -1572
rect 1908 -1584 1914 -1578
rect 1908 -1590 1914 -1584
rect 1908 -1596 1914 -1590
rect 1908 -1602 1914 -1596
rect 1908 -1608 1914 -1602
rect 1908 -1614 1914 -1608
rect 1908 -1620 1914 -1614
rect 1908 -1626 1914 -1620
rect 1908 -1632 1914 -1626
rect 1908 -1638 1914 -1632
rect 1908 -1644 1914 -1638
rect 1908 -1650 1914 -1644
rect 1908 -1656 1914 -1650
rect 1908 -1662 1914 -1656
rect 1908 -1668 1914 -1662
rect 1908 -1674 1914 -1668
rect 1908 -1680 1914 -1674
rect 1908 -1686 1914 -1680
rect 1908 -1692 1914 -1686
rect 1908 -1698 1914 -1692
rect 1908 -1704 1914 -1698
rect 1908 -1710 1914 -1704
rect 1908 -1716 1914 -1710
rect 1908 -1722 1914 -1716
rect 1908 -1728 1914 -1722
rect 1908 -1734 1914 -1728
rect 1908 -1740 1914 -1734
rect 1908 -1818 1914 -1812
rect 1908 -1824 1914 -1818
rect 1908 -1830 1914 -1824
rect 1908 -1836 1914 -1830
rect 1908 -1842 1914 -1836
rect 1908 -1848 1914 -1842
rect 1908 -1854 1914 -1848
rect 1908 -1860 1914 -1854
rect 1908 -1866 1914 -1860
rect 1908 -1872 1914 -1866
rect 1908 -1878 1914 -1872
rect 1908 -1884 1914 -1878
rect 1908 -1890 1914 -1884
rect 1908 -1896 1914 -1890
rect 1908 -1902 1914 -1896
rect 1908 -1908 1914 -1902
rect 1908 -1914 1914 -1908
rect 1908 -1920 1914 -1914
rect 1908 -1926 1914 -1920
rect 1908 -1932 1914 -1926
rect 1908 -1938 1914 -1932
rect 1908 -1944 1914 -1938
rect 1908 -1950 1914 -1944
rect 1908 -1956 1914 -1950
rect 1908 -1962 1914 -1956
rect 1908 -1968 1914 -1962
rect 1908 -1974 1914 -1968
rect 1908 -1980 1914 -1974
rect 1908 -1986 1914 -1980
rect 1908 -1992 1914 -1986
rect 1908 -1998 1914 -1992
rect 1908 -2004 1914 -1998
rect 1908 -2010 1914 -2004
rect 1908 -2016 1914 -2010
rect 1908 -2022 1914 -2016
rect 1908 -2028 1914 -2022
rect 1908 -2034 1914 -2028
rect 1908 -2040 1914 -2034
rect 1908 -2046 1914 -2040
rect 1908 -2052 1914 -2046
rect 1908 -2058 1914 -2052
rect 1908 -2064 1914 -2058
rect 1908 -2070 1914 -2064
rect 1908 -2076 1914 -2070
rect 1908 -2082 1914 -2076
rect 1908 -2088 1914 -2082
rect 1908 -2094 1914 -2088
rect 1908 -2100 1914 -2094
rect 1908 -2106 1914 -2100
rect 1908 -2112 1914 -2106
rect 1908 -2118 1914 -2112
rect 1908 -2124 1914 -2118
rect 1908 -2130 1914 -2124
rect 1908 -2136 1914 -2130
rect 1908 -2142 1914 -2136
rect 1908 -2148 1914 -2142
rect 1908 -2154 1914 -2148
rect 1908 -2160 1914 -2154
rect 1908 -2166 1914 -2160
rect 1908 -2172 1914 -2166
rect 1908 -2178 1914 -2172
rect 1908 -2184 1914 -2178
rect 1908 -2190 1914 -2184
rect 1908 -2196 1914 -2190
rect 1908 -2202 1914 -2196
rect 1908 -2208 1914 -2202
rect 1908 -2214 1914 -2208
rect 1908 -2220 1914 -2214
rect 1908 -2226 1914 -2220
rect 1908 -2232 1914 -2226
rect 1908 -2238 1914 -2232
rect 1908 -2244 1914 -2238
rect 1908 -2250 1914 -2244
rect 1908 -2256 1914 -2250
rect 1908 -2262 1914 -2256
rect 1908 -2268 1914 -2262
rect 1908 -2274 1914 -2268
rect 1908 -2280 1914 -2274
rect 1908 -2286 1914 -2280
rect 1908 -2292 1914 -2286
rect 1908 -2298 1914 -2292
rect 1908 -2304 1914 -2298
rect 1908 -2310 1914 -2304
rect 1908 -2316 1914 -2310
rect 1908 -2322 1914 -2316
rect 1908 -2328 1914 -2322
rect 1908 -2334 1914 -2328
rect 1908 -2340 1914 -2334
rect 1908 -2346 1914 -2340
rect 1908 -2352 1914 -2346
rect 1908 -2358 1914 -2352
rect 1908 -2364 1914 -2358
rect 1908 -2370 1914 -2364
rect 1908 -2376 1914 -2370
rect 1908 -2382 1914 -2376
rect 1908 -2388 1914 -2382
rect 1908 -2394 1914 -2388
rect 1908 -2400 1914 -2394
rect 1908 -2406 1914 -2400
rect 1908 -2412 1914 -2406
rect 1908 -2418 1914 -2412
rect 1908 -2424 1914 -2418
rect 1908 -2430 1914 -2424
rect 1908 -2436 1914 -2430
rect 1908 -2442 1914 -2436
rect 1908 -2448 1914 -2442
rect 1908 -2454 1914 -2448
rect 1908 -2460 1914 -2454
rect 1908 -2466 1914 -2460
rect 1908 -2472 1914 -2466
rect 1908 -2478 1914 -2472
rect 1908 -2484 1914 -2478
rect 1908 -2490 1914 -2484
rect 1908 -2496 1914 -2490
rect 1908 -2502 1914 -2496
rect 1908 -2508 1914 -2502
rect 1908 -2514 1914 -2508
rect 1908 -2520 1914 -2514
rect 1908 -2526 1914 -2520
rect 1908 -2532 1914 -2526
rect 1908 -2538 1914 -2532
rect 1908 -2544 1914 -2538
rect 1908 -2550 1914 -2544
rect 1908 -2556 1914 -2550
rect 1908 -2562 1914 -2556
rect 1908 -2568 1914 -2562
rect 1908 -2574 1914 -2568
rect 1908 -2652 1914 -2646
rect 1908 -2658 1914 -2652
rect 1908 -2664 1914 -2658
rect 1908 -2670 1914 -2664
rect 1908 -2676 1914 -2670
rect 1908 -2682 1914 -2676
rect 1908 -2688 1914 -2682
rect 1908 -2694 1914 -2688
rect 1908 -2700 1914 -2694
rect 1908 -2706 1914 -2700
rect 1908 -2712 1914 -2706
rect 1908 -2718 1914 -2712
rect 1908 -2724 1914 -2718
rect 1908 -2730 1914 -2724
rect 1908 -2736 1914 -2730
rect 1908 -2742 1914 -2736
rect 1908 -2748 1914 -2742
rect 1908 -2754 1914 -2748
rect 1908 -2760 1914 -2754
rect 1908 -2766 1914 -2760
rect 1908 -2772 1914 -2766
rect 1908 -2778 1914 -2772
rect 1908 -2784 1914 -2778
rect 1908 -2790 1914 -2784
rect 1908 -2796 1914 -2790
rect 1908 -2802 1914 -2796
rect 1908 -2808 1914 -2802
rect 1908 -2814 1914 -2808
rect 1908 -2820 1914 -2814
rect 1908 -2826 1914 -2820
rect 1908 -2832 1914 -2826
rect 1908 -2838 1914 -2832
rect 1908 -2844 1914 -2838
rect 1908 -2850 1914 -2844
rect 1908 -2856 1914 -2850
rect 1908 -2862 1914 -2856
rect 1908 -2868 1914 -2862
rect 1908 -2874 1914 -2868
rect 1908 -2880 1914 -2874
rect 1908 -2886 1914 -2880
rect 1908 -2892 1914 -2886
rect 1908 -2898 1914 -2892
rect 1908 -2904 1914 -2898
rect 1908 -2910 1914 -2904
rect 1908 -2916 1914 -2910
rect 1908 -2922 1914 -2916
rect 1908 -2928 1914 -2922
rect 1908 -2934 1914 -2928
rect 1908 -2940 1914 -2934
rect 1908 -2946 1914 -2940
rect 1908 -2952 1914 -2946
rect 1908 -2958 1914 -2952
rect 1908 -2964 1914 -2958
rect 1908 -2970 1914 -2964
rect 1908 -2976 1914 -2970
rect 1908 -2982 1914 -2976
rect 1908 -2988 1914 -2982
rect 1908 -2994 1914 -2988
rect 1908 -3000 1914 -2994
rect 1908 -3006 1914 -3000
rect 1908 -3012 1914 -3006
rect 1908 -3018 1914 -3012
rect 1908 -3024 1914 -3018
rect 1908 -3030 1914 -3024
rect 1908 -3036 1914 -3030
rect 1908 -3042 1914 -3036
rect 1908 -3048 1914 -3042
rect 1908 -3054 1914 -3048
rect 1908 -3060 1914 -3054
rect 1908 -3066 1914 -3060
rect 1908 -3072 1914 -3066
rect 1908 -3078 1914 -3072
rect 1908 -3084 1914 -3078
rect 1908 -3090 1914 -3084
rect 1908 -3096 1914 -3090
rect 1908 -3102 1914 -3096
rect 1908 -3108 1914 -3102
rect 1908 -3114 1914 -3108
rect 1908 -3120 1914 -3114
rect 1908 -3126 1914 -3120
rect 1908 -3132 1914 -3126
rect 1908 -3138 1914 -3132
rect 1908 -3192 1914 -3186
rect 1908 -3198 1914 -3192
rect 1908 -3204 1914 -3198
rect 1908 -3210 1914 -3204
rect 1908 -3216 1914 -3210
rect 1908 -3222 1914 -3216
rect 1908 -3228 1914 -3222
rect 1908 -3234 1914 -3228
rect 1908 -3240 1914 -3234
rect 1908 -3246 1914 -3240
rect 1908 -3252 1914 -3246
rect 1908 -3258 1914 -3252
rect 1908 -3264 1914 -3258
rect 1908 -3270 1914 -3264
rect 1908 -3276 1914 -3270
rect 1908 -3282 1914 -3276
rect 1908 -3288 1914 -3282
rect 1908 -3294 1914 -3288
rect 1914 -564 1920 -558
rect 1914 -570 1920 -564
rect 1914 -576 1920 -570
rect 1914 -582 1920 -576
rect 1914 -588 1920 -582
rect 1914 -594 1920 -588
rect 1914 -600 1920 -594
rect 1914 -606 1920 -600
rect 1914 -612 1920 -606
rect 1914 -618 1920 -612
rect 1914 -624 1920 -618
rect 1914 -630 1920 -624
rect 1914 -636 1920 -630
rect 1914 -642 1920 -636
rect 1914 -648 1920 -642
rect 1914 -654 1920 -648
rect 1914 -660 1920 -654
rect 1914 -666 1920 -660
rect 1914 -672 1920 -666
rect 1914 -678 1920 -672
rect 1914 -684 1920 -678
rect 1914 -690 1920 -684
rect 1914 -696 1920 -690
rect 1914 -702 1920 -696
rect 1914 -708 1920 -702
rect 1914 -714 1920 -708
rect 1914 -720 1920 -714
rect 1914 -726 1920 -720
rect 1914 -732 1920 -726
rect 1914 -738 1920 -732
rect 1914 -744 1920 -738
rect 1914 -750 1920 -744
rect 1914 -756 1920 -750
rect 1914 -762 1920 -756
rect 1914 -768 1920 -762
rect 1914 -774 1920 -768
rect 1914 -780 1920 -774
rect 1914 -786 1920 -780
rect 1914 -792 1920 -786
rect 1914 -798 1920 -792
rect 1914 -804 1920 -798
rect 1914 -810 1920 -804
rect 1914 -816 1920 -810
rect 1914 -822 1920 -816
rect 1914 -828 1920 -822
rect 1914 -834 1920 -828
rect 1914 -840 1920 -834
rect 1914 -846 1920 -840
rect 1914 -852 1920 -846
rect 1914 -858 1920 -852
rect 1914 -864 1920 -858
rect 1914 -870 1920 -864
rect 1914 -876 1920 -870
rect 1914 -882 1920 -876
rect 1914 -888 1920 -882
rect 1914 -894 1920 -888
rect 1914 -900 1920 -894
rect 1914 -906 1920 -900
rect 1914 -912 1920 -906
rect 1914 -918 1920 -912
rect 1914 -924 1920 -918
rect 1914 -930 1920 -924
rect 1914 -936 1920 -930
rect 1914 -942 1920 -936
rect 1914 -948 1920 -942
rect 1914 -954 1920 -948
rect 1914 -960 1920 -954
rect 1914 -966 1920 -960
rect 1914 -972 1920 -966
rect 1914 -978 1920 -972
rect 1914 -984 1920 -978
rect 1914 -990 1920 -984
rect 1914 -996 1920 -990
rect 1914 -1002 1920 -996
rect 1914 -1008 1920 -1002
rect 1914 -1014 1920 -1008
rect 1914 -1020 1920 -1014
rect 1914 -1026 1920 -1020
rect 1914 -1032 1920 -1026
rect 1914 -1038 1920 -1032
rect 1914 -1044 1920 -1038
rect 1914 -1050 1920 -1044
rect 1914 -1056 1920 -1050
rect 1914 -1062 1920 -1056
rect 1914 -1068 1920 -1062
rect 1914 -1074 1920 -1068
rect 1914 -1080 1920 -1074
rect 1914 -1086 1920 -1080
rect 1914 -1092 1920 -1086
rect 1914 -1098 1920 -1092
rect 1914 -1104 1920 -1098
rect 1914 -1110 1920 -1104
rect 1914 -1116 1920 -1110
rect 1914 -1122 1920 -1116
rect 1914 -1128 1920 -1122
rect 1914 -1134 1920 -1128
rect 1914 -1140 1920 -1134
rect 1914 -1146 1920 -1140
rect 1914 -1152 1920 -1146
rect 1914 -1158 1920 -1152
rect 1914 -1164 1920 -1158
rect 1914 -1170 1920 -1164
rect 1914 -1176 1920 -1170
rect 1914 -1182 1920 -1176
rect 1914 -1188 1920 -1182
rect 1914 -1194 1920 -1188
rect 1914 -1200 1920 -1194
rect 1914 -1206 1920 -1200
rect 1914 -1212 1920 -1206
rect 1914 -1218 1920 -1212
rect 1914 -1224 1920 -1218
rect 1914 -1230 1920 -1224
rect 1914 -1236 1920 -1230
rect 1914 -1242 1920 -1236
rect 1914 -1248 1920 -1242
rect 1914 -1254 1920 -1248
rect 1914 -1260 1920 -1254
rect 1914 -1266 1920 -1260
rect 1914 -1272 1920 -1266
rect 1914 -1278 1920 -1272
rect 1914 -1284 1920 -1278
rect 1914 -1290 1920 -1284
rect 1914 -1296 1920 -1290
rect 1914 -1302 1920 -1296
rect 1914 -1308 1920 -1302
rect 1914 -1314 1920 -1308
rect 1914 -1320 1920 -1314
rect 1914 -1326 1920 -1320
rect 1914 -1332 1920 -1326
rect 1914 -1338 1920 -1332
rect 1914 -1344 1920 -1338
rect 1914 -1350 1920 -1344
rect 1914 -1356 1920 -1350
rect 1914 -1362 1920 -1356
rect 1914 -1368 1920 -1362
rect 1914 -1374 1920 -1368
rect 1914 -1380 1920 -1374
rect 1914 -1386 1920 -1380
rect 1914 -1392 1920 -1386
rect 1914 -1398 1920 -1392
rect 1914 -1404 1920 -1398
rect 1914 -1410 1920 -1404
rect 1914 -1416 1920 -1410
rect 1914 -1422 1920 -1416
rect 1914 -1428 1920 -1422
rect 1914 -1434 1920 -1428
rect 1914 -1440 1920 -1434
rect 1914 -1446 1920 -1440
rect 1914 -1452 1920 -1446
rect 1914 -1458 1920 -1452
rect 1914 -1464 1920 -1458
rect 1914 -1470 1920 -1464
rect 1914 -1476 1920 -1470
rect 1914 -1482 1920 -1476
rect 1914 -1488 1920 -1482
rect 1914 -1494 1920 -1488
rect 1914 -1500 1920 -1494
rect 1914 -1506 1920 -1500
rect 1914 -1512 1920 -1506
rect 1914 -1518 1920 -1512
rect 1914 -1524 1920 -1518
rect 1914 -1530 1920 -1524
rect 1914 -1536 1920 -1530
rect 1914 -1542 1920 -1536
rect 1914 -1548 1920 -1542
rect 1914 -1554 1920 -1548
rect 1914 -1560 1920 -1554
rect 1914 -1566 1920 -1560
rect 1914 -1572 1920 -1566
rect 1914 -1578 1920 -1572
rect 1914 -1584 1920 -1578
rect 1914 -1590 1920 -1584
rect 1914 -1596 1920 -1590
rect 1914 -1602 1920 -1596
rect 1914 -1608 1920 -1602
rect 1914 -1614 1920 -1608
rect 1914 -1620 1920 -1614
rect 1914 -1626 1920 -1620
rect 1914 -1632 1920 -1626
rect 1914 -1638 1920 -1632
rect 1914 -1644 1920 -1638
rect 1914 -1650 1920 -1644
rect 1914 -1656 1920 -1650
rect 1914 -1662 1920 -1656
rect 1914 -1668 1920 -1662
rect 1914 -1674 1920 -1668
rect 1914 -1680 1920 -1674
rect 1914 -1686 1920 -1680
rect 1914 -1692 1920 -1686
rect 1914 -1698 1920 -1692
rect 1914 -1704 1920 -1698
rect 1914 -1710 1920 -1704
rect 1914 -1716 1920 -1710
rect 1914 -1722 1920 -1716
rect 1914 -1728 1920 -1722
rect 1914 -1734 1920 -1728
rect 1914 -1818 1920 -1812
rect 1914 -1824 1920 -1818
rect 1914 -1830 1920 -1824
rect 1914 -1836 1920 -1830
rect 1914 -1842 1920 -1836
rect 1914 -1848 1920 -1842
rect 1914 -1854 1920 -1848
rect 1914 -1860 1920 -1854
rect 1914 -1866 1920 -1860
rect 1914 -1872 1920 -1866
rect 1914 -1878 1920 -1872
rect 1914 -1884 1920 -1878
rect 1914 -1890 1920 -1884
rect 1914 -1896 1920 -1890
rect 1914 -1902 1920 -1896
rect 1914 -1908 1920 -1902
rect 1914 -1914 1920 -1908
rect 1914 -1920 1920 -1914
rect 1914 -1926 1920 -1920
rect 1914 -1932 1920 -1926
rect 1914 -1938 1920 -1932
rect 1914 -1944 1920 -1938
rect 1914 -1950 1920 -1944
rect 1914 -1956 1920 -1950
rect 1914 -1962 1920 -1956
rect 1914 -1968 1920 -1962
rect 1914 -1974 1920 -1968
rect 1914 -1980 1920 -1974
rect 1914 -1986 1920 -1980
rect 1914 -1992 1920 -1986
rect 1914 -1998 1920 -1992
rect 1914 -2004 1920 -1998
rect 1914 -2010 1920 -2004
rect 1914 -2016 1920 -2010
rect 1914 -2022 1920 -2016
rect 1914 -2028 1920 -2022
rect 1914 -2034 1920 -2028
rect 1914 -2040 1920 -2034
rect 1914 -2046 1920 -2040
rect 1914 -2052 1920 -2046
rect 1914 -2058 1920 -2052
rect 1914 -2064 1920 -2058
rect 1914 -2070 1920 -2064
rect 1914 -2076 1920 -2070
rect 1914 -2082 1920 -2076
rect 1914 -2088 1920 -2082
rect 1914 -2094 1920 -2088
rect 1914 -2100 1920 -2094
rect 1914 -2106 1920 -2100
rect 1914 -2112 1920 -2106
rect 1914 -2118 1920 -2112
rect 1914 -2124 1920 -2118
rect 1914 -2130 1920 -2124
rect 1914 -2136 1920 -2130
rect 1914 -2142 1920 -2136
rect 1914 -2148 1920 -2142
rect 1914 -2154 1920 -2148
rect 1914 -2160 1920 -2154
rect 1914 -2166 1920 -2160
rect 1914 -2172 1920 -2166
rect 1914 -2178 1920 -2172
rect 1914 -2184 1920 -2178
rect 1914 -2190 1920 -2184
rect 1914 -2196 1920 -2190
rect 1914 -2202 1920 -2196
rect 1914 -2208 1920 -2202
rect 1914 -2214 1920 -2208
rect 1914 -2220 1920 -2214
rect 1914 -2226 1920 -2220
rect 1914 -2232 1920 -2226
rect 1914 -2238 1920 -2232
rect 1914 -2244 1920 -2238
rect 1914 -2250 1920 -2244
rect 1914 -2256 1920 -2250
rect 1914 -2262 1920 -2256
rect 1914 -2268 1920 -2262
rect 1914 -2274 1920 -2268
rect 1914 -2280 1920 -2274
rect 1914 -2286 1920 -2280
rect 1914 -2292 1920 -2286
rect 1914 -2298 1920 -2292
rect 1914 -2304 1920 -2298
rect 1914 -2310 1920 -2304
rect 1914 -2316 1920 -2310
rect 1914 -2322 1920 -2316
rect 1914 -2328 1920 -2322
rect 1914 -2334 1920 -2328
rect 1914 -2340 1920 -2334
rect 1914 -2346 1920 -2340
rect 1914 -2352 1920 -2346
rect 1914 -2358 1920 -2352
rect 1914 -2364 1920 -2358
rect 1914 -2370 1920 -2364
rect 1914 -2376 1920 -2370
rect 1914 -2382 1920 -2376
rect 1914 -2388 1920 -2382
rect 1914 -2394 1920 -2388
rect 1914 -2400 1920 -2394
rect 1914 -2406 1920 -2400
rect 1914 -2412 1920 -2406
rect 1914 -2418 1920 -2412
rect 1914 -2424 1920 -2418
rect 1914 -2430 1920 -2424
rect 1914 -2436 1920 -2430
rect 1914 -2442 1920 -2436
rect 1914 -2448 1920 -2442
rect 1914 -2454 1920 -2448
rect 1914 -2460 1920 -2454
rect 1914 -2466 1920 -2460
rect 1914 -2472 1920 -2466
rect 1914 -2478 1920 -2472
rect 1914 -2484 1920 -2478
rect 1914 -2490 1920 -2484
rect 1914 -2496 1920 -2490
rect 1914 -2502 1920 -2496
rect 1914 -2508 1920 -2502
rect 1914 -2514 1920 -2508
rect 1914 -2520 1920 -2514
rect 1914 -2526 1920 -2520
rect 1914 -2532 1920 -2526
rect 1914 -2538 1920 -2532
rect 1914 -2544 1920 -2538
rect 1914 -2550 1920 -2544
rect 1914 -2556 1920 -2550
rect 1914 -2562 1920 -2556
rect 1914 -2568 1920 -2562
rect 1914 -2574 1920 -2568
rect 1914 -2652 1920 -2646
rect 1914 -2658 1920 -2652
rect 1914 -2664 1920 -2658
rect 1914 -2670 1920 -2664
rect 1914 -2676 1920 -2670
rect 1914 -2682 1920 -2676
rect 1914 -2688 1920 -2682
rect 1914 -2694 1920 -2688
rect 1914 -2700 1920 -2694
rect 1914 -2706 1920 -2700
rect 1914 -2712 1920 -2706
rect 1914 -2718 1920 -2712
rect 1914 -2724 1920 -2718
rect 1914 -2730 1920 -2724
rect 1914 -2736 1920 -2730
rect 1914 -2742 1920 -2736
rect 1914 -2748 1920 -2742
rect 1914 -2754 1920 -2748
rect 1914 -2760 1920 -2754
rect 1914 -2766 1920 -2760
rect 1914 -2772 1920 -2766
rect 1914 -2778 1920 -2772
rect 1914 -2784 1920 -2778
rect 1914 -2790 1920 -2784
rect 1914 -2796 1920 -2790
rect 1914 -2802 1920 -2796
rect 1914 -2808 1920 -2802
rect 1914 -2814 1920 -2808
rect 1914 -2820 1920 -2814
rect 1914 -2826 1920 -2820
rect 1914 -2832 1920 -2826
rect 1914 -2838 1920 -2832
rect 1914 -2844 1920 -2838
rect 1914 -2850 1920 -2844
rect 1914 -2856 1920 -2850
rect 1914 -2862 1920 -2856
rect 1914 -2868 1920 -2862
rect 1914 -2874 1920 -2868
rect 1914 -2880 1920 -2874
rect 1914 -2886 1920 -2880
rect 1914 -2892 1920 -2886
rect 1914 -2898 1920 -2892
rect 1914 -2904 1920 -2898
rect 1914 -2910 1920 -2904
rect 1914 -2916 1920 -2910
rect 1914 -2922 1920 -2916
rect 1914 -2928 1920 -2922
rect 1914 -2934 1920 -2928
rect 1914 -2940 1920 -2934
rect 1914 -2946 1920 -2940
rect 1914 -2952 1920 -2946
rect 1914 -2958 1920 -2952
rect 1914 -2964 1920 -2958
rect 1914 -2970 1920 -2964
rect 1914 -2976 1920 -2970
rect 1914 -2982 1920 -2976
rect 1914 -2988 1920 -2982
rect 1914 -2994 1920 -2988
rect 1914 -3000 1920 -2994
rect 1914 -3006 1920 -3000
rect 1914 -3012 1920 -3006
rect 1914 -3018 1920 -3012
rect 1914 -3024 1920 -3018
rect 1914 -3030 1920 -3024
rect 1914 -3036 1920 -3030
rect 1914 -3042 1920 -3036
rect 1914 -3048 1920 -3042
rect 1914 -3054 1920 -3048
rect 1914 -3060 1920 -3054
rect 1914 -3066 1920 -3060
rect 1914 -3072 1920 -3066
rect 1914 -3078 1920 -3072
rect 1914 -3084 1920 -3078
rect 1914 -3090 1920 -3084
rect 1914 -3096 1920 -3090
rect 1914 -3102 1920 -3096
rect 1914 -3108 1920 -3102
rect 1914 -3114 1920 -3108
rect 1914 -3120 1920 -3114
rect 1914 -3126 1920 -3120
rect 1914 -3132 1920 -3126
rect 1914 -3138 1920 -3132
rect 1914 -3192 1920 -3186
rect 1914 -3198 1920 -3192
rect 1914 -3204 1920 -3198
rect 1914 -3210 1920 -3204
rect 1914 -3216 1920 -3210
rect 1914 -3222 1920 -3216
rect 1914 -3228 1920 -3222
rect 1914 -3234 1920 -3228
rect 1914 -3240 1920 -3234
rect 1914 -3246 1920 -3240
rect 1914 -3252 1920 -3246
rect 1914 -3258 1920 -3252
rect 1914 -3264 1920 -3258
rect 1914 -3270 1920 -3264
rect 1914 -3276 1920 -3270
rect 1914 -3282 1920 -3276
rect 1914 -3288 1920 -3282
rect 1920 -558 1926 -552
rect 1920 -564 1926 -558
rect 1920 -570 1926 -564
rect 1920 -576 1926 -570
rect 1920 -582 1926 -576
rect 1920 -588 1926 -582
rect 1920 -594 1926 -588
rect 1920 -600 1926 -594
rect 1920 -606 1926 -600
rect 1920 -612 1926 -606
rect 1920 -618 1926 -612
rect 1920 -624 1926 -618
rect 1920 -630 1926 -624
rect 1920 -636 1926 -630
rect 1920 -642 1926 -636
rect 1920 -648 1926 -642
rect 1920 -654 1926 -648
rect 1920 -660 1926 -654
rect 1920 -666 1926 -660
rect 1920 -672 1926 -666
rect 1920 -678 1926 -672
rect 1920 -684 1926 -678
rect 1920 -690 1926 -684
rect 1920 -696 1926 -690
rect 1920 -702 1926 -696
rect 1920 -708 1926 -702
rect 1920 -714 1926 -708
rect 1920 -720 1926 -714
rect 1920 -726 1926 -720
rect 1920 -732 1926 -726
rect 1920 -738 1926 -732
rect 1920 -744 1926 -738
rect 1920 -750 1926 -744
rect 1920 -756 1926 -750
rect 1920 -762 1926 -756
rect 1920 -768 1926 -762
rect 1920 -774 1926 -768
rect 1920 -780 1926 -774
rect 1920 -786 1926 -780
rect 1920 -792 1926 -786
rect 1920 -798 1926 -792
rect 1920 -804 1926 -798
rect 1920 -810 1926 -804
rect 1920 -816 1926 -810
rect 1920 -822 1926 -816
rect 1920 -828 1926 -822
rect 1920 -834 1926 -828
rect 1920 -840 1926 -834
rect 1920 -846 1926 -840
rect 1920 -852 1926 -846
rect 1920 -858 1926 -852
rect 1920 -864 1926 -858
rect 1920 -870 1926 -864
rect 1920 -876 1926 -870
rect 1920 -882 1926 -876
rect 1920 -888 1926 -882
rect 1920 -894 1926 -888
rect 1920 -900 1926 -894
rect 1920 -906 1926 -900
rect 1920 -912 1926 -906
rect 1920 -918 1926 -912
rect 1920 -924 1926 -918
rect 1920 -930 1926 -924
rect 1920 -936 1926 -930
rect 1920 -942 1926 -936
rect 1920 -948 1926 -942
rect 1920 -954 1926 -948
rect 1920 -960 1926 -954
rect 1920 -966 1926 -960
rect 1920 -972 1926 -966
rect 1920 -978 1926 -972
rect 1920 -984 1926 -978
rect 1920 -990 1926 -984
rect 1920 -996 1926 -990
rect 1920 -1002 1926 -996
rect 1920 -1008 1926 -1002
rect 1920 -1014 1926 -1008
rect 1920 -1020 1926 -1014
rect 1920 -1026 1926 -1020
rect 1920 -1032 1926 -1026
rect 1920 -1038 1926 -1032
rect 1920 -1044 1926 -1038
rect 1920 -1050 1926 -1044
rect 1920 -1056 1926 -1050
rect 1920 -1062 1926 -1056
rect 1920 -1068 1926 -1062
rect 1920 -1074 1926 -1068
rect 1920 -1080 1926 -1074
rect 1920 -1086 1926 -1080
rect 1920 -1092 1926 -1086
rect 1920 -1098 1926 -1092
rect 1920 -1104 1926 -1098
rect 1920 -1110 1926 -1104
rect 1920 -1116 1926 -1110
rect 1920 -1122 1926 -1116
rect 1920 -1128 1926 -1122
rect 1920 -1134 1926 -1128
rect 1920 -1140 1926 -1134
rect 1920 -1146 1926 -1140
rect 1920 -1152 1926 -1146
rect 1920 -1158 1926 -1152
rect 1920 -1164 1926 -1158
rect 1920 -1170 1926 -1164
rect 1920 -1176 1926 -1170
rect 1920 -1182 1926 -1176
rect 1920 -1188 1926 -1182
rect 1920 -1194 1926 -1188
rect 1920 -1200 1926 -1194
rect 1920 -1206 1926 -1200
rect 1920 -1212 1926 -1206
rect 1920 -1218 1926 -1212
rect 1920 -1224 1926 -1218
rect 1920 -1230 1926 -1224
rect 1920 -1236 1926 -1230
rect 1920 -1242 1926 -1236
rect 1920 -1248 1926 -1242
rect 1920 -1254 1926 -1248
rect 1920 -1260 1926 -1254
rect 1920 -1266 1926 -1260
rect 1920 -1272 1926 -1266
rect 1920 -1278 1926 -1272
rect 1920 -1284 1926 -1278
rect 1920 -1290 1926 -1284
rect 1920 -1296 1926 -1290
rect 1920 -1302 1926 -1296
rect 1920 -1308 1926 -1302
rect 1920 -1314 1926 -1308
rect 1920 -1320 1926 -1314
rect 1920 -1326 1926 -1320
rect 1920 -1332 1926 -1326
rect 1920 -1338 1926 -1332
rect 1920 -1344 1926 -1338
rect 1920 -1350 1926 -1344
rect 1920 -1356 1926 -1350
rect 1920 -1362 1926 -1356
rect 1920 -1368 1926 -1362
rect 1920 -1374 1926 -1368
rect 1920 -1380 1926 -1374
rect 1920 -1386 1926 -1380
rect 1920 -1392 1926 -1386
rect 1920 -1398 1926 -1392
rect 1920 -1404 1926 -1398
rect 1920 -1410 1926 -1404
rect 1920 -1416 1926 -1410
rect 1920 -1422 1926 -1416
rect 1920 -1428 1926 -1422
rect 1920 -1434 1926 -1428
rect 1920 -1440 1926 -1434
rect 1920 -1446 1926 -1440
rect 1920 -1452 1926 -1446
rect 1920 -1458 1926 -1452
rect 1920 -1464 1926 -1458
rect 1920 -1470 1926 -1464
rect 1920 -1476 1926 -1470
rect 1920 -1482 1926 -1476
rect 1920 -1488 1926 -1482
rect 1920 -1494 1926 -1488
rect 1920 -1500 1926 -1494
rect 1920 -1506 1926 -1500
rect 1920 -1512 1926 -1506
rect 1920 -1518 1926 -1512
rect 1920 -1524 1926 -1518
rect 1920 -1530 1926 -1524
rect 1920 -1536 1926 -1530
rect 1920 -1542 1926 -1536
rect 1920 -1548 1926 -1542
rect 1920 -1554 1926 -1548
rect 1920 -1560 1926 -1554
rect 1920 -1566 1926 -1560
rect 1920 -1572 1926 -1566
rect 1920 -1578 1926 -1572
rect 1920 -1584 1926 -1578
rect 1920 -1590 1926 -1584
rect 1920 -1596 1926 -1590
rect 1920 -1602 1926 -1596
rect 1920 -1608 1926 -1602
rect 1920 -1614 1926 -1608
rect 1920 -1620 1926 -1614
rect 1920 -1626 1926 -1620
rect 1920 -1632 1926 -1626
rect 1920 -1638 1926 -1632
rect 1920 -1644 1926 -1638
rect 1920 -1650 1926 -1644
rect 1920 -1656 1926 -1650
rect 1920 -1662 1926 -1656
rect 1920 -1668 1926 -1662
rect 1920 -1674 1926 -1668
rect 1920 -1680 1926 -1674
rect 1920 -1686 1926 -1680
rect 1920 -1692 1926 -1686
rect 1920 -1698 1926 -1692
rect 1920 -1704 1926 -1698
rect 1920 -1710 1926 -1704
rect 1920 -1716 1926 -1710
rect 1920 -1722 1926 -1716
rect 1920 -1728 1926 -1722
rect 1920 -1812 1926 -1806
rect 1920 -1818 1926 -1812
rect 1920 -1824 1926 -1818
rect 1920 -1830 1926 -1824
rect 1920 -1836 1926 -1830
rect 1920 -1842 1926 -1836
rect 1920 -1848 1926 -1842
rect 1920 -1854 1926 -1848
rect 1920 -1860 1926 -1854
rect 1920 -1866 1926 -1860
rect 1920 -1872 1926 -1866
rect 1920 -1878 1926 -1872
rect 1920 -1884 1926 -1878
rect 1920 -1890 1926 -1884
rect 1920 -1896 1926 -1890
rect 1920 -1902 1926 -1896
rect 1920 -1908 1926 -1902
rect 1920 -1914 1926 -1908
rect 1920 -1920 1926 -1914
rect 1920 -1926 1926 -1920
rect 1920 -1932 1926 -1926
rect 1920 -1938 1926 -1932
rect 1920 -1944 1926 -1938
rect 1920 -1950 1926 -1944
rect 1920 -1956 1926 -1950
rect 1920 -1962 1926 -1956
rect 1920 -1968 1926 -1962
rect 1920 -1974 1926 -1968
rect 1920 -1980 1926 -1974
rect 1920 -1986 1926 -1980
rect 1920 -1992 1926 -1986
rect 1920 -1998 1926 -1992
rect 1920 -2004 1926 -1998
rect 1920 -2010 1926 -2004
rect 1920 -2016 1926 -2010
rect 1920 -2022 1926 -2016
rect 1920 -2028 1926 -2022
rect 1920 -2034 1926 -2028
rect 1920 -2040 1926 -2034
rect 1920 -2046 1926 -2040
rect 1920 -2052 1926 -2046
rect 1920 -2058 1926 -2052
rect 1920 -2064 1926 -2058
rect 1920 -2070 1926 -2064
rect 1920 -2076 1926 -2070
rect 1920 -2082 1926 -2076
rect 1920 -2088 1926 -2082
rect 1920 -2094 1926 -2088
rect 1920 -2100 1926 -2094
rect 1920 -2106 1926 -2100
rect 1920 -2112 1926 -2106
rect 1920 -2118 1926 -2112
rect 1920 -2124 1926 -2118
rect 1920 -2130 1926 -2124
rect 1920 -2136 1926 -2130
rect 1920 -2142 1926 -2136
rect 1920 -2148 1926 -2142
rect 1920 -2154 1926 -2148
rect 1920 -2160 1926 -2154
rect 1920 -2166 1926 -2160
rect 1920 -2172 1926 -2166
rect 1920 -2178 1926 -2172
rect 1920 -2184 1926 -2178
rect 1920 -2190 1926 -2184
rect 1920 -2196 1926 -2190
rect 1920 -2202 1926 -2196
rect 1920 -2208 1926 -2202
rect 1920 -2214 1926 -2208
rect 1920 -2220 1926 -2214
rect 1920 -2226 1926 -2220
rect 1920 -2232 1926 -2226
rect 1920 -2238 1926 -2232
rect 1920 -2244 1926 -2238
rect 1920 -2250 1926 -2244
rect 1920 -2256 1926 -2250
rect 1920 -2262 1926 -2256
rect 1920 -2268 1926 -2262
rect 1920 -2274 1926 -2268
rect 1920 -2280 1926 -2274
rect 1920 -2286 1926 -2280
rect 1920 -2292 1926 -2286
rect 1920 -2298 1926 -2292
rect 1920 -2304 1926 -2298
rect 1920 -2310 1926 -2304
rect 1920 -2316 1926 -2310
rect 1920 -2322 1926 -2316
rect 1920 -2328 1926 -2322
rect 1920 -2334 1926 -2328
rect 1920 -2340 1926 -2334
rect 1920 -2346 1926 -2340
rect 1920 -2352 1926 -2346
rect 1920 -2358 1926 -2352
rect 1920 -2364 1926 -2358
rect 1920 -2370 1926 -2364
rect 1920 -2376 1926 -2370
rect 1920 -2382 1926 -2376
rect 1920 -2388 1926 -2382
rect 1920 -2394 1926 -2388
rect 1920 -2400 1926 -2394
rect 1920 -2406 1926 -2400
rect 1920 -2412 1926 -2406
rect 1920 -2418 1926 -2412
rect 1920 -2424 1926 -2418
rect 1920 -2430 1926 -2424
rect 1920 -2436 1926 -2430
rect 1920 -2442 1926 -2436
rect 1920 -2448 1926 -2442
rect 1920 -2454 1926 -2448
rect 1920 -2460 1926 -2454
rect 1920 -2466 1926 -2460
rect 1920 -2472 1926 -2466
rect 1920 -2478 1926 -2472
rect 1920 -2484 1926 -2478
rect 1920 -2490 1926 -2484
rect 1920 -2496 1926 -2490
rect 1920 -2502 1926 -2496
rect 1920 -2508 1926 -2502
rect 1920 -2514 1926 -2508
rect 1920 -2520 1926 -2514
rect 1920 -2526 1926 -2520
rect 1920 -2532 1926 -2526
rect 1920 -2538 1926 -2532
rect 1920 -2544 1926 -2538
rect 1920 -2550 1926 -2544
rect 1920 -2556 1926 -2550
rect 1920 -2562 1926 -2556
rect 1920 -2568 1926 -2562
rect 1920 -2646 1926 -2640
rect 1920 -2652 1926 -2646
rect 1920 -2658 1926 -2652
rect 1920 -2664 1926 -2658
rect 1920 -2670 1926 -2664
rect 1920 -2676 1926 -2670
rect 1920 -2682 1926 -2676
rect 1920 -2688 1926 -2682
rect 1920 -2694 1926 -2688
rect 1920 -2700 1926 -2694
rect 1920 -2706 1926 -2700
rect 1920 -2712 1926 -2706
rect 1920 -2718 1926 -2712
rect 1920 -2724 1926 -2718
rect 1920 -2730 1926 -2724
rect 1920 -2736 1926 -2730
rect 1920 -2742 1926 -2736
rect 1920 -2748 1926 -2742
rect 1920 -2754 1926 -2748
rect 1920 -2760 1926 -2754
rect 1920 -2766 1926 -2760
rect 1920 -2772 1926 -2766
rect 1920 -2778 1926 -2772
rect 1920 -2784 1926 -2778
rect 1920 -2790 1926 -2784
rect 1920 -2796 1926 -2790
rect 1920 -2802 1926 -2796
rect 1920 -2808 1926 -2802
rect 1920 -2814 1926 -2808
rect 1920 -2820 1926 -2814
rect 1920 -2826 1926 -2820
rect 1920 -2832 1926 -2826
rect 1920 -2838 1926 -2832
rect 1920 -2844 1926 -2838
rect 1920 -2850 1926 -2844
rect 1920 -2856 1926 -2850
rect 1920 -2862 1926 -2856
rect 1920 -2868 1926 -2862
rect 1920 -2874 1926 -2868
rect 1920 -2880 1926 -2874
rect 1920 -2886 1926 -2880
rect 1920 -2892 1926 -2886
rect 1920 -2898 1926 -2892
rect 1920 -2904 1926 -2898
rect 1920 -2910 1926 -2904
rect 1920 -2916 1926 -2910
rect 1920 -2922 1926 -2916
rect 1920 -2928 1926 -2922
rect 1920 -2934 1926 -2928
rect 1920 -2940 1926 -2934
rect 1920 -2946 1926 -2940
rect 1920 -2952 1926 -2946
rect 1920 -2958 1926 -2952
rect 1920 -2964 1926 -2958
rect 1920 -2970 1926 -2964
rect 1920 -2976 1926 -2970
rect 1920 -2982 1926 -2976
rect 1920 -2988 1926 -2982
rect 1920 -2994 1926 -2988
rect 1920 -3000 1926 -2994
rect 1920 -3006 1926 -3000
rect 1920 -3012 1926 -3006
rect 1920 -3018 1926 -3012
rect 1920 -3024 1926 -3018
rect 1920 -3030 1926 -3024
rect 1920 -3036 1926 -3030
rect 1920 -3042 1926 -3036
rect 1920 -3048 1926 -3042
rect 1920 -3054 1926 -3048
rect 1920 -3060 1926 -3054
rect 1920 -3066 1926 -3060
rect 1920 -3072 1926 -3066
rect 1920 -3078 1926 -3072
rect 1920 -3084 1926 -3078
rect 1920 -3090 1926 -3084
rect 1920 -3096 1926 -3090
rect 1920 -3102 1926 -3096
rect 1920 -3108 1926 -3102
rect 1920 -3114 1926 -3108
rect 1920 -3120 1926 -3114
rect 1920 -3126 1926 -3120
rect 1920 -3132 1926 -3126
rect 1920 -3138 1926 -3132
rect 1920 -3186 1926 -3180
rect 1920 -3192 1926 -3186
rect 1920 -3198 1926 -3192
rect 1920 -3204 1926 -3198
rect 1920 -3210 1926 -3204
rect 1920 -3216 1926 -3210
rect 1920 -3222 1926 -3216
rect 1920 -3228 1926 -3222
rect 1920 -3234 1926 -3228
rect 1920 -3240 1926 -3234
rect 1920 -3246 1926 -3240
rect 1920 -3252 1926 -3246
rect 1920 -3258 1926 -3252
rect 1920 -3264 1926 -3258
rect 1920 -3270 1926 -3264
rect 1920 -3276 1926 -3270
rect 1920 -3282 1926 -3276
rect 1920 -3288 1926 -3282
rect 1926 -546 1932 -540
rect 1926 -552 1932 -546
rect 1926 -558 1932 -552
rect 1926 -564 1932 -558
rect 1926 -570 1932 -564
rect 1926 -576 1932 -570
rect 1926 -582 1932 -576
rect 1926 -588 1932 -582
rect 1926 -594 1932 -588
rect 1926 -600 1932 -594
rect 1926 -606 1932 -600
rect 1926 -612 1932 -606
rect 1926 -618 1932 -612
rect 1926 -624 1932 -618
rect 1926 -630 1932 -624
rect 1926 -636 1932 -630
rect 1926 -642 1932 -636
rect 1926 -648 1932 -642
rect 1926 -654 1932 -648
rect 1926 -660 1932 -654
rect 1926 -666 1932 -660
rect 1926 -672 1932 -666
rect 1926 -678 1932 -672
rect 1926 -684 1932 -678
rect 1926 -690 1932 -684
rect 1926 -696 1932 -690
rect 1926 -702 1932 -696
rect 1926 -708 1932 -702
rect 1926 -714 1932 -708
rect 1926 -720 1932 -714
rect 1926 -726 1932 -720
rect 1926 -732 1932 -726
rect 1926 -738 1932 -732
rect 1926 -744 1932 -738
rect 1926 -750 1932 -744
rect 1926 -756 1932 -750
rect 1926 -762 1932 -756
rect 1926 -768 1932 -762
rect 1926 -774 1932 -768
rect 1926 -780 1932 -774
rect 1926 -786 1932 -780
rect 1926 -792 1932 -786
rect 1926 -798 1932 -792
rect 1926 -804 1932 -798
rect 1926 -810 1932 -804
rect 1926 -816 1932 -810
rect 1926 -822 1932 -816
rect 1926 -828 1932 -822
rect 1926 -834 1932 -828
rect 1926 -840 1932 -834
rect 1926 -846 1932 -840
rect 1926 -852 1932 -846
rect 1926 -858 1932 -852
rect 1926 -864 1932 -858
rect 1926 -870 1932 -864
rect 1926 -876 1932 -870
rect 1926 -882 1932 -876
rect 1926 -888 1932 -882
rect 1926 -894 1932 -888
rect 1926 -900 1932 -894
rect 1926 -906 1932 -900
rect 1926 -912 1932 -906
rect 1926 -918 1932 -912
rect 1926 -924 1932 -918
rect 1926 -930 1932 -924
rect 1926 -936 1932 -930
rect 1926 -942 1932 -936
rect 1926 -948 1932 -942
rect 1926 -954 1932 -948
rect 1926 -960 1932 -954
rect 1926 -966 1932 -960
rect 1926 -972 1932 -966
rect 1926 -978 1932 -972
rect 1926 -984 1932 -978
rect 1926 -990 1932 -984
rect 1926 -996 1932 -990
rect 1926 -1002 1932 -996
rect 1926 -1008 1932 -1002
rect 1926 -1014 1932 -1008
rect 1926 -1020 1932 -1014
rect 1926 -1026 1932 -1020
rect 1926 -1032 1932 -1026
rect 1926 -1038 1932 -1032
rect 1926 -1044 1932 -1038
rect 1926 -1050 1932 -1044
rect 1926 -1056 1932 -1050
rect 1926 -1062 1932 -1056
rect 1926 -1068 1932 -1062
rect 1926 -1074 1932 -1068
rect 1926 -1080 1932 -1074
rect 1926 -1086 1932 -1080
rect 1926 -1092 1932 -1086
rect 1926 -1098 1932 -1092
rect 1926 -1104 1932 -1098
rect 1926 -1110 1932 -1104
rect 1926 -1116 1932 -1110
rect 1926 -1122 1932 -1116
rect 1926 -1128 1932 -1122
rect 1926 -1134 1932 -1128
rect 1926 -1140 1932 -1134
rect 1926 -1146 1932 -1140
rect 1926 -1152 1932 -1146
rect 1926 -1158 1932 -1152
rect 1926 -1164 1932 -1158
rect 1926 -1170 1932 -1164
rect 1926 -1176 1932 -1170
rect 1926 -1182 1932 -1176
rect 1926 -1188 1932 -1182
rect 1926 -1194 1932 -1188
rect 1926 -1200 1932 -1194
rect 1926 -1206 1932 -1200
rect 1926 -1212 1932 -1206
rect 1926 -1218 1932 -1212
rect 1926 -1224 1932 -1218
rect 1926 -1230 1932 -1224
rect 1926 -1236 1932 -1230
rect 1926 -1242 1932 -1236
rect 1926 -1248 1932 -1242
rect 1926 -1254 1932 -1248
rect 1926 -1260 1932 -1254
rect 1926 -1266 1932 -1260
rect 1926 -1272 1932 -1266
rect 1926 -1278 1932 -1272
rect 1926 -1284 1932 -1278
rect 1926 -1290 1932 -1284
rect 1926 -1296 1932 -1290
rect 1926 -1302 1932 -1296
rect 1926 -1308 1932 -1302
rect 1926 -1314 1932 -1308
rect 1926 -1320 1932 -1314
rect 1926 -1326 1932 -1320
rect 1926 -1332 1932 -1326
rect 1926 -1338 1932 -1332
rect 1926 -1344 1932 -1338
rect 1926 -1350 1932 -1344
rect 1926 -1356 1932 -1350
rect 1926 -1362 1932 -1356
rect 1926 -1368 1932 -1362
rect 1926 -1374 1932 -1368
rect 1926 -1380 1932 -1374
rect 1926 -1386 1932 -1380
rect 1926 -1392 1932 -1386
rect 1926 -1398 1932 -1392
rect 1926 -1404 1932 -1398
rect 1926 -1410 1932 -1404
rect 1926 -1416 1932 -1410
rect 1926 -1422 1932 -1416
rect 1926 -1428 1932 -1422
rect 1926 -1434 1932 -1428
rect 1926 -1440 1932 -1434
rect 1926 -1446 1932 -1440
rect 1926 -1452 1932 -1446
rect 1926 -1458 1932 -1452
rect 1926 -1464 1932 -1458
rect 1926 -1470 1932 -1464
rect 1926 -1476 1932 -1470
rect 1926 -1482 1932 -1476
rect 1926 -1488 1932 -1482
rect 1926 -1494 1932 -1488
rect 1926 -1500 1932 -1494
rect 1926 -1506 1932 -1500
rect 1926 -1512 1932 -1506
rect 1926 -1518 1932 -1512
rect 1926 -1524 1932 -1518
rect 1926 -1530 1932 -1524
rect 1926 -1536 1932 -1530
rect 1926 -1542 1932 -1536
rect 1926 -1548 1932 -1542
rect 1926 -1554 1932 -1548
rect 1926 -1560 1932 -1554
rect 1926 -1566 1932 -1560
rect 1926 -1572 1932 -1566
rect 1926 -1578 1932 -1572
rect 1926 -1584 1932 -1578
rect 1926 -1590 1932 -1584
rect 1926 -1596 1932 -1590
rect 1926 -1602 1932 -1596
rect 1926 -1608 1932 -1602
rect 1926 -1614 1932 -1608
rect 1926 -1620 1932 -1614
rect 1926 -1626 1932 -1620
rect 1926 -1632 1932 -1626
rect 1926 -1638 1932 -1632
rect 1926 -1644 1932 -1638
rect 1926 -1650 1932 -1644
rect 1926 -1656 1932 -1650
rect 1926 -1662 1932 -1656
rect 1926 -1668 1932 -1662
rect 1926 -1674 1932 -1668
rect 1926 -1680 1932 -1674
rect 1926 -1686 1932 -1680
rect 1926 -1692 1932 -1686
rect 1926 -1698 1932 -1692
rect 1926 -1704 1932 -1698
rect 1926 -1710 1932 -1704
rect 1926 -1716 1932 -1710
rect 1926 -1806 1932 -1800
rect 1926 -1812 1932 -1806
rect 1926 -1818 1932 -1812
rect 1926 -1824 1932 -1818
rect 1926 -1830 1932 -1824
rect 1926 -1836 1932 -1830
rect 1926 -1842 1932 -1836
rect 1926 -1848 1932 -1842
rect 1926 -1854 1932 -1848
rect 1926 -1860 1932 -1854
rect 1926 -1866 1932 -1860
rect 1926 -1872 1932 -1866
rect 1926 -1878 1932 -1872
rect 1926 -1884 1932 -1878
rect 1926 -1890 1932 -1884
rect 1926 -1896 1932 -1890
rect 1926 -1902 1932 -1896
rect 1926 -1908 1932 -1902
rect 1926 -1914 1932 -1908
rect 1926 -1920 1932 -1914
rect 1926 -1926 1932 -1920
rect 1926 -1932 1932 -1926
rect 1926 -1938 1932 -1932
rect 1926 -1944 1932 -1938
rect 1926 -1950 1932 -1944
rect 1926 -1956 1932 -1950
rect 1926 -1962 1932 -1956
rect 1926 -1968 1932 -1962
rect 1926 -1974 1932 -1968
rect 1926 -1980 1932 -1974
rect 1926 -1986 1932 -1980
rect 1926 -1992 1932 -1986
rect 1926 -1998 1932 -1992
rect 1926 -2004 1932 -1998
rect 1926 -2010 1932 -2004
rect 1926 -2016 1932 -2010
rect 1926 -2022 1932 -2016
rect 1926 -2028 1932 -2022
rect 1926 -2034 1932 -2028
rect 1926 -2040 1932 -2034
rect 1926 -2046 1932 -2040
rect 1926 -2052 1932 -2046
rect 1926 -2058 1932 -2052
rect 1926 -2064 1932 -2058
rect 1926 -2070 1932 -2064
rect 1926 -2076 1932 -2070
rect 1926 -2082 1932 -2076
rect 1926 -2088 1932 -2082
rect 1926 -2094 1932 -2088
rect 1926 -2100 1932 -2094
rect 1926 -2106 1932 -2100
rect 1926 -2112 1932 -2106
rect 1926 -2118 1932 -2112
rect 1926 -2124 1932 -2118
rect 1926 -2130 1932 -2124
rect 1926 -2136 1932 -2130
rect 1926 -2142 1932 -2136
rect 1926 -2148 1932 -2142
rect 1926 -2154 1932 -2148
rect 1926 -2160 1932 -2154
rect 1926 -2166 1932 -2160
rect 1926 -2172 1932 -2166
rect 1926 -2178 1932 -2172
rect 1926 -2184 1932 -2178
rect 1926 -2190 1932 -2184
rect 1926 -2196 1932 -2190
rect 1926 -2202 1932 -2196
rect 1926 -2208 1932 -2202
rect 1926 -2214 1932 -2208
rect 1926 -2220 1932 -2214
rect 1926 -2226 1932 -2220
rect 1926 -2232 1932 -2226
rect 1926 -2238 1932 -2232
rect 1926 -2244 1932 -2238
rect 1926 -2250 1932 -2244
rect 1926 -2256 1932 -2250
rect 1926 -2262 1932 -2256
rect 1926 -2268 1932 -2262
rect 1926 -2274 1932 -2268
rect 1926 -2280 1932 -2274
rect 1926 -2286 1932 -2280
rect 1926 -2292 1932 -2286
rect 1926 -2298 1932 -2292
rect 1926 -2304 1932 -2298
rect 1926 -2310 1932 -2304
rect 1926 -2316 1932 -2310
rect 1926 -2322 1932 -2316
rect 1926 -2328 1932 -2322
rect 1926 -2334 1932 -2328
rect 1926 -2340 1932 -2334
rect 1926 -2346 1932 -2340
rect 1926 -2352 1932 -2346
rect 1926 -2358 1932 -2352
rect 1926 -2364 1932 -2358
rect 1926 -2370 1932 -2364
rect 1926 -2376 1932 -2370
rect 1926 -2382 1932 -2376
rect 1926 -2388 1932 -2382
rect 1926 -2394 1932 -2388
rect 1926 -2400 1932 -2394
rect 1926 -2406 1932 -2400
rect 1926 -2412 1932 -2406
rect 1926 -2418 1932 -2412
rect 1926 -2424 1932 -2418
rect 1926 -2430 1932 -2424
rect 1926 -2436 1932 -2430
rect 1926 -2442 1932 -2436
rect 1926 -2448 1932 -2442
rect 1926 -2454 1932 -2448
rect 1926 -2460 1932 -2454
rect 1926 -2466 1932 -2460
rect 1926 -2472 1932 -2466
rect 1926 -2478 1932 -2472
rect 1926 -2484 1932 -2478
rect 1926 -2490 1932 -2484
rect 1926 -2496 1932 -2490
rect 1926 -2502 1932 -2496
rect 1926 -2508 1932 -2502
rect 1926 -2514 1932 -2508
rect 1926 -2520 1932 -2514
rect 1926 -2526 1932 -2520
rect 1926 -2532 1932 -2526
rect 1926 -2538 1932 -2532
rect 1926 -2544 1932 -2538
rect 1926 -2550 1932 -2544
rect 1926 -2556 1932 -2550
rect 1926 -2562 1932 -2556
rect 1926 -2646 1932 -2640
rect 1926 -2652 1932 -2646
rect 1926 -2658 1932 -2652
rect 1926 -2664 1932 -2658
rect 1926 -2670 1932 -2664
rect 1926 -2676 1932 -2670
rect 1926 -2682 1932 -2676
rect 1926 -2688 1932 -2682
rect 1926 -2694 1932 -2688
rect 1926 -2700 1932 -2694
rect 1926 -2706 1932 -2700
rect 1926 -2712 1932 -2706
rect 1926 -2718 1932 -2712
rect 1926 -2724 1932 -2718
rect 1926 -2730 1932 -2724
rect 1926 -2736 1932 -2730
rect 1926 -2742 1932 -2736
rect 1926 -2748 1932 -2742
rect 1926 -2754 1932 -2748
rect 1926 -2760 1932 -2754
rect 1926 -2766 1932 -2760
rect 1926 -2772 1932 -2766
rect 1926 -2778 1932 -2772
rect 1926 -2784 1932 -2778
rect 1926 -2790 1932 -2784
rect 1926 -2796 1932 -2790
rect 1926 -2802 1932 -2796
rect 1926 -2808 1932 -2802
rect 1926 -2814 1932 -2808
rect 1926 -2820 1932 -2814
rect 1926 -2826 1932 -2820
rect 1926 -2832 1932 -2826
rect 1926 -2838 1932 -2832
rect 1926 -2844 1932 -2838
rect 1926 -2850 1932 -2844
rect 1926 -2856 1932 -2850
rect 1926 -2862 1932 -2856
rect 1926 -2868 1932 -2862
rect 1926 -2874 1932 -2868
rect 1926 -2880 1932 -2874
rect 1926 -2886 1932 -2880
rect 1926 -2892 1932 -2886
rect 1926 -2898 1932 -2892
rect 1926 -2904 1932 -2898
rect 1926 -2910 1932 -2904
rect 1926 -2916 1932 -2910
rect 1926 -2922 1932 -2916
rect 1926 -2928 1932 -2922
rect 1926 -2934 1932 -2928
rect 1926 -2940 1932 -2934
rect 1926 -2946 1932 -2940
rect 1926 -2952 1932 -2946
rect 1926 -2958 1932 -2952
rect 1926 -2964 1932 -2958
rect 1926 -2970 1932 -2964
rect 1926 -2976 1932 -2970
rect 1926 -2982 1932 -2976
rect 1926 -2988 1932 -2982
rect 1926 -2994 1932 -2988
rect 1926 -3000 1932 -2994
rect 1926 -3006 1932 -3000
rect 1926 -3012 1932 -3006
rect 1926 -3018 1932 -3012
rect 1926 -3024 1932 -3018
rect 1926 -3030 1932 -3024
rect 1926 -3036 1932 -3030
rect 1926 -3042 1932 -3036
rect 1926 -3048 1932 -3042
rect 1926 -3054 1932 -3048
rect 1926 -3060 1932 -3054
rect 1926 -3066 1932 -3060
rect 1926 -3072 1932 -3066
rect 1926 -3078 1932 -3072
rect 1926 -3084 1932 -3078
rect 1926 -3090 1932 -3084
rect 1926 -3096 1932 -3090
rect 1926 -3102 1932 -3096
rect 1926 -3108 1932 -3102
rect 1926 -3114 1932 -3108
rect 1926 -3120 1932 -3114
rect 1926 -3126 1932 -3120
rect 1926 -3132 1932 -3126
rect 1926 -3186 1932 -3180
rect 1926 -3192 1932 -3186
rect 1926 -3198 1932 -3192
rect 1926 -3204 1932 -3198
rect 1926 -3210 1932 -3204
rect 1926 -3216 1932 -3210
rect 1926 -3222 1932 -3216
rect 1926 -3228 1932 -3222
rect 1926 -3234 1932 -3228
rect 1926 -3240 1932 -3234
rect 1926 -3246 1932 -3240
rect 1926 -3252 1932 -3246
rect 1926 -3258 1932 -3252
rect 1926 -3264 1932 -3258
rect 1926 -3270 1932 -3264
rect 1926 -3276 1932 -3270
rect 1926 -3282 1932 -3276
rect 1932 -540 1938 -534
rect 1932 -546 1938 -540
rect 1932 -552 1938 -546
rect 1932 -558 1938 -552
rect 1932 -564 1938 -558
rect 1932 -570 1938 -564
rect 1932 -576 1938 -570
rect 1932 -582 1938 -576
rect 1932 -588 1938 -582
rect 1932 -594 1938 -588
rect 1932 -600 1938 -594
rect 1932 -606 1938 -600
rect 1932 -612 1938 -606
rect 1932 -618 1938 -612
rect 1932 -624 1938 -618
rect 1932 -630 1938 -624
rect 1932 -636 1938 -630
rect 1932 -642 1938 -636
rect 1932 -648 1938 -642
rect 1932 -654 1938 -648
rect 1932 -660 1938 -654
rect 1932 -666 1938 -660
rect 1932 -672 1938 -666
rect 1932 -678 1938 -672
rect 1932 -684 1938 -678
rect 1932 -690 1938 -684
rect 1932 -696 1938 -690
rect 1932 -702 1938 -696
rect 1932 -708 1938 -702
rect 1932 -714 1938 -708
rect 1932 -720 1938 -714
rect 1932 -726 1938 -720
rect 1932 -732 1938 -726
rect 1932 -738 1938 -732
rect 1932 -744 1938 -738
rect 1932 -750 1938 -744
rect 1932 -756 1938 -750
rect 1932 -762 1938 -756
rect 1932 -768 1938 -762
rect 1932 -774 1938 -768
rect 1932 -780 1938 -774
rect 1932 -786 1938 -780
rect 1932 -792 1938 -786
rect 1932 -798 1938 -792
rect 1932 -804 1938 -798
rect 1932 -810 1938 -804
rect 1932 -816 1938 -810
rect 1932 -822 1938 -816
rect 1932 -828 1938 -822
rect 1932 -834 1938 -828
rect 1932 -840 1938 -834
rect 1932 -846 1938 -840
rect 1932 -852 1938 -846
rect 1932 -858 1938 -852
rect 1932 -864 1938 -858
rect 1932 -870 1938 -864
rect 1932 -876 1938 -870
rect 1932 -882 1938 -876
rect 1932 -888 1938 -882
rect 1932 -894 1938 -888
rect 1932 -900 1938 -894
rect 1932 -906 1938 -900
rect 1932 -912 1938 -906
rect 1932 -918 1938 -912
rect 1932 -924 1938 -918
rect 1932 -930 1938 -924
rect 1932 -936 1938 -930
rect 1932 -942 1938 -936
rect 1932 -948 1938 -942
rect 1932 -954 1938 -948
rect 1932 -960 1938 -954
rect 1932 -966 1938 -960
rect 1932 -972 1938 -966
rect 1932 -978 1938 -972
rect 1932 -984 1938 -978
rect 1932 -990 1938 -984
rect 1932 -996 1938 -990
rect 1932 -1002 1938 -996
rect 1932 -1008 1938 -1002
rect 1932 -1014 1938 -1008
rect 1932 -1020 1938 -1014
rect 1932 -1026 1938 -1020
rect 1932 -1032 1938 -1026
rect 1932 -1038 1938 -1032
rect 1932 -1044 1938 -1038
rect 1932 -1050 1938 -1044
rect 1932 -1056 1938 -1050
rect 1932 -1062 1938 -1056
rect 1932 -1068 1938 -1062
rect 1932 -1074 1938 -1068
rect 1932 -1080 1938 -1074
rect 1932 -1086 1938 -1080
rect 1932 -1092 1938 -1086
rect 1932 -1098 1938 -1092
rect 1932 -1104 1938 -1098
rect 1932 -1110 1938 -1104
rect 1932 -1116 1938 -1110
rect 1932 -1122 1938 -1116
rect 1932 -1128 1938 -1122
rect 1932 -1134 1938 -1128
rect 1932 -1140 1938 -1134
rect 1932 -1146 1938 -1140
rect 1932 -1152 1938 -1146
rect 1932 -1158 1938 -1152
rect 1932 -1164 1938 -1158
rect 1932 -1170 1938 -1164
rect 1932 -1176 1938 -1170
rect 1932 -1182 1938 -1176
rect 1932 -1188 1938 -1182
rect 1932 -1194 1938 -1188
rect 1932 -1200 1938 -1194
rect 1932 -1206 1938 -1200
rect 1932 -1212 1938 -1206
rect 1932 -1218 1938 -1212
rect 1932 -1224 1938 -1218
rect 1932 -1230 1938 -1224
rect 1932 -1236 1938 -1230
rect 1932 -1242 1938 -1236
rect 1932 -1248 1938 -1242
rect 1932 -1254 1938 -1248
rect 1932 -1260 1938 -1254
rect 1932 -1266 1938 -1260
rect 1932 -1272 1938 -1266
rect 1932 -1278 1938 -1272
rect 1932 -1284 1938 -1278
rect 1932 -1290 1938 -1284
rect 1932 -1296 1938 -1290
rect 1932 -1302 1938 -1296
rect 1932 -1308 1938 -1302
rect 1932 -1314 1938 -1308
rect 1932 -1320 1938 -1314
rect 1932 -1326 1938 -1320
rect 1932 -1332 1938 -1326
rect 1932 -1338 1938 -1332
rect 1932 -1344 1938 -1338
rect 1932 -1350 1938 -1344
rect 1932 -1356 1938 -1350
rect 1932 -1362 1938 -1356
rect 1932 -1368 1938 -1362
rect 1932 -1374 1938 -1368
rect 1932 -1380 1938 -1374
rect 1932 -1386 1938 -1380
rect 1932 -1392 1938 -1386
rect 1932 -1398 1938 -1392
rect 1932 -1404 1938 -1398
rect 1932 -1410 1938 -1404
rect 1932 -1416 1938 -1410
rect 1932 -1422 1938 -1416
rect 1932 -1428 1938 -1422
rect 1932 -1434 1938 -1428
rect 1932 -1440 1938 -1434
rect 1932 -1446 1938 -1440
rect 1932 -1452 1938 -1446
rect 1932 -1458 1938 -1452
rect 1932 -1464 1938 -1458
rect 1932 -1470 1938 -1464
rect 1932 -1476 1938 -1470
rect 1932 -1482 1938 -1476
rect 1932 -1488 1938 -1482
rect 1932 -1494 1938 -1488
rect 1932 -1500 1938 -1494
rect 1932 -1506 1938 -1500
rect 1932 -1512 1938 -1506
rect 1932 -1518 1938 -1512
rect 1932 -1524 1938 -1518
rect 1932 -1530 1938 -1524
rect 1932 -1536 1938 -1530
rect 1932 -1542 1938 -1536
rect 1932 -1548 1938 -1542
rect 1932 -1554 1938 -1548
rect 1932 -1560 1938 -1554
rect 1932 -1566 1938 -1560
rect 1932 -1572 1938 -1566
rect 1932 -1578 1938 -1572
rect 1932 -1584 1938 -1578
rect 1932 -1590 1938 -1584
rect 1932 -1596 1938 -1590
rect 1932 -1602 1938 -1596
rect 1932 -1608 1938 -1602
rect 1932 -1614 1938 -1608
rect 1932 -1620 1938 -1614
rect 1932 -1626 1938 -1620
rect 1932 -1632 1938 -1626
rect 1932 -1638 1938 -1632
rect 1932 -1644 1938 -1638
rect 1932 -1650 1938 -1644
rect 1932 -1656 1938 -1650
rect 1932 -1662 1938 -1656
rect 1932 -1668 1938 -1662
rect 1932 -1674 1938 -1668
rect 1932 -1680 1938 -1674
rect 1932 -1686 1938 -1680
rect 1932 -1692 1938 -1686
rect 1932 -1698 1938 -1692
rect 1932 -1704 1938 -1698
rect 1932 -1710 1938 -1704
rect 1932 -1800 1938 -1794
rect 1932 -1806 1938 -1800
rect 1932 -1812 1938 -1806
rect 1932 -1818 1938 -1812
rect 1932 -1824 1938 -1818
rect 1932 -1830 1938 -1824
rect 1932 -1836 1938 -1830
rect 1932 -1842 1938 -1836
rect 1932 -1848 1938 -1842
rect 1932 -1854 1938 -1848
rect 1932 -1860 1938 -1854
rect 1932 -1866 1938 -1860
rect 1932 -1872 1938 -1866
rect 1932 -1878 1938 -1872
rect 1932 -1884 1938 -1878
rect 1932 -1890 1938 -1884
rect 1932 -1896 1938 -1890
rect 1932 -1902 1938 -1896
rect 1932 -1908 1938 -1902
rect 1932 -1914 1938 -1908
rect 1932 -1920 1938 -1914
rect 1932 -1926 1938 -1920
rect 1932 -1932 1938 -1926
rect 1932 -1938 1938 -1932
rect 1932 -1944 1938 -1938
rect 1932 -1950 1938 -1944
rect 1932 -1956 1938 -1950
rect 1932 -1962 1938 -1956
rect 1932 -1968 1938 -1962
rect 1932 -1974 1938 -1968
rect 1932 -1980 1938 -1974
rect 1932 -1986 1938 -1980
rect 1932 -1992 1938 -1986
rect 1932 -1998 1938 -1992
rect 1932 -2004 1938 -1998
rect 1932 -2010 1938 -2004
rect 1932 -2016 1938 -2010
rect 1932 -2022 1938 -2016
rect 1932 -2028 1938 -2022
rect 1932 -2034 1938 -2028
rect 1932 -2040 1938 -2034
rect 1932 -2046 1938 -2040
rect 1932 -2052 1938 -2046
rect 1932 -2058 1938 -2052
rect 1932 -2064 1938 -2058
rect 1932 -2070 1938 -2064
rect 1932 -2076 1938 -2070
rect 1932 -2082 1938 -2076
rect 1932 -2088 1938 -2082
rect 1932 -2094 1938 -2088
rect 1932 -2100 1938 -2094
rect 1932 -2106 1938 -2100
rect 1932 -2112 1938 -2106
rect 1932 -2118 1938 -2112
rect 1932 -2124 1938 -2118
rect 1932 -2130 1938 -2124
rect 1932 -2136 1938 -2130
rect 1932 -2142 1938 -2136
rect 1932 -2148 1938 -2142
rect 1932 -2154 1938 -2148
rect 1932 -2160 1938 -2154
rect 1932 -2166 1938 -2160
rect 1932 -2172 1938 -2166
rect 1932 -2178 1938 -2172
rect 1932 -2184 1938 -2178
rect 1932 -2190 1938 -2184
rect 1932 -2196 1938 -2190
rect 1932 -2202 1938 -2196
rect 1932 -2208 1938 -2202
rect 1932 -2214 1938 -2208
rect 1932 -2220 1938 -2214
rect 1932 -2226 1938 -2220
rect 1932 -2232 1938 -2226
rect 1932 -2238 1938 -2232
rect 1932 -2244 1938 -2238
rect 1932 -2250 1938 -2244
rect 1932 -2256 1938 -2250
rect 1932 -2262 1938 -2256
rect 1932 -2268 1938 -2262
rect 1932 -2274 1938 -2268
rect 1932 -2280 1938 -2274
rect 1932 -2286 1938 -2280
rect 1932 -2292 1938 -2286
rect 1932 -2298 1938 -2292
rect 1932 -2304 1938 -2298
rect 1932 -2310 1938 -2304
rect 1932 -2316 1938 -2310
rect 1932 -2322 1938 -2316
rect 1932 -2328 1938 -2322
rect 1932 -2334 1938 -2328
rect 1932 -2340 1938 -2334
rect 1932 -2346 1938 -2340
rect 1932 -2352 1938 -2346
rect 1932 -2358 1938 -2352
rect 1932 -2364 1938 -2358
rect 1932 -2370 1938 -2364
rect 1932 -2376 1938 -2370
rect 1932 -2382 1938 -2376
rect 1932 -2388 1938 -2382
rect 1932 -2394 1938 -2388
rect 1932 -2400 1938 -2394
rect 1932 -2406 1938 -2400
rect 1932 -2412 1938 -2406
rect 1932 -2418 1938 -2412
rect 1932 -2424 1938 -2418
rect 1932 -2430 1938 -2424
rect 1932 -2436 1938 -2430
rect 1932 -2442 1938 -2436
rect 1932 -2448 1938 -2442
rect 1932 -2454 1938 -2448
rect 1932 -2460 1938 -2454
rect 1932 -2466 1938 -2460
rect 1932 -2472 1938 -2466
rect 1932 -2478 1938 -2472
rect 1932 -2484 1938 -2478
rect 1932 -2490 1938 -2484
rect 1932 -2496 1938 -2490
rect 1932 -2502 1938 -2496
rect 1932 -2508 1938 -2502
rect 1932 -2514 1938 -2508
rect 1932 -2520 1938 -2514
rect 1932 -2526 1938 -2520
rect 1932 -2532 1938 -2526
rect 1932 -2538 1938 -2532
rect 1932 -2544 1938 -2538
rect 1932 -2550 1938 -2544
rect 1932 -2556 1938 -2550
rect 1932 -2562 1938 -2556
rect 1932 -2640 1938 -2634
rect 1932 -2646 1938 -2640
rect 1932 -2652 1938 -2646
rect 1932 -2658 1938 -2652
rect 1932 -2664 1938 -2658
rect 1932 -2670 1938 -2664
rect 1932 -2676 1938 -2670
rect 1932 -2682 1938 -2676
rect 1932 -2688 1938 -2682
rect 1932 -2694 1938 -2688
rect 1932 -2700 1938 -2694
rect 1932 -2706 1938 -2700
rect 1932 -2712 1938 -2706
rect 1932 -2718 1938 -2712
rect 1932 -2724 1938 -2718
rect 1932 -2730 1938 -2724
rect 1932 -2736 1938 -2730
rect 1932 -2742 1938 -2736
rect 1932 -2748 1938 -2742
rect 1932 -2754 1938 -2748
rect 1932 -2760 1938 -2754
rect 1932 -2766 1938 -2760
rect 1932 -2772 1938 -2766
rect 1932 -2778 1938 -2772
rect 1932 -2784 1938 -2778
rect 1932 -2790 1938 -2784
rect 1932 -2796 1938 -2790
rect 1932 -2802 1938 -2796
rect 1932 -2808 1938 -2802
rect 1932 -2814 1938 -2808
rect 1932 -2820 1938 -2814
rect 1932 -2826 1938 -2820
rect 1932 -2832 1938 -2826
rect 1932 -2838 1938 -2832
rect 1932 -2844 1938 -2838
rect 1932 -2850 1938 -2844
rect 1932 -2856 1938 -2850
rect 1932 -2862 1938 -2856
rect 1932 -2868 1938 -2862
rect 1932 -2874 1938 -2868
rect 1932 -2880 1938 -2874
rect 1932 -2886 1938 -2880
rect 1932 -2892 1938 -2886
rect 1932 -2898 1938 -2892
rect 1932 -2904 1938 -2898
rect 1932 -2910 1938 -2904
rect 1932 -2916 1938 -2910
rect 1932 -2922 1938 -2916
rect 1932 -2928 1938 -2922
rect 1932 -2934 1938 -2928
rect 1932 -2940 1938 -2934
rect 1932 -2946 1938 -2940
rect 1932 -2952 1938 -2946
rect 1932 -2958 1938 -2952
rect 1932 -2964 1938 -2958
rect 1932 -2970 1938 -2964
rect 1932 -2976 1938 -2970
rect 1932 -2982 1938 -2976
rect 1932 -2988 1938 -2982
rect 1932 -2994 1938 -2988
rect 1932 -3000 1938 -2994
rect 1932 -3006 1938 -3000
rect 1932 -3012 1938 -3006
rect 1932 -3018 1938 -3012
rect 1932 -3024 1938 -3018
rect 1932 -3030 1938 -3024
rect 1932 -3036 1938 -3030
rect 1932 -3042 1938 -3036
rect 1932 -3048 1938 -3042
rect 1932 -3054 1938 -3048
rect 1932 -3060 1938 -3054
rect 1932 -3066 1938 -3060
rect 1932 -3072 1938 -3066
rect 1932 -3078 1938 -3072
rect 1932 -3084 1938 -3078
rect 1932 -3090 1938 -3084
rect 1932 -3096 1938 -3090
rect 1932 -3102 1938 -3096
rect 1932 -3108 1938 -3102
rect 1932 -3114 1938 -3108
rect 1932 -3120 1938 -3114
rect 1932 -3126 1938 -3120
rect 1932 -3132 1938 -3126
rect 1932 -3186 1938 -3180
rect 1932 -3192 1938 -3186
rect 1932 -3198 1938 -3192
rect 1932 -3204 1938 -3198
rect 1932 -3210 1938 -3204
rect 1932 -3216 1938 -3210
rect 1932 -3222 1938 -3216
rect 1932 -3228 1938 -3222
rect 1932 -3234 1938 -3228
rect 1932 -3240 1938 -3234
rect 1932 -3246 1938 -3240
rect 1932 -3252 1938 -3246
rect 1932 -3258 1938 -3252
rect 1932 -3264 1938 -3258
rect 1932 -3270 1938 -3264
rect 1932 -3276 1938 -3270
rect 1938 -534 1944 -528
rect 1938 -540 1944 -534
rect 1938 -546 1944 -540
rect 1938 -552 1944 -546
rect 1938 -558 1944 -552
rect 1938 -564 1944 -558
rect 1938 -570 1944 -564
rect 1938 -576 1944 -570
rect 1938 -582 1944 -576
rect 1938 -588 1944 -582
rect 1938 -594 1944 -588
rect 1938 -600 1944 -594
rect 1938 -606 1944 -600
rect 1938 -612 1944 -606
rect 1938 -618 1944 -612
rect 1938 -624 1944 -618
rect 1938 -630 1944 -624
rect 1938 -636 1944 -630
rect 1938 -642 1944 -636
rect 1938 -648 1944 -642
rect 1938 -654 1944 -648
rect 1938 -660 1944 -654
rect 1938 -666 1944 -660
rect 1938 -672 1944 -666
rect 1938 -678 1944 -672
rect 1938 -684 1944 -678
rect 1938 -690 1944 -684
rect 1938 -696 1944 -690
rect 1938 -702 1944 -696
rect 1938 -708 1944 -702
rect 1938 -714 1944 -708
rect 1938 -720 1944 -714
rect 1938 -726 1944 -720
rect 1938 -732 1944 -726
rect 1938 -738 1944 -732
rect 1938 -744 1944 -738
rect 1938 -750 1944 -744
rect 1938 -756 1944 -750
rect 1938 -762 1944 -756
rect 1938 -768 1944 -762
rect 1938 -774 1944 -768
rect 1938 -780 1944 -774
rect 1938 -786 1944 -780
rect 1938 -792 1944 -786
rect 1938 -798 1944 -792
rect 1938 -804 1944 -798
rect 1938 -810 1944 -804
rect 1938 -816 1944 -810
rect 1938 -822 1944 -816
rect 1938 -828 1944 -822
rect 1938 -834 1944 -828
rect 1938 -840 1944 -834
rect 1938 -846 1944 -840
rect 1938 -852 1944 -846
rect 1938 -858 1944 -852
rect 1938 -864 1944 -858
rect 1938 -870 1944 -864
rect 1938 -876 1944 -870
rect 1938 -882 1944 -876
rect 1938 -888 1944 -882
rect 1938 -894 1944 -888
rect 1938 -900 1944 -894
rect 1938 -906 1944 -900
rect 1938 -912 1944 -906
rect 1938 -918 1944 -912
rect 1938 -924 1944 -918
rect 1938 -930 1944 -924
rect 1938 -936 1944 -930
rect 1938 -942 1944 -936
rect 1938 -948 1944 -942
rect 1938 -954 1944 -948
rect 1938 -960 1944 -954
rect 1938 -966 1944 -960
rect 1938 -972 1944 -966
rect 1938 -978 1944 -972
rect 1938 -984 1944 -978
rect 1938 -990 1944 -984
rect 1938 -996 1944 -990
rect 1938 -1002 1944 -996
rect 1938 -1008 1944 -1002
rect 1938 -1014 1944 -1008
rect 1938 -1020 1944 -1014
rect 1938 -1026 1944 -1020
rect 1938 -1032 1944 -1026
rect 1938 -1038 1944 -1032
rect 1938 -1044 1944 -1038
rect 1938 -1050 1944 -1044
rect 1938 -1056 1944 -1050
rect 1938 -1062 1944 -1056
rect 1938 -1068 1944 -1062
rect 1938 -1074 1944 -1068
rect 1938 -1080 1944 -1074
rect 1938 -1086 1944 -1080
rect 1938 -1092 1944 -1086
rect 1938 -1098 1944 -1092
rect 1938 -1104 1944 -1098
rect 1938 -1110 1944 -1104
rect 1938 -1116 1944 -1110
rect 1938 -1122 1944 -1116
rect 1938 -1128 1944 -1122
rect 1938 -1134 1944 -1128
rect 1938 -1140 1944 -1134
rect 1938 -1146 1944 -1140
rect 1938 -1152 1944 -1146
rect 1938 -1158 1944 -1152
rect 1938 -1164 1944 -1158
rect 1938 -1170 1944 -1164
rect 1938 -1176 1944 -1170
rect 1938 -1182 1944 -1176
rect 1938 -1188 1944 -1182
rect 1938 -1194 1944 -1188
rect 1938 -1200 1944 -1194
rect 1938 -1206 1944 -1200
rect 1938 -1212 1944 -1206
rect 1938 -1218 1944 -1212
rect 1938 -1224 1944 -1218
rect 1938 -1230 1944 -1224
rect 1938 -1236 1944 -1230
rect 1938 -1242 1944 -1236
rect 1938 -1248 1944 -1242
rect 1938 -1254 1944 -1248
rect 1938 -1260 1944 -1254
rect 1938 -1266 1944 -1260
rect 1938 -1272 1944 -1266
rect 1938 -1278 1944 -1272
rect 1938 -1284 1944 -1278
rect 1938 -1290 1944 -1284
rect 1938 -1296 1944 -1290
rect 1938 -1302 1944 -1296
rect 1938 -1308 1944 -1302
rect 1938 -1314 1944 -1308
rect 1938 -1320 1944 -1314
rect 1938 -1326 1944 -1320
rect 1938 -1332 1944 -1326
rect 1938 -1338 1944 -1332
rect 1938 -1344 1944 -1338
rect 1938 -1350 1944 -1344
rect 1938 -1356 1944 -1350
rect 1938 -1362 1944 -1356
rect 1938 -1368 1944 -1362
rect 1938 -1374 1944 -1368
rect 1938 -1380 1944 -1374
rect 1938 -1386 1944 -1380
rect 1938 -1392 1944 -1386
rect 1938 -1398 1944 -1392
rect 1938 -1404 1944 -1398
rect 1938 -1410 1944 -1404
rect 1938 -1416 1944 -1410
rect 1938 -1422 1944 -1416
rect 1938 -1428 1944 -1422
rect 1938 -1434 1944 -1428
rect 1938 -1440 1944 -1434
rect 1938 -1446 1944 -1440
rect 1938 -1452 1944 -1446
rect 1938 -1458 1944 -1452
rect 1938 -1464 1944 -1458
rect 1938 -1470 1944 -1464
rect 1938 -1476 1944 -1470
rect 1938 -1482 1944 -1476
rect 1938 -1488 1944 -1482
rect 1938 -1494 1944 -1488
rect 1938 -1500 1944 -1494
rect 1938 -1506 1944 -1500
rect 1938 -1512 1944 -1506
rect 1938 -1518 1944 -1512
rect 1938 -1524 1944 -1518
rect 1938 -1530 1944 -1524
rect 1938 -1536 1944 -1530
rect 1938 -1542 1944 -1536
rect 1938 -1548 1944 -1542
rect 1938 -1554 1944 -1548
rect 1938 -1560 1944 -1554
rect 1938 -1566 1944 -1560
rect 1938 -1572 1944 -1566
rect 1938 -1578 1944 -1572
rect 1938 -1584 1944 -1578
rect 1938 -1590 1944 -1584
rect 1938 -1596 1944 -1590
rect 1938 -1602 1944 -1596
rect 1938 -1608 1944 -1602
rect 1938 -1614 1944 -1608
rect 1938 -1620 1944 -1614
rect 1938 -1626 1944 -1620
rect 1938 -1632 1944 -1626
rect 1938 -1638 1944 -1632
rect 1938 -1644 1944 -1638
rect 1938 -1650 1944 -1644
rect 1938 -1656 1944 -1650
rect 1938 -1662 1944 -1656
rect 1938 -1668 1944 -1662
rect 1938 -1674 1944 -1668
rect 1938 -1680 1944 -1674
rect 1938 -1686 1944 -1680
rect 1938 -1692 1944 -1686
rect 1938 -1698 1944 -1692
rect 1938 -1704 1944 -1698
rect 1938 -1794 1944 -1788
rect 1938 -1800 1944 -1794
rect 1938 -1806 1944 -1800
rect 1938 -1812 1944 -1806
rect 1938 -1818 1944 -1812
rect 1938 -1824 1944 -1818
rect 1938 -1830 1944 -1824
rect 1938 -1836 1944 -1830
rect 1938 -1842 1944 -1836
rect 1938 -1848 1944 -1842
rect 1938 -1854 1944 -1848
rect 1938 -1860 1944 -1854
rect 1938 -1866 1944 -1860
rect 1938 -1872 1944 -1866
rect 1938 -1878 1944 -1872
rect 1938 -1884 1944 -1878
rect 1938 -1890 1944 -1884
rect 1938 -1896 1944 -1890
rect 1938 -1902 1944 -1896
rect 1938 -1908 1944 -1902
rect 1938 -1914 1944 -1908
rect 1938 -1920 1944 -1914
rect 1938 -1926 1944 -1920
rect 1938 -1932 1944 -1926
rect 1938 -1938 1944 -1932
rect 1938 -1944 1944 -1938
rect 1938 -1950 1944 -1944
rect 1938 -1956 1944 -1950
rect 1938 -1962 1944 -1956
rect 1938 -1968 1944 -1962
rect 1938 -1974 1944 -1968
rect 1938 -1980 1944 -1974
rect 1938 -1986 1944 -1980
rect 1938 -1992 1944 -1986
rect 1938 -1998 1944 -1992
rect 1938 -2004 1944 -1998
rect 1938 -2010 1944 -2004
rect 1938 -2016 1944 -2010
rect 1938 -2022 1944 -2016
rect 1938 -2028 1944 -2022
rect 1938 -2034 1944 -2028
rect 1938 -2040 1944 -2034
rect 1938 -2046 1944 -2040
rect 1938 -2052 1944 -2046
rect 1938 -2058 1944 -2052
rect 1938 -2064 1944 -2058
rect 1938 -2070 1944 -2064
rect 1938 -2076 1944 -2070
rect 1938 -2082 1944 -2076
rect 1938 -2088 1944 -2082
rect 1938 -2094 1944 -2088
rect 1938 -2100 1944 -2094
rect 1938 -2106 1944 -2100
rect 1938 -2112 1944 -2106
rect 1938 -2118 1944 -2112
rect 1938 -2124 1944 -2118
rect 1938 -2130 1944 -2124
rect 1938 -2136 1944 -2130
rect 1938 -2142 1944 -2136
rect 1938 -2148 1944 -2142
rect 1938 -2154 1944 -2148
rect 1938 -2160 1944 -2154
rect 1938 -2166 1944 -2160
rect 1938 -2172 1944 -2166
rect 1938 -2178 1944 -2172
rect 1938 -2184 1944 -2178
rect 1938 -2190 1944 -2184
rect 1938 -2196 1944 -2190
rect 1938 -2202 1944 -2196
rect 1938 -2208 1944 -2202
rect 1938 -2214 1944 -2208
rect 1938 -2220 1944 -2214
rect 1938 -2226 1944 -2220
rect 1938 -2232 1944 -2226
rect 1938 -2238 1944 -2232
rect 1938 -2244 1944 -2238
rect 1938 -2250 1944 -2244
rect 1938 -2256 1944 -2250
rect 1938 -2262 1944 -2256
rect 1938 -2268 1944 -2262
rect 1938 -2274 1944 -2268
rect 1938 -2280 1944 -2274
rect 1938 -2286 1944 -2280
rect 1938 -2292 1944 -2286
rect 1938 -2298 1944 -2292
rect 1938 -2304 1944 -2298
rect 1938 -2310 1944 -2304
rect 1938 -2316 1944 -2310
rect 1938 -2322 1944 -2316
rect 1938 -2328 1944 -2322
rect 1938 -2334 1944 -2328
rect 1938 -2340 1944 -2334
rect 1938 -2346 1944 -2340
rect 1938 -2352 1944 -2346
rect 1938 -2358 1944 -2352
rect 1938 -2364 1944 -2358
rect 1938 -2370 1944 -2364
rect 1938 -2376 1944 -2370
rect 1938 -2382 1944 -2376
rect 1938 -2388 1944 -2382
rect 1938 -2394 1944 -2388
rect 1938 -2400 1944 -2394
rect 1938 -2406 1944 -2400
rect 1938 -2412 1944 -2406
rect 1938 -2418 1944 -2412
rect 1938 -2424 1944 -2418
rect 1938 -2430 1944 -2424
rect 1938 -2436 1944 -2430
rect 1938 -2442 1944 -2436
rect 1938 -2448 1944 -2442
rect 1938 -2454 1944 -2448
rect 1938 -2460 1944 -2454
rect 1938 -2466 1944 -2460
rect 1938 -2472 1944 -2466
rect 1938 -2478 1944 -2472
rect 1938 -2484 1944 -2478
rect 1938 -2490 1944 -2484
rect 1938 -2496 1944 -2490
rect 1938 -2502 1944 -2496
rect 1938 -2508 1944 -2502
rect 1938 -2514 1944 -2508
rect 1938 -2520 1944 -2514
rect 1938 -2526 1944 -2520
rect 1938 -2532 1944 -2526
rect 1938 -2538 1944 -2532
rect 1938 -2544 1944 -2538
rect 1938 -2550 1944 -2544
rect 1938 -2556 1944 -2550
rect 1938 -2640 1944 -2634
rect 1938 -2646 1944 -2640
rect 1938 -2652 1944 -2646
rect 1938 -2658 1944 -2652
rect 1938 -2664 1944 -2658
rect 1938 -2670 1944 -2664
rect 1938 -2676 1944 -2670
rect 1938 -2682 1944 -2676
rect 1938 -2688 1944 -2682
rect 1938 -2694 1944 -2688
rect 1938 -2700 1944 -2694
rect 1938 -2706 1944 -2700
rect 1938 -2712 1944 -2706
rect 1938 -2718 1944 -2712
rect 1938 -2724 1944 -2718
rect 1938 -2730 1944 -2724
rect 1938 -2736 1944 -2730
rect 1938 -2742 1944 -2736
rect 1938 -2748 1944 -2742
rect 1938 -2754 1944 -2748
rect 1938 -2760 1944 -2754
rect 1938 -2766 1944 -2760
rect 1938 -2772 1944 -2766
rect 1938 -2778 1944 -2772
rect 1938 -2784 1944 -2778
rect 1938 -2790 1944 -2784
rect 1938 -2796 1944 -2790
rect 1938 -2802 1944 -2796
rect 1938 -2808 1944 -2802
rect 1938 -2814 1944 -2808
rect 1938 -2820 1944 -2814
rect 1938 -2826 1944 -2820
rect 1938 -2832 1944 -2826
rect 1938 -2838 1944 -2832
rect 1938 -2844 1944 -2838
rect 1938 -2850 1944 -2844
rect 1938 -2856 1944 -2850
rect 1938 -2862 1944 -2856
rect 1938 -2868 1944 -2862
rect 1938 -2874 1944 -2868
rect 1938 -2880 1944 -2874
rect 1938 -2886 1944 -2880
rect 1938 -2892 1944 -2886
rect 1938 -2898 1944 -2892
rect 1938 -2904 1944 -2898
rect 1938 -2910 1944 -2904
rect 1938 -2916 1944 -2910
rect 1938 -2922 1944 -2916
rect 1938 -2928 1944 -2922
rect 1938 -2934 1944 -2928
rect 1938 -2940 1944 -2934
rect 1938 -2946 1944 -2940
rect 1938 -2952 1944 -2946
rect 1938 -2958 1944 -2952
rect 1938 -2964 1944 -2958
rect 1938 -2970 1944 -2964
rect 1938 -2976 1944 -2970
rect 1938 -2982 1944 -2976
rect 1938 -2988 1944 -2982
rect 1938 -2994 1944 -2988
rect 1938 -3000 1944 -2994
rect 1938 -3006 1944 -3000
rect 1938 -3012 1944 -3006
rect 1938 -3018 1944 -3012
rect 1938 -3024 1944 -3018
rect 1938 -3030 1944 -3024
rect 1938 -3036 1944 -3030
rect 1938 -3042 1944 -3036
rect 1938 -3048 1944 -3042
rect 1938 -3054 1944 -3048
rect 1938 -3060 1944 -3054
rect 1938 -3066 1944 -3060
rect 1938 -3072 1944 -3066
rect 1938 -3078 1944 -3072
rect 1938 -3084 1944 -3078
rect 1938 -3090 1944 -3084
rect 1938 -3096 1944 -3090
rect 1938 -3102 1944 -3096
rect 1938 -3108 1944 -3102
rect 1938 -3114 1944 -3108
rect 1938 -3120 1944 -3114
rect 1938 -3126 1944 -3120
rect 1938 -3180 1944 -3174
rect 1938 -3186 1944 -3180
rect 1938 -3192 1944 -3186
rect 1938 -3198 1944 -3192
rect 1938 -3204 1944 -3198
rect 1938 -3210 1944 -3204
rect 1938 -3216 1944 -3210
rect 1938 -3222 1944 -3216
rect 1938 -3228 1944 -3222
rect 1938 -3234 1944 -3228
rect 1938 -3240 1944 -3234
rect 1938 -3246 1944 -3240
rect 1938 -3252 1944 -3246
rect 1938 -3258 1944 -3252
rect 1938 -3264 1944 -3258
rect 1938 -3270 1944 -3264
rect 1944 -522 1950 -516
rect 1944 -528 1950 -522
rect 1944 -534 1950 -528
rect 1944 -540 1950 -534
rect 1944 -546 1950 -540
rect 1944 -552 1950 -546
rect 1944 -558 1950 -552
rect 1944 -564 1950 -558
rect 1944 -570 1950 -564
rect 1944 -576 1950 -570
rect 1944 -582 1950 -576
rect 1944 -588 1950 -582
rect 1944 -594 1950 -588
rect 1944 -600 1950 -594
rect 1944 -606 1950 -600
rect 1944 -612 1950 -606
rect 1944 -618 1950 -612
rect 1944 -624 1950 -618
rect 1944 -630 1950 -624
rect 1944 -636 1950 -630
rect 1944 -642 1950 -636
rect 1944 -648 1950 -642
rect 1944 -654 1950 -648
rect 1944 -660 1950 -654
rect 1944 -666 1950 -660
rect 1944 -672 1950 -666
rect 1944 -678 1950 -672
rect 1944 -684 1950 -678
rect 1944 -690 1950 -684
rect 1944 -696 1950 -690
rect 1944 -702 1950 -696
rect 1944 -708 1950 -702
rect 1944 -714 1950 -708
rect 1944 -720 1950 -714
rect 1944 -726 1950 -720
rect 1944 -732 1950 -726
rect 1944 -738 1950 -732
rect 1944 -744 1950 -738
rect 1944 -750 1950 -744
rect 1944 -756 1950 -750
rect 1944 -762 1950 -756
rect 1944 -768 1950 -762
rect 1944 -774 1950 -768
rect 1944 -780 1950 -774
rect 1944 -786 1950 -780
rect 1944 -792 1950 -786
rect 1944 -798 1950 -792
rect 1944 -804 1950 -798
rect 1944 -810 1950 -804
rect 1944 -816 1950 -810
rect 1944 -822 1950 -816
rect 1944 -828 1950 -822
rect 1944 -834 1950 -828
rect 1944 -840 1950 -834
rect 1944 -846 1950 -840
rect 1944 -852 1950 -846
rect 1944 -858 1950 -852
rect 1944 -864 1950 -858
rect 1944 -870 1950 -864
rect 1944 -876 1950 -870
rect 1944 -882 1950 -876
rect 1944 -888 1950 -882
rect 1944 -894 1950 -888
rect 1944 -900 1950 -894
rect 1944 -906 1950 -900
rect 1944 -912 1950 -906
rect 1944 -918 1950 -912
rect 1944 -924 1950 -918
rect 1944 -930 1950 -924
rect 1944 -936 1950 -930
rect 1944 -942 1950 -936
rect 1944 -948 1950 -942
rect 1944 -954 1950 -948
rect 1944 -960 1950 -954
rect 1944 -966 1950 -960
rect 1944 -972 1950 -966
rect 1944 -978 1950 -972
rect 1944 -984 1950 -978
rect 1944 -990 1950 -984
rect 1944 -996 1950 -990
rect 1944 -1002 1950 -996
rect 1944 -1008 1950 -1002
rect 1944 -1014 1950 -1008
rect 1944 -1020 1950 -1014
rect 1944 -1026 1950 -1020
rect 1944 -1032 1950 -1026
rect 1944 -1038 1950 -1032
rect 1944 -1044 1950 -1038
rect 1944 -1050 1950 -1044
rect 1944 -1056 1950 -1050
rect 1944 -1062 1950 -1056
rect 1944 -1068 1950 -1062
rect 1944 -1074 1950 -1068
rect 1944 -1080 1950 -1074
rect 1944 -1086 1950 -1080
rect 1944 -1092 1950 -1086
rect 1944 -1098 1950 -1092
rect 1944 -1104 1950 -1098
rect 1944 -1110 1950 -1104
rect 1944 -1116 1950 -1110
rect 1944 -1122 1950 -1116
rect 1944 -1128 1950 -1122
rect 1944 -1134 1950 -1128
rect 1944 -1140 1950 -1134
rect 1944 -1146 1950 -1140
rect 1944 -1152 1950 -1146
rect 1944 -1158 1950 -1152
rect 1944 -1164 1950 -1158
rect 1944 -1170 1950 -1164
rect 1944 -1176 1950 -1170
rect 1944 -1182 1950 -1176
rect 1944 -1188 1950 -1182
rect 1944 -1194 1950 -1188
rect 1944 -1200 1950 -1194
rect 1944 -1206 1950 -1200
rect 1944 -1212 1950 -1206
rect 1944 -1218 1950 -1212
rect 1944 -1224 1950 -1218
rect 1944 -1230 1950 -1224
rect 1944 -1236 1950 -1230
rect 1944 -1242 1950 -1236
rect 1944 -1248 1950 -1242
rect 1944 -1254 1950 -1248
rect 1944 -1260 1950 -1254
rect 1944 -1266 1950 -1260
rect 1944 -1272 1950 -1266
rect 1944 -1278 1950 -1272
rect 1944 -1284 1950 -1278
rect 1944 -1290 1950 -1284
rect 1944 -1296 1950 -1290
rect 1944 -1302 1950 -1296
rect 1944 -1308 1950 -1302
rect 1944 -1314 1950 -1308
rect 1944 -1320 1950 -1314
rect 1944 -1326 1950 -1320
rect 1944 -1332 1950 -1326
rect 1944 -1338 1950 -1332
rect 1944 -1344 1950 -1338
rect 1944 -1350 1950 -1344
rect 1944 -1356 1950 -1350
rect 1944 -1362 1950 -1356
rect 1944 -1368 1950 -1362
rect 1944 -1374 1950 -1368
rect 1944 -1380 1950 -1374
rect 1944 -1386 1950 -1380
rect 1944 -1392 1950 -1386
rect 1944 -1398 1950 -1392
rect 1944 -1404 1950 -1398
rect 1944 -1410 1950 -1404
rect 1944 -1416 1950 -1410
rect 1944 -1422 1950 -1416
rect 1944 -1428 1950 -1422
rect 1944 -1434 1950 -1428
rect 1944 -1440 1950 -1434
rect 1944 -1446 1950 -1440
rect 1944 -1452 1950 -1446
rect 1944 -1458 1950 -1452
rect 1944 -1464 1950 -1458
rect 1944 -1470 1950 -1464
rect 1944 -1476 1950 -1470
rect 1944 -1482 1950 -1476
rect 1944 -1488 1950 -1482
rect 1944 -1494 1950 -1488
rect 1944 -1500 1950 -1494
rect 1944 -1506 1950 -1500
rect 1944 -1512 1950 -1506
rect 1944 -1518 1950 -1512
rect 1944 -1524 1950 -1518
rect 1944 -1530 1950 -1524
rect 1944 -1536 1950 -1530
rect 1944 -1542 1950 -1536
rect 1944 -1548 1950 -1542
rect 1944 -1554 1950 -1548
rect 1944 -1560 1950 -1554
rect 1944 -1566 1950 -1560
rect 1944 -1572 1950 -1566
rect 1944 -1578 1950 -1572
rect 1944 -1584 1950 -1578
rect 1944 -1590 1950 -1584
rect 1944 -1596 1950 -1590
rect 1944 -1602 1950 -1596
rect 1944 -1608 1950 -1602
rect 1944 -1614 1950 -1608
rect 1944 -1620 1950 -1614
rect 1944 -1626 1950 -1620
rect 1944 -1632 1950 -1626
rect 1944 -1638 1950 -1632
rect 1944 -1644 1950 -1638
rect 1944 -1650 1950 -1644
rect 1944 -1656 1950 -1650
rect 1944 -1662 1950 -1656
rect 1944 -1668 1950 -1662
rect 1944 -1674 1950 -1668
rect 1944 -1680 1950 -1674
rect 1944 -1686 1950 -1680
rect 1944 -1692 1950 -1686
rect 1944 -1698 1950 -1692
rect 1944 -1788 1950 -1782
rect 1944 -1794 1950 -1788
rect 1944 -1800 1950 -1794
rect 1944 -1806 1950 -1800
rect 1944 -1812 1950 -1806
rect 1944 -1818 1950 -1812
rect 1944 -1824 1950 -1818
rect 1944 -1830 1950 -1824
rect 1944 -1836 1950 -1830
rect 1944 -1842 1950 -1836
rect 1944 -1848 1950 -1842
rect 1944 -1854 1950 -1848
rect 1944 -1860 1950 -1854
rect 1944 -1866 1950 -1860
rect 1944 -1872 1950 -1866
rect 1944 -1878 1950 -1872
rect 1944 -1884 1950 -1878
rect 1944 -1890 1950 -1884
rect 1944 -1896 1950 -1890
rect 1944 -1902 1950 -1896
rect 1944 -1908 1950 -1902
rect 1944 -1914 1950 -1908
rect 1944 -1920 1950 -1914
rect 1944 -1926 1950 -1920
rect 1944 -1932 1950 -1926
rect 1944 -1938 1950 -1932
rect 1944 -1944 1950 -1938
rect 1944 -1950 1950 -1944
rect 1944 -1956 1950 -1950
rect 1944 -1962 1950 -1956
rect 1944 -1968 1950 -1962
rect 1944 -1974 1950 -1968
rect 1944 -1980 1950 -1974
rect 1944 -1986 1950 -1980
rect 1944 -1992 1950 -1986
rect 1944 -1998 1950 -1992
rect 1944 -2004 1950 -1998
rect 1944 -2010 1950 -2004
rect 1944 -2016 1950 -2010
rect 1944 -2022 1950 -2016
rect 1944 -2028 1950 -2022
rect 1944 -2034 1950 -2028
rect 1944 -2040 1950 -2034
rect 1944 -2046 1950 -2040
rect 1944 -2052 1950 -2046
rect 1944 -2058 1950 -2052
rect 1944 -2064 1950 -2058
rect 1944 -2070 1950 -2064
rect 1944 -2076 1950 -2070
rect 1944 -2082 1950 -2076
rect 1944 -2088 1950 -2082
rect 1944 -2094 1950 -2088
rect 1944 -2100 1950 -2094
rect 1944 -2106 1950 -2100
rect 1944 -2112 1950 -2106
rect 1944 -2118 1950 -2112
rect 1944 -2124 1950 -2118
rect 1944 -2130 1950 -2124
rect 1944 -2136 1950 -2130
rect 1944 -2142 1950 -2136
rect 1944 -2148 1950 -2142
rect 1944 -2154 1950 -2148
rect 1944 -2160 1950 -2154
rect 1944 -2166 1950 -2160
rect 1944 -2172 1950 -2166
rect 1944 -2178 1950 -2172
rect 1944 -2184 1950 -2178
rect 1944 -2190 1950 -2184
rect 1944 -2196 1950 -2190
rect 1944 -2202 1950 -2196
rect 1944 -2208 1950 -2202
rect 1944 -2214 1950 -2208
rect 1944 -2220 1950 -2214
rect 1944 -2226 1950 -2220
rect 1944 -2232 1950 -2226
rect 1944 -2238 1950 -2232
rect 1944 -2244 1950 -2238
rect 1944 -2250 1950 -2244
rect 1944 -2256 1950 -2250
rect 1944 -2262 1950 -2256
rect 1944 -2268 1950 -2262
rect 1944 -2274 1950 -2268
rect 1944 -2280 1950 -2274
rect 1944 -2286 1950 -2280
rect 1944 -2292 1950 -2286
rect 1944 -2298 1950 -2292
rect 1944 -2304 1950 -2298
rect 1944 -2310 1950 -2304
rect 1944 -2316 1950 -2310
rect 1944 -2322 1950 -2316
rect 1944 -2328 1950 -2322
rect 1944 -2334 1950 -2328
rect 1944 -2340 1950 -2334
rect 1944 -2346 1950 -2340
rect 1944 -2352 1950 -2346
rect 1944 -2358 1950 -2352
rect 1944 -2364 1950 -2358
rect 1944 -2370 1950 -2364
rect 1944 -2376 1950 -2370
rect 1944 -2382 1950 -2376
rect 1944 -2388 1950 -2382
rect 1944 -2394 1950 -2388
rect 1944 -2400 1950 -2394
rect 1944 -2406 1950 -2400
rect 1944 -2412 1950 -2406
rect 1944 -2418 1950 -2412
rect 1944 -2424 1950 -2418
rect 1944 -2430 1950 -2424
rect 1944 -2436 1950 -2430
rect 1944 -2442 1950 -2436
rect 1944 -2448 1950 -2442
rect 1944 -2454 1950 -2448
rect 1944 -2460 1950 -2454
rect 1944 -2466 1950 -2460
rect 1944 -2472 1950 -2466
rect 1944 -2478 1950 -2472
rect 1944 -2484 1950 -2478
rect 1944 -2490 1950 -2484
rect 1944 -2496 1950 -2490
rect 1944 -2502 1950 -2496
rect 1944 -2508 1950 -2502
rect 1944 -2514 1950 -2508
rect 1944 -2520 1950 -2514
rect 1944 -2526 1950 -2520
rect 1944 -2532 1950 -2526
rect 1944 -2538 1950 -2532
rect 1944 -2544 1950 -2538
rect 1944 -2550 1950 -2544
rect 1944 -2556 1950 -2550
rect 1944 -2634 1950 -2628
rect 1944 -2640 1950 -2634
rect 1944 -2646 1950 -2640
rect 1944 -2652 1950 -2646
rect 1944 -2658 1950 -2652
rect 1944 -2664 1950 -2658
rect 1944 -2670 1950 -2664
rect 1944 -2676 1950 -2670
rect 1944 -2682 1950 -2676
rect 1944 -2688 1950 -2682
rect 1944 -2694 1950 -2688
rect 1944 -2700 1950 -2694
rect 1944 -2706 1950 -2700
rect 1944 -2712 1950 -2706
rect 1944 -2718 1950 -2712
rect 1944 -2724 1950 -2718
rect 1944 -2730 1950 -2724
rect 1944 -2736 1950 -2730
rect 1944 -2742 1950 -2736
rect 1944 -2748 1950 -2742
rect 1944 -2754 1950 -2748
rect 1944 -2760 1950 -2754
rect 1944 -2766 1950 -2760
rect 1944 -2772 1950 -2766
rect 1944 -2778 1950 -2772
rect 1944 -2784 1950 -2778
rect 1944 -2790 1950 -2784
rect 1944 -2796 1950 -2790
rect 1944 -2802 1950 -2796
rect 1944 -2808 1950 -2802
rect 1944 -2814 1950 -2808
rect 1944 -2820 1950 -2814
rect 1944 -2826 1950 -2820
rect 1944 -2832 1950 -2826
rect 1944 -2838 1950 -2832
rect 1944 -2844 1950 -2838
rect 1944 -2850 1950 -2844
rect 1944 -2856 1950 -2850
rect 1944 -2862 1950 -2856
rect 1944 -2868 1950 -2862
rect 1944 -2874 1950 -2868
rect 1944 -2880 1950 -2874
rect 1944 -2886 1950 -2880
rect 1944 -2892 1950 -2886
rect 1944 -2898 1950 -2892
rect 1944 -2904 1950 -2898
rect 1944 -2910 1950 -2904
rect 1944 -2916 1950 -2910
rect 1944 -2922 1950 -2916
rect 1944 -2928 1950 -2922
rect 1944 -2934 1950 -2928
rect 1944 -2940 1950 -2934
rect 1944 -2946 1950 -2940
rect 1944 -2952 1950 -2946
rect 1944 -2958 1950 -2952
rect 1944 -2964 1950 -2958
rect 1944 -2970 1950 -2964
rect 1944 -2976 1950 -2970
rect 1944 -2982 1950 -2976
rect 1944 -2988 1950 -2982
rect 1944 -2994 1950 -2988
rect 1944 -3000 1950 -2994
rect 1944 -3006 1950 -3000
rect 1944 -3012 1950 -3006
rect 1944 -3018 1950 -3012
rect 1944 -3024 1950 -3018
rect 1944 -3030 1950 -3024
rect 1944 -3036 1950 -3030
rect 1944 -3042 1950 -3036
rect 1944 -3048 1950 -3042
rect 1944 -3054 1950 -3048
rect 1944 -3060 1950 -3054
rect 1944 -3066 1950 -3060
rect 1944 -3072 1950 -3066
rect 1944 -3078 1950 -3072
rect 1944 -3084 1950 -3078
rect 1944 -3090 1950 -3084
rect 1944 -3096 1950 -3090
rect 1944 -3102 1950 -3096
rect 1944 -3108 1950 -3102
rect 1944 -3114 1950 -3108
rect 1944 -3120 1950 -3114
rect 1944 -3126 1950 -3120
rect 1944 -3180 1950 -3174
rect 1944 -3186 1950 -3180
rect 1944 -3192 1950 -3186
rect 1944 -3198 1950 -3192
rect 1944 -3204 1950 -3198
rect 1944 -3210 1950 -3204
rect 1944 -3216 1950 -3210
rect 1944 -3222 1950 -3216
rect 1944 -3228 1950 -3222
rect 1944 -3234 1950 -3228
rect 1944 -3240 1950 -3234
rect 1944 -3246 1950 -3240
rect 1944 -3252 1950 -3246
rect 1944 -3258 1950 -3252
rect 1944 -3264 1950 -3258
rect 1944 -3270 1950 -3264
rect 1950 -516 1956 -510
rect 1950 -522 1956 -516
rect 1950 -528 1956 -522
rect 1950 -534 1956 -528
rect 1950 -540 1956 -534
rect 1950 -546 1956 -540
rect 1950 -552 1956 -546
rect 1950 -558 1956 -552
rect 1950 -564 1956 -558
rect 1950 -570 1956 -564
rect 1950 -576 1956 -570
rect 1950 -582 1956 -576
rect 1950 -588 1956 -582
rect 1950 -594 1956 -588
rect 1950 -600 1956 -594
rect 1950 -606 1956 -600
rect 1950 -612 1956 -606
rect 1950 -618 1956 -612
rect 1950 -624 1956 -618
rect 1950 -630 1956 -624
rect 1950 -636 1956 -630
rect 1950 -642 1956 -636
rect 1950 -648 1956 -642
rect 1950 -654 1956 -648
rect 1950 -660 1956 -654
rect 1950 -666 1956 -660
rect 1950 -672 1956 -666
rect 1950 -678 1956 -672
rect 1950 -684 1956 -678
rect 1950 -690 1956 -684
rect 1950 -696 1956 -690
rect 1950 -702 1956 -696
rect 1950 -708 1956 -702
rect 1950 -714 1956 -708
rect 1950 -720 1956 -714
rect 1950 -726 1956 -720
rect 1950 -732 1956 -726
rect 1950 -738 1956 -732
rect 1950 -744 1956 -738
rect 1950 -750 1956 -744
rect 1950 -756 1956 -750
rect 1950 -762 1956 -756
rect 1950 -768 1956 -762
rect 1950 -774 1956 -768
rect 1950 -780 1956 -774
rect 1950 -786 1956 -780
rect 1950 -792 1956 -786
rect 1950 -798 1956 -792
rect 1950 -804 1956 -798
rect 1950 -810 1956 -804
rect 1950 -816 1956 -810
rect 1950 -822 1956 -816
rect 1950 -828 1956 -822
rect 1950 -834 1956 -828
rect 1950 -840 1956 -834
rect 1950 -846 1956 -840
rect 1950 -852 1956 -846
rect 1950 -858 1956 -852
rect 1950 -864 1956 -858
rect 1950 -870 1956 -864
rect 1950 -876 1956 -870
rect 1950 -882 1956 -876
rect 1950 -888 1956 -882
rect 1950 -894 1956 -888
rect 1950 -900 1956 -894
rect 1950 -906 1956 -900
rect 1950 -912 1956 -906
rect 1950 -918 1956 -912
rect 1950 -924 1956 -918
rect 1950 -930 1956 -924
rect 1950 -936 1956 -930
rect 1950 -942 1956 -936
rect 1950 -948 1956 -942
rect 1950 -954 1956 -948
rect 1950 -960 1956 -954
rect 1950 -966 1956 -960
rect 1950 -972 1956 -966
rect 1950 -978 1956 -972
rect 1950 -984 1956 -978
rect 1950 -990 1956 -984
rect 1950 -996 1956 -990
rect 1950 -1002 1956 -996
rect 1950 -1008 1956 -1002
rect 1950 -1014 1956 -1008
rect 1950 -1020 1956 -1014
rect 1950 -1026 1956 -1020
rect 1950 -1032 1956 -1026
rect 1950 -1038 1956 -1032
rect 1950 -1044 1956 -1038
rect 1950 -1050 1956 -1044
rect 1950 -1056 1956 -1050
rect 1950 -1062 1956 -1056
rect 1950 -1068 1956 -1062
rect 1950 -1074 1956 -1068
rect 1950 -1080 1956 -1074
rect 1950 -1086 1956 -1080
rect 1950 -1092 1956 -1086
rect 1950 -1098 1956 -1092
rect 1950 -1104 1956 -1098
rect 1950 -1110 1956 -1104
rect 1950 -1116 1956 -1110
rect 1950 -1122 1956 -1116
rect 1950 -1128 1956 -1122
rect 1950 -1134 1956 -1128
rect 1950 -1140 1956 -1134
rect 1950 -1146 1956 -1140
rect 1950 -1152 1956 -1146
rect 1950 -1158 1956 -1152
rect 1950 -1164 1956 -1158
rect 1950 -1170 1956 -1164
rect 1950 -1176 1956 -1170
rect 1950 -1182 1956 -1176
rect 1950 -1188 1956 -1182
rect 1950 -1194 1956 -1188
rect 1950 -1200 1956 -1194
rect 1950 -1206 1956 -1200
rect 1950 -1212 1956 -1206
rect 1950 -1218 1956 -1212
rect 1950 -1224 1956 -1218
rect 1950 -1230 1956 -1224
rect 1950 -1236 1956 -1230
rect 1950 -1242 1956 -1236
rect 1950 -1248 1956 -1242
rect 1950 -1254 1956 -1248
rect 1950 -1260 1956 -1254
rect 1950 -1266 1956 -1260
rect 1950 -1272 1956 -1266
rect 1950 -1278 1956 -1272
rect 1950 -1284 1956 -1278
rect 1950 -1290 1956 -1284
rect 1950 -1296 1956 -1290
rect 1950 -1302 1956 -1296
rect 1950 -1308 1956 -1302
rect 1950 -1314 1956 -1308
rect 1950 -1320 1956 -1314
rect 1950 -1326 1956 -1320
rect 1950 -1332 1956 -1326
rect 1950 -1338 1956 -1332
rect 1950 -1344 1956 -1338
rect 1950 -1350 1956 -1344
rect 1950 -1356 1956 -1350
rect 1950 -1362 1956 -1356
rect 1950 -1368 1956 -1362
rect 1950 -1374 1956 -1368
rect 1950 -1380 1956 -1374
rect 1950 -1386 1956 -1380
rect 1950 -1392 1956 -1386
rect 1950 -1398 1956 -1392
rect 1950 -1404 1956 -1398
rect 1950 -1410 1956 -1404
rect 1950 -1416 1956 -1410
rect 1950 -1422 1956 -1416
rect 1950 -1428 1956 -1422
rect 1950 -1434 1956 -1428
rect 1950 -1440 1956 -1434
rect 1950 -1446 1956 -1440
rect 1950 -1452 1956 -1446
rect 1950 -1458 1956 -1452
rect 1950 -1464 1956 -1458
rect 1950 -1470 1956 -1464
rect 1950 -1476 1956 -1470
rect 1950 -1482 1956 -1476
rect 1950 -1488 1956 -1482
rect 1950 -1494 1956 -1488
rect 1950 -1500 1956 -1494
rect 1950 -1506 1956 -1500
rect 1950 -1512 1956 -1506
rect 1950 -1518 1956 -1512
rect 1950 -1524 1956 -1518
rect 1950 -1530 1956 -1524
rect 1950 -1536 1956 -1530
rect 1950 -1542 1956 -1536
rect 1950 -1548 1956 -1542
rect 1950 -1554 1956 -1548
rect 1950 -1560 1956 -1554
rect 1950 -1566 1956 -1560
rect 1950 -1572 1956 -1566
rect 1950 -1578 1956 -1572
rect 1950 -1584 1956 -1578
rect 1950 -1590 1956 -1584
rect 1950 -1596 1956 -1590
rect 1950 -1602 1956 -1596
rect 1950 -1608 1956 -1602
rect 1950 -1614 1956 -1608
rect 1950 -1620 1956 -1614
rect 1950 -1626 1956 -1620
rect 1950 -1632 1956 -1626
rect 1950 -1638 1956 -1632
rect 1950 -1644 1956 -1638
rect 1950 -1650 1956 -1644
rect 1950 -1656 1956 -1650
rect 1950 -1662 1956 -1656
rect 1950 -1668 1956 -1662
rect 1950 -1674 1956 -1668
rect 1950 -1680 1956 -1674
rect 1950 -1686 1956 -1680
rect 1950 -1692 1956 -1686
rect 1950 -1782 1956 -1776
rect 1950 -1788 1956 -1782
rect 1950 -1794 1956 -1788
rect 1950 -1800 1956 -1794
rect 1950 -1806 1956 -1800
rect 1950 -1812 1956 -1806
rect 1950 -1818 1956 -1812
rect 1950 -1824 1956 -1818
rect 1950 -1830 1956 -1824
rect 1950 -1836 1956 -1830
rect 1950 -1842 1956 -1836
rect 1950 -1848 1956 -1842
rect 1950 -1854 1956 -1848
rect 1950 -1860 1956 -1854
rect 1950 -1866 1956 -1860
rect 1950 -1872 1956 -1866
rect 1950 -1878 1956 -1872
rect 1950 -1884 1956 -1878
rect 1950 -1890 1956 -1884
rect 1950 -1896 1956 -1890
rect 1950 -1902 1956 -1896
rect 1950 -1908 1956 -1902
rect 1950 -1914 1956 -1908
rect 1950 -1920 1956 -1914
rect 1950 -1926 1956 -1920
rect 1950 -1932 1956 -1926
rect 1950 -1938 1956 -1932
rect 1950 -1944 1956 -1938
rect 1950 -1950 1956 -1944
rect 1950 -1956 1956 -1950
rect 1950 -1962 1956 -1956
rect 1950 -1968 1956 -1962
rect 1950 -1974 1956 -1968
rect 1950 -1980 1956 -1974
rect 1950 -1986 1956 -1980
rect 1950 -1992 1956 -1986
rect 1950 -1998 1956 -1992
rect 1950 -2004 1956 -1998
rect 1950 -2010 1956 -2004
rect 1950 -2016 1956 -2010
rect 1950 -2022 1956 -2016
rect 1950 -2028 1956 -2022
rect 1950 -2034 1956 -2028
rect 1950 -2040 1956 -2034
rect 1950 -2046 1956 -2040
rect 1950 -2052 1956 -2046
rect 1950 -2058 1956 -2052
rect 1950 -2064 1956 -2058
rect 1950 -2070 1956 -2064
rect 1950 -2076 1956 -2070
rect 1950 -2082 1956 -2076
rect 1950 -2088 1956 -2082
rect 1950 -2094 1956 -2088
rect 1950 -2100 1956 -2094
rect 1950 -2106 1956 -2100
rect 1950 -2112 1956 -2106
rect 1950 -2118 1956 -2112
rect 1950 -2124 1956 -2118
rect 1950 -2130 1956 -2124
rect 1950 -2136 1956 -2130
rect 1950 -2142 1956 -2136
rect 1950 -2148 1956 -2142
rect 1950 -2154 1956 -2148
rect 1950 -2160 1956 -2154
rect 1950 -2166 1956 -2160
rect 1950 -2172 1956 -2166
rect 1950 -2178 1956 -2172
rect 1950 -2184 1956 -2178
rect 1950 -2190 1956 -2184
rect 1950 -2196 1956 -2190
rect 1950 -2202 1956 -2196
rect 1950 -2208 1956 -2202
rect 1950 -2214 1956 -2208
rect 1950 -2220 1956 -2214
rect 1950 -2226 1956 -2220
rect 1950 -2232 1956 -2226
rect 1950 -2238 1956 -2232
rect 1950 -2244 1956 -2238
rect 1950 -2250 1956 -2244
rect 1950 -2256 1956 -2250
rect 1950 -2262 1956 -2256
rect 1950 -2268 1956 -2262
rect 1950 -2274 1956 -2268
rect 1950 -2280 1956 -2274
rect 1950 -2286 1956 -2280
rect 1950 -2292 1956 -2286
rect 1950 -2298 1956 -2292
rect 1950 -2304 1956 -2298
rect 1950 -2310 1956 -2304
rect 1950 -2316 1956 -2310
rect 1950 -2322 1956 -2316
rect 1950 -2328 1956 -2322
rect 1950 -2334 1956 -2328
rect 1950 -2340 1956 -2334
rect 1950 -2346 1956 -2340
rect 1950 -2352 1956 -2346
rect 1950 -2358 1956 -2352
rect 1950 -2364 1956 -2358
rect 1950 -2370 1956 -2364
rect 1950 -2376 1956 -2370
rect 1950 -2382 1956 -2376
rect 1950 -2388 1956 -2382
rect 1950 -2394 1956 -2388
rect 1950 -2400 1956 -2394
rect 1950 -2406 1956 -2400
rect 1950 -2412 1956 -2406
rect 1950 -2418 1956 -2412
rect 1950 -2424 1956 -2418
rect 1950 -2430 1956 -2424
rect 1950 -2436 1956 -2430
rect 1950 -2442 1956 -2436
rect 1950 -2448 1956 -2442
rect 1950 -2454 1956 -2448
rect 1950 -2460 1956 -2454
rect 1950 -2466 1956 -2460
rect 1950 -2472 1956 -2466
rect 1950 -2478 1956 -2472
rect 1950 -2484 1956 -2478
rect 1950 -2490 1956 -2484
rect 1950 -2496 1956 -2490
rect 1950 -2502 1956 -2496
rect 1950 -2508 1956 -2502
rect 1950 -2514 1956 -2508
rect 1950 -2520 1956 -2514
rect 1950 -2526 1956 -2520
rect 1950 -2532 1956 -2526
rect 1950 -2538 1956 -2532
rect 1950 -2544 1956 -2538
rect 1950 -2550 1956 -2544
rect 1950 -2634 1956 -2628
rect 1950 -2640 1956 -2634
rect 1950 -2646 1956 -2640
rect 1950 -2652 1956 -2646
rect 1950 -2658 1956 -2652
rect 1950 -2664 1956 -2658
rect 1950 -2670 1956 -2664
rect 1950 -2676 1956 -2670
rect 1950 -2682 1956 -2676
rect 1950 -2688 1956 -2682
rect 1950 -2694 1956 -2688
rect 1950 -2700 1956 -2694
rect 1950 -2706 1956 -2700
rect 1950 -2712 1956 -2706
rect 1950 -2718 1956 -2712
rect 1950 -2724 1956 -2718
rect 1950 -2730 1956 -2724
rect 1950 -2736 1956 -2730
rect 1950 -2742 1956 -2736
rect 1950 -2748 1956 -2742
rect 1950 -2754 1956 -2748
rect 1950 -2760 1956 -2754
rect 1950 -2766 1956 -2760
rect 1950 -2772 1956 -2766
rect 1950 -2778 1956 -2772
rect 1950 -2784 1956 -2778
rect 1950 -2790 1956 -2784
rect 1950 -2796 1956 -2790
rect 1950 -2802 1956 -2796
rect 1950 -2808 1956 -2802
rect 1950 -2814 1956 -2808
rect 1950 -2820 1956 -2814
rect 1950 -2826 1956 -2820
rect 1950 -2832 1956 -2826
rect 1950 -2838 1956 -2832
rect 1950 -2844 1956 -2838
rect 1950 -2850 1956 -2844
rect 1950 -2856 1956 -2850
rect 1950 -2862 1956 -2856
rect 1950 -2868 1956 -2862
rect 1950 -2874 1956 -2868
rect 1950 -2880 1956 -2874
rect 1950 -2886 1956 -2880
rect 1950 -2892 1956 -2886
rect 1950 -2898 1956 -2892
rect 1950 -2904 1956 -2898
rect 1950 -2910 1956 -2904
rect 1950 -2916 1956 -2910
rect 1950 -2922 1956 -2916
rect 1950 -2928 1956 -2922
rect 1950 -2934 1956 -2928
rect 1950 -2940 1956 -2934
rect 1950 -2946 1956 -2940
rect 1950 -2952 1956 -2946
rect 1950 -2958 1956 -2952
rect 1950 -2964 1956 -2958
rect 1950 -2970 1956 -2964
rect 1950 -2976 1956 -2970
rect 1950 -2982 1956 -2976
rect 1950 -2988 1956 -2982
rect 1950 -2994 1956 -2988
rect 1950 -3000 1956 -2994
rect 1950 -3006 1956 -3000
rect 1950 -3012 1956 -3006
rect 1950 -3018 1956 -3012
rect 1950 -3024 1956 -3018
rect 1950 -3030 1956 -3024
rect 1950 -3036 1956 -3030
rect 1950 -3042 1956 -3036
rect 1950 -3048 1956 -3042
rect 1950 -3054 1956 -3048
rect 1950 -3060 1956 -3054
rect 1950 -3066 1956 -3060
rect 1950 -3072 1956 -3066
rect 1950 -3078 1956 -3072
rect 1950 -3084 1956 -3078
rect 1950 -3090 1956 -3084
rect 1950 -3096 1956 -3090
rect 1950 -3102 1956 -3096
rect 1950 -3108 1956 -3102
rect 1950 -3114 1956 -3108
rect 1950 -3120 1956 -3114
rect 1950 -3126 1956 -3120
rect 1950 -3180 1956 -3174
rect 1950 -3186 1956 -3180
rect 1950 -3192 1956 -3186
rect 1950 -3198 1956 -3192
rect 1950 -3204 1956 -3198
rect 1950 -3210 1956 -3204
rect 1950 -3216 1956 -3210
rect 1950 -3222 1956 -3216
rect 1950 -3228 1956 -3222
rect 1950 -3234 1956 -3228
rect 1950 -3240 1956 -3234
rect 1950 -3246 1956 -3240
rect 1950 -3252 1956 -3246
rect 1950 -3258 1956 -3252
rect 1950 -3264 1956 -3258
rect 1956 -510 1962 -504
rect 1956 -516 1962 -510
rect 1956 -522 1962 -516
rect 1956 -528 1962 -522
rect 1956 -534 1962 -528
rect 1956 -540 1962 -534
rect 1956 -546 1962 -540
rect 1956 -552 1962 -546
rect 1956 -558 1962 -552
rect 1956 -564 1962 -558
rect 1956 -570 1962 -564
rect 1956 -576 1962 -570
rect 1956 -582 1962 -576
rect 1956 -588 1962 -582
rect 1956 -594 1962 -588
rect 1956 -600 1962 -594
rect 1956 -606 1962 -600
rect 1956 -612 1962 -606
rect 1956 -618 1962 -612
rect 1956 -624 1962 -618
rect 1956 -630 1962 -624
rect 1956 -636 1962 -630
rect 1956 -642 1962 -636
rect 1956 -648 1962 -642
rect 1956 -654 1962 -648
rect 1956 -660 1962 -654
rect 1956 -666 1962 -660
rect 1956 -672 1962 -666
rect 1956 -678 1962 -672
rect 1956 -684 1962 -678
rect 1956 -690 1962 -684
rect 1956 -696 1962 -690
rect 1956 -702 1962 -696
rect 1956 -708 1962 -702
rect 1956 -714 1962 -708
rect 1956 -720 1962 -714
rect 1956 -726 1962 -720
rect 1956 -732 1962 -726
rect 1956 -738 1962 -732
rect 1956 -744 1962 -738
rect 1956 -750 1962 -744
rect 1956 -756 1962 -750
rect 1956 -762 1962 -756
rect 1956 -768 1962 -762
rect 1956 -774 1962 -768
rect 1956 -780 1962 -774
rect 1956 -786 1962 -780
rect 1956 -792 1962 -786
rect 1956 -798 1962 -792
rect 1956 -804 1962 -798
rect 1956 -810 1962 -804
rect 1956 -816 1962 -810
rect 1956 -822 1962 -816
rect 1956 -828 1962 -822
rect 1956 -834 1962 -828
rect 1956 -840 1962 -834
rect 1956 -846 1962 -840
rect 1956 -852 1962 -846
rect 1956 -858 1962 -852
rect 1956 -864 1962 -858
rect 1956 -870 1962 -864
rect 1956 -876 1962 -870
rect 1956 -882 1962 -876
rect 1956 -888 1962 -882
rect 1956 -894 1962 -888
rect 1956 -900 1962 -894
rect 1956 -906 1962 -900
rect 1956 -912 1962 -906
rect 1956 -918 1962 -912
rect 1956 -924 1962 -918
rect 1956 -930 1962 -924
rect 1956 -936 1962 -930
rect 1956 -942 1962 -936
rect 1956 -948 1962 -942
rect 1956 -954 1962 -948
rect 1956 -960 1962 -954
rect 1956 -966 1962 -960
rect 1956 -972 1962 -966
rect 1956 -978 1962 -972
rect 1956 -984 1962 -978
rect 1956 -990 1962 -984
rect 1956 -996 1962 -990
rect 1956 -1002 1962 -996
rect 1956 -1008 1962 -1002
rect 1956 -1014 1962 -1008
rect 1956 -1020 1962 -1014
rect 1956 -1026 1962 -1020
rect 1956 -1032 1962 -1026
rect 1956 -1038 1962 -1032
rect 1956 -1044 1962 -1038
rect 1956 -1050 1962 -1044
rect 1956 -1056 1962 -1050
rect 1956 -1062 1962 -1056
rect 1956 -1068 1962 -1062
rect 1956 -1074 1962 -1068
rect 1956 -1080 1962 -1074
rect 1956 -1086 1962 -1080
rect 1956 -1092 1962 -1086
rect 1956 -1098 1962 -1092
rect 1956 -1104 1962 -1098
rect 1956 -1110 1962 -1104
rect 1956 -1116 1962 -1110
rect 1956 -1122 1962 -1116
rect 1956 -1128 1962 -1122
rect 1956 -1134 1962 -1128
rect 1956 -1140 1962 -1134
rect 1956 -1146 1962 -1140
rect 1956 -1152 1962 -1146
rect 1956 -1158 1962 -1152
rect 1956 -1164 1962 -1158
rect 1956 -1170 1962 -1164
rect 1956 -1176 1962 -1170
rect 1956 -1182 1962 -1176
rect 1956 -1188 1962 -1182
rect 1956 -1194 1962 -1188
rect 1956 -1200 1962 -1194
rect 1956 -1206 1962 -1200
rect 1956 -1212 1962 -1206
rect 1956 -1218 1962 -1212
rect 1956 -1224 1962 -1218
rect 1956 -1230 1962 -1224
rect 1956 -1236 1962 -1230
rect 1956 -1242 1962 -1236
rect 1956 -1248 1962 -1242
rect 1956 -1254 1962 -1248
rect 1956 -1260 1962 -1254
rect 1956 -1266 1962 -1260
rect 1956 -1272 1962 -1266
rect 1956 -1278 1962 -1272
rect 1956 -1284 1962 -1278
rect 1956 -1290 1962 -1284
rect 1956 -1296 1962 -1290
rect 1956 -1302 1962 -1296
rect 1956 -1308 1962 -1302
rect 1956 -1314 1962 -1308
rect 1956 -1320 1962 -1314
rect 1956 -1326 1962 -1320
rect 1956 -1332 1962 -1326
rect 1956 -1338 1962 -1332
rect 1956 -1344 1962 -1338
rect 1956 -1350 1962 -1344
rect 1956 -1356 1962 -1350
rect 1956 -1362 1962 -1356
rect 1956 -1368 1962 -1362
rect 1956 -1374 1962 -1368
rect 1956 -1380 1962 -1374
rect 1956 -1386 1962 -1380
rect 1956 -1392 1962 -1386
rect 1956 -1398 1962 -1392
rect 1956 -1404 1962 -1398
rect 1956 -1410 1962 -1404
rect 1956 -1416 1962 -1410
rect 1956 -1422 1962 -1416
rect 1956 -1428 1962 -1422
rect 1956 -1434 1962 -1428
rect 1956 -1440 1962 -1434
rect 1956 -1446 1962 -1440
rect 1956 -1452 1962 -1446
rect 1956 -1458 1962 -1452
rect 1956 -1464 1962 -1458
rect 1956 -1470 1962 -1464
rect 1956 -1476 1962 -1470
rect 1956 -1482 1962 -1476
rect 1956 -1488 1962 -1482
rect 1956 -1494 1962 -1488
rect 1956 -1500 1962 -1494
rect 1956 -1506 1962 -1500
rect 1956 -1512 1962 -1506
rect 1956 -1518 1962 -1512
rect 1956 -1524 1962 -1518
rect 1956 -1530 1962 -1524
rect 1956 -1536 1962 -1530
rect 1956 -1542 1962 -1536
rect 1956 -1548 1962 -1542
rect 1956 -1554 1962 -1548
rect 1956 -1560 1962 -1554
rect 1956 -1566 1962 -1560
rect 1956 -1572 1962 -1566
rect 1956 -1578 1962 -1572
rect 1956 -1584 1962 -1578
rect 1956 -1590 1962 -1584
rect 1956 -1596 1962 -1590
rect 1956 -1602 1962 -1596
rect 1956 -1608 1962 -1602
rect 1956 -1614 1962 -1608
rect 1956 -1620 1962 -1614
rect 1956 -1626 1962 -1620
rect 1956 -1632 1962 -1626
rect 1956 -1638 1962 -1632
rect 1956 -1644 1962 -1638
rect 1956 -1650 1962 -1644
rect 1956 -1656 1962 -1650
rect 1956 -1662 1962 -1656
rect 1956 -1668 1962 -1662
rect 1956 -1674 1962 -1668
rect 1956 -1680 1962 -1674
rect 1956 -1686 1962 -1680
rect 1956 -1776 1962 -1770
rect 1956 -1782 1962 -1776
rect 1956 -1788 1962 -1782
rect 1956 -1794 1962 -1788
rect 1956 -1800 1962 -1794
rect 1956 -1806 1962 -1800
rect 1956 -1812 1962 -1806
rect 1956 -1818 1962 -1812
rect 1956 -1824 1962 -1818
rect 1956 -1830 1962 -1824
rect 1956 -1836 1962 -1830
rect 1956 -1842 1962 -1836
rect 1956 -1848 1962 -1842
rect 1956 -1854 1962 -1848
rect 1956 -1860 1962 -1854
rect 1956 -1866 1962 -1860
rect 1956 -1872 1962 -1866
rect 1956 -1878 1962 -1872
rect 1956 -1884 1962 -1878
rect 1956 -1890 1962 -1884
rect 1956 -1896 1962 -1890
rect 1956 -1902 1962 -1896
rect 1956 -1908 1962 -1902
rect 1956 -1914 1962 -1908
rect 1956 -1920 1962 -1914
rect 1956 -1926 1962 -1920
rect 1956 -1932 1962 -1926
rect 1956 -1938 1962 -1932
rect 1956 -1944 1962 -1938
rect 1956 -1950 1962 -1944
rect 1956 -1956 1962 -1950
rect 1956 -1962 1962 -1956
rect 1956 -1968 1962 -1962
rect 1956 -1974 1962 -1968
rect 1956 -1980 1962 -1974
rect 1956 -1986 1962 -1980
rect 1956 -1992 1962 -1986
rect 1956 -1998 1962 -1992
rect 1956 -2004 1962 -1998
rect 1956 -2010 1962 -2004
rect 1956 -2016 1962 -2010
rect 1956 -2022 1962 -2016
rect 1956 -2028 1962 -2022
rect 1956 -2034 1962 -2028
rect 1956 -2040 1962 -2034
rect 1956 -2046 1962 -2040
rect 1956 -2052 1962 -2046
rect 1956 -2058 1962 -2052
rect 1956 -2064 1962 -2058
rect 1956 -2070 1962 -2064
rect 1956 -2076 1962 -2070
rect 1956 -2082 1962 -2076
rect 1956 -2088 1962 -2082
rect 1956 -2094 1962 -2088
rect 1956 -2100 1962 -2094
rect 1956 -2106 1962 -2100
rect 1956 -2112 1962 -2106
rect 1956 -2118 1962 -2112
rect 1956 -2124 1962 -2118
rect 1956 -2130 1962 -2124
rect 1956 -2136 1962 -2130
rect 1956 -2142 1962 -2136
rect 1956 -2148 1962 -2142
rect 1956 -2154 1962 -2148
rect 1956 -2160 1962 -2154
rect 1956 -2166 1962 -2160
rect 1956 -2172 1962 -2166
rect 1956 -2178 1962 -2172
rect 1956 -2184 1962 -2178
rect 1956 -2190 1962 -2184
rect 1956 -2196 1962 -2190
rect 1956 -2202 1962 -2196
rect 1956 -2208 1962 -2202
rect 1956 -2214 1962 -2208
rect 1956 -2220 1962 -2214
rect 1956 -2226 1962 -2220
rect 1956 -2232 1962 -2226
rect 1956 -2238 1962 -2232
rect 1956 -2244 1962 -2238
rect 1956 -2250 1962 -2244
rect 1956 -2256 1962 -2250
rect 1956 -2262 1962 -2256
rect 1956 -2268 1962 -2262
rect 1956 -2274 1962 -2268
rect 1956 -2280 1962 -2274
rect 1956 -2286 1962 -2280
rect 1956 -2292 1962 -2286
rect 1956 -2298 1962 -2292
rect 1956 -2304 1962 -2298
rect 1956 -2310 1962 -2304
rect 1956 -2316 1962 -2310
rect 1956 -2322 1962 -2316
rect 1956 -2328 1962 -2322
rect 1956 -2334 1962 -2328
rect 1956 -2340 1962 -2334
rect 1956 -2346 1962 -2340
rect 1956 -2352 1962 -2346
rect 1956 -2358 1962 -2352
rect 1956 -2364 1962 -2358
rect 1956 -2370 1962 -2364
rect 1956 -2376 1962 -2370
rect 1956 -2382 1962 -2376
rect 1956 -2388 1962 -2382
rect 1956 -2394 1962 -2388
rect 1956 -2400 1962 -2394
rect 1956 -2406 1962 -2400
rect 1956 -2412 1962 -2406
rect 1956 -2418 1962 -2412
rect 1956 -2424 1962 -2418
rect 1956 -2430 1962 -2424
rect 1956 -2436 1962 -2430
rect 1956 -2442 1962 -2436
rect 1956 -2448 1962 -2442
rect 1956 -2454 1962 -2448
rect 1956 -2460 1962 -2454
rect 1956 -2466 1962 -2460
rect 1956 -2472 1962 -2466
rect 1956 -2478 1962 -2472
rect 1956 -2484 1962 -2478
rect 1956 -2490 1962 -2484
rect 1956 -2496 1962 -2490
rect 1956 -2502 1962 -2496
rect 1956 -2508 1962 -2502
rect 1956 -2514 1962 -2508
rect 1956 -2520 1962 -2514
rect 1956 -2526 1962 -2520
rect 1956 -2532 1962 -2526
rect 1956 -2538 1962 -2532
rect 1956 -2544 1962 -2538
rect 1956 -2550 1962 -2544
rect 1956 -2628 1962 -2622
rect 1956 -2634 1962 -2628
rect 1956 -2640 1962 -2634
rect 1956 -2646 1962 -2640
rect 1956 -2652 1962 -2646
rect 1956 -2658 1962 -2652
rect 1956 -2664 1962 -2658
rect 1956 -2670 1962 -2664
rect 1956 -2676 1962 -2670
rect 1956 -2682 1962 -2676
rect 1956 -2688 1962 -2682
rect 1956 -2694 1962 -2688
rect 1956 -2700 1962 -2694
rect 1956 -2706 1962 -2700
rect 1956 -2712 1962 -2706
rect 1956 -2718 1962 -2712
rect 1956 -2724 1962 -2718
rect 1956 -2730 1962 -2724
rect 1956 -2736 1962 -2730
rect 1956 -2742 1962 -2736
rect 1956 -2748 1962 -2742
rect 1956 -2754 1962 -2748
rect 1956 -2760 1962 -2754
rect 1956 -2766 1962 -2760
rect 1956 -2772 1962 -2766
rect 1956 -2778 1962 -2772
rect 1956 -2784 1962 -2778
rect 1956 -2790 1962 -2784
rect 1956 -2796 1962 -2790
rect 1956 -2802 1962 -2796
rect 1956 -2808 1962 -2802
rect 1956 -2814 1962 -2808
rect 1956 -2820 1962 -2814
rect 1956 -2826 1962 -2820
rect 1956 -2832 1962 -2826
rect 1956 -2838 1962 -2832
rect 1956 -2844 1962 -2838
rect 1956 -2850 1962 -2844
rect 1956 -2856 1962 -2850
rect 1956 -2862 1962 -2856
rect 1956 -2868 1962 -2862
rect 1956 -2874 1962 -2868
rect 1956 -2880 1962 -2874
rect 1956 -2886 1962 -2880
rect 1956 -2892 1962 -2886
rect 1956 -2898 1962 -2892
rect 1956 -2904 1962 -2898
rect 1956 -2910 1962 -2904
rect 1956 -2916 1962 -2910
rect 1956 -2922 1962 -2916
rect 1956 -2928 1962 -2922
rect 1956 -2934 1962 -2928
rect 1956 -2940 1962 -2934
rect 1956 -2946 1962 -2940
rect 1956 -2952 1962 -2946
rect 1956 -2958 1962 -2952
rect 1956 -2964 1962 -2958
rect 1956 -2970 1962 -2964
rect 1956 -2976 1962 -2970
rect 1956 -2982 1962 -2976
rect 1956 -2988 1962 -2982
rect 1956 -2994 1962 -2988
rect 1956 -3000 1962 -2994
rect 1956 -3006 1962 -3000
rect 1956 -3012 1962 -3006
rect 1956 -3018 1962 -3012
rect 1956 -3024 1962 -3018
rect 1956 -3030 1962 -3024
rect 1956 -3036 1962 -3030
rect 1956 -3042 1962 -3036
rect 1956 -3048 1962 -3042
rect 1956 -3054 1962 -3048
rect 1956 -3060 1962 -3054
rect 1956 -3066 1962 -3060
rect 1956 -3072 1962 -3066
rect 1956 -3078 1962 -3072
rect 1956 -3084 1962 -3078
rect 1956 -3090 1962 -3084
rect 1956 -3096 1962 -3090
rect 1956 -3102 1962 -3096
rect 1956 -3108 1962 -3102
rect 1956 -3114 1962 -3108
rect 1956 -3120 1962 -3114
rect 1956 -3174 1962 -3168
rect 1956 -3180 1962 -3174
rect 1956 -3186 1962 -3180
rect 1956 -3192 1962 -3186
rect 1956 -3198 1962 -3192
rect 1956 -3204 1962 -3198
rect 1956 -3210 1962 -3204
rect 1956 -3216 1962 -3210
rect 1956 -3222 1962 -3216
rect 1956 -3228 1962 -3222
rect 1956 -3234 1962 -3228
rect 1956 -3240 1962 -3234
rect 1956 -3246 1962 -3240
rect 1956 -3252 1962 -3246
rect 1956 -3258 1962 -3252
rect 1962 -498 1968 -492
rect 1962 -504 1968 -498
rect 1962 -510 1968 -504
rect 1962 -516 1968 -510
rect 1962 -522 1968 -516
rect 1962 -528 1968 -522
rect 1962 -534 1968 -528
rect 1962 -540 1968 -534
rect 1962 -546 1968 -540
rect 1962 -552 1968 -546
rect 1962 -558 1968 -552
rect 1962 -564 1968 -558
rect 1962 -570 1968 -564
rect 1962 -576 1968 -570
rect 1962 -582 1968 -576
rect 1962 -588 1968 -582
rect 1962 -594 1968 -588
rect 1962 -600 1968 -594
rect 1962 -606 1968 -600
rect 1962 -612 1968 -606
rect 1962 -618 1968 -612
rect 1962 -624 1968 -618
rect 1962 -630 1968 -624
rect 1962 -636 1968 -630
rect 1962 -642 1968 -636
rect 1962 -648 1968 -642
rect 1962 -654 1968 -648
rect 1962 -660 1968 -654
rect 1962 -666 1968 -660
rect 1962 -672 1968 -666
rect 1962 -678 1968 -672
rect 1962 -684 1968 -678
rect 1962 -690 1968 -684
rect 1962 -696 1968 -690
rect 1962 -702 1968 -696
rect 1962 -708 1968 -702
rect 1962 -714 1968 -708
rect 1962 -720 1968 -714
rect 1962 -726 1968 -720
rect 1962 -732 1968 -726
rect 1962 -738 1968 -732
rect 1962 -744 1968 -738
rect 1962 -750 1968 -744
rect 1962 -756 1968 -750
rect 1962 -762 1968 -756
rect 1962 -768 1968 -762
rect 1962 -774 1968 -768
rect 1962 -780 1968 -774
rect 1962 -786 1968 -780
rect 1962 -792 1968 -786
rect 1962 -798 1968 -792
rect 1962 -804 1968 -798
rect 1962 -810 1968 -804
rect 1962 -816 1968 -810
rect 1962 -822 1968 -816
rect 1962 -828 1968 -822
rect 1962 -834 1968 -828
rect 1962 -840 1968 -834
rect 1962 -846 1968 -840
rect 1962 -852 1968 -846
rect 1962 -858 1968 -852
rect 1962 -864 1968 -858
rect 1962 -870 1968 -864
rect 1962 -876 1968 -870
rect 1962 -882 1968 -876
rect 1962 -888 1968 -882
rect 1962 -894 1968 -888
rect 1962 -900 1968 -894
rect 1962 -906 1968 -900
rect 1962 -912 1968 -906
rect 1962 -918 1968 -912
rect 1962 -924 1968 -918
rect 1962 -930 1968 -924
rect 1962 -936 1968 -930
rect 1962 -942 1968 -936
rect 1962 -948 1968 -942
rect 1962 -954 1968 -948
rect 1962 -960 1968 -954
rect 1962 -966 1968 -960
rect 1962 -972 1968 -966
rect 1962 -978 1968 -972
rect 1962 -984 1968 -978
rect 1962 -990 1968 -984
rect 1962 -996 1968 -990
rect 1962 -1002 1968 -996
rect 1962 -1008 1968 -1002
rect 1962 -1014 1968 -1008
rect 1962 -1020 1968 -1014
rect 1962 -1026 1968 -1020
rect 1962 -1032 1968 -1026
rect 1962 -1038 1968 -1032
rect 1962 -1044 1968 -1038
rect 1962 -1050 1968 -1044
rect 1962 -1056 1968 -1050
rect 1962 -1062 1968 -1056
rect 1962 -1068 1968 -1062
rect 1962 -1074 1968 -1068
rect 1962 -1080 1968 -1074
rect 1962 -1086 1968 -1080
rect 1962 -1092 1968 -1086
rect 1962 -1098 1968 -1092
rect 1962 -1104 1968 -1098
rect 1962 -1110 1968 -1104
rect 1962 -1116 1968 -1110
rect 1962 -1122 1968 -1116
rect 1962 -1128 1968 -1122
rect 1962 -1134 1968 -1128
rect 1962 -1140 1968 -1134
rect 1962 -1146 1968 -1140
rect 1962 -1152 1968 -1146
rect 1962 -1158 1968 -1152
rect 1962 -1164 1968 -1158
rect 1962 -1170 1968 -1164
rect 1962 -1176 1968 -1170
rect 1962 -1182 1968 -1176
rect 1962 -1188 1968 -1182
rect 1962 -1194 1968 -1188
rect 1962 -1200 1968 -1194
rect 1962 -1206 1968 -1200
rect 1962 -1212 1968 -1206
rect 1962 -1218 1968 -1212
rect 1962 -1224 1968 -1218
rect 1962 -1230 1968 -1224
rect 1962 -1236 1968 -1230
rect 1962 -1242 1968 -1236
rect 1962 -1248 1968 -1242
rect 1962 -1254 1968 -1248
rect 1962 -1260 1968 -1254
rect 1962 -1266 1968 -1260
rect 1962 -1272 1968 -1266
rect 1962 -1278 1968 -1272
rect 1962 -1284 1968 -1278
rect 1962 -1290 1968 -1284
rect 1962 -1296 1968 -1290
rect 1962 -1302 1968 -1296
rect 1962 -1308 1968 -1302
rect 1962 -1314 1968 -1308
rect 1962 -1320 1968 -1314
rect 1962 -1326 1968 -1320
rect 1962 -1332 1968 -1326
rect 1962 -1338 1968 -1332
rect 1962 -1344 1968 -1338
rect 1962 -1350 1968 -1344
rect 1962 -1356 1968 -1350
rect 1962 -1362 1968 -1356
rect 1962 -1368 1968 -1362
rect 1962 -1374 1968 -1368
rect 1962 -1380 1968 -1374
rect 1962 -1386 1968 -1380
rect 1962 -1392 1968 -1386
rect 1962 -1398 1968 -1392
rect 1962 -1404 1968 -1398
rect 1962 -1410 1968 -1404
rect 1962 -1416 1968 -1410
rect 1962 -1422 1968 -1416
rect 1962 -1428 1968 -1422
rect 1962 -1434 1968 -1428
rect 1962 -1440 1968 -1434
rect 1962 -1446 1968 -1440
rect 1962 -1452 1968 -1446
rect 1962 -1458 1968 -1452
rect 1962 -1464 1968 -1458
rect 1962 -1470 1968 -1464
rect 1962 -1476 1968 -1470
rect 1962 -1482 1968 -1476
rect 1962 -1488 1968 -1482
rect 1962 -1494 1968 -1488
rect 1962 -1500 1968 -1494
rect 1962 -1506 1968 -1500
rect 1962 -1512 1968 -1506
rect 1962 -1518 1968 -1512
rect 1962 -1524 1968 -1518
rect 1962 -1530 1968 -1524
rect 1962 -1536 1968 -1530
rect 1962 -1542 1968 -1536
rect 1962 -1548 1968 -1542
rect 1962 -1554 1968 -1548
rect 1962 -1560 1968 -1554
rect 1962 -1566 1968 -1560
rect 1962 -1572 1968 -1566
rect 1962 -1578 1968 -1572
rect 1962 -1584 1968 -1578
rect 1962 -1590 1968 -1584
rect 1962 -1596 1968 -1590
rect 1962 -1602 1968 -1596
rect 1962 -1608 1968 -1602
rect 1962 -1614 1968 -1608
rect 1962 -1620 1968 -1614
rect 1962 -1626 1968 -1620
rect 1962 -1632 1968 -1626
rect 1962 -1638 1968 -1632
rect 1962 -1644 1968 -1638
rect 1962 -1650 1968 -1644
rect 1962 -1656 1968 -1650
rect 1962 -1662 1968 -1656
rect 1962 -1668 1968 -1662
rect 1962 -1674 1968 -1668
rect 1962 -1680 1968 -1674
rect 1962 -1770 1968 -1764
rect 1962 -1776 1968 -1770
rect 1962 -1782 1968 -1776
rect 1962 -1788 1968 -1782
rect 1962 -1794 1968 -1788
rect 1962 -1800 1968 -1794
rect 1962 -1806 1968 -1800
rect 1962 -1812 1968 -1806
rect 1962 -1818 1968 -1812
rect 1962 -1824 1968 -1818
rect 1962 -1830 1968 -1824
rect 1962 -1836 1968 -1830
rect 1962 -1842 1968 -1836
rect 1962 -1848 1968 -1842
rect 1962 -1854 1968 -1848
rect 1962 -1860 1968 -1854
rect 1962 -1866 1968 -1860
rect 1962 -1872 1968 -1866
rect 1962 -1878 1968 -1872
rect 1962 -1884 1968 -1878
rect 1962 -1890 1968 -1884
rect 1962 -1896 1968 -1890
rect 1962 -1902 1968 -1896
rect 1962 -1908 1968 -1902
rect 1962 -1914 1968 -1908
rect 1962 -1920 1968 -1914
rect 1962 -1926 1968 -1920
rect 1962 -1932 1968 -1926
rect 1962 -1938 1968 -1932
rect 1962 -1944 1968 -1938
rect 1962 -1950 1968 -1944
rect 1962 -1956 1968 -1950
rect 1962 -1962 1968 -1956
rect 1962 -1968 1968 -1962
rect 1962 -1974 1968 -1968
rect 1962 -1980 1968 -1974
rect 1962 -1986 1968 -1980
rect 1962 -1992 1968 -1986
rect 1962 -1998 1968 -1992
rect 1962 -2004 1968 -1998
rect 1962 -2010 1968 -2004
rect 1962 -2016 1968 -2010
rect 1962 -2022 1968 -2016
rect 1962 -2028 1968 -2022
rect 1962 -2034 1968 -2028
rect 1962 -2040 1968 -2034
rect 1962 -2046 1968 -2040
rect 1962 -2052 1968 -2046
rect 1962 -2058 1968 -2052
rect 1962 -2064 1968 -2058
rect 1962 -2070 1968 -2064
rect 1962 -2076 1968 -2070
rect 1962 -2082 1968 -2076
rect 1962 -2088 1968 -2082
rect 1962 -2094 1968 -2088
rect 1962 -2100 1968 -2094
rect 1962 -2106 1968 -2100
rect 1962 -2112 1968 -2106
rect 1962 -2118 1968 -2112
rect 1962 -2124 1968 -2118
rect 1962 -2130 1968 -2124
rect 1962 -2136 1968 -2130
rect 1962 -2142 1968 -2136
rect 1962 -2148 1968 -2142
rect 1962 -2154 1968 -2148
rect 1962 -2160 1968 -2154
rect 1962 -2166 1968 -2160
rect 1962 -2172 1968 -2166
rect 1962 -2178 1968 -2172
rect 1962 -2184 1968 -2178
rect 1962 -2190 1968 -2184
rect 1962 -2196 1968 -2190
rect 1962 -2202 1968 -2196
rect 1962 -2208 1968 -2202
rect 1962 -2214 1968 -2208
rect 1962 -2220 1968 -2214
rect 1962 -2226 1968 -2220
rect 1962 -2232 1968 -2226
rect 1962 -2238 1968 -2232
rect 1962 -2244 1968 -2238
rect 1962 -2250 1968 -2244
rect 1962 -2256 1968 -2250
rect 1962 -2262 1968 -2256
rect 1962 -2268 1968 -2262
rect 1962 -2274 1968 -2268
rect 1962 -2280 1968 -2274
rect 1962 -2286 1968 -2280
rect 1962 -2292 1968 -2286
rect 1962 -2298 1968 -2292
rect 1962 -2304 1968 -2298
rect 1962 -2310 1968 -2304
rect 1962 -2316 1968 -2310
rect 1962 -2322 1968 -2316
rect 1962 -2328 1968 -2322
rect 1962 -2334 1968 -2328
rect 1962 -2340 1968 -2334
rect 1962 -2346 1968 -2340
rect 1962 -2352 1968 -2346
rect 1962 -2358 1968 -2352
rect 1962 -2364 1968 -2358
rect 1962 -2370 1968 -2364
rect 1962 -2376 1968 -2370
rect 1962 -2382 1968 -2376
rect 1962 -2388 1968 -2382
rect 1962 -2394 1968 -2388
rect 1962 -2400 1968 -2394
rect 1962 -2406 1968 -2400
rect 1962 -2412 1968 -2406
rect 1962 -2418 1968 -2412
rect 1962 -2424 1968 -2418
rect 1962 -2430 1968 -2424
rect 1962 -2436 1968 -2430
rect 1962 -2442 1968 -2436
rect 1962 -2448 1968 -2442
rect 1962 -2454 1968 -2448
rect 1962 -2460 1968 -2454
rect 1962 -2466 1968 -2460
rect 1962 -2472 1968 -2466
rect 1962 -2478 1968 -2472
rect 1962 -2484 1968 -2478
rect 1962 -2490 1968 -2484
rect 1962 -2496 1968 -2490
rect 1962 -2502 1968 -2496
rect 1962 -2508 1968 -2502
rect 1962 -2514 1968 -2508
rect 1962 -2520 1968 -2514
rect 1962 -2526 1968 -2520
rect 1962 -2532 1968 -2526
rect 1962 -2538 1968 -2532
rect 1962 -2544 1968 -2538
rect 1962 -2628 1968 -2622
rect 1962 -2634 1968 -2628
rect 1962 -2640 1968 -2634
rect 1962 -2646 1968 -2640
rect 1962 -2652 1968 -2646
rect 1962 -2658 1968 -2652
rect 1962 -2664 1968 -2658
rect 1962 -2670 1968 -2664
rect 1962 -2676 1968 -2670
rect 1962 -2682 1968 -2676
rect 1962 -2688 1968 -2682
rect 1962 -2694 1968 -2688
rect 1962 -2700 1968 -2694
rect 1962 -2706 1968 -2700
rect 1962 -2712 1968 -2706
rect 1962 -2718 1968 -2712
rect 1962 -2724 1968 -2718
rect 1962 -2730 1968 -2724
rect 1962 -2736 1968 -2730
rect 1962 -2742 1968 -2736
rect 1962 -2748 1968 -2742
rect 1962 -2754 1968 -2748
rect 1962 -2760 1968 -2754
rect 1962 -2766 1968 -2760
rect 1962 -2772 1968 -2766
rect 1962 -2778 1968 -2772
rect 1962 -2784 1968 -2778
rect 1962 -2790 1968 -2784
rect 1962 -2796 1968 -2790
rect 1962 -2802 1968 -2796
rect 1962 -2808 1968 -2802
rect 1962 -2814 1968 -2808
rect 1962 -2820 1968 -2814
rect 1962 -2826 1968 -2820
rect 1962 -2832 1968 -2826
rect 1962 -2838 1968 -2832
rect 1962 -2844 1968 -2838
rect 1962 -2850 1968 -2844
rect 1962 -2856 1968 -2850
rect 1962 -2862 1968 -2856
rect 1962 -2868 1968 -2862
rect 1962 -2874 1968 -2868
rect 1962 -2880 1968 -2874
rect 1962 -2886 1968 -2880
rect 1962 -2892 1968 -2886
rect 1962 -2898 1968 -2892
rect 1962 -2904 1968 -2898
rect 1962 -2910 1968 -2904
rect 1962 -2916 1968 -2910
rect 1962 -2922 1968 -2916
rect 1962 -2928 1968 -2922
rect 1962 -2934 1968 -2928
rect 1962 -2940 1968 -2934
rect 1962 -2946 1968 -2940
rect 1962 -2952 1968 -2946
rect 1962 -2958 1968 -2952
rect 1962 -2964 1968 -2958
rect 1962 -2970 1968 -2964
rect 1962 -2976 1968 -2970
rect 1962 -2982 1968 -2976
rect 1962 -2988 1968 -2982
rect 1962 -2994 1968 -2988
rect 1962 -3000 1968 -2994
rect 1962 -3006 1968 -3000
rect 1962 -3012 1968 -3006
rect 1962 -3018 1968 -3012
rect 1962 -3024 1968 -3018
rect 1962 -3030 1968 -3024
rect 1962 -3036 1968 -3030
rect 1962 -3042 1968 -3036
rect 1962 -3048 1968 -3042
rect 1962 -3054 1968 -3048
rect 1962 -3060 1968 -3054
rect 1962 -3066 1968 -3060
rect 1962 -3072 1968 -3066
rect 1962 -3078 1968 -3072
rect 1962 -3084 1968 -3078
rect 1962 -3090 1968 -3084
rect 1962 -3096 1968 -3090
rect 1962 -3102 1968 -3096
rect 1962 -3108 1968 -3102
rect 1962 -3114 1968 -3108
rect 1962 -3120 1968 -3114
rect 1962 -3174 1968 -3168
rect 1962 -3180 1968 -3174
rect 1962 -3186 1968 -3180
rect 1962 -3192 1968 -3186
rect 1962 -3198 1968 -3192
rect 1962 -3204 1968 -3198
rect 1962 -3210 1968 -3204
rect 1962 -3216 1968 -3210
rect 1962 -3222 1968 -3216
rect 1962 -3228 1968 -3222
rect 1962 -3234 1968 -3228
rect 1962 -3240 1968 -3234
rect 1962 -3246 1968 -3240
rect 1962 -3252 1968 -3246
rect 1968 -492 1974 -486
rect 1968 -498 1974 -492
rect 1968 -504 1974 -498
rect 1968 -510 1974 -504
rect 1968 -516 1974 -510
rect 1968 -522 1974 -516
rect 1968 -528 1974 -522
rect 1968 -534 1974 -528
rect 1968 -540 1974 -534
rect 1968 -546 1974 -540
rect 1968 -552 1974 -546
rect 1968 -558 1974 -552
rect 1968 -564 1974 -558
rect 1968 -570 1974 -564
rect 1968 -576 1974 -570
rect 1968 -582 1974 -576
rect 1968 -588 1974 -582
rect 1968 -594 1974 -588
rect 1968 -600 1974 -594
rect 1968 -606 1974 -600
rect 1968 -612 1974 -606
rect 1968 -618 1974 -612
rect 1968 -624 1974 -618
rect 1968 -630 1974 -624
rect 1968 -636 1974 -630
rect 1968 -642 1974 -636
rect 1968 -648 1974 -642
rect 1968 -654 1974 -648
rect 1968 -660 1974 -654
rect 1968 -666 1974 -660
rect 1968 -672 1974 -666
rect 1968 -678 1974 -672
rect 1968 -684 1974 -678
rect 1968 -690 1974 -684
rect 1968 -696 1974 -690
rect 1968 -702 1974 -696
rect 1968 -708 1974 -702
rect 1968 -714 1974 -708
rect 1968 -720 1974 -714
rect 1968 -726 1974 -720
rect 1968 -732 1974 -726
rect 1968 -738 1974 -732
rect 1968 -744 1974 -738
rect 1968 -750 1974 -744
rect 1968 -756 1974 -750
rect 1968 -762 1974 -756
rect 1968 -768 1974 -762
rect 1968 -774 1974 -768
rect 1968 -780 1974 -774
rect 1968 -786 1974 -780
rect 1968 -792 1974 -786
rect 1968 -798 1974 -792
rect 1968 -804 1974 -798
rect 1968 -810 1974 -804
rect 1968 -816 1974 -810
rect 1968 -822 1974 -816
rect 1968 -828 1974 -822
rect 1968 -834 1974 -828
rect 1968 -840 1974 -834
rect 1968 -846 1974 -840
rect 1968 -852 1974 -846
rect 1968 -858 1974 -852
rect 1968 -864 1974 -858
rect 1968 -870 1974 -864
rect 1968 -876 1974 -870
rect 1968 -882 1974 -876
rect 1968 -888 1974 -882
rect 1968 -894 1974 -888
rect 1968 -900 1974 -894
rect 1968 -906 1974 -900
rect 1968 -912 1974 -906
rect 1968 -918 1974 -912
rect 1968 -924 1974 -918
rect 1968 -930 1974 -924
rect 1968 -936 1974 -930
rect 1968 -942 1974 -936
rect 1968 -948 1974 -942
rect 1968 -954 1974 -948
rect 1968 -960 1974 -954
rect 1968 -966 1974 -960
rect 1968 -972 1974 -966
rect 1968 -978 1974 -972
rect 1968 -984 1974 -978
rect 1968 -990 1974 -984
rect 1968 -996 1974 -990
rect 1968 -1002 1974 -996
rect 1968 -1008 1974 -1002
rect 1968 -1014 1974 -1008
rect 1968 -1020 1974 -1014
rect 1968 -1026 1974 -1020
rect 1968 -1032 1974 -1026
rect 1968 -1038 1974 -1032
rect 1968 -1044 1974 -1038
rect 1968 -1050 1974 -1044
rect 1968 -1056 1974 -1050
rect 1968 -1062 1974 -1056
rect 1968 -1068 1974 -1062
rect 1968 -1074 1974 -1068
rect 1968 -1080 1974 -1074
rect 1968 -1086 1974 -1080
rect 1968 -1092 1974 -1086
rect 1968 -1098 1974 -1092
rect 1968 -1104 1974 -1098
rect 1968 -1110 1974 -1104
rect 1968 -1116 1974 -1110
rect 1968 -1122 1974 -1116
rect 1968 -1128 1974 -1122
rect 1968 -1134 1974 -1128
rect 1968 -1140 1974 -1134
rect 1968 -1146 1974 -1140
rect 1968 -1152 1974 -1146
rect 1968 -1158 1974 -1152
rect 1968 -1164 1974 -1158
rect 1968 -1170 1974 -1164
rect 1968 -1176 1974 -1170
rect 1968 -1182 1974 -1176
rect 1968 -1188 1974 -1182
rect 1968 -1194 1974 -1188
rect 1968 -1200 1974 -1194
rect 1968 -1206 1974 -1200
rect 1968 -1212 1974 -1206
rect 1968 -1218 1974 -1212
rect 1968 -1224 1974 -1218
rect 1968 -1230 1974 -1224
rect 1968 -1236 1974 -1230
rect 1968 -1242 1974 -1236
rect 1968 -1248 1974 -1242
rect 1968 -1254 1974 -1248
rect 1968 -1260 1974 -1254
rect 1968 -1266 1974 -1260
rect 1968 -1272 1974 -1266
rect 1968 -1278 1974 -1272
rect 1968 -1284 1974 -1278
rect 1968 -1290 1974 -1284
rect 1968 -1296 1974 -1290
rect 1968 -1302 1974 -1296
rect 1968 -1308 1974 -1302
rect 1968 -1314 1974 -1308
rect 1968 -1320 1974 -1314
rect 1968 -1326 1974 -1320
rect 1968 -1332 1974 -1326
rect 1968 -1338 1974 -1332
rect 1968 -1344 1974 -1338
rect 1968 -1350 1974 -1344
rect 1968 -1356 1974 -1350
rect 1968 -1362 1974 -1356
rect 1968 -1368 1974 -1362
rect 1968 -1374 1974 -1368
rect 1968 -1380 1974 -1374
rect 1968 -1386 1974 -1380
rect 1968 -1392 1974 -1386
rect 1968 -1398 1974 -1392
rect 1968 -1404 1974 -1398
rect 1968 -1410 1974 -1404
rect 1968 -1416 1974 -1410
rect 1968 -1422 1974 -1416
rect 1968 -1428 1974 -1422
rect 1968 -1434 1974 -1428
rect 1968 -1440 1974 -1434
rect 1968 -1446 1974 -1440
rect 1968 -1452 1974 -1446
rect 1968 -1458 1974 -1452
rect 1968 -1464 1974 -1458
rect 1968 -1470 1974 -1464
rect 1968 -1476 1974 -1470
rect 1968 -1482 1974 -1476
rect 1968 -1488 1974 -1482
rect 1968 -1494 1974 -1488
rect 1968 -1500 1974 -1494
rect 1968 -1506 1974 -1500
rect 1968 -1512 1974 -1506
rect 1968 -1518 1974 -1512
rect 1968 -1524 1974 -1518
rect 1968 -1530 1974 -1524
rect 1968 -1536 1974 -1530
rect 1968 -1542 1974 -1536
rect 1968 -1548 1974 -1542
rect 1968 -1554 1974 -1548
rect 1968 -1560 1974 -1554
rect 1968 -1566 1974 -1560
rect 1968 -1572 1974 -1566
rect 1968 -1578 1974 -1572
rect 1968 -1584 1974 -1578
rect 1968 -1590 1974 -1584
rect 1968 -1596 1974 -1590
rect 1968 -1602 1974 -1596
rect 1968 -1608 1974 -1602
rect 1968 -1614 1974 -1608
rect 1968 -1620 1974 -1614
rect 1968 -1626 1974 -1620
rect 1968 -1632 1974 -1626
rect 1968 -1638 1974 -1632
rect 1968 -1644 1974 -1638
rect 1968 -1650 1974 -1644
rect 1968 -1656 1974 -1650
rect 1968 -1662 1974 -1656
rect 1968 -1668 1974 -1662
rect 1968 -1674 1974 -1668
rect 1968 -1764 1974 -1758
rect 1968 -1770 1974 -1764
rect 1968 -1776 1974 -1770
rect 1968 -1782 1974 -1776
rect 1968 -1788 1974 -1782
rect 1968 -1794 1974 -1788
rect 1968 -1800 1974 -1794
rect 1968 -1806 1974 -1800
rect 1968 -1812 1974 -1806
rect 1968 -1818 1974 -1812
rect 1968 -1824 1974 -1818
rect 1968 -1830 1974 -1824
rect 1968 -1836 1974 -1830
rect 1968 -1842 1974 -1836
rect 1968 -1848 1974 -1842
rect 1968 -1854 1974 -1848
rect 1968 -1860 1974 -1854
rect 1968 -1866 1974 -1860
rect 1968 -1872 1974 -1866
rect 1968 -1878 1974 -1872
rect 1968 -1884 1974 -1878
rect 1968 -1890 1974 -1884
rect 1968 -1896 1974 -1890
rect 1968 -1902 1974 -1896
rect 1968 -1908 1974 -1902
rect 1968 -1914 1974 -1908
rect 1968 -1920 1974 -1914
rect 1968 -1926 1974 -1920
rect 1968 -1932 1974 -1926
rect 1968 -1938 1974 -1932
rect 1968 -1944 1974 -1938
rect 1968 -1950 1974 -1944
rect 1968 -1956 1974 -1950
rect 1968 -1962 1974 -1956
rect 1968 -1968 1974 -1962
rect 1968 -1974 1974 -1968
rect 1968 -1980 1974 -1974
rect 1968 -1986 1974 -1980
rect 1968 -1992 1974 -1986
rect 1968 -1998 1974 -1992
rect 1968 -2004 1974 -1998
rect 1968 -2010 1974 -2004
rect 1968 -2016 1974 -2010
rect 1968 -2022 1974 -2016
rect 1968 -2028 1974 -2022
rect 1968 -2034 1974 -2028
rect 1968 -2040 1974 -2034
rect 1968 -2046 1974 -2040
rect 1968 -2052 1974 -2046
rect 1968 -2058 1974 -2052
rect 1968 -2064 1974 -2058
rect 1968 -2070 1974 -2064
rect 1968 -2076 1974 -2070
rect 1968 -2082 1974 -2076
rect 1968 -2088 1974 -2082
rect 1968 -2094 1974 -2088
rect 1968 -2100 1974 -2094
rect 1968 -2106 1974 -2100
rect 1968 -2112 1974 -2106
rect 1968 -2118 1974 -2112
rect 1968 -2124 1974 -2118
rect 1968 -2130 1974 -2124
rect 1968 -2136 1974 -2130
rect 1968 -2142 1974 -2136
rect 1968 -2148 1974 -2142
rect 1968 -2154 1974 -2148
rect 1968 -2160 1974 -2154
rect 1968 -2166 1974 -2160
rect 1968 -2172 1974 -2166
rect 1968 -2178 1974 -2172
rect 1968 -2184 1974 -2178
rect 1968 -2190 1974 -2184
rect 1968 -2196 1974 -2190
rect 1968 -2202 1974 -2196
rect 1968 -2208 1974 -2202
rect 1968 -2214 1974 -2208
rect 1968 -2220 1974 -2214
rect 1968 -2226 1974 -2220
rect 1968 -2232 1974 -2226
rect 1968 -2238 1974 -2232
rect 1968 -2244 1974 -2238
rect 1968 -2250 1974 -2244
rect 1968 -2256 1974 -2250
rect 1968 -2262 1974 -2256
rect 1968 -2268 1974 -2262
rect 1968 -2274 1974 -2268
rect 1968 -2280 1974 -2274
rect 1968 -2286 1974 -2280
rect 1968 -2292 1974 -2286
rect 1968 -2298 1974 -2292
rect 1968 -2304 1974 -2298
rect 1968 -2310 1974 -2304
rect 1968 -2316 1974 -2310
rect 1968 -2322 1974 -2316
rect 1968 -2328 1974 -2322
rect 1968 -2334 1974 -2328
rect 1968 -2340 1974 -2334
rect 1968 -2346 1974 -2340
rect 1968 -2352 1974 -2346
rect 1968 -2358 1974 -2352
rect 1968 -2364 1974 -2358
rect 1968 -2370 1974 -2364
rect 1968 -2376 1974 -2370
rect 1968 -2382 1974 -2376
rect 1968 -2388 1974 -2382
rect 1968 -2394 1974 -2388
rect 1968 -2400 1974 -2394
rect 1968 -2406 1974 -2400
rect 1968 -2412 1974 -2406
rect 1968 -2418 1974 -2412
rect 1968 -2424 1974 -2418
rect 1968 -2430 1974 -2424
rect 1968 -2436 1974 -2430
rect 1968 -2442 1974 -2436
rect 1968 -2448 1974 -2442
rect 1968 -2454 1974 -2448
rect 1968 -2460 1974 -2454
rect 1968 -2466 1974 -2460
rect 1968 -2472 1974 -2466
rect 1968 -2478 1974 -2472
rect 1968 -2484 1974 -2478
rect 1968 -2490 1974 -2484
rect 1968 -2496 1974 -2490
rect 1968 -2502 1974 -2496
rect 1968 -2508 1974 -2502
rect 1968 -2514 1974 -2508
rect 1968 -2520 1974 -2514
rect 1968 -2526 1974 -2520
rect 1968 -2532 1974 -2526
rect 1968 -2538 1974 -2532
rect 1968 -2544 1974 -2538
rect 1968 -2622 1974 -2616
rect 1968 -2628 1974 -2622
rect 1968 -2634 1974 -2628
rect 1968 -2640 1974 -2634
rect 1968 -2646 1974 -2640
rect 1968 -2652 1974 -2646
rect 1968 -2658 1974 -2652
rect 1968 -2664 1974 -2658
rect 1968 -2670 1974 -2664
rect 1968 -2676 1974 -2670
rect 1968 -2682 1974 -2676
rect 1968 -2688 1974 -2682
rect 1968 -2694 1974 -2688
rect 1968 -2700 1974 -2694
rect 1968 -2706 1974 -2700
rect 1968 -2712 1974 -2706
rect 1968 -2718 1974 -2712
rect 1968 -2724 1974 -2718
rect 1968 -2730 1974 -2724
rect 1968 -2736 1974 -2730
rect 1968 -2742 1974 -2736
rect 1968 -2748 1974 -2742
rect 1968 -2754 1974 -2748
rect 1968 -2760 1974 -2754
rect 1968 -2766 1974 -2760
rect 1968 -2772 1974 -2766
rect 1968 -2778 1974 -2772
rect 1968 -2784 1974 -2778
rect 1968 -2790 1974 -2784
rect 1968 -2796 1974 -2790
rect 1968 -2802 1974 -2796
rect 1968 -2808 1974 -2802
rect 1968 -2814 1974 -2808
rect 1968 -2820 1974 -2814
rect 1968 -2826 1974 -2820
rect 1968 -2832 1974 -2826
rect 1968 -2838 1974 -2832
rect 1968 -2844 1974 -2838
rect 1968 -2850 1974 -2844
rect 1968 -2856 1974 -2850
rect 1968 -2862 1974 -2856
rect 1968 -2868 1974 -2862
rect 1968 -2874 1974 -2868
rect 1968 -2880 1974 -2874
rect 1968 -2886 1974 -2880
rect 1968 -2892 1974 -2886
rect 1968 -2898 1974 -2892
rect 1968 -2904 1974 -2898
rect 1968 -2910 1974 -2904
rect 1968 -2916 1974 -2910
rect 1968 -2922 1974 -2916
rect 1968 -2928 1974 -2922
rect 1968 -2934 1974 -2928
rect 1968 -2940 1974 -2934
rect 1968 -2946 1974 -2940
rect 1968 -2952 1974 -2946
rect 1968 -2958 1974 -2952
rect 1968 -2964 1974 -2958
rect 1968 -2970 1974 -2964
rect 1968 -2976 1974 -2970
rect 1968 -2982 1974 -2976
rect 1968 -2988 1974 -2982
rect 1968 -2994 1974 -2988
rect 1968 -3000 1974 -2994
rect 1968 -3006 1974 -3000
rect 1968 -3012 1974 -3006
rect 1968 -3018 1974 -3012
rect 1968 -3024 1974 -3018
rect 1968 -3030 1974 -3024
rect 1968 -3036 1974 -3030
rect 1968 -3042 1974 -3036
rect 1968 -3048 1974 -3042
rect 1968 -3054 1974 -3048
rect 1968 -3060 1974 -3054
rect 1968 -3066 1974 -3060
rect 1968 -3072 1974 -3066
rect 1968 -3078 1974 -3072
rect 1968 -3084 1974 -3078
rect 1968 -3090 1974 -3084
rect 1968 -3096 1974 -3090
rect 1968 -3102 1974 -3096
rect 1968 -3108 1974 -3102
rect 1968 -3114 1974 -3108
rect 1968 -3174 1974 -3168
rect 1968 -3180 1974 -3174
rect 1968 -3186 1974 -3180
rect 1968 -3192 1974 -3186
rect 1968 -3198 1974 -3192
rect 1968 -3204 1974 -3198
rect 1968 -3210 1974 -3204
rect 1968 -3216 1974 -3210
rect 1968 -3222 1974 -3216
rect 1968 -3228 1974 -3222
rect 1968 -3234 1974 -3228
rect 1968 -3240 1974 -3234
rect 1968 -3246 1974 -3240
rect 1974 -486 1980 -480
rect 1974 -492 1980 -486
rect 1974 -498 1980 -492
rect 1974 -504 1980 -498
rect 1974 -510 1980 -504
rect 1974 -516 1980 -510
rect 1974 -522 1980 -516
rect 1974 -528 1980 -522
rect 1974 -534 1980 -528
rect 1974 -540 1980 -534
rect 1974 -546 1980 -540
rect 1974 -552 1980 -546
rect 1974 -558 1980 -552
rect 1974 -564 1980 -558
rect 1974 -570 1980 -564
rect 1974 -576 1980 -570
rect 1974 -582 1980 -576
rect 1974 -588 1980 -582
rect 1974 -594 1980 -588
rect 1974 -600 1980 -594
rect 1974 -606 1980 -600
rect 1974 -612 1980 -606
rect 1974 -618 1980 -612
rect 1974 -624 1980 -618
rect 1974 -630 1980 -624
rect 1974 -636 1980 -630
rect 1974 -642 1980 -636
rect 1974 -648 1980 -642
rect 1974 -654 1980 -648
rect 1974 -660 1980 -654
rect 1974 -666 1980 -660
rect 1974 -672 1980 -666
rect 1974 -678 1980 -672
rect 1974 -684 1980 -678
rect 1974 -690 1980 -684
rect 1974 -696 1980 -690
rect 1974 -702 1980 -696
rect 1974 -708 1980 -702
rect 1974 -714 1980 -708
rect 1974 -720 1980 -714
rect 1974 -726 1980 -720
rect 1974 -732 1980 -726
rect 1974 -738 1980 -732
rect 1974 -744 1980 -738
rect 1974 -750 1980 -744
rect 1974 -756 1980 -750
rect 1974 -762 1980 -756
rect 1974 -768 1980 -762
rect 1974 -774 1980 -768
rect 1974 -780 1980 -774
rect 1974 -786 1980 -780
rect 1974 -792 1980 -786
rect 1974 -798 1980 -792
rect 1974 -804 1980 -798
rect 1974 -810 1980 -804
rect 1974 -816 1980 -810
rect 1974 -822 1980 -816
rect 1974 -828 1980 -822
rect 1974 -834 1980 -828
rect 1974 -840 1980 -834
rect 1974 -846 1980 -840
rect 1974 -852 1980 -846
rect 1974 -858 1980 -852
rect 1974 -864 1980 -858
rect 1974 -870 1980 -864
rect 1974 -876 1980 -870
rect 1974 -882 1980 -876
rect 1974 -888 1980 -882
rect 1974 -894 1980 -888
rect 1974 -900 1980 -894
rect 1974 -906 1980 -900
rect 1974 -912 1980 -906
rect 1974 -918 1980 -912
rect 1974 -924 1980 -918
rect 1974 -930 1980 -924
rect 1974 -936 1980 -930
rect 1974 -942 1980 -936
rect 1974 -948 1980 -942
rect 1974 -954 1980 -948
rect 1974 -960 1980 -954
rect 1974 -966 1980 -960
rect 1974 -972 1980 -966
rect 1974 -978 1980 -972
rect 1974 -984 1980 -978
rect 1974 -990 1980 -984
rect 1974 -996 1980 -990
rect 1974 -1002 1980 -996
rect 1974 -1008 1980 -1002
rect 1974 -1014 1980 -1008
rect 1974 -1020 1980 -1014
rect 1974 -1026 1980 -1020
rect 1974 -1032 1980 -1026
rect 1974 -1038 1980 -1032
rect 1974 -1044 1980 -1038
rect 1974 -1050 1980 -1044
rect 1974 -1056 1980 -1050
rect 1974 -1062 1980 -1056
rect 1974 -1068 1980 -1062
rect 1974 -1074 1980 -1068
rect 1974 -1080 1980 -1074
rect 1974 -1086 1980 -1080
rect 1974 -1092 1980 -1086
rect 1974 -1098 1980 -1092
rect 1974 -1104 1980 -1098
rect 1974 -1110 1980 -1104
rect 1974 -1116 1980 -1110
rect 1974 -1122 1980 -1116
rect 1974 -1128 1980 -1122
rect 1974 -1134 1980 -1128
rect 1974 -1140 1980 -1134
rect 1974 -1146 1980 -1140
rect 1974 -1152 1980 -1146
rect 1974 -1158 1980 -1152
rect 1974 -1164 1980 -1158
rect 1974 -1170 1980 -1164
rect 1974 -1176 1980 -1170
rect 1974 -1182 1980 -1176
rect 1974 -1188 1980 -1182
rect 1974 -1194 1980 -1188
rect 1974 -1200 1980 -1194
rect 1974 -1206 1980 -1200
rect 1974 -1212 1980 -1206
rect 1974 -1218 1980 -1212
rect 1974 -1224 1980 -1218
rect 1974 -1230 1980 -1224
rect 1974 -1236 1980 -1230
rect 1974 -1242 1980 -1236
rect 1974 -1248 1980 -1242
rect 1974 -1254 1980 -1248
rect 1974 -1260 1980 -1254
rect 1974 -1266 1980 -1260
rect 1974 -1272 1980 -1266
rect 1974 -1278 1980 -1272
rect 1974 -1284 1980 -1278
rect 1974 -1290 1980 -1284
rect 1974 -1296 1980 -1290
rect 1974 -1302 1980 -1296
rect 1974 -1308 1980 -1302
rect 1974 -1314 1980 -1308
rect 1974 -1320 1980 -1314
rect 1974 -1326 1980 -1320
rect 1974 -1332 1980 -1326
rect 1974 -1338 1980 -1332
rect 1974 -1344 1980 -1338
rect 1974 -1350 1980 -1344
rect 1974 -1356 1980 -1350
rect 1974 -1362 1980 -1356
rect 1974 -1368 1980 -1362
rect 1974 -1374 1980 -1368
rect 1974 -1380 1980 -1374
rect 1974 -1386 1980 -1380
rect 1974 -1392 1980 -1386
rect 1974 -1398 1980 -1392
rect 1974 -1404 1980 -1398
rect 1974 -1410 1980 -1404
rect 1974 -1416 1980 -1410
rect 1974 -1422 1980 -1416
rect 1974 -1428 1980 -1422
rect 1974 -1434 1980 -1428
rect 1974 -1440 1980 -1434
rect 1974 -1446 1980 -1440
rect 1974 -1452 1980 -1446
rect 1974 -1458 1980 -1452
rect 1974 -1464 1980 -1458
rect 1974 -1470 1980 -1464
rect 1974 -1476 1980 -1470
rect 1974 -1482 1980 -1476
rect 1974 -1488 1980 -1482
rect 1974 -1494 1980 -1488
rect 1974 -1500 1980 -1494
rect 1974 -1506 1980 -1500
rect 1974 -1512 1980 -1506
rect 1974 -1518 1980 -1512
rect 1974 -1524 1980 -1518
rect 1974 -1530 1980 -1524
rect 1974 -1536 1980 -1530
rect 1974 -1542 1980 -1536
rect 1974 -1548 1980 -1542
rect 1974 -1554 1980 -1548
rect 1974 -1560 1980 -1554
rect 1974 -1566 1980 -1560
rect 1974 -1572 1980 -1566
rect 1974 -1578 1980 -1572
rect 1974 -1584 1980 -1578
rect 1974 -1590 1980 -1584
rect 1974 -1596 1980 -1590
rect 1974 -1602 1980 -1596
rect 1974 -1608 1980 -1602
rect 1974 -1614 1980 -1608
rect 1974 -1620 1980 -1614
rect 1974 -1626 1980 -1620
rect 1974 -1632 1980 -1626
rect 1974 -1638 1980 -1632
rect 1974 -1644 1980 -1638
rect 1974 -1650 1980 -1644
rect 1974 -1656 1980 -1650
rect 1974 -1662 1980 -1656
rect 1974 -1668 1980 -1662
rect 1974 -1758 1980 -1752
rect 1974 -1764 1980 -1758
rect 1974 -1770 1980 -1764
rect 1974 -1776 1980 -1770
rect 1974 -1782 1980 -1776
rect 1974 -1788 1980 -1782
rect 1974 -1794 1980 -1788
rect 1974 -1800 1980 -1794
rect 1974 -1806 1980 -1800
rect 1974 -1812 1980 -1806
rect 1974 -1818 1980 -1812
rect 1974 -1824 1980 -1818
rect 1974 -1830 1980 -1824
rect 1974 -1836 1980 -1830
rect 1974 -1842 1980 -1836
rect 1974 -1848 1980 -1842
rect 1974 -1854 1980 -1848
rect 1974 -1860 1980 -1854
rect 1974 -1866 1980 -1860
rect 1974 -1872 1980 -1866
rect 1974 -1878 1980 -1872
rect 1974 -1884 1980 -1878
rect 1974 -1890 1980 -1884
rect 1974 -1896 1980 -1890
rect 1974 -1902 1980 -1896
rect 1974 -1908 1980 -1902
rect 1974 -1914 1980 -1908
rect 1974 -1920 1980 -1914
rect 1974 -1926 1980 -1920
rect 1974 -1932 1980 -1926
rect 1974 -1938 1980 -1932
rect 1974 -1944 1980 -1938
rect 1974 -1950 1980 -1944
rect 1974 -1956 1980 -1950
rect 1974 -1962 1980 -1956
rect 1974 -1968 1980 -1962
rect 1974 -1974 1980 -1968
rect 1974 -1980 1980 -1974
rect 1974 -1986 1980 -1980
rect 1974 -1992 1980 -1986
rect 1974 -1998 1980 -1992
rect 1974 -2004 1980 -1998
rect 1974 -2010 1980 -2004
rect 1974 -2016 1980 -2010
rect 1974 -2022 1980 -2016
rect 1974 -2028 1980 -2022
rect 1974 -2034 1980 -2028
rect 1974 -2040 1980 -2034
rect 1974 -2046 1980 -2040
rect 1974 -2052 1980 -2046
rect 1974 -2058 1980 -2052
rect 1974 -2064 1980 -2058
rect 1974 -2070 1980 -2064
rect 1974 -2076 1980 -2070
rect 1974 -2082 1980 -2076
rect 1974 -2088 1980 -2082
rect 1974 -2094 1980 -2088
rect 1974 -2100 1980 -2094
rect 1974 -2106 1980 -2100
rect 1974 -2112 1980 -2106
rect 1974 -2118 1980 -2112
rect 1974 -2124 1980 -2118
rect 1974 -2130 1980 -2124
rect 1974 -2136 1980 -2130
rect 1974 -2142 1980 -2136
rect 1974 -2148 1980 -2142
rect 1974 -2154 1980 -2148
rect 1974 -2160 1980 -2154
rect 1974 -2166 1980 -2160
rect 1974 -2172 1980 -2166
rect 1974 -2178 1980 -2172
rect 1974 -2184 1980 -2178
rect 1974 -2190 1980 -2184
rect 1974 -2196 1980 -2190
rect 1974 -2202 1980 -2196
rect 1974 -2208 1980 -2202
rect 1974 -2214 1980 -2208
rect 1974 -2220 1980 -2214
rect 1974 -2226 1980 -2220
rect 1974 -2232 1980 -2226
rect 1974 -2238 1980 -2232
rect 1974 -2244 1980 -2238
rect 1974 -2250 1980 -2244
rect 1974 -2256 1980 -2250
rect 1974 -2262 1980 -2256
rect 1974 -2268 1980 -2262
rect 1974 -2274 1980 -2268
rect 1974 -2280 1980 -2274
rect 1974 -2286 1980 -2280
rect 1974 -2292 1980 -2286
rect 1974 -2298 1980 -2292
rect 1974 -2304 1980 -2298
rect 1974 -2310 1980 -2304
rect 1974 -2316 1980 -2310
rect 1974 -2322 1980 -2316
rect 1974 -2328 1980 -2322
rect 1974 -2334 1980 -2328
rect 1974 -2340 1980 -2334
rect 1974 -2346 1980 -2340
rect 1974 -2352 1980 -2346
rect 1974 -2358 1980 -2352
rect 1974 -2364 1980 -2358
rect 1974 -2370 1980 -2364
rect 1974 -2376 1980 -2370
rect 1974 -2382 1980 -2376
rect 1974 -2388 1980 -2382
rect 1974 -2394 1980 -2388
rect 1974 -2400 1980 -2394
rect 1974 -2406 1980 -2400
rect 1974 -2412 1980 -2406
rect 1974 -2418 1980 -2412
rect 1974 -2424 1980 -2418
rect 1974 -2430 1980 -2424
rect 1974 -2436 1980 -2430
rect 1974 -2442 1980 -2436
rect 1974 -2448 1980 -2442
rect 1974 -2454 1980 -2448
rect 1974 -2460 1980 -2454
rect 1974 -2466 1980 -2460
rect 1974 -2472 1980 -2466
rect 1974 -2478 1980 -2472
rect 1974 -2484 1980 -2478
rect 1974 -2490 1980 -2484
rect 1974 -2496 1980 -2490
rect 1974 -2502 1980 -2496
rect 1974 -2508 1980 -2502
rect 1974 -2514 1980 -2508
rect 1974 -2520 1980 -2514
rect 1974 -2526 1980 -2520
rect 1974 -2532 1980 -2526
rect 1974 -2538 1980 -2532
rect 1974 -2622 1980 -2616
rect 1974 -2628 1980 -2622
rect 1974 -2634 1980 -2628
rect 1974 -2640 1980 -2634
rect 1974 -2646 1980 -2640
rect 1974 -2652 1980 -2646
rect 1974 -2658 1980 -2652
rect 1974 -2664 1980 -2658
rect 1974 -2670 1980 -2664
rect 1974 -2676 1980 -2670
rect 1974 -2682 1980 -2676
rect 1974 -2688 1980 -2682
rect 1974 -2694 1980 -2688
rect 1974 -2700 1980 -2694
rect 1974 -2706 1980 -2700
rect 1974 -2712 1980 -2706
rect 1974 -2718 1980 -2712
rect 1974 -2724 1980 -2718
rect 1974 -2730 1980 -2724
rect 1974 -2736 1980 -2730
rect 1974 -2742 1980 -2736
rect 1974 -2748 1980 -2742
rect 1974 -2754 1980 -2748
rect 1974 -2760 1980 -2754
rect 1974 -2766 1980 -2760
rect 1974 -2772 1980 -2766
rect 1974 -2778 1980 -2772
rect 1974 -2784 1980 -2778
rect 1974 -2790 1980 -2784
rect 1974 -2796 1980 -2790
rect 1974 -2802 1980 -2796
rect 1974 -2808 1980 -2802
rect 1974 -2814 1980 -2808
rect 1974 -2820 1980 -2814
rect 1974 -2826 1980 -2820
rect 1974 -2832 1980 -2826
rect 1974 -2838 1980 -2832
rect 1974 -2844 1980 -2838
rect 1974 -2850 1980 -2844
rect 1974 -2856 1980 -2850
rect 1974 -2862 1980 -2856
rect 1974 -2868 1980 -2862
rect 1974 -2874 1980 -2868
rect 1974 -2880 1980 -2874
rect 1974 -2886 1980 -2880
rect 1974 -2892 1980 -2886
rect 1974 -2898 1980 -2892
rect 1974 -2904 1980 -2898
rect 1974 -2910 1980 -2904
rect 1974 -2916 1980 -2910
rect 1974 -2922 1980 -2916
rect 1974 -2928 1980 -2922
rect 1974 -2934 1980 -2928
rect 1974 -2940 1980 -2934
rect 1974 -2946 1980 -2940
rect 1974 -2952 1980 -2946
rect 1974 -2958 1980 -2952
rect 1974 -2964 1980 -2958
rect 1974 -2970 1980 -2964
rect 1974 -2976 1980 -2970
rect 1974 -2982 1980 -2976
rect 1974 -2988 1980 -2982
rect 1974 -2994 1980 -2988
rect 1974 -3000 1980 -2994
rect 1974 -3006 1980 -3000
rect 1974 -3012 1980 -3006
rect 1974 -3018 1980 -3012
rect 1974 -3024 1980 -3018
rect 1974 -3030 1980 -3024
rect 1974 -3036 1980 -3030
rect 1974 -3042 1980 -3036
rect 1974 -3048 1980 -3042
rect 1974 -3054 1980 -3048
rect 1974 -3060 1980 -3054
rect 1974 -3066 1980 -3060
rect 1974 -3072 1980 -3066
rect 1974 -3078 1980 -3072
rect 1974 -3084 1980 -3078
rect 1974 -3090 1980 -3084
rect 1974 -3096 1980 -3090
rect 1974 -3102 1980 -3096
rect 1974 -3108 1980 -3102
rect 1974 -3114 1980 -3108
rect 1974 -3168 1980 -3162
rect 1974 -3174 1980 -3168
rect 1974 -3180 1980 -3174
rect 1974 -3186 1980 -3180
rect 1974 -3192 1980 -3186
rect 1974 -3198 1980 -3192
rect 1974 -3204 1980 -3198
rect 1974 -3210 1980 -3204
rect 1974 -3216 1980 -3210
rect 1974 -3222 1980 -3216
rect 1974 -3228 1980 -3222
rect 1974 -3234 1980 -3228
rect 1974 -3240 1980 -3234
rect 1980 -480 1986 -474
rect 1980 -486 1986 -480
rect 1980 -492 1986 -486
rect 1980 -498 1986 -492
rect 1980 -504 1986 -498
rect 1980 -510 1986 -504
rect 1980 -516 1986 -510
rect 1980 -522 1986 -516
rect 1980 -528 1986 -522
rect 1980 -534 1986 -528
rect 1980 -540 1986 -534
rect 1980 -546 1986 -540
rect 1980 -552 1986 -546
rect 1980 -558 1986 -552
rect 1980 -564 1986 -558
rect 1980 -570 1986 -564
rect 1980 -576 1986 -570
rect 1980 -582 1986 -576
rect 1980 -588 1986 -582
rect 1980 -594 1986 -588
rect 1980 -600 1986 -594
rect 1980 -606 1986 -600
rect 1980 -612 1986 -606
rect 1980 -618 1986 -612
rect 1980 -624 1986 -618
rect 1980 -630 1986 -624
rect 1980 -636 1986 -630
rect 1980 -642 1986 -636
rect 1980 -648 1986 -642
rect 1980 -654 1986 -648
rect 1980 -660 1986 -654
rect 1980 -666 1986 -660
rect 1980 -672 1986 -666
rect 1980 -678 1986 -672
rect 1980 -684 1986 -678
rect 1980 -690 1986 -684
rect 1980 -696 1986 -690
rect 1980 -702 1986 -696
rect 1980 -708 1986 -702
rect 1980 -714 1986 -708
rect 1980 -720 1986 -714
rect 1980 -726 1986 -720
rect 1980 -732 1986 -726
rect 1980 -738 1986 -732
rect 1980 -744 1986 -738
rect 1980 -750 1986 -744
rect 1980 -756 1986 -750
rect 1980 -762 1986 -756
rect 1980 -768 1986 -762
rect 1980 -774 1986 -768
rect 1980 -780 1986 -774
rect 1980 -786 1986 -780
rect 1980 -792 1986 -786
rect 1980 -798 1986 -792
rect 1980 -804 1986 -798
rect 1980 -810 1986 -804
rect 1980 -816 1986 -810
rect 1980 -822 1986 -816
rect 1980 -828 1986 -822
rect 1980 -834 1986 -828
rect 1980 -840 1986 -834
rect 1980 -846 1986 -840
rect 1980 -852 1986 -846
rect 1980 -858 1986 -852
rect 1980 -864 1986 -858
rect 1980 -870 1986 -864
rect 1980 -876 1986 -870
rect 1980 -882 1986 -876
rect 1980 -888 1986 -882
rect 1980 -894 1986 -888
rect 1980 -900 1986 -894
rect 1980 -906 1986 -900
rect 1980 -912 1986 -906
rect 1980 -918 1986 -912
rect 1980 -924 1986 -918
rect 1980 -930 1986 -924
rect 1980 -936 1986 -930
rect 1980 -942 1986 -936
rect 1980 -948 1986 -942
rect 1980 -954 1986 -948
rect 1980 -960 1986 -954
rect 1980 -966 1986 -960
rect 1980 -972 1986 -966
rect 1980 -978 1986 -972
rect 1980 -984 1986 -978
rect 1980 -990 1986 -984
rect 1980 -996 1986 -990
rect 1980 -1002 1986 -996
rect 1980 -1008 1986 -1002
rect 1980 -1014 1986 -1008
rect 1980 -1020 1986 -1014
rect 1980 -1026 1986 -1020
rect 1980 -1032 1986 -1026
rect 1980 -1038 1986 -1032
rect 1980 -1044 1986 -1038
rect 1980 -1050 1986 -1044
rect 1980 -1056 1986 -1050
rect 1980 -1062 1986 -1056
rect 1980 -1068 1986 -1062
rect 1980 -1074 1986 -1068
rect 1980 -1080 1986 -1074
rect 1980 -1086 1986 -1080
rect 1980 -1092 1986 -1086
rect 1980 -1098 1986 -1092
rect 1980 -1104 1986 -1098
rect 1980 -1110 1986 -1104
rect 1980 -1116 1986 -1110
rect 1980 -1122 1986 -1116
rect 1980 -1128 1986 -1122
rect 1980 -1134 1986 -1128
rect 1980 -1140 1986 -1134
rect 1980 -1146 1986 -1140
rect 1980 -1152 1986 -1146
rect 1980 -1158 1986 -1152
rect 1980 -1164 1986 -1158
rect 1980 -1170 1986 -1164
rect 1980 -1176 1986 -1170
rect 1980 -1182 1986 -1176
rect 1980 -1188 1986 -1182
rect 1980 -1194 1986 -1188
rect 1980 -1200 1986 -1194
rect 1980 -1206 1986 -1200
rect 1980 -1212 1986 -1206
rect 1980 -1218 1986 -1212
rect 1980 -1224 1986 -1218
rect 1980 -1230 1986 -1224
rect 1980 -1236 1986 -1230
rect 1980 -1242 1986 -1236
rect 1980 -1248 1986 -1242
rect 1980 -1254 1986 -1248
rect 1980 -1260 1986 -1254
rect 1980 -1266 1986 -1260
rect 1980 -1272 1986 -1266
rect 1980 -1278 1986 -1272
rect 1980 -1284 1986 -1278
rect 1980 -1290 1986 -1284
rect 1980 -1296 1986 -1290
rect 1980 -1302 1986 -1296
rect 1980 -1308 1986 -1302
rect 1980 -1314 1986 -1308
rect 1980 -1320 1986 -1314
rect 1980 -1326 1986 -1320
rect 1980 -1332 1986 -1326
rect 1980 -1338 1986 -1332
rect 1980 -1344 1986 -1338
rect 1980 -1350 1986 -1344
rect 1980 -1356 1986 -1350
rect 1980 -1362 1986 -1356
rect 1980 -1368 1986 -1362
rect 1980 -1374 1986 -1368
rect 1980 -1380 1986 -1374
rect 1980 -1386 1986 -1380
rect 1980 -1392 1986 -1386
rect 1980 -1398 1986 -1392
rect 1980 -1404 1986 -1398
rect 1980 -1410 1986 -1404
rect 1980 -1416 1986 -1410
rect 1980 -1422 1986 -1416
rect 1980 -1428 1986 -1422
rect 1980 -1434 1986 -1428
rect 1980 -1440 1986 -1434
rect 1980 -1446 1986 -1440
rect 1980 -1452 1986 -1446
rect 1980 -1458 1986 -1452
rect 1980 -1464 1986 -1458
rect 1980 -1470 1986 -1464
rect 1980 -1476 1986 -1470
rect 1980 -1482 1986 -1476
rect 1980 -1488 1986 -1482
rect 1980 -1494 1986 -1488
rect 1980 -1500 1986 -1494
rect 1980 -1506 1986 -1500
rect 1980 -1512 1986 -1506
rect 1980 -1518 1986 -1512
rect 1980 -1524 1986 -1518
rect 1980 -1530 1986 -1524
rect 1980 -1536 1986 -1530
rect 1980 -1542 1986 -1536
rect 1980 -1548 1986 -1542
rect 1980 -1554 1986 -1548
rect 1980 -1560 1986 -1554
rect 1980 -1566 1986 -1560
rect 1980 -1572 1986 -1566
rect 1980 -1578 1986 -1572
rect 1980 -1584 1986 -1578
rect 1980 -1590 1986 -1584
rect 1980 -1596 1986 -1590
rect 1980 -1602 1986 -1596
rect 1980 -1608 1986 -1602
rect 1980 -1614 1986 -1608
rect 1980 -1620 1986 -1614
rect 1980 -1626 1986 -1620
rect 1980 -1632 1986 -1626
rect 1980 -1638 1986 -1632
rect 1980 -1644 1986 -1638
rect 1980 -1650 1986 -1644
rect 1980 -1656 1986 -1650
rect 1980 -1662 1986 -1656
rect 1980 -1752 1986 -1746
rect 1980 -1758 1986 -1752
rect 1980 -1764 1986 -1758
rect 1980 -1770 1986 -1764
rect 1980 -1776 1986 -1770
rect 1980 -1782 1986 -1776
rect 1980 -1788 1986 -1782
rect 1980 -1794 1986 -1788
rect 1980 -1800 1986 -1794
rect 1980 -1806 1986 -1800
rect 1980 -1812 1986 -1806
rect 1980 -1818 1986 -1812
rect 1980 -1824 1986 -1818
rect 1980 -1830 1986 -1824
rect 1980 -1836 1986 -1830
rect 1980 -1842 1986 -1836
rect 1980 -1848 1986 -1842
rect 1980 -1854 1986 -1848
rect 1980 -1860 1986 -1854
rect 1980 -1866 1986 -1860
rect 1980 -1872 1986 -1866
rect 1980 -1878 1986 -1872
rect 1980 -1884 1986 -1878
rect 1980 -1890 1986 -1884
rect 1980 -1896 1986 -1890
rect 1980 -1902 1986 -1896
rect 1980 -1908 1986 -1902
rect 1980 -1914 1986 -1908
rect 1980 -1920 1986 -1914
rect 1980 -1926 1986 -1920
rect 1980 -1932 1986 -1926
rect 1980 -1938 1986 -1932
rect 1980 -1944 1986 -1938
rect 1980 -1950 1986 -1944
rect 1980 -1956 1986 -1950
rect 1980 -1962 1986 -1956
rect 1980 -1968 1986 -1962
rect 1980 -1974 1986 -1968
rect 1980 -1980 1986 -1974
rect 1980 -1986 1986 -1980
rect 1980 -1992 1986 -1986
rect 1980 -1998 1986 -1992
rect 1980 -2004 1986 -1998
rect 1980 -2010 1986 -2004
rect 1980 -2016 1986 -2010
rect 1980 -2022 1986 -2016
rect 1980 -2028 1986 -2022
rect 1980 -2034 1986 -2028
rect 1980 -2040 1986 -2034
rect 1980 -2046 1986 -2040
rect 1980 -2052 1986 -2046
rect 1980 -2058 1986 -2052
rect 1980 -2064 1986 -2058
rect 1980 -2070 1986 -2064
rect 1980 -2076 1986 -2070
rect 1980 -2082 1986 -2076
rect 1980 -2088 1986 -2082
rect 1980 -2094 1986 -2088
rect 1980 -2100 1986 -2094
rect 1980 -2106 1986 -2100
rect 1980 -2112 1986 -2106
rect 1980 -2118 1986 -2112
rect 1980 -2124 1986 -2118
rect 1980 -2130 1986 -2124
rect 1980 -2136 1986 -2130
rect 1980 -2142 1986 -2136
rect 1980 -2148 1986 -2142
rect 1980 -2154 1986 -2148
rect 1980 -2160 1986 -2154
rect 1980 -2166 1986 -2160
rect 1980 -2172 1986 -2166
rect 1980 -2178 1986 -2172
rect 1980 -2184 1986 -2178
rect 1980 -2190 1986 -2184
rect 1980 -2196 1986 -2190
rect 1980 -2202 1986 -2196
rect 1980 -2208 1986 -2202
rect 1980 -2214 1986 -2208
rect 1980 -2220 1986 -2214
rect 1980 -2226 1986 -2220
rect 1980 -2232 1986 -2226
rect 1980 -2238 1986 -2232
rect 1980 -2244 1986 -2238
rect 1980 -2250 1986 -2244
rect 1980 -2256 1986 -2250
rect 1980 -2262 1986 -2256
rect 1980 -2268 1986 -2262
rect 1980 -2274 1986 -2268
rect 1980 -2280 1986 -2274
rect 1980 -2286 1986 -2280
rect 1980 -2292 1986 -2286
rect 1980 -2298 1986 -2292
rect 1980 -2304 1986 -2298
rect 1980 -2310 1986 -2304
rect 1980 -2316 1986 -2310
rect 1980 -2322 1986 -2316
rect 1980 -2328 1986 -2322
rect 1980 -2334 1986 -2328
rect 1980 -2340 1986 -2334
rect 1980 -2346 1986 -2340
rect 1980 -2352 1986 -2346
rect 1980 -2358 1986 -2352
rect 1980 -2364 1986 -2358
rect 1980 -2370 1986 -2364
rect 1980 -2376 1986 -2370
rect 1980 -2382 1986 -2376
rect 1980 -2388 1986 -2382
rect 1980 -2394 1986 -2388
rect 1980 -2400 1986 -2394
rect 1980 -2406 1986 -2400
rect 1980 -2412 1986 -2406
rect 1980 -2418 1986 -2412
rect 1980 -2424 1986 -2418
rect 1980 -2430 1986 -2424
rect 1980 -2436 1986 -2430
rect 1980 -2442 1986 -2436
rect 1980 -2448 1986 -2442
rect 1980 -2454 1986 -2448
rect 1980 -2460 1986 -2454
rect 1980 -2466 1986 -2460
rect 1980 -2472 1986 -2466
rect 1980 -2478 1986 -2472
rect 1980 -2484 1986 -2478
rect 1980 -2490 1986 -2484
rect 1980 -2496 1986 -2490
rect 1980 -2502 1986 -2496
rect 1980 -2508 1986 -2502
rect 1980 -2514 1986 -2508
rect 1980 -2520 1986 -2514
rect 1980 -2526 1986 -2520
rect 1980 -2532 1986 -2526
rect 1980 -2538 1986 -2532
rect 1980 -2622 1986 -2616
rect 1980 -2628 1986 -2622
rect 1980 -2634 1986 -2628
rect 1980 -2640 1986 -2634
rect 1980 -2646 1986 -2640
rect 1980 -2652 1986 -2646
rect 1980 -2658 1986 -2652
rect 1980 -2664 1986 -2658
rect 1980 -2670 1986 -2664
rect 1980 -2676 1986 -2670
rect 1980 -2682 1986 -2676
rect 1980 -2688 1986 -2682
rect 1980 -2694 1986 -2688
rect 1980 -2700 1986 -2694
rect 1980 -2706 1986 -2700
rect 1980 -2712 1986 -2706
rect 1980 -2718 1986 -2712
rect 1980 -2724 1986 -2718
rect 1980 -2730 1986 -2724
rect 1980 -2736 1986 -2730
rect 1980 -2742 1986 -2736
rect 1980 -2748 1986 -2742
rect 1980 -2754 1986 -2748
rect 1980 -2760 1986 -2754
rect 1980 -2766 1986 -2760
rect 1980 -2772 1986 -2766
rect 1980 -2778 1986 -2772
rect 1980 -2784 1986 -2778
rect 1980 -2790 1986 -2784
rect 1980 -2796 1986 -2790
rect 1980 -2802 1986 -2796
rect 1980 -2808 1986 -2802
rect 1980 -2814 1986 -2808
rect 1980 -2820 1986 -2814
rect 1980 -2826 1986 -2820
rect 1980 -2832 1986 -2826
rect 1980 -2838 1986 -2832
rect 1980 -2844 1986 -2838
rect 1980 -2850 1986 -2844
rect 1980 -2856 1986 -2850
rect 1980 -2862 1986 -2856
rect 1980 -2868 1986 -2862
rect 1980 -2874 1986 -2868
rect 1980 -2880 1986 -2874
rect 1980 -2886 1986 -2880
rect 1980 -2892 1986 -2886
rect 1980 -2898 1986 -2892
rect 1980 -2904 1986 -2898
rect 1980 -2910 1986 -2904
rect 1980 -2916 1986 -2910
rect 1980 -2922 1986 -2916
rect 1980 -2928 1986 -2922
rect 1980 -2934 1986 -2928
rect 1980 -2940 1986 -2934
rect 1980 -2946 1986 -2940
rect 1980 -2952 1986 -2946
rect 1980 -2958 1986 -2952
rect 1980 -2964 1986 -2958
rect 1980 -2970 1986 -2964
rect 1980 -2976 1986 -2970
rect 1980 -2982 1986 -2976
rect 1980 -2988 1986 -2982
rect 1980 -2994 1986 -2988
rect 1980 -3000 1986 -2994
rect 1980 -3006 1986 -3000
rect 1980 -3012 1986 -3006
rect 1980 -3018 1986 -3012
rect 1980 -3024 1986 -3018
rect 1980 -3030 1986 -3024
rect 1980 -3036 1986 -3030
rect 1980 -3042 1986 -3036
rect 1980 -3048 1986 -3042
rect 1980 -3054 1986 -3048
rect 1980 -3060 1986 -3054
rect 1980 -3066 1986 -3060
rect 1980 -3072 1986 -3066
rect 1980 -3078 1986 -3072
rect 1980 -3084 1986 -3078
rect 1980 -3090 1986 -3084
rect 1980 -3096 1986 -3090
rect 1980 -3102 1986 -3096
rect 1980 -3108 1986 -3102
rect 1980 -3114 1986 -3108
rect 1980 -3168 1986 -3162
rect 1980 -3174 1986 -3168
rect 1980 -3180 1986 -3174
rect 1980 -3186 1986 -3180
rect 1980 -3192 1986 -3186
rect 1980 -3198 1986 -3192
rect 1980 -3204 1986 -3198
rect 1980 -3210 1986 -3204
rect 1980 -3216 1986 -3210
rect 1980 -3222 1986 -3216
rect 1980 -3228 1986 -3222
rect 1980 -3234 1986 -3228
rect 1986 -468 1992 -462
rect 1986 -474 1992 -468
rect 1986 -480 1992 -474
rect 1986 -486 1992 -480
rect 1986 -492 1992 -486
rect 1986 -498 1992 -492
rect 1986 -504 1992 -498
rect 1986 -510 1992 -504
rect 1986 -516 1992 -510
rect 1986 -522 1992 -516
rect 1986 -528 1992 -522
rect 1986 -534 1992 -528
rect 1986 -540 1992 -534
rect 1986 -546 1992 -540
rect 1986 -552 1992 -546
rect 1986 -558 1992 -552
rect 1986 -564 1992 -558
rect 1986 -570 1992 -564
rect 1986 -576 1992 -570
rect 1986 -582 1992 -576
rect 1986 -588 1992 -582
rect 1986 -594 1992 -588
rect 1986 -600 1992 -594
rect 1986 -606 1992 -600
rect 1986 -612 1992 -606
rect 1986 -618 1992 -612
rect 1986 -624 1992 -618
rect 1986 -630 1992 -624
rect 1986 -636 1992 -630
rect 1986 -642 1992 -636
rect 1986 -648 1992 -642
rect 1986 -654 1992 -648
rect 1986 -660 1992 -654
rect 1986 -666 1992 -660
rect 1986 -672 1992 -666
rect 1986 -678 1992 -672
rect 1986 -684 1992 -678
rect 1986 -690 1992 -684
rect 1986 -696 1992 -690
rect 1986 -702 1992 -696
rect 1986 -708 1992 -702
rect 1986 -714 1992 -708
rect 1986 -720 1992 -714
rect 1986 -726 1992 -720
rect 1986 -732 1992 -726
rect 1986 -738 1992 -732
rect 1986 -744 1992 -738
rect 1986 -750 1992 -744
rect 1986 -756 1992 -750
rect 1986 -762 1992 -756
rect 1986 -768 1992 -762
rect 1986 -774 1992 -768
rect 1986 -780 1992 -774
rect 1986 -786 1992 -780
rect 1986 -792 1992 -786
rect 1986 -798 1992 -792
rect 1986 -804 1992 -798
rect 1986 -810 1992 -804
rect 1986 -816 1992 -810
rect 1986 -822 1992 -816
rect 1986 -828 1992 -822
rect 1986 -834 1992 -828
rect 1986 -840 1992 -834
rect 1986 -846 1992 -840
rect 1986 -852 1992 -846
rect 1986 -858 1992 -852
rect 1986 -864 1992 -858
rect 1986 -870 1992 -864
rect 1986 -876 1992 -870
rect 1986 -882 1992 -876
rect 1986 -888 1992 -882
rect 1986 -894 1992 -888
rect 1986 -900 1992 -894
rect 1986 -906 1992 -900
rect 1986 -912 1992 -906
rect 1986 -918 1992 -912
rect 1986 -924 1992 -918
rect 1986 -930 1992 -924
rect 1986 -936 1992 -930
rect 1986 -942 1992 -936
rect 1986 -948 1992 -942
rect 1986 -954 1992 -948
rect 1986 -960 1992 -954
rect 1986 -966 1992 -960
rect 1986 -972 1992 -966
rect 1986 -978 1992 -972
rect 1986 -984 1992 -978
rect 1986 -990 1992 -984
rect 1986 -996 1992 -990
rect 1986 -1002 1992 -996
rect 1986 -1008 1992 -1002
rect 1986 -1014 1992 -1008
rect 1986 -1020 1992 -1014
rect 1986 -1026 1992 -1020
rect 1986 -1032 1992 -1026
rect 1986 -1038 1992 -1032
rect 1986 -1044 1992 -1038
rect 1986 -1050 1992 -1044
rect 1986 -1056 1992 -1050
rect 1986 -1062 1992 -1056
rect 1986 -1068 1992 -1062
rect 1986 -1074 1992 -1068
rect 1986 -1080 1992 -1074
rect 1986 -1086 1992 -1080
rect 1986 -1092 1992 -1086
rect 1986 -1098 1992 -1092
rect 1986 -1104 1992 -1098
rect 1986 -1110 1992 -1104
rect 1986 -1116 1992 -1110
rect 1986 -1122 1992 -1116
rect 1986 -1128 1992 -1122
rect 1986 -1134 1992 -1128
rect 1986 -1140 1992 -1134
rect 1986 -1146 1992 -1140
rect 1986 -1152 1992 -1146
rect 1986 -1158 1992 -1152
rect 1986 -1164 1992 -1158
rect 1986 -1170 1992 -1164
rect 1986 -1176 1992 -1170
rect 1986 -1182 1992 -1176
rect 1986 -1188 1992 -1182
rect 1986 -1194 1992 -1188
rect 1986 -1200 1992 -1194
rect 1986 -1206 1992 -1200
rect 1986 -1212 1992 -1206
rect 1986 -1218 1992 -1212
rect 1986 -1224 1992 -1218
rect 1986 -1230 1992 -1224
rect 1986 -1236 1992 -1230
rect 1986 -1242 1992 -1236
rect 1986 -1248 1992 -1242
rect 1986 -1254 1992 -1248
rect 1986 -1260 1992 -1254
rect 1986 -1266 1992 -1260
rect 1986 -1272 1992 -1266
rect 1986 -1278 1992 -1272
rect 1986 -1284 1992 -1278
rect 1986 -1290 1992 -1284
rect 1986 -1296 1992 -1290
rect 1986 -1302 1992 -1296
rect 1986 -1308 1992 -1302
rect 1986 -1314 1992 -1308
rect 1986 -1320 1992 -1314
rect 1986 -1326 1992 -1320
rect 1986 -1332 1992 -1326
rect 1986 -1338 1992 -1332
rect 1986 -1344 1992 -1338
rect 1986 -1350 1992 -1344
rect 1986 -1356 1992 -1350
rect 1986 -1362 1992 -1356
rect 1986 -1368 1992 -1362
rect 1986 -1374 1992 -1368
rect 1986 -1380 1992 -1374
rect 1986 -1386 1992 -1380
rect 1986 -1392 1992 -1386
rect 1986 -1398 1992 -1392
rect 1986 -1404 1992 -1398
rect 1986 -1410 1992 -1404
rect 1986 -1416 1992 -1410
rect 1986 -1422 1992 -1416
rect 1986 -1428 1992 -1422
rect 1986 -1434 1992 -1428
rect 1986 -1440 1992 -1434
rect 1986 -1446 1992 -1440
rect 1986 -1452 1992 -1446
rect 1986 -1458 1992 -1452
rect 1986 -1464 1992 -1458
rect 1986 -1470 1992 -1464
rect 1986 -1476 1992 -1470
rect 1986 -1482 1992 -1476
rect 1986 -1488 1992 -1482
rect 1986 -1494 1992 -1488
rect 1986 -1500 1992 -1494
rect 1986 -1506 1992 -1500
rect 1986 -1512 1992 -1506
rect 1986 -1518 1992 -1512
rect 1986 -1524 1992 -1518
rect 1986 -1530 1992 -1524
rect 1986 -1536 1992 -1530
rect 1986 -1542 1992 -1536
rect 1986 -1548 1992 -1542
rect 1986 -1554 1992 -1548
rect 1986 -1560 1992 -1554
rect 1986 -1566 1992 -1560
rect 1986 -1572 1992 -1566
rect 1986 -1578 1992 -1572
rect 1986 -1584 1992 -1578
rect 1986 -1590 1992 -1584
rect 1986 -1596 1992 -1590
rect 1986 -1602 1992 -1596
rect 1986 -1608 1992 -1602
rect 1986 -1614 1992 -1608
rect 1986 -1620 1992 -1614
rect 1986 -1626 1992 -1620
rect 1986 -1632 1992 -1626
rect 1986 -1638 1992 -1632
rect 1986 -1644 1992 -1638
rect 1986 -1650 1992 -1644
rect 1986 -1656 1992 -1650
rect 1986 -1746 1992 -1740
rect 1986 -1752 1992 -1746
rect 1986 -1758 1992 -1752
rect 1986 -1764 1992 -1758
rect 1986 -1770 1992 -1764
rect 1986 -1776 1992 -1770
rect 1986 -1782 1992 -1776
rect 1986 -1788 1992 -1782
rect 1986 -1794 1992 -1788
rect 1986 -1800 1992 -1794
rect 1986 -1806 1992 -1800
rect 1986 -1812 1992 -1806
rect 1986 -1818 1992 -1812
rect 1986 -1824 1992 -1818
rect 1986 -1830 1992 -1824
rect 1986 -1836 1992 -1830
rect 1986 -1842 1992 -1836
rect 1986 -1848 1992 -1842
rect 1986 -1854 1992 -1848
rect 1986 -1860 1992 -1854
rect 1986 -1866 1992 -1860
rect 1986 -1872 1992 -1866
rect 1986 -1878 1992 -1872
rect 1986 -1884 1992 -1878
rect 1986 -1890 1992 -1884
rect 1986 -1896 1992 -1890
rect 1986 -1902 1992 -1896
rect 1986 -1908 1992 -1902
rect 1986 -1914 1992 -1908
rect 1986 -1920 1992 -1914
rect 1986 -1926 1992 -1920
rect 1986 -1932 1992 -1926
rect 1986 -1938 1992 -1932
rect 1986 -1944 1992 -1938
rect 1986 -1950 1992 -1944
rect 1986 -1956 1992 -1950
rect 1986 -1962 1992 -1956
rect 1986 -1968 1992 -1962
rect 1986 -1974 1992 -1968
rect 1986 -1980 1992 -1974
rect 1986 -1986 1992 -1980
rect 1986 -1992 1992 -1986
rect 1986 -1998 1992 -1992
rect 1986 -2004 1992 -1998
rect 1986 -2010 1992 -2004
rect 1986 -2016 1992 -2010
rect 1986 -2022 1992 -2016
rect 1986 -2028 1992 -2022
rect 1986 -2034 1992 -2028
rect 1986 -2040 1992 -2034
rect 1986 -2046 1992 -2040
rect 1986 -2052 1992 -2046
rect 1986 -2058 1992 -2052
rect 1986 -2064 1992 -2058
rect 1986 -2070 1992 -2064
rect 1986 -2076 1992 -2070
rect 1986 -2082 1992 -2076
rect 1986 -2088 1992 -2082
rect 1986 -2094 1992 -2088
rect 1986 -2100 1992 -2094
rect 1986 -2106 1992 -2100
rect 1986 -2112 1992 -2106
rect 1986 -2118 1992 -2112
rect 1986 -2124 1992 -2118
rect 1986 -2130 1992 -2124
rect 1986 -2136 1992 -2130
rect 1986 -2142 1992 -2136
rect 1986 -2148 1992 -2142
rect 1986 -2154 1992 -2148
rect 1986 -2160 1992 -2154
rect 1986 -2166 1992 -2160
rect 1986 -2172 1992 -2166
rect 1986 -2178 1992 -2172
rect 1986 -2184 1992 -2178
rect 1986 -2190 1992 -2184
rect 1986 -2196 1992 -2190
rect 1986 -2202 1992 -2196
rect 1986 -2208 1992 -2202
rect 1986 -2214 1992 -2208
rect 1986 -2220 1992 -2214
rect 1986 -2226 1992 -2220
rect 1986 -2232 1992 -2226
rect 1986 -2238 1992 -2232
rect 1986 -2244 1992 -2238
rect 1986 -2250 1992 -2244
rect 1986 -2256 1992 -2250
rect 1986 -2262 1992 -2256
rect 1986 -2268 1992 -2262
rect 1986 -2274 1992 -2268
rect 1986 -2280 1992 -2274
rect 1986 -2286 1992 -2280
rect 1986 -2292 1992 -2286
rect 1986 -2298 1992 -2292
rect 1986 -2304 1992 -2298
rect 1986 -2310 1992 -2304
rect 1986 -2316 1992 -2310
rect 1986 -2322 1992 -2316
rect 1986 -2328 1992 -2322
rect 1986 -2334 1992 -2328
rect 1986 -2340 1992 -2334
rect 1986 -2346 1992 -2340
rect 1986 -2352 1992 -2346
rect 1986 -2358 1992 -2352
rect 1986 -2364 1992 -2358
rect 1986 -2370 1992 -2364
rect 1986 -2376 1992 -2370
rect 1986 -2382 1992 -2376
rect 1986 -2388 1992 -2382
rect 1986 -2394 1992 -2388
rect 1986 -2400 1992 -2394
rect 1986 -2406 1992 -2400
rect 1986 -2412 1992 -2406
rect 1986 -2418 1992 -2412
rect 1986 -2424 1992 -2418
rect 1986 -2430 1992 -2424
rect 1986 -2436 1992 -2430
rect 1986 -2442 1992 -2436
rect 1986 -2448 1992 -2442
rect 1986 -2454 1992 -2448
rect 1986 -2460 1992 -2454
rect 1986 -2466 1992 -2460
rect 1986 -2472 1992 -2466
rect 1986 -2478 1992 -2472
rect 1986 -2484 1992 -2478
rect 1986 -2490 1992 -2484
rect 1986 -2496 1992 -2490
rect 1986 -2502 1992 -2496
rect 1986 -2508 1992 -2502
rect 1986 -2514 1992 -2508
rect 1986 -2520 1992 -2514
rect 1986 -2526 1992 -2520
rect 1986 -2532 1992 -2526
rect 1986 -2616 1992 -2610
rect 1986 -2622 1992 -2616
rect 1986 -2628 1992 -2622
rect 1986 -2634 1992 -2628
rect 1986 -2640 1992 -2634
rect 1986 -2646 1992 -2640
rect 1986 -2652 1992 -2646
rect 1986 -2658 1992 -2652
rect 1986 -2664 1992 -2658
rect 1986 -2670 1992 -2664
rect 1986 -2676 1992 -2670
rect 1986 -2682 1992 -2676
rect 1986 -2688 1992 -2682
rect 1986 -2694 1992 -2688
rect 1986 -2700 1992 -2694
rect 1986 -2706 1992 -2700
rect 1986 -2712 1992 -2706
rect 1986 -2718 1992 -2712
rect 1986 -2724 1992 -2718
rect 1986 -2730 1992 -2724
rect 1986 -2736 1992 -2730
rect 1986 -2742 1992 -2736
rect 1986 -2748 1992 -2742
rect 1986 -2754 1992 -2748
rect 1986 -2760 1992 -2754
rect 1986 -2766 1992 -2760
rect 1986 -2772 1992 -2766
rect 1986 -2778 1992 -2772
rect 1986 -2784 1992 -2778
rect 1986 -2790 1992 -2784
rect 1986 -2796 1992 -2790
rect 1986 -2802 1992 -2796
rect 1986 -2808 1992 -2802
rect 1986 -2814 1992 -2808
rect 1986 -2820 1992 -2814
rect 1986 -2826 1992 -2820
rect 1986 -2832 1992 -2826
rect 1986 -2838 1992 -2832
rect 1986 -2844 1992 -2838
rect 1986 -2850 1992 -2844
rect 1986 -2856 1992 -2850
rect 1986 -2862 1992 -2856
rect 1986 -2868 1992 -2862
rect 1986 -2874 1992 -2868
rect 1986 -2880 1992 -2874
rect 1986 -2886 1992 -2880
rect 1986 -2892 1992 -2886
rect 1986 -2898 1992 -2892
rect 1986 -2904 1992 -2898
rect 1986 -2910 1992 -2904
rect 1986 -2916 1992 -2910
rect 1986 -2922 1992 -2916
rect 1986 -2928 1992 -2922
rect 1986 -2934 1992 -2928
rect 1986 -2940 1992 -2934
rect 1986 -2946 1992 -2940
rect 1986 -2952 1992 -2946
rect 1986 -2958 1992 -2952
rect 1986 -2964 1992 -2958
rect 1986 -2970 1992 -2964
rect 1986 -2976 1992 -2970
rect 1986 -2982 1992 -2976
rect 1986 -2988 1992 -2982
rect 1986 -2994 1992 -2988
rect 1986 -3000 1992 -2994
rect 1986 -3006 1992 -3000
rect 1986 -3012 1992 -3006
rect 1986 -3018 1992 -3012
rect 1986 -3024 1992 -3018
rect 1986 -3030 1992 -3024
rect 1986 -3036 1992 -3030
rect 1986 -3042 1992 -3036
rect 1986 -3048 1992 -3042
rect 1986 -3054 1992 -3048
rect 1986 -3060 1992 -3054
rect 1986 -3066 1992 -3060
rect 1986 -3072 1992 -3066
rect 1986 -3078 1992 -3072
rect 1986 -3084 1992 -3078
rect 1986 -3090 1992 -3084
rect 1986 -3096 1992 -3090
rect 1986 -3102 1992 -3096
rect 1986 -3108 1992 -3102
rect 1986 -3162 1992 -3156
rect 1986 -3168 1992 -3162
rect 1986 -3174 1992 -3168
rect 1986 -3180 1992 -3174
rect 1986 -3186 1992 -3180
rect 1986 -3192 1992 -3186
rect 1986 -3198 1992 -3192
rect 1986 -3204 1992 -3198
rect 1986 -3210 1992 -3204
rect 1986 -3216 1992 -3210
rect 1986 -3222 1992 -3216
rect 1986 -3228 1992 -3222
rect 1992 -462 1998 -456
rect 1992 -468 1998 -462
rect 1992 -474 1998 -468
rect 1992 -480 1998 -474
rect 1992 -486 1998 -480
rect 1992 -492 1998 -486
rect 1992 -498 1998 -492
rect 1992 -504 1998 -498
rect 1992 -510 1998 -504
rect 1992 -516 1998 -510
rect 1992 -522 1998 -516
rect 1992 -528 1998 -522
rect 1992 -534 1998 -528
rect 1992 -540 1998 -534
rect 1992 -546 1998 -540
rect 1992 -552 1998 -546
rect 1992 -558 1998 -552
rect 1992 -564 1998 -558
rect 1992 -570 1998 -564
rect 1992 -576 1998 -570
rect 1992 -582 1998 -576
rect 1992 -588 1998 -582
rect 1992 -594 1998 -588
rect 1992 -600 1998 -594
rect 1992 -606 1998 -600
rect 1992 -612 1998 -606
rect 1992 -618 1998 -612
rect 1992 -624 1998 -618
rect 1992 -630 1998 -624
rect 1992 -636 1998 -630
rect 1992 -642 1998 -636
rect 1992 -648 1998 -642
rect 1992 -654 1998 -648
rect 1992 -660 1998 -654
rect 1992 -666 1998 -660
rect 1992 -672 1998 -666
rect 1992 -678 1998 -672
rect 1992 -684 1998 -678
rect 1992 -690 1998 -684
rect 1992 -696 1998 -690
rect 1992 -702 1998 -696
rect 1992 -708 1998 -702
rect 1992 -714 1998 -708
rect 1992 -720 1998 -714
rect 1992 -726 1998 -720
rect 1992 -732 1998 -726
rect 1992 -738 1998 -732
rect 1992 -744 1998 -738
rect 1992 -750 1998 -744
rect 1992 -756 1998 -750
rect 1992 -762 1998 -756
rect 1992 -768 1998 -762
rect 1992 -774 1998 -768
rect 1992 -780 1998 -774
rect 1992 -786 1998 -780
rect 1992 -792 1998 -786
rect 1992 -798 1998 -792
rect 1992 -804 1998 -798
rect 1992 -810 1998 -804
rect 1992 -816 1998 -810
rect 1992 -822 1998 -816
rect 1992 -828 1998 -822
rect 1992 -834 1998 -828
rect 1992 -840 1998 -834
rect 1992 -846 1998 -840
rect 1992 -852 1998 -846
rect 1992 -858 1998 -852
rect 1992 -864 1998 -858
rect 1992 -870 1998 -864
rect 1992 -876 1998 -870
rect 1992 -882 1998 -876
rect 1992 -888 1998 -882
rect 1992 -894 1998 -888
rect 1992 -900 1998 -894
rect 1992 -906 1998 -900
rect 1992 -912 1998 -906
rect 1992 -918 1998 -912
rect 1992 -924 1998 -918
rect 1992 -930 1998 -924
rect 1992 -936 1998 -930
rect 1992 -942 1998 -936
rect 1992 -948 1998 -942
rect 1992 -954 1998 -948
rect 1992 -960 1998 -954
rect 1992 -966 1998 -960
rect 1992 -972 1998 -966
rect 1992 -978 1998 -972
rect 1992 -984 1998 -978
rect 1992 -990 1998 -984
rect 1992 -996 1998 -990
rect 1992 -1002 1998 -996
rect 1992 -1008 1998 -1002
rect 1992 -1014 1998 -1008
rect 1992 -1020 1998 -1014
rect 1992 -1026 1998 -1020
rect 1992 -1032 1998 -1026
rect 1992 -1038 1998 -1032
rect 1992 -1044 1998 -1038
rect 1992 -1050 1998 -1044
rect 1992 -1056 1998 -1050
rect 1992 -1062 1998 -1056
rect 1992 -1068 1998 -1062
rect 1992 -1074 1998 -1068
rect 1992 -1080 1998 -1074
rect 1992 -1086 1998 -1080
rect 1992 -1092 1998 -1086
rect 1992 -1098 1998 -1092
rect 1992 -1104 1998 -1098
rect 1992 -1110 1998 -1104
rect 1992 -1116 1998 -1110
rect 1992 -1122 1998 -1116
rect 1992 -1128 1998 -1122
rect 1992 -1134 1998 -1128
rect 1992 -1140 1998 -1134
rect 1992 -1146 1998 -1140
rect 1992 -1152 1998 -1146
rect 1992 -1158 1998 -1152
rect 1992 -1164 1998 -1158
rect 1992 -1170 1998 -1164
rect 1992 -1176 1998 -1170
rect 1992 -1182 1998 -1176
rect 1992 -1188 1998 -1182
rect 1992 -1194 1998 -1188
rect 1992 -1200 1998 -1194
rect 1992 -1206 1998 -1200
rect 1992 -1212 1998 -1206
rect 1992 -1218 1998 -1212
rect 1992 -1224 1998 -1218
rect 1992 -1230 1998 -1224
rect 1992 -1236 1998 -1230
rect 1992 -1242 1998 -1236
rect 1992 -1248 1998 -1242
rect 1992 -1254 1998 -1248
rect 1992 -1260 1998 -1254
rect 1992 -1266 1998 -1260
rect 1992 -1272 1998 -1266
rect 1992 -1278 1998 -1272
rect 1992 -1284 1998 -1278
rect 1992 -1290 1998 -1284
rect 1992 -1296 1998 -1290
rect 1992 -1302 1998 -1296
rect 1992 -1308 1998 -1302
rect 1992 -1314 1998 -1308
rect 1992 -1320 1998 -1314
rect 1992 -1326 1998 -1320
rect 1992 -1332 1998 -1326
rect 1992 -1338 1998 -1332
rect 1992 -1344 1998 -1338
rect 1992 -1350 1998 -1344
rect 1992 -1356 1998 -1350
rect 1992 -1362 1998 -1356
rect 1992 -1368 1998 -1362
rect 1992 -1374 1998 -1368
rect 1992 -1380 1998 -1374
rect 1992 -1386 1998 -1380
rect 1992 -1392 1998 -1386
rect 1992 -1398 1998 -1392
rect 1992 -1404 1998 -1398
rect 1992 -1410 1998 -1404
rect 1992 -1416 1998 -1410
rect 1992 -1422 1998 -1416
rect 1992 -1428 1998 -1422
rect 1992 -1434 1998 -1428
rect 1992 -1440 1998 -1434
rect 1992 -1446 1998 -1440
rect 1992 -1452 1998 -1446
rect 1992 -1458 1998 -1452
rect 1992 -1464 1998 -1458
rect 1992 -1470 1998 -1464
rect 1992 -1476 1998 -1470
rect 1992 -1482 1998 -1476
rect 1992 -1488 1998 -1482
rect 1992 -1494 1998 -1488
rect 1992 -1500 1998 -1494
rect 1992 -1506 1998 -1500
rect 1992 -1512 1998 -1506
rect 1992 -1518 1998 -1512
rect 1992 -1524 1998 -1518
rect 1992 -1530 1998 -1524
rect 1992 -1536 1998 -1530
rect 1992 -1542 1998 -1536
rect 1992 -1548 1998 -1542
rect 1992 -1554 1998 -1548
rect 1992 -1560 1998 -1554
rect 1992 -1566 1998 -1560
rect 1992 -1572 1998 -1566
rect 1992 -1578 1998 -1572
rect 1992 -1584 1998 -1578
rect 1992 -1590 1998 -1584
rect 1992 -1596 1998 -1590
rect 1992 -1602 1998 -1596
rect 1992 -1608 1998 -1602
rect 1992 -1614 1998 -1608
rect 1992 -1620 1998 -1614
rect 1992 -1626 1998 -1620
rect 1992 -1632 1998 -1626
rect 1992 -1638 1998 -1632
rect 1992 -1644 1998 -1638
rect 1992 -1650 1998 -1644
rect 1992 -1740 1998 -1734
rect 1992 -1746 1998 -1740
rect 1992 -1752 1998 -1746
rect 1992 -1758 1998 -1752
rect 1992 -1764 1998 -1758
rect 1992 -1770 1998 -1764
rect 1992 -1776 1998 -1770
rect 1992 -1782 1998 -1776
rect 1992 -1788 1998 -1782
rect 1992 -1794 1998 -1788
rect 1992 -1800 1998 -1794
rect 1992 -1806 1998 -1800
rect 1992 -1812 1998 -1806
rect 1992 -1818 1998 -1812
rect 1992 -1824 1998 -1818
rect 1992 -1830 1998 -1824
rect 1992 -1836 1998 -1830
rect 1992 -1842 1998 -1836
rect 1992 -1848 1998 -1842
rect 1992 -1854 1998 -1848
rect 1992 -1860 1998 -1854
rect 1992 -1866 1998 -1860
rect 1992 -1872 1998 -1866
rect 1992 -1878 1998 -1872
rect 1992 -1884 1998 -1878
rect 1992 -1890 1998 -1884
rect 1992 -1896 1998 -1890
rect 1992 -1902 1998 -1896
rect 1992 -1908 1998 -1902
rect 1992 -1914 1998 -1908
rect 1992 -1920 1998 -1914
rect 1992 -1926 1998 -1920
rect 1992 -1932 1998 -1926
rect 1992 -1938 1998 -1932
rect 1992 -1944 1998 -1938
rect 1992 -1950 1998 -1944
rect 1992 -1956 1998 -1950
rect 1992 -1962 1998 -1956
rect 1992 -1968 1998 -1962
rect 1992 -1974 1998 -1968
rect 1992 -1980 1998 -1974
rect 1992 -1986 1998 -1980
rect 1992 -1992 1998 -1986
rect 1992 -1998 1998 -1992
rect 1992 -2004 1998 -1998
rect 1992 -2010 1998 -2004
rect 1992 -2016 1998 -2010
rect 1992 -2022 1998 -2016
rect 1992 -2028 1998 -2022
rect 1992 -2034 1998 -2028
rect 1992 -2040 1998 -2034
rect 1992 -2046 1998 -2040
rect 1992 -2052 1998 -2046
rect 1992 -2058 1998 -2052
rect 1992 -2064 1998 -2058
rect 1992 -2070 1998 -2064
rect 1992 -2076 1998 -2070
rect 1992 -2082 1998 -2076
rect 1992 -2088 1998 -2082
rect 1992 -2094 1998 -2088
rect 1992 -2100 1998 -2094
rect 1992 -2106 1998 -2100
rect 1992 -2112 1998 -2106
rect 1992 -2118 1998 -2112
rect 1992 -2124 1998 -2118
rect 1992 -2130 1998 -2124
rect 1992 -2136 1998 -2130
rect 1992 -2142 1998 -2136
rect 1992 -2148 1998 -2142
rect 1992 -2154 1998 -2148
rect 1992 -2160 1998 -2154
rect 1992 -2166 1998 -2160
rect 1992 -2172 1998 -2166
rect 1992 -2178 1998 -2172
rect 1992 -2184 1998 -2178
rect 1992 -2190 1998 -2184
rect 1992 -2196 1998 -2190
rect 1992 -2202 1998 -2196
rect 1992 -2208 1998 -2202
rect 1992 -2214 1998 -2208
rect 1992 -2220 1998 -2214
rect 1992 -2226 1998 -2220
rect 1992 -2232 1998 -2226
rect 1992 -2238 1998 -2232
rect 1992 -2244 1998 -2238
rect 1992 -2250 1998 -2244
rect 1992 -2256 1998 -2250
rect 1992 -2262 1998 -2256
rect 1992 -2268 1998 -2262
rect 1992 -2274 1998 -2268
rect 1992 -2280 1998 -2274
rect 1992 -2286 1998 -2280
rect 1992 -2292 1998 -2286
rect 1992 -2298 1998 -2292
rect 1992 -2304 1998 -2298
rect 1992 -2310 1998 -2304
rect 1992 -2316 1998 -2310
rect 1992 -2322 1998 -2316
rect 1992 -2328 1998 -2322
rect 1992 -2334 1998 -2328
rect 1992 -2340 1998 -2334
rect 1992 -2346 1998 -2340
rect 1992 -2352 1998 -2346
rect 1992 -2358 1998 -2352
rect 1992 -2364 1998 -2358
rect 1992 -2370 1998 -2364
rect 1992 -2376 1998 -2370
rect 1992 -2382 1998 -2376
rect 1992 -2388 1998 -2382
rect 1992 -2394 1998 -2388
rect 1992 -2400 1998 -2394
rect 1992 -2406 1998 -2400
rect 1992 -2412 1998 -2406
rect 1992 -2418 1998 -2412
rect 1992 -2424 1998 -2418
rect 1992 -2430 1998 -2424
rect 1992 -2436 1998 -2430
rect 1992 -2442 1998 -2436
rect 1992 -2448 1998 -2442
rect 1992 -2454 1998 -2448
rect 1992 -2460 1998 -2454
rect 1992 -2466 1998 -2460
rect 1992 -2472 1998 -2466
rect 1992 -2478 1998 -2472
rect 1992 -2484 1998 -2478
rect 1992 -2490 1998 -2484
rect 1992 -2496 1998 -2490
rect 1992 -2502 1998 -2496
rect 1992 -2508 1998 -2502
rect 1992 -2514 1998 -2508
rect 1992 -2520 1998 -2514
rect 1992 -2526 1998 -2520
rect 1992 -2532 1998 -2526
rect 1992 -2616 1998 -2610
rect 1992 -2622 1998 -2616
rect 1992 -2628 1998 -2622
rect 1992 -2634 1998 -2628
rect 1992 -2640 1998 -2634
rect 1992 -2646 1998 -2640
rect 1992 -2652 1998 -2646
rect 1992 -2658 1998 -2652
rect 1992 -2664 1998 -2658
rect 1992 -2670 1998 -2664
rect 1992 -2676 1998 -2670
rect 1992 -2682 1998 -2676
rect 1992 -2688 1998 -2682
rect 1992 -2694 1998 -2688
rect 1992 -2700 1998 -2694
rect 1992 -2706 1998 -2700
rect 1992 -2712 1998 -2706
rect 1992 -2718 1998 -2712
rect 1992 -2724 1998 -2718
rect 1992 -2730 1998 -2724
rect 1992 -2736 1998 -2730
rect 1992 -2742 1998 -2736
rect 1992 -2748 1998 -2742
rect 1992 -2754 1998 -2748
rect 1992 -2760 1998 -2754
rect 1992 -2766 1998 -2760
rect 1992 -2772 1998 -2766
rect 1992 -2778 1998 -2772
rect 1992 -2784 1998 -2778
rect 1992 -2790 1998 -2784
rect 1992 -2796 1998 -2790
rect 1992 -2802 1998 -2796
rect 1992 -2808 1998 -2802
rect 1992 -2814 1998 -2808
rect 1992 -2820 1998 -2814
rect 1992 -2826 1998 -2820
rect 1992 -2832 1998 -2826
rect 1992 -2838 1998 -2832
rect 1992 -2844 1998 -2838
rect 1992 -2850 1998 -2844
rect 1992 -2856 1998 -2850
rect 1992 -2862 1998 -2856
rect 1992 -2868 1998 -2862
rect 1992 -2874 1998 -2868
rect 1992 -2880 1998 -2874
rect 1992 -2886 1998 -2880
rect 1992 -2892 1998 -2886
rect 1992 -2898 1998 -2892
rect 1992 -2904 1998 -2898
rect 1992 -2910 1998 -2904
rect 1992 -2916 1998 -2910
rect 1992 -2922 1998 -2916
rect 1992 -2928 1998 -2922
rect 1992 -2934 1998 -2928
rect 1992 -2940 1998 -2934
rect 1992 -2946 1998 -2940
rect 1992 -2952 1998 -2946
rect 1992 -2958 1998 -2952
rect 1992 -2964 1998 -2958
rect 1992 -2970 1998 -2964
rect 1992 -2976 1998 -2970
rect 1992 -2982 1998 -2976
rect 1992 -2988 1998 -2982
rect 1992 -2994 1998 -2988
rect 1992 -3000 1998 -2994
rect 1992 -3006 1998 -3000
rect 1992 -3012 1998 -3006
rect 1992 -3018 1998 -3012
rect 1992 -3024 1998 -3018
rect 1992 -3030 1998 -3024
rect 1992 -3036 1998 -3030
rect 1992 -3042 1998 -3036
rect 1992 -3048 1998 -3042
rect 1992 -3054 1998 -3048
rect 1992 -3060 1998 -3054
rect 1992 -3066 1998 -3060
rect 1992 -3072 1998 -3066
rect 1992 -3078 1998 -3072
rect 1992 -3084 1998 -3078
rect 1992 -3090 1998 -3084
rect 1992 -3096 1998 -3090
rect 1992 -3102 1998 -3096
rect 1992 -3108 1998 -3102
rect 1992 -3162 1998 -3156
rect 1992 -3168 1998 -3162
rect 1992 -3174 1998 -3168
rect 1992 -3180 1998 -3174
rect 1992 -3186 1998 -3180
rect 1992 -3192 1998 -3186
rect 1992 -3198 1998 -3192
rect 1992 -3204 1998 -3198
rect 1992 -3210 1998 -3204
rect 1992 -3216 1998 -3210
rect 1992 -3222 1998 -3216
rect 1992 -3228 1998 -3222
rect 1998 -456 2004 -450
rect 1998 -462 2004 -456
rect 1998 -468 2004 -462
rect 1998 -474 2004 -468
rect 1998 -480 2004 -474
rect 1998 -486 2004 -480
rect 1998 -492 2004 -486
rect 1998 -498 2004 -492
rect 1998 -504 2004 -498
rect 1998 -510 2004 -504
rect 1998 -516 2004 -510
rect 1998 -522 2004 -516
rect 1998 -528 2004 -522
rect 1998 -534 2004 -528
rect 1998 -540 2004 -534
rect 1998 -546 2004 -540
rect 1998 -552 2004 -546
rect 1998 -558 2004 -552
rect 1998 -564 2004 -558
rect 1998 -570 2004 -564
rect 1998 -576 2004 -570
rect 1998 -582 2004 -576
rect 1998 -588 2004 -582
rect 1998 -594 2004 -588
rect 1998 -600 2004 -594
rect 1998 -606 2004 -600
rect 1998 -612 2004 -606
rect 1998 -618 2004 -612
rect 1998 -624 2004 -618
rect 1998 -630 2004 -624
rect 1998 -636 2004 -630
rect 1998 -642 2004 -636
rect 1998 -648 2004 -642
rect 1998 -654 2004 -648
rect 1998 -660 2004 -654
rect 1998 -666 2004 -660
rect 1998 -672 2004 -666
rect 1998 -678 2004 -672
rect 1998 -684 2004 -678
rect 1998 -690 2004 -684
rect 1998 -696 2004 -690
rect 1998 -702 2004 -696
rect 1998 -708 2004 -702
rect 1998 -714 2004 -708
rect 1998 -720 2004 -714
rect 1998 -726 2004 -720
rect 1998 -732 2004 -726
rect 1998 -738 2004 -732
rect 1998 -744 2004 -738
rect 1998 -750 2004 -744
rect 1998 -756 2004 -750
rect 1998 -762 2004 -756
rect 1998 -768 2004 -762
rect 1998 -774 2004 -768
rect 1998 -780 2004 -774
rect 1998 -786 2004 -780
rect 1998 -792 2004 -786
rect 1998 -798 2004 -792
rect 1998 -804 2004 -798
rect 1998 -810 2004 -804
rect 1998 -816 2004 -810
rect 1998 -822 2004 -816
rect 1998 -828 2004 -822
rect 1998 -834 2004 -828
rect 1998 -840 2004 -834
rect 1998 -846 2004 -840
rect 1998 -852 2004 -846
rect 1998 -858 2004 -852
rect 1998 -864 2004 -858
rect 1998 -870 2004 -864
rect 1998 -876 2004 -870
rect 1998 -882 2004 -876
rect 1998 -888 2004 -882
rect 1998 -894 2004 -888
rect 1998 -900 2004 -894
rect 1998 -906 2004 -900
rect 1998 -912 2004 -906
rect 1998 -918 2004 -912
rect 1998 -924 2004 -918
rect 1998 -930 2004 -924
rect 1998 -936 2004 -930
rect 1998 -942 2004 -936
rect 1998 -948 2004 -942
rect 1998 -954 2004 -948
rect 1998 -960 2004 -954
rect 1998 -966 2004 -960
rect 1998 -972 2004 -966
rect 1998 -978 2004 -972
rect 1998 -984 2004 -978
rect 1998 -990 2004 -984
rect 1998 -996 2004 -990
rect 1998 -1002 2004 -996
rect 1998 -1008 2004 -1002
rect 1998 -1014 2004 -1008
rect 1998 -1020 2004 -1014
rect 1998 -1026 2004 -1020
rect 1998 -1032 2004 -1026
rect 1998 -1038 2004 -1032
rect 1998 -1044 2004 -1038
rect 1998 -1050 2004 -1044
rect 1998 -1056 2004 -1050
rect 1998 -1062 2004 -1056
rect 1998 -1068 2004 -1062
rect 1998 -1074 2004 -1068
rect 1998 -1080 2004 -1074
rect 1998 -1086 2004 -1080
rect 1998 -1092 2004 -1086
rect 1998 -1098 2004 -1092
rect 1998 -1104 2004 -1098
rect 1998 -1110 2004 -1104
rect 1998 -1116 2004 -1110
rect 1998 -1122 2004 -1116
rect 1998 -1128 2004 -1122
rect 1998 -1134 2004 -1128
rect 1998 -1140 2004 -1134
rect 1998 -1146 2004 -1140
rect 1998 -1152 2004 -1146
rect 1998 -1158 2004 -1152
rect 1998 -1164 2004 -1158
rect 1998 -1170 2004 -1164
rect 1998 -1176 2004 -1170
rect 1998 -1182 2004 -1176
rect 1998 -1188 2004 -1182
rect 1998 -1194 2004 -1188
rect 1998 -1200 2004 -1194
rect 1998 -1206 2004 -1200
rect 1998 -1212 2004 -1206
rect 1998 -1218 2004 -1212
rect 1998 -1224 2004 -1218
rect 1998 -1230 2004 -1224
rect 1998 -1236 2004 -1230
rect 1998 -1242 2004 -1236
rect 1998 -1248 2004 -1242
rect 1998 -1254 2004 -1248
rect 1998 -1260 2004 -1254
rect 1998 -1266 2004 -1260
rect 1998 -1272 2004 -1266
rect 1998 -1278 2004 -1272
rect 1998 -1284 2004 -1278
rect 1998 -1290 2004 -1284
rect 1998 -1296 2004 -1290
rect 1998 -1302 2004 -1296
rect 1998 -1308 2004 -1302
rect 1998 -1314 2004 -1308
rect 1998 -1320 2004 -1314
rect 1998 -1326 2004 -1320
rect 1998 -1332 2004 -1326
rect 1998 -1338 2004 -1332
rect 1998 -1344 2004 -1338
rect 1998 -1350 2004 -1344
rect 1998 -1356 2004 -1350
rect 1998 -1362 2004 -1356
rect 1998 -1368 2004 -1362
rect 1998 -1374 2004 -1368
rect 1998 -1380 2004 -1374
rect 1998 -1386 2004 -1380
rect 1998 -1392 2004 -1386
rect 1998 -1398 2004 -1392
rect 1998 -1404 2004 -1398
rect 1998 -1410 2004 -1404
rect 1998 -1416 2004 -1410
rect 1998 -1422 2004 -1416
rect 1998 -1428 2004 -1422
rect 1998 -1434 2004 -1428
rect 1998 -1440 2004 -1434
rect 1998 -1446 2004 -1440
rect 1998 -1452 2004 -1446
rect 1998 -1458 2004 -1452
rect 1998 -1464 2004 -1458
rect 1998 -1470 2004 -1464
rect 1998 -1476 2004 -1470
rect 1998 -1482 2004 -1476
rect 1998 -1488 2004 -1482
rect 1998 -1494 2004 -1488
rect 1998 -1500 2004 -1494
rect 1998 -1506 2004 -1500
rect 1998 -1512 2004 -1506
rect 1998 -1518 2004 -1512
rect 1998 -1524 2004 -1518
rect 1998 -1530 2004 -1524
rect 1998 -1536 2004 -1530
rect 1998 -1542 2004 -1536
rect 1998 -1548 2004 -1542
rect 1998 -1554 2004 -1548
rect 1998 -1560 2004 -1554
rect 1998 -1566 2004 -1560
rect 1998 -1572 2004 -1566
rect 1998 -1578 2004 -1572
rect 1998 -1584 2004 -1578
rect 1998 -1590 2004 -1584
rect 1998 -1596 2004 -1590
rect 1998 -1602 2004 -1596
rect 1998 -1608 2004 -1602
rect 1998 -1614 2004 -1608
rect 1998 -1620 2004 -1614
rect 1998 -1626 2004 -1620
rect 1998 -1632 2004 -1626
rect 1998 -1638 2004 -1632
rect 1998 -1644 2004 -1638
rect 1998 -1734 2004 -1728
rect 1998 -1740 2004 -1734
rect 1998 -1746 2004 -1740
rect 1998 -1752 2004 -1746
rect 1998 -1758 2004 -1752
rect 1998 -1764 2004 -1758
rect 1998 -1770 2004 -1764
rect 1998 -1776 2004 -1770
rect 1998 -1782 2004 -1776
rect 1998 -1788 2004 -1782
rect 1998 -1794 2004 -1788
rect 1998 -1800 2004 -1794
rect 1998 -1806 2004 -1800
rect 1998 -1812 2004 -1806
rect 1998 -1818 2004 -1812
rect 1998 -1824 2004 -1818
rect 1998 -1830 2004 -1824
rect 1998 -1836 2004 -1830
rect 1998 -1842 2004 -1836
rect 1998 -1848 2004 -1842
rect 1998 -1854 2004 -1848
rect 1998 -1860 2004 -1854
rect 1998 -1866 2004 -1860
rect 1998 -1872 2004 -1866
rect 1998 -1878 2004 -1872
rect 1998 -1884 2004 -1878
rect 1998 -1890 2004 -1884
rect 1998 -1896 2004 -1890
rect 1998 -1902 2004 -1896
rect 1998 -1908 2004 -1902
rect 1998 -1914 2004 -1908
rect 1998 -1920 2004 -1914
rect 1998 -1926 2004 -1920
rect 1998 -1932 2004 -1926
rect 1998 -1938 2004 -1932
rect 1998 -1944 2004 -1938
rect 1998 -1950 2004 -1944
rect 1998 -1956 2004 -1950
rect 1998 -1962 2004 -1956
rect 1998 -1968 2004 -1962
rect 1998 -1974 2004 -1968
rect 1998 -1980 2004 -1974
rect 1998 -1986 2004 -1980
rect 1998 -1992 2004 -1986
rect 1998 -1998 2004 -1992
rect 1998 -2004 2004 -1998
rect 1998 -2010 2004 -2004
rect 1998 -2016 2004 -2010
rect 1998 -2022 2004 -2016
rect 1998 -2028 2004 -2022
rect 1998 -2034 2004 -2028
rect 1998 -2040 2004 -2034
rect 1998 -2046 2004 -2040
rect 1998 -2052 2004 -2046
rect 1998 -2058 2004 -2052
rect 1998 -2064 2004 -2058
rect 1998 -2070 2004 -2064
rect 1998 -2076 2004 -2070
rect 1998 -2082 2004 -2076
rect 1998 -2088 2004 -2082
rect 1998 -2094 2004 -2088
rect 1998 -2100 2004 -2094
rect 1998 -2106 2004 -2100
rect 1998 -2112 2004 -2106
rect 1998 -2118 2004 -2112
rect 1998 -2124 2004 -2118
rect 1998 -2130 2004 -2124
rect 1998 -2136 2004 -2130
rect 1998 -2142 2004 -2136
rect 1998 -2148 2004 -2142
rect 1998 -2154 2004 -2148
rect 1998 -2160 2004 -2154
rect 1998 -2166 2004 -2160
rect 1998 -2172 2004 -2166
rect 1998 -2178 2004 -2172
rect 1998 -2184 2004 -2178
rect 1998 -2190 2004 -2184
rect 1998 -2196 2004 -2190
rect 1998 -2202 2004 -2196
rect 1998 -2208 2004 -2202
rect 1998 -2214 2004 -2208
rect 1998 -2220 2004 -2214
rect 1998 -2226 2004 -2220
rect 1998 -2232 2004 -2226
rect 1998 -2238 2004 -2232
rect 1998 -2244 2004 -2238
rect 1998 -2250 2004 -2244
rect 1998 -2256 2004 -2250
rect 1998 -2262 2004 -2256
rect 1998 -2268 2004 -2262
rect 1998 -2274 2004 -2268
rect 1998 -2280 2004 -2274
rect 1998 -2286 2004 -2280
rect 1998 -2292 2004 -2286
rect 1998 -2298 2004 -2292
rect 1998 -2304 2004 -2298
rect 1998 -2310 2004 -2304
rect 1998 -2316 2004 -2310
rect 1998 -2322 2004 -2316
rect 1998 -2328 2004 -2322
rect 1998 -2334 2004 -2328
rect 1998 -2340 2004 -2334
rect 1998 -2346 2004 -2340
rect 1998 -2352 2004 -2346
rect 1998 -2358 2004 -2352
rect 1998 -2364 2004 -2358
rect 1998 -2370 2004 -2364
rect 1998 -2376 2004 -2370
rect 1998 -2382 2004 -2376
rect 1998 -2388 2004 -2382
rect 1998 -2394 2004 -2388
rect 1998 -2400 2004 -2394
rect 1998 -2406 2004 -2400
rect 1998 -2412 2004 -2406
rect 1998 -2418 2004 -2412
rect 1998 -2424 2004 -2418
rect 1998 -2430 2004 -2424
rect 1998 -2436 2004 -2430
rect 1998 -2442 2004 -2436
rect 1998 -2448 2004 -2442
rect 1998 -2454 2004 -2448
rect 1998 -2460 2004 -2454
rect 1998 -2466 2004 -2460
rect 1998 -2472 2004 -2466
rect 1998 -2478 2004 -2472
rect 1998 -2484 2004 -2478
rect 1998 -2490 2004 -2484
rect 1998 -2496 2004 -2490
rect 1998 -2502 2004 -2496
rect 1998 -2508 2004 -2502
rect 1998 -2514 2004 -2508
rect 1998 -2520 2004 -2514
rect 1998 -2526 2004 -2520
rect 1998 -2610 2004 -2604
rect 1998 -2616 2004 -2610
rect 1998 -2622 2004 -2616
rect 1998 -2628 2004 -2622
rect 1998 -2634 2004 -2628
rect 1998 -2640 2004 -2634
rect 1998 -2646 2004 -2640
rect 1998 -2652 2004 -2646
rect 1998 -2658 2004 -2652
rect 1998 -2664 2004 -2658
rect 1998 -2670 2004 -2664
rect 1998 -2676 2004 -2670
rect 1998 -2682 2004 -2676
rect 1998 -2688 2004 -2682
rect 1998 -2694 2004 -2688
rect 1998 -2700 2004 -2694
rect 1998 -2706 2004 -2700
rect 1998 -2712 2004 -2706
rect 1998 -2718 2004 -2712
rect 1998 -2724 2004 -2718
rect 1998 -2730 2004 -2724
rect 1998 -2736 2004 -2730
rect 1998 -2742 2004 -2736
rect 1998 -2748 2004 -2742
rect 1998 -2754 2004 -2748
rect 1998 -2760 2004 -2754
rect 1998 -2766 2004 -2760
rect 1998 -2772 2004 -2766
rect 1998 -2778 2004 -2772
rect 1998 -2784 2004 -2778
rect 1998 -2790 2004 -2784
rect 1998 -2796 2004 -2790
rect 1998 -2802 2004 -2796
rect 1998 -2808 2004 -2802
rect 1998 -2814 2004 -2808
rect 1998 -2820 2004 -2814
rect 1998 -2826 2004 -2820
rect 1998 -2832 2004 -2826
rect 1998 -2838 2004 -2832
rect 1998 -2844 2004 -2838
rect 1998 -2850 2004 -2844
rect 1998 -2856 2004 -2850
rect 1998 -2862 2004 -2856
rect 1998 -2868 2004 -2862
rect 1998 -2874 2004 -2868
rect 1998 -2880 2004 -2874
rect 1998 -2886 2004 -2880
rect 1998 -2892 2004 -2886
rect 1998 -2898 2004 -2892
rect 1998 -2904 2004 -2898
rect 1998 -2910 2004 -2904
rect 1998 -2916 2004 -2910
rect 1998 -2922 2004 -2916
rect 1998 -2928 2004 -2922
rect 1998 -2934 2004 -2928
rect 1998 -2940 2004 -2934
rect 1998 -2946 2004 -2940
rect 1998 -2952 2004 -2946
rect 1998 -2958 2004 -2952
rect 1998 -2964 2004 -2958
rect 1998 -2970 2004 -2964
rect 1998 -2976 2004 -2970
rect 1998 -2982 2004 -2976
rect 1998 -2988 2004 -2982
rect 1998 -2994 2004 -2988
rect 1998 -3000 2004 -2994
rect 1998 -3006 2004 -3000
rect 1998 -3012 2004 -3006
rect 1998 -3018 2004 -3012
rect 1998 -3024 2004 -3018
rect 1998 -3030 2004 -3024
rect 1998 -3036 2004 -3030
rect 1998 -3042 2004 -3036
rect 1998 -3048 2004 -3042
rect 1998 -3054 2004 -3048
rect 1998 -3060 2004 -3054
rect 1998 -3066 2004 -3060
rect 1998 -3072 2004 -3066
rect 1998 -3078 2004 -3072
rect 1998 -3084 2004 -3078
rect 1998 -3090 2004 -3084
rect 1998 -3096 2004 -3090
rect 1998 -3102 2004 -3096
rect 1998 -3162 2004 -3156
rect 1998 -3168 2004 -3162
rect 1998 -3174 2004 -3168
rect 1998 -3180 2004 -3174
rect 1998 -3186 2004 -3180
rect 1998 -3192 2004 -3186
rect 1998 -3198 2004 -3192
rect 1998 -3204 2004 -3198
rect 1998 -3210 2004 -3204
rect 1998 -3216 2004 -3210
rect 1998 -3222 2004 -3216
rect 2004 -444 2010 -438
rect 2004 -450 2010 -444
rect 2004 -456 2010 -450
rect 2004 -462 2010 -456
rect 2004 -468 2010 -462
rect 2004 -474 2010 -468
rect 2004 -480 2010 -474
rect 2004 -486 2010 -480
rect 2004 -492 2010 -486
rect 2004 -498 2010 -492
rect 2004 -504 2010 -498
rect 2004 -510 2010 -504
rect 2004 -516 2010 -510
rect 2004 -522 2010 -516
rect 2004 -528 2010 -522
rect 2004 -534 2010 -528
rect 2004 -540 2010 -534
rect 2004 -546 2010 -540
rect 2004 -552 2010 -546
rect 2004 -558 2010 -552
rect 2004 -564 2010 -558
rect 2004 -570 2010 -564
rect 2004 -576 2010 -570
rect 2004 -582 2010 -576
rect 2004 -588 2010 -582
rect 2004 -594 2010 -588
rect 2004 -600 2010 -594
rect 2004 -606 2010 -600
rect 2004 -612 2010 -606
rect 2004 -618 2010 -612
rect 2004 -624 2010 -618
rect 2004 -630 2010 -624
rect 2004 -636 2010 -630
rect 2004 -642 2010 -636
rect 2004 -648 2010 -642
rect 2004 -654 2010 -648
rect 2004 -660 2010 -654
rect 2004 -666 2010 -660
rect 2004 -672 2010 -666
rect 2004 -678 2010 -672
rect 2004 -684 2010 -678
rect 2004 -690 2010 -684
rect 2004 -696 2010 -690
rect 2004 -702 2010 -696
rect 2004 -708 2010 -702
rect 2004 -714 2010 -708
rect 2004 -720 2010 -714
rect 2004 -726 2010 -720
rect 2004 -732 2010 -726
rect 2004 -738 2010 -732
rect 2004 -744 2010 -738
rect 2004 -750 2010 -744
rect 2004 -756 2010 -750
rect 2004 -762 2010 -756
rect 2004 -768 2010 -762
rect 2004 -774 2010 -768
rect 2004 -780 2010 -774
rect 2004 -786 2010 -780
rect 2004 -792 2010 -786
rect 2004 -798 2010 -792
rect 2004 -804 2010 -798
rect 2004 -810 2010 -804
rect 2004 -816 2010 -810
rect 2004 -822 2010 -816
rect 2004 -828 2010 -822
rect 2004 -834 2010 -828
rect 2004 -840 2010 -834
rect 2004 -846 2010 -840
rect 2004 -852 2010 -846
rect 2004 -858 2010 -852
rect 2004 -864 2010 -858
rect 2004 -870 2010 -864
rect 2004 -876 2010 -870
rect 2004 -882 2010 -876
rect 2004 -888 2010 -882
rect 2004 -894 2010 -888
rect 2004 -900 2010 -894
rect 2004 -906 2010 -900
rect 2004 -912 2010 -906
rect 2004 -918 2010 -912
rect 2004 -924 2010 -918
rect 2004 -930 2010 -924
rect 2004 -936 2010 -930
rect 2004 -942 2010 -936
rect 2004 -948 2010 -942
rect 2004 -954 2010 -948
rect 2004 -960 2010 -954
rect 2004 -966 2010 -960
rect 2004 -972 2010 -966
rect 2004 -978 2010 -972
rect 2004 -984 2010 -978
rect 2004 -990 2010 -984
rect 2004 -996 2010 -990
rect 2004 -1002 2010 -996
rect 2004 -1008 2010 -1002
rect 2004 -1014 2010 -1008
rect 2004 -1020 2010 -1014
rect 2004 -1026 2010 -1020
rect 2004 -1032 2010 -1026
rect 2004 -1038 2010 -1032
rect 2004 -1044 2010 -1038
rect 2004 -1050 2010 -1044
rect 2004 -1056 2010 -1050
rect 2004 -1062 2010 -1056
rect 2004 -1068 2010 -1062
rect 2004 -1074 2010 -1068
rect 2004 -1080 2010 -1074
rect 2004 -1086 2010 -1080
rect 2004 -1092 2010 -1086
rect 2004 -1098 2010 -1092
rect 2004 -1104 2010 -1098
rect 2004 -1110 2010 -1104
rect 2004 -1116 2010 -1110
rect 2004 -1122 2010 -1116
rect 2004 -1128 2010 -1122
rect 2004 -1134 2010 -1128
rect 2004 -1140 2010 -1134
rect 2004 -1146 2010 -1140
rect 2004 -1152 2010 -1146
rect 2004 -1158 2010 -1152
rect 2004 -1164 2010 -1158
rect 2004 -1170 2010 -1164
rect 2004 -1176 2010 -1170
rect 2004 -1182 2010 -1176
rect 2004 -1188 2010 -1182
rect 2004 -1194 2010 -1188
rect 2004 -1200 2010 -1194
rect 2004 -1206 2010 -1200
rect 2004 -1212 2010 -1206
rect 2004 -1218 2010 -1212
rect 2004 -1224 2010 -1218
rect 2004 -1230 2010 -1224
rect 2004 -1236 2010 -1230
rect 2004 -1242 2010 -1236
rect 2004 -1248 2010 -1242
rect 2004 -1254 2010 -1248
rect 2004 -1260 2010 -1254
rect 2004 -1266 2010 -1260
rect 2004 -1272 2010 -1266
rect 2004 -1278 2010 -1272
rect 2004 -1284 2010 -1278
rect 2004 -1290 2010 -1284
rect 2004 -1296 2010 -1290
rect 2004 -1302 2010 -1296
rect 2004 -1308 2010 -1302
rect 2004 -1314 2010 -1308
rect 2004 -1320 2010 -1314
rect 2004 -1326 2010 -1320
rect 2004 -1332 2010 -1326
rect 2004 -1338 2010 -1332
rect 2004 -1344 2010 -1338
rect 2004 -1350 2010 -1344
rect 2004 -1356 2010 -1350
rect 2004 -1362 2010 -1356
rect 2004 -1368 2010 -1362
rect 2004 -1374 2010 -1368
rect 2004 -1380 2010 -1374
rect 2004 -1386 2010 -1380
rect 2004 -1392 2010 -1386
rect 2004 -1398 2010 -1392
rect 2004 -1404 2010 -1398
rect 2004 -1410 2010 -1404
rect 2004 -1416 2010 -1410
rect 2004 -1422 2010 -1416
rect 2004 -1428 2010 -1422
rect 2004 -1434 2010 -1428
rect 2004 -1440 2010 -1434
rect 2004 -1446 2010 -1440
rect 2004 -1452 2010 -1446
rect 2004 -1458 2010 -1452
rect 2004 -1464 2010 -1458
rect 2004 -1470 2010 -1464
rect 2004 -1476 2010 -1470
rect 2004 -1482 2010 -1476
rect 2004 -1488 2010 -1482
rect 2004 -1494 2010 -1488
rect 2004 -1500 2010 -1494
rect 2004 -1506 2010 -1500
rect 2004 -1512 2010 -1506
rect 2004 -1518 2010 -1512
rect 2004 -1524 2010 -1518
rect 2004 -1530 2010 -1524
rect 2004 -1536 2010 -1530
rect 2004 -1542 2010 -1536
rect 2004 -1548 2010 -1542
rect 2004 -1554 2010 -1548
rect 2004 -1560 2010 -1554
rect 2004 -1566 2010 -1560
rect 2004 -1572 2010 -1566
rect 2004 -1578 2010 -1572
rect 2004 -1584 2010 -1578
rect 2004 -1590 2010 -1584
rect 2004 -1596 2010 -1590
rect 2004 -1602 2010 -1596
rect 2004 -1608 2010 -1602
rect 2004 -1614 2010 -1608
rect 2004 -1620 2010 -1614
rect 2004 -1626 2010 -1620
rect 2004 -1632 2010 -1626
rect 2004 -1638 2010 -1632
rect 2004 -1728 2010 -1722
rect 2004 -1734 2010 -1728
rect 2004 -1740 2010 -1734
rect 2004 -1746 2010 -1740
rect 2004 -1752 2010 -1746
rect 2004 -1758 2010 -1752
rect 2004 -1764 2010 -1758
rect 2004 -1770 2010 -1764
rect 2004 -1776 2010 -1770
rect 2004 -1782 2010 -1776
rect 2004 -1788 2010 -1782
rect 2004 -1794 2010 -1788
rect 2004 -1800 2010 -1794
rect 2004 -1806 2010 -1800
rect 2004 -1812 2010 -1806
rect 2004 -1818 2010 -1812
rect 2004 -1824 2010 -1818
rect 2004 -1830 2010 -1824
rect 2004 -1836 2010 -1830
rect 2004 -1842 2010 -1836
rect 2004 -1848 2010 -1842
rect 2004 -1854 2010 -1848
rect 2004 -1860 2010 -1854
rect 2004 -1866 2010 -1860
rect 2004 -1872 2010 -1866
rect 2004 -1878 2010 -1872
rect 2004 -1884 2010 -1878
rect 2004 -1890 2010 -1884
rect 2004 -1896 2010 -1890
rect 2004 -1902 2010 -1896
rect 2004 -1908 2010 -1902
rect 2004 -1914 2010 -1908
rect 2004 -1920 2010 -1914
rect 2004 -1926 2010 -1920
rect 2004 -1932 2010 -1926
rect 2004 -1938 2010 -1932
rect 2004 -1944 2010 -1938
rect 2004 -1950 2010 -1944
rect 2004 -1956 2010 -1950
rect 2004 -1962 2010 -1956
rect 2004 -1968 2010 -1962
rect 2004 -1974 2010 -1968
rect 2004 -1980 2010 -1974
rect 2004 -1986 2010 -1980
rect 2004 -1992 2010 -1986
rect 2004 -1998 2010 -1992
rect 2004 -2004 2010 -1998
rect 2004 -2010 2010 -2004
rect 2004 -2016 2010 -2010
rect 2004 -2022 2010 -2016
rect 2004 -2028 2010 -2022
rect 2004 -2034 2010 -2028
rect 2004 -2040 2010 -2034
rect 2004 -2046 2010 -2040
rect 2004 -2052 2010 -2046
rect 2004 -2058 2010 -2052
rect 2004 -2064 2010 -2058
rect 2004 -2070 2010 -2064
rect 2004 -2076 2010 -2070
rect 2004 -2082 2010 -2076
rect 2004 -2088 2010 -2082
rect 2004 -2094 2010 -2088
rect 2004 -2100 2010 -2094
rect 2004 -2106 2010 -2100
rect 2004 -2112 2010 -2106
rect 2004 -2118 2010 -2112
rect 2004 -2124 2010 -2118
rect 2004 -2130 2010 -2124
rect 2004 -2136 2010 -2130
rect 2004 -2142 2010 -2136
rect 2004 -2148 2010 -2142
rect 2004 -2154 2010 -2148
rect 2004 -2160 2010 -2154
rect 2004 -2166 2010 -2160
rect 2004 -2172 2010 -2166
rect 2004 -2178 2010 -2172
rect 2004 -2184 2010 -2178
rect 2004 -2190 2010 -2184
rect 2004 -2196 2010 -2190
rect 2004 -2202 2010 -2196
rect 2004 -2208 2010 -2202
rect 2004 -2214 2010 -2208
rect 2004 -2220 2010 -2214
rect 2004 -2226 2010 -2220
rect 2004 -2232 2010 -2226
rect 2004 -2238 2010 -2232
rect 2004 -2244 2010 -2238
rect 2004 -2250 2010 -2244
rect 2004 -2256 2010 -2250
rect 2004 -2262 2010 -2256
rect 2004 -2268 2010 -2262
rect 2004 -2274 2010 -2268
rect 2004 -2280 2010 -2274
rect 2004 -2286 2010 -2280
rect 2004 -2292 2010 -2286
rect 2004 -2298 2010 -2292
rect 2004 -2304 2010 -2298
rect 2004 -2310 2010 -2304
rect 2004 -2316 2010 -2310
rect 2004 -2322 2010 -2316
rect 2004 -2328 2010 -2322
rect 2004 -2334 2010 -2328
rect 2004 -2340 2010 -2334
rect 2004 -2346 2010 -2340
rect 2004 -2352 2010 -2346
rect 2004 -2358 2010 -2352
rect 2004 -2364 2010 -2358
rect 2004 -2370 2010 -2364
rect 2004 -2376 2010 -2370
rect 2004 -2382 2010 -2376
rect 2004 -2388 2010 -2382
rect 2004 -2394 2010 -2388
rect 2004 -2400 2010 -2394
rect 2004 -2406 2010 -2400
rect 2004 -2412 2010 -2406
rect 2004 -2418 2010 -2412
rect 2004 -2424 2010 -2418
rect 2004 -2430 2010 -2424
rect 2004 -2436 2010 -2430
rect 2004 -2442 2010 -2436
rect 2004 -2448 2010 -2442
rect 2004 -2454 2010 -2448
rect 2004 -2460 2010 -2454
rect 2004 -2466 2010 -2460
rect 2004 -2472 2010 -2466
rect 2004 -2478 2010 -2472
rect 2004 -2484 2010 -2478
rect 2004 -2490 2010 -2484
rect 2004 -2496 2010 -2490
rect 2004 -2502 2010 -2496
rect 2004 -2508 2010 -2502
rect 2004 -2514 2010 -2508
rect 2004 -2520 2010 -2514
rect 2004 -2526 2010 -2520
rect 2004 -2610 2010 -2604
rect 2004 -2616 2010 -2610
rect 2004 -2622 2010 -2616
rect 2004 -2628 2010 -2622
rect 2004 -2634 2010 -2628
rect 2004 -2640 2010 -2634
rect 2004 -2646 2010 -2640
rect 2004 -2652 2010 -2646
rect 2004 -2658 2010 -2652
rect 2004 -2664 2010 -2658
rect 2004 -2670 2010 -2664
rect 2004 -2676 2010 -2670
rect 2004 -2682 2010 -2676
rect 2004 -2688 2010 -2682
rect 2004 -2694 2010 -2688
rect 2004 -2700 2010 -2694
rect 2004 -2706 2010 -2700
rect 2004 -2712 2010 -2706
rect 2004 -2718 2010 -2712
rect 2004 -2724 2010 -2718
rect 2004 -2730 2010 -2724
rect 2004 -2736 2010 -2730
rect 2004 -2742 2010 -2736
rect 2004 -2748 2010 -2742
rect 2004 -2754 2010 -2748
rect 2004 -2760 2010 -2754
rect 2004 -2766 2010 -2760
rect 2004 -2772 2010 -2766
rect 2004 -2778 2010 -2772
rect 2004 -2784 2010 -2778
rect 2004 -2790 2010 -2784
rect 2004 -2796 2010 -2790
rect 2004 -2802 2010 -2796
rect 2004 -2808 2010 -2802
rect 2004 -2814 2010 -2808
rect 2004 -2820 2010 -2814
rect 2004 -2826 2010 -2820
rect 2004 -2832 2010 -2826
rect 2004 -2838 2010 -2832
rect 2004 -2844 2010 -2838
rect 2004 -2850 2010 -2844
rect 2004 -2856 2010 -2850
rect 2004 -2862 2010 -2856
rect 2004 -2868 2010 -2862
rect 2004 -2874 2010 -2868
rect 2004 -2880 2010 -2874
rect 2004 -2886 2010 -2880
rect 2004 -2892 2010 -2886
rect 2004 -2898 2010 -2892
rect 2004 -2904 2010 -2898
rect 2004 -2910 2010 -2904
rect 2004 -2916 2010 -2910
rect 2004 -2922 2010 -2916
rect 2004 -2928 2010 -2922
rect 2004 -2934 2010 -2928
rect 2004 -2940 2010 -2934
rect 2004 -2946 2010 -2940
rect 2004 -2952 2010 -2946
rect 2004 -2958 2010 -2952
rect 2004 -2964 2010 -2958
rect 2004 -2970 2010 -2964
rect 2004 -2976 2010 -2970
rect 2004 -2982 2010 -2976
rect 2004 -2988 2010 -2982
rect 2004 -2994 2010 -2988
rect 2004 -3000 2010 -2994
rect 2004 -3006 2010 -3000
rect 2004 -3012 2010 -3006
rect 2004 -3018 2010 -3012
rect 2004 -3024 2010 -3018
rect 2004 -3030 2010 -3024
rect 2004 -3036 2010 -3030
rect 2004 -3042 2010 -3036
rect 2004 -3048 2010 -3042
rect 2004 -3054 2010 -3048
rect 2004 -3060 2010 -3054
rect 2004 -3066 2010 -3060
rect 2004 -3072 2010 -3066
rect 2004 -3078 2010 -3072
rect 2004 -3084 2010 -3078
rect 2004 -3090 2010 -3084
rect 2004 -3096 2010 -3090
rect 2004 -3102 2010 -3096
rect 2004 -3156 2010 -3150
rect 2004 -3162 2010 -3156
rect 2004 -3168 2010 -3162
rect 2004 -3174 2010 -3168
rect 2004 -3180 2010 -3174
rect 2004 -3186 2010 -3180
rect 2004 -3192 2010 -3186
rect 2004 -3198 2010 -3192
rect 2004 -3204 2010 -3198
rect 2004 -3210 2010 -3204
rect 2004 -3216 2010 -3210
rect 2010 -438 2016 -432
rect 2010 -444 2016 -438
rect 2010 -450 2016 -444
rect 2010 -456 2016 -450
rect 2010 -462 2016 -456
rect 2010 -468 2016 -462
rect 2010 -474 2016 -468
rect 2010 -480 2016 -474
rect 2010 -486 2016 -480
rect 2010 -492 2016 -486
rect 2010 -498 2016 -492
rect 2010 -504 2016 -498
rect 2010 -510 2016 -504
rect 2010 -516 2016 -510
rect 2010 -522 2016 -516
rect 2010 -528 2016 -522
rect 2010 -534 2016 -528
rect 2010 -540 2016 -534
rect 2010 -546 2016 -540
rect 2010 -552 2016 -546
rect 2010 -558 2016 -552
rect 2010 -564 2016 -558
rect 2010 -570 2016 -564
rect 2010 -576 2016 -570
rect 2010 -582 2016 -576
rect 2010 -588 2016 -582
rect 2010 -594 2016 -588
rect 2010 -600 2016 -594
rect 2010 -606 2016 -600
rect 2010 -612 2016 -606
rect 2010 -618 2016 -612
rect 2010 -624 2016 -618
rect 2010 -630 2016 -624
rect 2010 -636 2016 -630
rect 2010 -642 2016 -636
rect 2010 -648 2016 -642
rect 2010 -654 2016 -648
rect 2010 -660 2016 -654
rect 2010 -666 2016 -660
rect 2010 -672 2016 -666
rect 2010 -678 2016 -672
rect 2010 -684 2016 -678
rect 2010 -690 2016 -684
rect 2010 -696 2016 -690
rect 2010 -702 2016 -696
rect 2010 -708 2016 -702
rect 2010 -714 2016 -708
rect 2010 -720 2016 -714
rect 2010 -726 2016 -720
rect 2010 -732 2016 -726
rect 2010 -738 2016 -732
rect 2010 -744 2016 -738
rect 2010 -750 2016 -744
rect 2010 -756 2016 -750
rect 2010 -762 2016 -756
rect 2010 -768 2016 -762
rect 2010 -774 2016 -768
rect 2010 -780 2016 -774
rect 2010 -786 2016 -780
rect 2010 -792 2016 -786
rect 2010 -798 2016 -792
rect 2010 -804 2016 -798
rect 2010 -810 2016 -804
rect 2010 -816 2016 -810
rect 2010 -822 2016 -816
rect 2010 -828 2016 -822
rect 2010 -834 2016 -828
rect 2010 -840 2016 -834
rect 2010 -846 2016 -840
rect 2010 -852 2016 -846
rect 2010 -858 2016 -852
rect 2010 -864 2016 -858
rect 2010 -870 2016 -864
rect 2010 -876 2016 -870
rect 2010 -882 2016 -876
rect 2010 -888 2016 -882
rect 2010 -894 2016 -888
rect 2010 -900 2016 -894
rect 2010 -906 2016 -900
rect 2010 -912 2016 -906
rect 2010 -918 2016 -912
rect 2010 -924 2016 -918
rect 2010 -930 2016 -924
rect 2010 -936 2016 -930
rect 2010 -942 2016 -936
rect 2010 -948 2016 -942
rect 2010 -954 2016 -948
rect 2010 -960 2016 -954
rect 2010 -966 2016 -960
rect 2010 -972 2016 -966
rect 2010 -978 2016 -972
rect 2010 -984 2016 -978
rect 2010 -990 2016 -984
rect 2010 -996 2016 -990
rect 2010 -1002 2016 -996
rect 2010 -1008 2016 -1002
rect 2010 -1014 2016 -1008
rect 2010 -1020 2016 -1014
rect 2010 -1026 2016 -1020
rect 2010 -1032 2016 -1026
rect 2010 -1038 2016 -1032
rect 2010 -1044 2016 -1038
rect 2010 -1050 2016 -1044
rect 2010 -1056 2016 -1050
rect 2010 -1062 2016 -1056
rect 2010 -1068 2016 -1062
rect 2010 -1074 2016 -1068
rect 2010 -1080 2016 -1074
rect 2010 -1086 2016 -1080
rect 2010 -1092 2016 -1086
rect 2010 -1098 2016 -1092
rect 2010 -1104 2016 -1098
rect 2010 -1110 2016 -1104
rect 2010 -1116 2016 -1110
rect 2010 -1122 2016 -1116
rect 2010 -1128 2016 -1122
rect 2010 -1134 2016 -1128
rect 2010 -1140 2016 -1134
rect 2010 -1146 2016 -1140
rect 2010 -1152 2016 -1146
rect 2010 -1158 2016 -1152
rect 2010 -1164 2016 -1158
rect 2010 -1170 2016 -1164
rect 2010 -1176 2016 -1170
rect 2010 -1182 2016 -1176
rect 2010 -1188 2016 -1182
rect 2010 -1194 2016 -1188
rect 2010 -1200 2016 -1194
rect 2010 -1206 2016 -1200
rect 2010 -1212 2016 -1206
rect 2010 -1218 2016 -1212
rect 2010 -1224 2016 -1218
rect 2010 -1230 2016 -1224
rect 2010 -1236 2016 -1230
rect 2010 -1242 2016 -1236
rect 2010 -1248 2016 -1242
rect 2010 -1254 2016 -1248
rect 2010 -1260 2016 -1254
rect 2010 -1266 2016 -1260
rect 2010 -1272 2016 -1266
rect 2010 -1278 2016 -1272
rect 2010 -1284 2016 -1278
rect 2010 -1290 2016 -1284
rect 2010 -1296 2016 -1290
rect 2010 -1302 2016 -1296
rect 2010 -1308 2016 -1302
rect 2010 -1314 2016 -1308
rect 2010 -1320 2016 -1314
rect 2010 -1326 2016 -1320
rect 2010 -1332 2016 -1326
rect 2010 -1338 2016 -1332
rect 2010 -1344 2016 -1338
rect 2010 -1350 2016 -1344
rect 2010 -1356 2016 -1350
rect 2010 -1362 2016 -1356
rect 2010 -1368 2016 -1362
rect 2010 -1374 2016 -1368
rect 2010 -1380 2016 -1374
rect 2010 -1386 2016 -1380
rect 2010 -1392 2016 -1386
rect 2010 -1398 2016 -1392
rect 2010 -1404 2016 -1398
rect 2010 -1410 2016 -1404
rect 2010 -1416 2016 -1410
rect 2010 -1422 2016 -1416
rect 2010 -1428 2016 -1422
rect 2010 -1434 2016 -1428
rect 2010 -1440 2016 -1434
rect 2010 -1446 2016 -1440
rect 2010 -1452 2016 -1446
rect 2010 -1458 2016 -1452
rect 2010 -1464 2016 -1458
rect 2010 -1470 2016 -1464
rect 2010 -1476 2016 -1470
rect 2010 -1482 2016 -1476
rect 2010 -1488 2016 -1482
rect 2010 -1494 2016 -1488
rect 2010 -1500 2016 -1494
rect 2010 -1506 2016 -1500
rect 2010 -1512 2016 -1506
rect 2010 -1518 2016 -1512
rect 2010 -1524 2016 -1518
rect 2010 -1530 2016 -1524
rect 2010 -1536 2016 -1530
rect 2010 -1542 2016 -1536
rect 2010 -1548 2016 -1542
rect 2010 -1554 2016 -1548
rect 2010 -1560 2016 -1554
rect 2010 -1566 2016 -1560
rect 2010 -1572 2016 -1566
rect 2010 -1578 2016 -1572
rect 2010 -1584 2016 -1578
rect 2010 -1590 2016 -1584
rect 2010 -1596 2016 -1590
rect 2010 -1602 2016 -1596
rect 2010 -1608 2016 -1602
rect 2010 -1614 2016 -1608
rect 2010 -1620 2016 -1614
rect 2010 -1626 2016 -1620
rect 2010 -1632 2016 -1626
rect 2010 -1722 2016 -1716
rect 2010 -1728 2016 -1722
rect 2010 -1734 2016 -1728
rect 2010 -1740 2016 -1734
rect 2010 -1746 2016 -1740
rect 2010 -1752 2016 -1746
rect 2010 -1758 2016 -1752
rect 2010 -1764 2016 -1758
rect 2010 -1770 2016 -1764
rect 2010 -1776 2016 -1770
rect 2010 -1782 2016 -1776
rect 2010 -1788 2016 -1782
rect 2010 -1794 2016 -1788
rect 2010 -1800 2016 -1794
rect 2010 -1806 2016 -1800
rect 2010 -1812 2016 -1806
rect 2010 -1818 2016 -1812
rect 2010 -1824 2016 -1818
rect 2010 -1830 2016 -1824
rect 2010 -1836 2016 -1830
rect 2010 -1842 2016 -1836
rect 2010 -1848 2016 -1842
rect 2010 -1854 2016 -1848
rect 2010 -1860 2016 -1854
rect 2010 -1866 2016 -1860
rect 2010 -1872 2016 -1866
rect 2010 -1878 2016 -1872
rect 2010 -1884 2016 -1878
rect 2010 -1890 2016 -1884
rect 2010 -1896 2016 -1890
rect 2010 -1902 2016 -1896
rect 2010 -1908 2016 -1902
rect 2010 -1914 2016 -1908
rect 2010 -1920 2016 -1914
rect 2010 -1926 2016 -1920
rect 2010 -1932 2016 -1926
rect 2010 -1938 2016 -1932
rect 2010 -1944 2016 -1938
rect 2010 -1950 2016 -1944
rect 2010 -1956 2016 -1950
rect 2010 -1962 2016 -1956
rect 2010 -1968 2016 -1962
rect 2010 -1974 2016 -1968
rect 2010 -1980 2016 -1974
rect 2010 -1986 2016 -1980
rect 2010 -1992 2016 -1986
rect 2010 -1998 2016 -1992
rect 2010 -2004 2016 -1998
rect 2010 -2010 2016 -2004
rect 2010 -2016 2016 -2010
rect 2010 -2022 2016 -2016
rect 2010 -2028 2016 -2022
rect 2010 -2034 2016 -2028
rect 2010 -2040 2016 -2034
rect 2010 -2046 2016 -2040
rect 2010 -2052 2016 -2046
rect 2010 -2058 2016 -2052
rect 2010 -2064 2016 -2058
rect 2010 -2070 2016 -2064
rect 2010 -2076 2016 -2070
rect 2010 -2082 2016 -2076
rect 2010 -2088 2016 -2082
rect 2010 -2094 2016 -2088
rect 2010 -2100 2016 -2094
rect 2010 -2106 2016 -2100
rect 2010 -2112 2016 -2106
rect 2010 -2118 2016 -2112
rect 2010 -2124 2016 -2118
rect 2010 -2130 2016 -2124
rect 2010 -2136 2016 -2130
rect 2010 -2142 2016 -2136
rect 2010 -2148 2016 -2142
rect 2010 -2154 2016 -2148
rect 2010 -2160 2016 -2154
rect 2010 -2166 2016 -2160
rect 2010 -2172 2016 -2166
rect 2010 -2178 2016 -2172
rect 2010 -2184 2016 -2178
rect 2010 -2190 2016 -2184
rect 2010 -2196 2016 -2190
rect 2010 -2202 2016 -2196
rect 2010 -2208 2016 -2202
rect 2010 -2214 2016 -2208
rect 2010 -2220 2016 -2214
rect 2010 -2226 2016 -2220
rect 2010 -2232 2016 -2226
rect 2010 -2238 2016 -2232
rect 2010 -2244 2016 -2238
rect 2010 -2250 2016 -2244
rect 2010 -2256 2016 -2250
rect 2010 -2262 2016 -2256
rect 2010 -2268 2016 -2262
rect 2010 -2274 2016 -2268
rect 2010 -2280 2016 -2274
rect 2010 -2286 2016 -2280
rect 2010 -2292 2016 -2286
rect 2010 -2298 2016 -2292
rect 2010 -2304 2016 -2298
rect 2010 -2310 2016 -2304
rect 2010 -2316 2016 -2310
rect 2010 -2322 2016 -2316
rect 2010 -2328 2016 -2322
rect 2010 -2334 2016 -2328
rect 2010 -2340 2016 -2334
rect 2010 -2346 2016 -2340
rect 2010 -2352 2016 -2346
rect 2010 -2358 2016 -2352
rect 2010 -2364 2016 -2358
rect 2010 -2370 2016 -2364
rect 2010 -2376 2016 -2370
rect 2010 -2382 2016 -2376
rect 2010 -2388 2016 -2382
rect 2010 -2394 2016 -2388
rect 2010 -2400 2016 -2394
rect 2010 -2406 2016 -2400
rect 2010 -2412 2016 -2406
rect 2010 -2418 2016 -2412
rect 2010 -2424 2016 -2418
rect 2010 -2430 2016 -2424
rect 2010 -2436 2016 -2430
rect 2010 -2442 2016 -2436
rect 2010 -2448 2016 -2442
rect 2010 -2454 2016 -2448
rect 2010 -2460 2016 -2454
rect 2010 -2466 2016 -2460
rect 2010 -2472 2016 -2466
rect 2010 -2478 2016 -2472
rect 2010 -2484 2016 -2478
rect 2010 -2490 2016 -2484
rect 2010 -2496 2016 -2490
rect 2010 -2502 2016 -2496
rect 2010 -2508 2016 -2502
rect 2010 -2514 2016 -2508
rect 2010 -2520 2016 -2514
rect 2010 -2610 2016 -2604
rect 2010 -2616 2016 -2610
rect 2010 -2622 2016 -2616
rect 2010 -2628 2016 -2622
rect 2010 -2634 2016 -2628
rect 2010 -2640 2016 -2634
rect 2010 -2646 2016 -2640
rect 2010 -2652 2016 -2646
rect 2010 -2658 2016 -2652
rect 2010 -2664 2016 -2658
rect 2010 -2670 2016 -2664
rect 2010 -2676 2016 -2670
rect 2010 -2682 2016 -2676
rect 2010 -2688 2016 -2682
rect 2010 -2694 2016 -2688
rect 2010 -2700 2016 -2694
rect 2010 -2706 2016 -2700
rect 2010 -2712 2016 -2706
rect 2010 -2718 2016 -2712
rect 2010 -2724 2016 -2718
rect 2010 -2730 2016 -2724
rect 2010 -2736 2016 -2730
rect 2010 -2742 2016 -2736
rect 2010 -2748 2016 -2742
rect 2010 -2754 2016 -2748
rect 2010 -2760 2016 -2754
rect 2010 -2766 2016 -2760
rect 2010 -2772 2016 -2766
rect 2010 -2778 2016 -2772
rect 2010 -2784 2016 -2778
rect 2010 -2790 2016 -2784
rect 2010 -2796 2016 -2790
rect 2010 -2802 2016 -2796
rect 2010 -2808 2016 -2802
rect 2010 -2814 2016 -2808
rect 2010 -2820 2016 -2814
rect 2010 -2826 2016 -2820
rect 2010 -2832 2016 -2826
rect 2010 -2838 2016 -2832
rect 2010 -2844 2016 -2838
rect 2010 -2850 2016 -2844
rect 2010 -2856 2016 -2850
rect 2010 -2862 2016 -2856
rect 2010 -2868 2016 -2862
rect 2010 -2874 2016 -2868
rect 2010 -2880 2016 -2874
rect 2010 -2886 2016 -2880
rect 2010 -2892 2016 -2886
rect 2010 -2898 2016 -2892
rect 2010 -2904 2016 -2898
rect 2010 -2910 2016 -2904
rect 2010 -2916 2016 -2910
rect 2010 -2922 2016 -2916
rect 2010 -2928 2016 -2922
rect 2010 -2934 2016 -2928
rect 2010 -2940 2016 -2934
rect 2010 -2946 2016 -2940
rect 2010 -2952 2016 -2946
rect 2010 -2958 2016 -2952
rect 2010 -2964 2016 -2958
rect 2010 -2970 2016 -2964
rect 2010 -2976 2016 -2970
rect 2010 -2982 2016 -2976
rect 2010 -2988 2016 -2982
rect 2010 -2994 2016 -2988
rect 2010 -3000 2016 -2994
rect 2010 -3006 2016 -3000
rect 2010 -3012 2016 -3006
rect 2010 -3018 2016 -3012
rect 2010 -3024 2016 -3018
rect 2010 -3030 2016 -3024
rect 2010 -3036 2016 -3030
rect 2010 -3042 2016 -3036
rect 2010 -3048 2016 -3042
rect 2010 -3054 2016 -3048
rect 2010 -3060 2016 -3054
rect 2010 -3066 2016 -3060
rect 2010 -3072 2016 -3066
rect 2010 -3078 2016 -3072
rect 2010 -3084 2016 -3078
rect 2010 -3090 2016 -3084
rect 2010 -3096 2016 -3090
rect 2010 -3102 2016 -3096
rect 2010 -3156 2016 -3150
rect 2010 -3162 2016 -3156
rect 2010 -3168 2016 -3162
rect 2010 -3174 2016 -3168
rect 2010 -3180 2016 -3174
rect 2010 -3186 2016 -3180
rect 2010 -3192 2016 -3186
rect 2010 -3198 2016 -3192
rect 2010 -3204 2016 -3198
rect 2010 -3210 2016 -3204
rect 2016 -432 2022 -426
rect 2016 -438 2022 -432
rect 2016 -444 2022 -438
rect 2016 -450 2022 -444
rect 2016 -456 2022 -450
rect 2016 -462 2022 -456
rect 2016 -468 2022 -462
rect 2016 -474 2022 -468
rect 2016 -480 2022 -474
rect 2016 -486 2022 -480
rect 2016 -492 2022 -486
rect 2016 -498 2022 -492
rect 2016 -504 2022 -498
rect 2016 -510 2022 -504
rect 2016 -516 2022 -510
rect 2016 -522 2022 -516
rect 2016 -528 2022 -522
rect 2016 -534 2022 -528
rect 2016 -540 2022 -534
rect 2016 -546 2022 -540
rect 2016 -552 2022 -546
rect 2016 -558 2022 -552
rect 2016 -564 2022 -558
rect 2016 -570 2022 -564
rect 2016 -576 2022 -570
rect 2016 -582 2022 -576
rect 2016 -588 2022 -582
rect 2016 -594 2022 -588
rect 2016 -600 2022 -594
rect 2016 -606 2022 -600
rect 2016 -612 2022 -606
rect 2016 -618 2022 -612
rect 2016 -624 2022 -618
rect 2016 -630 2022 -624
rect 2016 -636 2022 -630
rect 2016 -642 2022 -636
rect 2016 -648 2022 -642
rect 2016 -654 2022 -648
rect 2016 -660 2022 -654
rect 2016 -666 2022 -660
rect 2016 -672 2022 -666
rect 2016 -678 2022 -672
rect 2016 -684 2022 -678
rect 2016 -690 2022 -684
rect 2016 -696 2022 -690
rect 2016 -702 2022 -696
rect 2016 -708 2022 -702
rect 2016 -714 2022 -708
rect 2016 -720 2022 -714
rect 2016 -726 2022 -720
rect 2016 -732 2022 -726
rect 2016 -738 2022 -732
rect 2016 -744 2022 -738
rect 2016 -750 2022 -744
rect 2016 -756 2022 -750
rect 2016 -762 2022 -756
rect 2016 -768 2022 -762
rect 2016 -774 2022 -768
rect 2016 -780 2022 -774
rect 2016 -786 2022 -780
rect 2016 -792 2022 -786
rect 2016 -798 2022 -792
rect 2016 -804 2022 -798
rect 2016 -810 2022 -804
rect 2016 -816 2022 -810
rect 2016 -822 2022 -816
rect 2016 -828 2022 -822
rect 2016 -834 2022 -828
rect 2016 -840 2022 -834
rect 2016 -846 2022 -840
rect 2016 -852 2022 -846
rect 2016 -858 2022 -852
rect 2016 -864 2022 -858
rect 2016 -870 2022 -864
rect 2016 -876 2022 -870
rect 2016 -882 2022 -876
rect 2016 -888 2022 -882
rect 2016 -894 2022 -888
rect 2016 -900 2022 -894
rect 2016 -906 2022 -900
rect 2016 -912 2022 -906
rect 2016 -918 2022 -912
rect 2016 -924 2022 -918
rect 2016 -930 2022 -924
rect 2016 -936 2022 -930
rect 2016 -942 2022 -936
rect 2016 -948 2022 -942
rect 2016 -954 2022 -948
rect 2016 -960 2022 -954
rect 2016 -966 2022 -960
rect 2016 -972 2022 -966
rect 2016 -978 2022 -972
rect 2016 -984 2022 -978
rect 2016 -990 2022 -984
rect 2016 -996 2022 -990
rect 2016 -1002 2022 -996
rect 2016 -1008 2022 -1002
rect 2016 -1014 2022 -1008
rect 2016 -1020 2022 -1014
rect 2016 -1026 2022 -1020
rect 2016 -1032 2022 -1026
rect 2016 -1038 2022 -1032
rect 2016 -1044 2022 -1038
rect 2016 -1050 2022 -1044
rect 2016 -1056 2022 -1050
rect 2016 -1062 2022 -1056
rect 2016 -1068 2022 -1062
rect 2016 -1074 2022 -1068
rect 2016 -1080 2022 -1074
rect 2016 -1086 2022 -1080
rect 2016 -1092 2022 -1086
rect 2016 -1098 2022 -1092
rect 2016 -1104 2022 -1098
rect 2016 -1110 2022 -1104
rect 2016 -1116 2022 -1110
rect 2016 -1122 2022 -1116
rect 2016 -1128 2022 -1122
rect 2016 -1134 2022 -1128
rect 2016 -1140 2022 -1134
rect 2016 -1146 2022 -1140
rect 2016 -1152 2022 -1146
rect 2016 -1158 2022 -1152
rect 2016 -1164 2022 -1158
rect 2016 -1170 2022 -1164
rect 2016 -1176 2022 -1170
rect 2016 -1182 2022 -1176
rect 2016 -1188 2022 -1182
rect 2016 -1194 2022 -1188
rect 2016 -1200 2022 -1194
rect 2016 -1206 2022 -1200
rect 2016 -1212 2022 -1206
rect 2016 -1218 2022 -1212
rect 2016 -1224 2022 -1218
rect 2016 -1230 2022 -1224
rect 2016 -1236 2022 -1230
rect 2016 -1242 2022 -1236
rect 2016 -1248 2022 -1242
rect 2016 -1254 2022 -1248
rect 2016 -1260 2022 -1254
rect 2016 -1266 2022 -1260
rect 2016 -1272 2022 -1266
rect 2016 -1278 2022 -1272
rect 2016 -1284 2022 -1278
rect 2016 -1290 2022 -1284
rect 2016 -1296 2022 -1290
rect 2016 -1302 2022 -1296
rect 2016 -1308 2022 -1302
rect 2016 -1314 2022 -1308
rect 2016 -1320 2022 -1314
rect 2016 -1326 2022 -1320
rect 2016 -1332 2022 -1326
rect 2016 -1338 2022 -1332
rect 2016 -1344 2022 -1338
rect 2016 -1350 2022 -1344
rect 2016 -1356 2022 -1350
rect 2016 -1362 2022 -1356
rect 2016 -1368 2022 -1362
rect 2016 -1374 2022 -1368
rect 2016 -1380 2022 -1374
rect 2016 -1386 2022 -1380
rect 2016 -1392 2022 -1386
rect 2016 -1398 2022 -1392
rect 2016 -1404 2022 -1398
rect 2016 -1410 2022 -1404
rect 2016 -1416 2022 -1410
rect 2016 -1422 2022 -1416
rect 2016 -1428 2022 -1422
rect 2016 -1434 2022 -1428
rect 2016 -1440 2022 -1434
rect 2016 -1446 2022 -1440
rect 2016 -1452 2022 -1446
rect 2016 -1458 2022 -1452
rect 2016 -1464 2022 -1458
rect 2016 -1470 2022 -1464
rect 2016 -1476 2022 -1470
rect 2016 -1482 2022 -1476
rect 2016 -1488 2022 -1482
rect 2016 -1494 2022 -1488
rect 2016 -1500 2022 -1494
rect 2016 -1506 2022 -1500
rect 2016 -1512 2022 -1506
rect 2016 -1518 2022 -1512
rect 2016 -1524 2022 -1518
rect 2016 -1530 2022 -1524
rect 2016 -1536 2022 -1530
rect 2016 -1542 2022 -1536
rect 2016 -1548 2022 -1542
rect 2016 -1554 2022 -1548
rect 2016 -1560 2022 -1554
rect 2016 -1566 2022 -1560
rect 2016 -1572 2022 -1566
rect 2016 -1578 2022 -1572
rect 2016 -1584 2022 -1578
rect 2016 -1590 2022 -1584
rect 2016 -1596 2022 -1590
rect 2016 -1602 2022 -1596
rect 2016 -1608 2022 -1602
rect 2016 -1614 2022 -1608
rect 2016 -1620 2022 -1614
rect 2016 -1626 2022 -1620
rect 2016 -1716 2022 -1710
rect 2016 -1722 2022 -1716
rect 2016 -1728 2022 -1722
rect 2016 -1734 2022 -1728
rect 2016 -1740 2022 -1734
rect 2016 -1746 2022 -1740
rect 2016 -1752 2022 -1746
rect 2016 -1758 2022 -1752
rect 2016 -1764 2022 -1758
rect 2016 -1770 2022 -1764
rect 2016 -1776 2022 -1770
rect 2016 -1782 2022 -1776
rect 2016 -1788 2022 -1782
rect 2016 -1794 2022 -1788
rect 2016 -1800 2022 -1794
rect 2016 -1806 2022 -1800
rect 2016 -1812 2022 -1806
rect 2016 -1818 2022 -1812
rect 2016 -1824 2022 -1818
rect 2016 -1830 2022 -1824
rect 2016 -1836 2022 -1830
rect 2016 -1842 2022 -1836
rect 2016 -1848 2022 -1842
rect 2016 -1854 2022 -1848
rect 2016 -1860 2022 -1854
rect 2016 -1866 2022 -1860
rect 2016 -1872 2022 -1866
rect 2016 -1878 2022 -1872
rect 2016 -1884 2022 -1878
rect 2016 -1890 2022 -1884
rect 2016 -1896 2022 -1890
rect 2016 -1902 2022 -1896
rect 2016 -1908 2022 -1902
rect 2016 -1914 2022 -1908
rect 2016 -1920 2022 -1914
rect 2016 -1926 2022 -1920
rect 2016 -1932 2022 -1926
rect 2016 -1938 2022 -1932
rect 2016 -1944 2022 -1938
rect 2016 -1950 2022 -1944
rect 2016 -1956 2022 -1950
rect 2016 -1962 2022 -1956
rect 2016 -1968 2022 -1962
rect 2016 -1974 2022 -1968
rect 2016 -1980 2022 -1974
rect 2016 -1986 2022 -1980
rect 2016 -1992 2022 -1986
rect 2016 -1998 2022 -1992
rect 2016 -2004 2022 -1998
rect 2016 -2010 2022 -2004
rect 2016 -2016 2022 -2010
rect 2016 -2022 2022 -2016
rect 2016 -2028 2022 -2022
rect 2016 -2034 2022 -2028
rect 2016 -2040 2022 -2034
rect 2016 -2046 2022 -2040
rect 2016 -2052 2022 -2046
rect 2016 -2058 2022 -2052
rect 2016 -2064 2022 -2058
rect 2016 -2070 2022 -2064
rect 2016 -2076 2022 -2070
rect 2016 -2082 2022 -2076
rect 2016 -2088 2022 -2082
rect 2016 -2094 2022 -2088
rect 2016 -2100 2022 -2094
rect 2016 -2106 2022 -2100
rect 2016 -2112 2022 -2106
rect 2016 -2118 2022 -2112
rect 2016 -2124 2022 -2118
rect 2016 -2130 2022 -2124
rect 2016 -2136 2022 -2130
rect 2016 -2142 2022 -2136
rect 2016 -2148 2022 -2142
rect 2016 -2154 2022 -2148
rect 2016 -2160 2022 -2154
rect 2016 -2166 2022 -2160
rect 2016 -2172 2022 -2166
rect 2016 -2178 2022 -2172
rect 2016 -2184 2022 -2178
rect 2016 -2190 2022 -2184
rect 2016 -2196 2022 -2190
rect 2016 -2202 2022 -2196
rect 2016 -2208 2022 -2202
rect 2016 -2214 2022 -2208
rect 2016 -2220 2022 -2214
rect 2016 -2226 2022 -2220
rect 2016 -2232 2022 -2226
rect 2016 -2238 2022 -2232
rect 2016 -2244 2022 -2238
rect 2016 -2250 2022 -2244
rect 2016 -2256 2022 -2250
rect 2016 -2262 2022 -2256
rect 2016 -2268 2022 -2262
rect 2016 -2274 2022 -2268
rect 2016 -2280 2022 -2274
rect 2016 -2286 2022 -2280
rect 2016 -2292 2022 -2286
rect 2016 -2298 2022 -2292
rect 2016 -2304 2022 -2298
rect 2016 -2310 2022 -2304
rect 2016 -2316 2022 -2310
rect 2016 -2322 2022 -2316
rect 2016 -2328 2022 -2322
rect 2016 -2334 2022 -2328
rect 2016 -2340 2022 -2334
rect 2016 -2346 2022 -2340
rect 2016 -2352 2022 -2346
rect 2016 -2358 2022 -2352
rect 2016 -2364 2022 -2358
rect 2016 -2370 2022 -2364
rect 2016 -2376 2022 -2370
rect 2016 -2382 2022 -2376
rect 2016 -2388 2022 -2382
rect 2016 -2394 2022 -2388
rect 2016 -2400 2022 -2394
rect 2016 -2406 2022 -2400
rect 2016 -2412 2022 -2406
rect 2016 -2418 2022 -2412
rect 2016 -2424 2022 -2418
rect 2016 -2430 2022 -2424
rect 2016 -2436 2022 -2430
rect 2016 -2442 2022 -2436
rect 2016 -2448 2022 -2442
rect 2016 -2454 2022 -2448
rect 2016 -2460 2022 -2454
rect 2016 -2466 2022 -2460
rect 2016 -2472 2022 -2466
rect 2016 -2478 2022 -2472
rect 2016 -2484 2022 -2478
rect 2016 -2490 2022 -2484
rect 2016 -2496 2022 -2490
rect 2016 -2502 2022 -2496
rect 2016 -2508 2022 -2502
rect 2016 -2514 2022 -2508
rect 2016 -2520 2022 -2514
rect 2016 -2604 2022 -2598
rect 2016 -2610 2022 -2604
rect 2016 -2616 2022 -2610
rect 2016 -2622 2022 -2616
rect 2016 -2628 2022 -2622
rect 2016 -2634 2022 -2628
rect 2016 -2640 2022 -2634
rect 2016 -2646 2022 -2640
rect 2016 -2652 2022 -2646
rect 2016 -2658 2022 -2652
rect 2016 -2664 2022 -2658
rect 2016 -2670 2022 -2664
rect 2016 -2676 2022 -2670
rect 2016 -2682 2022 -2676
rect 2016 -2688 2022 -2682
rect 2016 -2694 2022 -2688
rect 2016 -2700 2022 -2694
rect 2016 -2706 2022 -2700
rect 2016 -2712 2022 -2706
rect 2016 -2718 2022 -2712
rect 2016 -2724 2022 -2718
rect 2016 -2730 2022 -2724
rect 2016 -2736 2022 -2730
rect 2016 -2742 2022 -2736
rect 2016 -2748 2022 -2742
rect 2016 -2754 2022 -2748
rect 2016 -2760 2022 -2754
rect 2016 -2766 2022 -2760
rect 2016 -2772 2022 -2766
rect 2016 -2778 2022 -2772
rect 2016 -2784 2022 -2778
rect 2016 -2790 2022 -2784
rect 2016 -2796 2022 -2790
rect 2016 -2802 2022 -2796
rect 2016 -2808 2022 -2802
rect 2016 -2814 2022 -2808
rect 2016 -2820 2022 -2814
rect 2016 -2826 2022 -2820
rect 2016 -2832 2022 -2826
rect 2016 -2838 2022 -2832
rect 2016 -2844 2022 -2838
rect 2016 -2850 2022 -2844
rect 2016 -2856 2022 -2850
rect 2016 -2862 2022 -2856
rect 2016 -2868 2022 -2862
rect 2016 -2874 2022 -2868
rect 2016 -2880 2022 -2874
rect 2016 -2886 2022 -2880
rect 2016 -2892 2022 -2886
rect 2016 -2898 2022 -2892
rect 2016 -2904 2022 -2898
rect 2016 -2910 2022 -2904
rect 2016 -2916 2022 -2910
rect 2016 -2922 2022 -2916
rect 2016 -2928 2022 -2922
rect 2016 -2934 2022 -2928
rect 2016 -2940 2022 -2934
rect 2016 -2946 2022 -2940
rect 2016 -2952 2022 -2946
rect 2016 -2958 2022 -2952
rect 2016 -2964 2022 -2958
rect 2016 -2970 2022 -2964
rect 2016 -2976 2022 -2970
rect 2016 -2982 2022 -2976
rect 2016 -2988 2022 -2982
rect 2016 -2994 2022 -2988
rect 2016 -3000 2022 -2994
rect 2016 -3006 2022 -3000
rect 2016 -3012 2022 -3006
rect 2016 -3018 2022 -3012
rect 2016 -3024 2022 -3018
rect 2016 -3030 2022 -3024
rect 2016 -3036 2022 -3030
rect 2016 -3042 2022 -3036
rect 2016 -3048 2022 -3042
rect 2016 -3054 2022 -3048
rect 2016 -3060 2022 -3054
rect 2016 -3066 2022 -3060
rect 2016 -3072 2022 -3066
rect 2016 -3078 2022 -3072
rect 2016 -3084 2022 -3078
rect 2016 -3090 2022 -3084
rect 2016 -3096 2022 -3090
rect 2016 -3156 2022 -3150
rect 2016 -3162 2022 -3156
rect 2016 -3168 2022 -3162
rect 2016 -3174 2022 -3168
rect 2016 -3180 2022 -3174
rect 2016 -3186 2022 -3180
rect 2016 -3192 2022 -3186
rect 2016 -3198 2022 -3192
rect 2016 -3204 2022 -3198
rect 2022 -420 2028 -414
rect 2022 -426 2028 -420
rect 2022 -432 2028 -426
rect 2022 -438 2028 -432
rect 2022 -444 2028 -438
rect 2022 -450 2028 -444
rect 2022 -456 2028 -450
rect 2022 -462 2028 -456
rect 2022 -468 2028 -462
rect 2022 -474 2028 -468
rect 2022 -480 2028 -474
rect 2022 -486 2028 -480
rect 2022 -492 2028 -486
rect 2022 -498 2028 -492
rect 2022 -504 2028 -498
rect 2022 -510 2028 -504
rect 2022 -516 2028 -510
rect 2022 -522 2028 -516
rect 2022 -528 2028 -522
rect 2022 -534 2028 -528
rect 2022 -540 2028 -534
rect 2022 -546 2028 -540
rect 2022 -552 2028 -546
rect 2022 -558 2028 -552
rect 2022 -564 2028 -558
rect 2022 -570 2028 -564
rect 2022 -576 2028 -570
rect 2022 -582 2028 -576
rect 2022 -588 2028 -582
rect 2022 -594 2028 -588
rect 2022 -600 2028 -594
rect 2022 -606 2028 -600
rect 2022 -612 2028 -606
rect 2022 -618 2028 -612
rect 2022 -624 2028 -618
rect 2022 -630 2028 -624
rect 2022 -636 2028 -630
rect 2022 -642 2028 -636
rect 2022 -648 2028 -642
rect 2022 -654 2028 -648
rect 2022 -660 2028 -654
rect 2022 -666 2028 -660
rect 2022 -672 2028 -666
rect 2022 -678 2028 -672
rect 2022 -684 2028 -678
rect 2022 -690 2028 -684
rect 2022 -696 2028 -690
rect 2022 -702 2028 -696
rect 2022 -708 2028 -702
rect 2022 -714 2028 -708
rect 2022 -720 2028 -714
rect 2022 -726 2028 -720
rect 2022 -732 2028 -726
rect 2022 -738 2028 -732
rect 2022 -744 2028 -738
rect 2022 -750 2028 -744
rect 2022 -756 2028 -750
rect 2022 -762 2028 -756
rect 2022 -768 2028 -762
rect 2022 -774 2028 -768
rect 2022 -780 2028 -774
rect 2022 -786 2028 -780
rect 2022 -792 2028 -786
rect 2022 -798 2028 -792
rect 2022 -804 2028 -798
rect 2022 -810 2028 -804
rect 2022 -816 2028 -810
rect 2022 -822 2028 -816
rect 2022 -828 2028 -822
rect 2022 -834 2028 -828
rect 2022 -840 2028 -834
rect 2022 -846 2028 -840
rect 2022 -852 2028 -846
rect 2022 -858 2028 -852
rect 2022 -864 2028 -858
rect 2022 -870 2028 -864
rect 2022 -876 2028 -870
rect 2022 -882 2028 -876
rect 2022 -888 2028 -882
rect 2022 -894 2028 -888
rect 2022 -900 2028 -894
rect 2022 -906 2028 -900
rect 2022 -912 2028 -906
rect 2022 -918 2028 -912
rect 2022 -924 2028 -918
rect 2022 -930 2028 -924
rect 2022 -936 2028 -930
rect 2022 -942 2028 -936
rect 2022 -948 2028 -942
rect 2022 -954 2028 -948
rect 2022 -960 2028 -954
rect 2022 -966 2028 -960
rect 2022 -972 2028 -966
rect 2022 -978 2028 -972
rect 2022 -984 2028 -978
rect 2022 -990 2028 -984
rect 2022 -996 2028 -990
rect 2022 -1002 2028 -996
rect 2022 -1008 2028 -1002
rect 2022 -1014 2028 -1008
rect 2022 -1020 2028 -1014
rect 2022 -1026 2028 -1020
rect 2022 -1032 2028 -1026
rect 2022 -1038 2028 -1032
rect 2022 -1044 2028 -1038
rect 2022 -1050 2028 -1044
rect 2022 -1056 2028 -1050
rect 2022 -1062 2028 -1056
rect 2022 -1068 2028 -1062
rect 2022 -1074 2028 -1068
rect 2022 -1080 2028 -1074
rect 2022 -1086 2028 -1080
rect 2022 -1092 2028 -1086
rect 2022 -1098 2028 -1092
rect 2022 -1104 2028 -1098
rect 2022 -1110 2028 -1104
rect 2022 -1116 2028 -1110
rect 2022 -1122 2028 -1116
rect 2022 -1128 2028 -1122
rect 2022 -1134 2028 -1128
rect 2022 -1140 2028 -1134
rect 2022 -1146 2028 -1140
rect 2022 -1152 2028 -1146
rect 2022 -1158 2028 -1152
rect 2022 -1164 2028 -1158
rect 2022 -1170 2028 -1164
rect 2022 -1176 2028 -1170
rect 2022 -1182 2028 -1176
rect 2022 -1188 2028 -1182
rect 2022 -1194 2028 -1188
rect 2022 -1200 2028 -1194
rect 2022 -1206 2028 -1200
rect 2022 -1212 2028 -1206
rect 2022 -1218 2028 -1212
rect 2022 -1224 2028 -1218
rect 2022 -1230 2028 -1224
rect 2022 -1236 2028 -1230
rect 2022 -1242 2028 -1236
rect 2022 -1248 2028 -1242
rect 2022 -1254 2028 -1248
rect 2022 -1260 2028 -1254
rect 2022 -1266 2028 -1260
rect 2022 -1272 2028 -1266
rect 2022 -1278 2028 -1272
rect 2022 -1284 2028 -1278
rect 2022 -1290 2028 -1284
rect 2022 -1296 2028 -1290
rect 2022 -1302 2028 -1296
rect 2022 -1308 2028 -1302
rect 2022 -1314 2028 -1308
rect 2022 -1320 2028 -1314
rect 2022 -1326 2028 -1320
rect 2022 -1332 2028 -1326
rect 2022 -1338 2028 -1332
rect 2022 -1344 2028 -1338
rect 2022 -1350 2028 -1344
rect 2022 -1356 2028 -1350
rect 2022 -1362 2028 -1356
rect 2022 -1368 2028 -1362
rect 2022 -1374 2028 -1368
rect 2022 -1380 2028 -1374
rect 2022 -1386 2028 -1380
rect 2022 -1392 2028 -1386
rect 2022 -1398 2028 -1392
rect 2022 -1404 2028 -1398
rect 2022 -1410 2028 -1404
rect 2022 -1416 2028 -1410
rect 2022 -1422 2028 -1416
rect 2022 -1428 2028 -1422
rect 2022 -1434 2028 -1428
rect 2022 -1440 2028 -1434
rect 2022 -1446 2028 -1440
rect 2022 -1452 2028 -1446
rect 2022 -1458 2028 -1452
rect 2022 -1464 2028 -1458
rect 2022 -1470 2028 -1464
rect 2022 -1476 2028 -1470
rect 2022 -1482 2028 -1476
rect 2022 -1488 2028 -1482
rect 2022 -1494 2028 -1488
rect 2022 -1500 2028 -1494
rect 2022 -1506 2028 -1500
rect 2022 -1512 2028 -1506
rect 2022 -1518 2028 -1512
rect 2022 -1524 2028 -1518
rect 2022 -1530 2028 -1524
rect 2022 -1536 2028 -1530
rect 2022 -1542 2028 -1536
rect 2022 -1548 2028 -1542
rect 2022 -1554 2028 -1548
rect 2022 -1560 2028 -1554
rect 2022 -1566 2028 -1560
rect 2022 -1572 2028 -1566
rect 2022 -1578 2028 -1572
rect 2022 -1584 2028 -1578
rect 2022 -1590 2028 -1584
rect 2022 -1596 2028 -1590
rect 2022 -1602 2028 -1596
rect 2022 -1608 2028 -1602
rect 2022 -1614 2028 -1608
rect 2022 -1620 2028 -1614
rect 2022 -1710 2028 -1704
rect 2022 -1716 2028 -1710
rect 2022 -1722 2028 -1716
rect 2022 -1728 2028 -1722
rect 2022 -1734 2028 -1728
rect 2022 -1740 2028 -1734
rect 2022 -1746 2028 -1740
rect 2022 -1752 2028 -1746
rect 2022 -1758 2028 -1752
rect 2022 -1764 2028 -1758
rect 2022 -1770 2028 -1764
rect 2022 -1776 2028 -1770
rect 2022 -1782 2028 -1776
rect 2022 -1788 2028 -1782
rect 2022 -1794 2028 -1788
rect 2022 -1800 2028 -1794
rect 2022 -1806 2028 -1800
rect 2022 -1812 2028 -1806
rect 2022 -1818 2028 -1812
rect 2022 -1824 2028 -1818
rect 2022 -1830 2028 -1824
rect 2022 -1836 2028 -1830
rect 2022 -1842 2028 -1836
rect 2022 -1848 2028 -1842
rect 2022 -1854 2028 -1848
rect 2022 -1860 2028 -1854
rect 2022 -1866 2028 -1860
rect 2022 -1872 2028 -1866
rect 2022 -1878 2028 -1872
rect 2022 -1884 2028 -1878
rect 2022 -1890 2028 -1884
rect 2022 -1896 2028 -1890
rect 2022 -1902 2028 -1896
rect 2022 -1908 2028 -1902
rect 2022 -1914 2028 -1908
rect 2022 -1920 2028 -1914
rect 2022 -1926 2028 -1920
rect 2022 -1932 2028 -1926
rect 2022 -1938 2028 -1932
rect 2022 -1944 2028 -1938
rect 2022 -1950 2028 -1944
rect 2022 -1956 2028 -1950
rect 2022 -1962 2028 -1956
rect 2022 -1968 2028 -1962
rect 2022 -1974 2028 -1968
rect 2022 -1980 2028 -1974
rect 2022 -1986 2028 -1980
rect 2022 -1992 2028 -1986
rect 2022 -1998 2028 -1992
rect 2022 -2004 2028 -1998
rect 2022 -2010 2028 -2004
rect 2022 -2016 2028 -2010
rect 2022 -2022 2028 -2016
rect 2022 -2028 2028 -2022
rect 2022 -2034 2028 -2028
rect 2022 -2040 2028 -2034
rect 2022 -2046 2028 -2040
rect 2022 -2052 2028 -2046
rect 2022 -2058 2028 -2052
rect 2022 -2064 2028 -2058
rect 2022 -2070 2028 -2064
rect 2022 -2076 2028 -2070
rect 2022 -2082 2028 -2076
rect 2022 -2088 2028 -2082
rect 2022 -2094 2028 -2088
rect 2022 -2100 2028 -2094
rect 2022 -2106 2028 -2100
rect 2022 -2112 2028 -2106
rect 2022 -2118 2028 -2112
rect 2022 -2124 2028 -2118
rect 2022 -2130 2028 -2124
rect 2022 -2136 2028 -2130
rect 2022 -2142 2028 -2136
rect 2022 -2148 2028 -2142
rect 2022 -2154 2028 -2148
rect 2022 -2160 2028 -2154
rect 2022 -2166 2028 -2160
rect 2022 -2172 2028 -2166
rect 2022 -2178 2028 -2172
rect 2022 -2184 2028 -2178
rect 2022 -2190 2028 -2184
rect 2022 -2196 2028 -2190
rect 2022 -2202 2028 -2196
rect 2022 -2208 2028 -2202
rect 2022 -2214 2028 -2208
rect 2022 -2220 2028 -2214
rect 2022 -2226 2028 -2220
rect 2022 -2232 2028 -2226
rect 2022 -2238 2028 -2232
rect 2022 -2244 2028 -2238
rect 2022 -2250 2028 -2244
rect 2022 -2256 2028 -2250
rect 2022 -2262 2028 -2256
rect 2022 -2268 2028 -2262
rect 2022 -2274 2028 -2268
rect 2022 -2280 2028 -2274
rect 2022 -2286 2028 -2280
rect 2022 -2292 2028 -2286
rect 2022 -2298 2028 -2292
rect 2022 -2304 2028 -2298
rect 2022 -2310 2028 -2304
rect 2022 -2316 2028 -2310
rect 2022 -2322 2028 -2316
rect 2022 -2328 2028 -2322
rect 2022 -2334 2028 -2328
rect 2022 -2340 2028 -2334
rect 2022 -2346 2028 -2340
rect 2022 -2352 2028 -2346
rect 2022 -2358 2028 -2352
rect 2022 -2364 2028 -2358
rect 2022 -2370 2028 -2364
rect 2022 -2376 2028 -2370
rect 2022 -2382 2028 -2376
rect 2022 -2388 2028 -2382
rect 2022 -2394 2028 -2388
rect 2022 -2400 2028 -2394
rect 2022 -2406 2028 -2400
rect 2022 -2412 2028 -2406
rect 2022 -2418 2028 -2412
rect 2022 -2424 2028 -2418
rect 2022 -2430 2028 -2424
rect 2022 -2436 2028 -2430
rect 2022 -2442 2028 -2436
rect 2022 -2448 2028 -2442
rect 2022 -2454 2028 -2448
rect 2022 -2460 2028 -2454
rect 2022 -2466 2028 -2460
rect 2022 -2472 2028 -2466
rect 2022 -2478 2028 -2472
rect 2022 -2484 2028 -2478
rect 2022 -2490 2028 -2484
rect 2022 -2496 2028 -2490
rect 2022 -2502 2028 -2496
rect 2022 -2508 2028 -2502
rect 2022 -2514 2028 -2508
rect 2022 -2604 2028 -2598
rect 2022 -2610 2028 -2604
rect 2022 -2616 2028 -2610
rect 2022 -2622 2028 -2616
rect 2022 -2628 2028 -2622
rect 2022 -2634 2028 -2628
rect 2022 -2640 2028 -2634
rect 2022 -2646 2028 -2640
rect 2022 -2652 2028 -2646
rect 2022 -2658 2028 -2652
rect 2022 -2664 2028 -2658
rect 2022 -2670 2028 -2664
rect 2022 -2676 2028 -2670
rect 2022 -2682 2028 -2676
rect 2022 -2688 2028 -2682
rect 2022 -2694 2028 -2688
rect 2022 -2700 2028 -2694
rect 2022 -2706 2028 -2700
rect 2022 -2712 2028 -2706
rect 2022 -2718 2028 -2712
rect 2022 -2724 2028 -2718
rect 2022 -2730 2028 -2724
rect 2022 -2736 2028 -2730
rect 2022 -2742 2028 -2736
rect 2022 -2748 2028 -2742
rect 2022 -2754 2028 -2748
rect 2022 -2760 2028 -2754
rect 2022 -2766 2028 -2760
rect 2022 -2772 2028 -2766
rect 2022 -2778 2028 -2772
rect 2022 -2784 2028 -2778
rect 2022 -2790 2028 -2784
rect 2022 -2796 2028 -2790
rect 2022 -2802 2028 -2796
rect 2022 -2808 2028 -2802
rect 2022 -2814 2028 -2808
rect 2022 -2820 2028 -2814
rect 2022 -2826 2028 -2820
rect 2022 -2832 2028 -2826
rect 2022 -2838 2028 -2832
rect 2022 -2844 2028 -2838
rect 2022 -2850 2028 -2844
rect 2022 -2856 2028 -2850
rect 2022 -2862 2028 -2856
rect 2022 -2868 2028 -2862
rect 2022 -2874 2028 -2868
rect 2022 -2880 2028 -2874
rect 2022 -2886 2028 -2880
rect 2022 -2892 2028 -2886
rect 2022 -2898 2028 -2892
rect 2022 -2904 2028 -2898
rect 2022 -2910 2028 -2904
rect 2022 -2916 2028 -2910
rect 2022 -2922 2028 -2916
rect 2022 -2928 2028 -2922
rect 2022 -2934 2028 -2928
rect 2022 -2940 2028 -2934
rect 2022 -2946 2028 -2940
rect 2022 -2952 2028 -2946
rect 2022 -2958 2028 -2952
rect 2022 -2964 2028 -2958
rect 2022 -2970 2028 -2964
rect 2022 -2976 2028 -2970
rect 2022 -2982 2028 -2976
rect 2022 -2988 2028 -2982
rect 2022 -2994 2028 -2988
rect 2022 -3000 2028 -2994
rect 2022 -3006 2028 -3000
rect 2022 -3012 2028 -3006
rect 2022 -3018 2028 -3012
rect 2022 -3024 2028 -3018
rect 2022 -3030 2028 -3024
rect 2022 -3036 2028 -3030
rect 2022 -3042 2028 -3036
rect 2022 -3048 2028 -3042
rect 2022 -3054 2028 -3048
rect 2022 -3060 2028 -3054
rect 2022 -3066 2028 -3060
rect 2022 -3072 2028 -3066
rect 2022 -3078 2028 -3072
rect 2022 -3084 2028 -3078
rect 2022 -3090 2028 -3084
rect 2022 -3096 2028 -3090
rect 2022 -3150 2028 -3144
rect 2022 -3156 2028 -3150
rect 2022 -3162 2028 -3156
rect 2022 -3168 2028 -3162
rect 2022 -3174 2028 -3168
rect 2022 -3180 2028 -3174
rect 2022 -3186 2028 -3180
rect 2022 -3192 2028 -3186
rect 2022 -3198 2028 -3192
rect 2028 -414 2034 -408
rect 2028 -420 2034 -414
rect 2028 -426 2034 -420
rect 2028 -432 2034 -426
rect 2028 -438 2034 -432
rect 2028 -444 2034 -438
rect 2028 -450 2034 -444
rect 2028 -456 2034 -450
rect 2028 -462 2034 -456
rect 2028 -468 2034 -462
rect 2028 -474 2034 -468
rect 2028 -480 2034 -474
rect 2028 -486 2034 -480
rect 2028 -492 2034 -486
rect 2028 -498 2034 -492
rect 2028 -504 2034 -498
rect 2028 -510 2034 -504
rect 2028 -516 2034 -510
rect 2028 -522 2034 -516
rect 2028 -528 2034 -522
rect 2028 -534 2034 -528
rect 2028 -540 2034 -534
rect 2028 -546 2034 -540
rect 2028 -552 2034 -546
rect 2028 -558 2034 -552
rect 2028 -564 2034 -558
rect 2028 -570 2034 -564
rect 2028 -576 2034 -570
rect 2028 -582 2034 -576
rect 2028 -588 2034 -582
rect 2028 -594 2034 -588
rect 2028 -600 2034 -594
rect 2028 -606 2034 -600
rect 2028 -612 2034 -606
rect 2028 -618 2034 -612
rect 2028 -624 2034 -618
rect 2028 -630 2034 -624
rect 2028 -636 2034 -630
rect 2028 -642 2034 -636
rect 2028 -648 2034 -642
rect 2028 -654 2034 -648
rect 2028 -660 2034 -654
rect 2028 -666 2034 -660
rect 2028 -672 2034 -666
rect 2028 -678 2034 -672
rect 2028 -684 2034 -678
rect 2028 -690 2034 -684
rect 2028 -696 2034 -690
rect 2028 -702 2034 -696
rect 2028 -708 2034 -702
rect 2028 -714 2034 -708
rect 2028 -720 2034 -714
rect 2028 -726 2034 -720
rect 2028 -732 2034 -726
rect 2028 -738 2034 -732
rect 2028 -744 2034 -738
rect 2028 -750 2034 -744
rect 2028 -756 2034 -750
rect 2028 -762 2034 -756
rect 2028 -768 2034 -762
rect 2028 -774 2034 -768
rect 2028 -780 2034 -774
rect 2028 -786 2034 -780
rect 2028 -792 2034 -786
rect 2028 -798 2034 -792
rect 2028 -804 2034 -798
rect 2028 -810 2034 -804
rect 2028 -816 2034 -810
rect 2028 -822 2034 -816
rect 2028 -828 2034 -822
rect 2028 -834 2034 -828
rect 2028 -840 2034 -834
rect 2028 -846 2034 -840
rect 2028 -852 2034 -846
rect 2028 -858 2034 -852
rect 2028 -864 2034 -858
rect 2028 -870 2034 -864
rect 2028 -876 2034 -870
rect 2028 -882 2034 -876
rect 2028 -888 2034 -882
rect 2028 -894 2034 -888
rect 2028 -900 2034 -894
rect 2028 -906 2034 -900
rect 2028 -912 2034 -906
rect 2028 -918 2034 -912
rect 2028 -924 2034 -918
rect 2028 -930 2034 -924
rect 2028 -936 2034 -930
rect 2028 -942 2034 -936
rect 2028 -948 2034 -942
rect 2028 -954 2034 -948
rect 2028 -960 2034 -954
rect 2028 -966 2034 -960
rect 2028 -972 2034 -966
rect 2028 -978 2034 -972
rect 2028 -984 2034 -978
rect 2028 -990 2034 -984
rect 2028 -996 2034 -990
rect 2028 -1002 2034 -996
rect 2028 -1008 2034 -1002
rect 2028 -1014 2034 -1008
rect 2028 -1020 2034 -1014
rect 2028 -1026 2034 -1020
rect 2028 -1032 2034 -1026
rect 2028 -1038 2034 -1032
rect 2028 -1044 2034 -1038
rect 2028 -1050 2034 -1044
rect 2028 -1056 2034 -1050
rect 2028 -1062 2034 -1056
rect 2028 -1068 2034 -1062
rect 2028 -1074 2034 -1068
rect 2028 -1080 2034 -1074
rect 2028 -1086 2034 -1080
rect 2028 -1092 2034 -1086
rect 2028 -1098 2034 -1092
rect 2028 -1104 2034 -1098
rect 2028 -1110 2034 -1104
rect 2028 -1116 2034 -1110
rect 2028 -1122 2034 -1116
rect 2028 -1128 2034 -1122
rect 2028 -1134 2034 -1128
rect 2028 -1140 2034 -1134
rect 2028 -1146 2034 -1140
rect 2028 -1152 2034 -1146
rect 2028 -1158 2034 -1152
rect 2028 -1164 2034 -1158
rect 2028 -1170 2034 -1164
rect 2028 -1176 2034 -1170
rect 2028 -1182 2034 -1176
rect 2028 -1188 2034 -1182
rect 2028 -1194 2034 -1188
rect 2028 -1200 2034 -1194
rect 2028 -1206 2034 -1200
rect 2028 -1212 2034 -1206
rect 2028 -1218 2034 -1212
rect 2028 -1224 2034 -1218
rect 2028 -1230 2034 -1224
rect 2028 -1236 2034 -1230
rect 2028 -1242 2034 -1236
rect 2028 -1248 2034 -1242
rect 2028 -1254 2034 -1248
rect 2028 -1260 2034 -1254
rect 2028 -1266 2034 -1260
rect 2028 -1272 2034 -1266
rect 2028 -1278 2034 -1272
rect 2028 -1284 2034 -1278
rect 2028 -1290 2034 -1284
rect 2028 -1296 2034 -1290
rect 2028 -1302 2034 -1296
rect 2028 -1308 2034 -1302
rect 2028 -1314 2034 -1308
rect 2028 -1320 2034 -1314
rect 2028 -1326 2034 -1320
rect 2028 -1332 2034 -1326
rect 2028 -1338 2034 -1332
rect 2028 -1344 2034 -1338
rect 2028 -1350 2034 -1344
rect 2028 -1356 2034 -1350
rect 2028 -1362 2034 -1356
rect 2028 -1368 2034 -1362
rect 2028 -1374 2034 -1368
rect 2028 -1380 2034 -1374
rect 2028 -1386 2034 -1380
rect 2028 -1392 2034 -1386
rect 2028 -1398 2034 -1392
rect 2028 -1404 2034 -1398
rect 2028 -1410 2034 -1404
rect 2028 -1416 2034 -1410
rect 2028 -1422 2034 -1416
rect 2028 -1428 2034 -1422
rect 2028 -1434 2034 -1428
rect 2028 -1440 2034 -1434
rect 2028 -1446 2034 -1440
rect 2028 -1452 2034 -1446
rect 2028 -1458 2034 -1452
rect 2028 -1464 2034 -1458
rect 2028 -1470 2034 -1464
rect 2028 -1476 2034 -1470
rect 2028 -1482 2034 -1476
rect 2028 -1488 2034 -1482
rect 2028 -1494 2034 -1488
rect 2028 -1500 2034 -1494
rect 2028 -1506 2034 -1500
rect 2028 -1512 2034 -1506
rect 2028 -1518 2034 -1512
rect 2028 -1524 2034 -1518
rect 2028 -1530 2034 -1524
rect 2028 -1536 2034 -1530
rect 2028 -1542 2034 -1536
rect 2028 -1548 2034 -1542
rect 2028 -1554 2034 -1548
rect 2028 -1560 2034 -1554
rect 2028 -1566 2034 -1560
rect 2028 -1572 2034 -1566
rect 2028 -1578 2034 -1572
rect 2028 -1584 2034 -1578
rect 2028 -1590 2034 -1584
rect 2028 -1596 2034 -1590
rect 2028 -1602 2034 -1596
rect 2028 -1608 2034 -1602
rect 2028 -1614 2034 -1608
rect 2028 -1710 2034 -1704
rect 2028 -1716 2034 -1710
rect 2028 -1722 2034 -1716
rect 2028 -1728 2034 -1722
rect 2028 -1734 2034 -1728
rect 2028 -1740 2034 -1734
rect 2028 -1746 2034 -1740
rect 2028 -1752 2034 -1746
rect 2028 -1758 2034 -1752
rect 2028 -1764 2034 -1758
rect 2028 -1770 2034 -1764
rect 2028 -1776 2034 -1770
rect 2028 -1782 2034 -1776
rect 2028 -1788 2034 -1782
rect 2028 -1794 2034 -1788
rect 2028 -1800 2034 -1794
rect 2028 -1806 2034 -1800
rect 2028 -1812 2034 -1806
rect 2028 -1818 2034 -1812
rect 2028 -1824 2034 -1818
rect 2028 -1830 2034 -1824
rect 2028 -1836 2034 -1830
rect 2028 -1842 2034 -1836
rect 2028 -1848 2034 -1842
rect 2028 -1854 2034 -1848
rect 2028 -1860 2034 -1854
rect 2028 -1866 2034 -1860
rect 2028 -1872 2034 -1866
rect 2028 -1878 2034 -1872
rect 2028 -1884 2034 -1878
rect 2028 -1890 2034 -1884
rect 2028 -1896 2034 -1890
rect 2028 -1902 2034 -1896
rect 2028 -1908 2034 -1902
rect 2028 -1914 2034 -1908
rect 2028 -1920 2034 -1914
rect 2028 -1926 2034 -1920
rect 2028 -1932 2034 -1926
rect 2028 -1938 2034 -1932
rect 2028 -1944 2034 -1938
rect 2028 -1950 2034 -1944
rect 2028 -1956 2034 -1950
rect 2028 -1962 2034 -1956
rect 2028 -1968 2034 -1962
rect 2028 -1974 2034 -1968
rect 2028 -1980 2034 -1974
rect 2028 -1986 2034 -1980
rect 2028 -1992 2034 -1986
rect 2028 -1998 2034 -1992
rect 2028 -2004 2034 -1998
rect 2028 -2010 2034 -2004
rect 2028 -2016 2034 -2010
rect 2028 -2022 2034 -2016
rect 2028 -2028 2034 -2022
rect 2028 -2034 2034 -2028
rect 2028 -2040 2034 -2034
rect 2028 -2046 2034 -2040
rect 2028 -2052 2034 -2046
rect 2028 -2058 2034 -2052
rect 2028 -2064 2034 -2058
rect 2028 -2070 2034 -2064
rect 2028 -2076 2034 -2070
rect 2028 -2082 2034 -2076
rect 2028 -2088 2034 -2082
rect 2028 -2094 2034 -2088
rect 2028 -2100 2034 -2094
rect 2028 -2106 2034 -2100
rect 2028 -2112 2034 -2106
rect 2028 -2118 2034 -2112
rect 2028 -2124 2034 -2118
rect 2028 -2130 2034 -2124
rect 2028 -2136 2034 -2130
rect 2028 -2142 2034 -2136
rect 2028 -2148 2034 -2142
rect 2028 -2154 2034 -2148
rect 2028 -2160 2034 -2154
rect 2028 -2166 2034 -2160
rect 2028 -2172 2034 -2166
rect 2028 -2178 2034 -2172
rect 2028 -2184 2034 -2178
rect 2028 -2190 2034 -2184
rect 2028 -2196 2034 -2190
rect 2028 -2202 2034 -2196
rect 2028 -2208 2034 -2202
rect 2028 -2214 2034 -2208
rect 2028 -2220 2034 -2214
rect 2028 -2226 2034 -2220
rect 2028 -2232 2034 -2226
rect 2028 -2238 2034 -2232
rect 2028 -2244 2034 -2238
rect 2028 -2250 2034 -2244
rect 2028 -2256 2034 -2250
rect 2028 -2262 2034 -2256
rect 2028 -2268 2034 -2262
rect 2028 -2274 2034 -2268
rect 2028 -2280 2034 -2274
rect 2028 -2286 2034 -2280
rect 2028 -2292 2034 -2286
rect 2028 -2298 2034 -2292
rect 2028 -2304 2034 -2298
rect 2028 -2310 2034 -2304
rect 2028 -2316 2034 -2310
rect 2028 -2322 2034 -2316
rect 2028 -2328 2034 -2322
rect 2028 -2334 2034 -2328
rect 2028 -2340 2034 -2334
rect 2028 -2346 2034 -2340
rect 2028 -2352 2034 -2346
rect 2028 -2358 2034 -2352
rect 2028 -2364 2034 -2358
rect 2028 -2370 2034 -2364
rect 2028 -2376 2034 -2370
rect 2028 -2382 2034 -2376
rect 2028 -2388 2034 -2382
rect 2028 -2394 2034 -2388
rect 2028 -2400 2034 -2394
rect 2028 -2406 2034 -2400
rect 2028 -2412 2034 -2406
rect 2028 -2418 2034 -2412
rect 2028 -2424 2034 -2418
rect 2028 -2430 2034 -2424
rect 2028 -2436 2034 -2430
rect 2028 -2442 2034 -2436
rect 2028 -2448 2034 -2442
rect 2028 -2454 2034 -2448
rect 2028 -2460 2034 -2454
rect 2028 -2466 2034 -2460
rect 2028 -2472 2034 -2466
rect 2028 -2478 2034 -2472
rect 2028 -2484 2034 -2478
rect 2028 -2490 2034 -2484
rect 2028 -2496 2034 -2490
rect 2028 -2502 2034 -2496
rect 2028 -2508 2034 -2502
rect 2028 -2514 2034 -2508
rect 2028 -2598 2034 -2592
rect 2028 -2604 2034 -2598
rect 2028 -2610 2034 -2604
rect 2028 -2616 2034 -2610
rect 2028 -2622 2034 -2616
rect 2028 -2628 2034 -2622
rect 2028 -2634 2034 -2628
rect 2028 -2640 2034 -2634
rect 2028 -2646 2034 -2640
rect 2028 -2652 2034 -2646
rect 2028 -2658 2034 -2652
rect 2028 -2664 2034 -2658
rect 2028 -2670 2034 -2664
rect 2028 -2676 2034 -2670
rect 2028 -2682 2034 -2676
rect 2028 -2688 2034 -2682
rect 2028 -2694 2034 -2688
rect 2028 -2700 2034 -2694
rect 2028 -2706 2034 -2700
rect 2028 -2712 2034 -2706
rect 2028 -2718 2034 -2712
rect 2028 -2724 2034 -2718
rect 2028 -2730 2034 -2724
rect 2028 -2736 2034 -2730
rect 2028 -2742 2034 -2736
rect 2028 -2748 2034 -2742
rect 2028 -2754 2034 -2748
rect 2028 -2760 2034 -2754
rect 2028 -2766 2034 -2760
rect 2028 -2772 2034 -2766
rect 2028 -2778 2034 -2772
rect 2028 -2784 2034 -2778
rect 2028 -2790 2034 -2784
rect 2028 -2796 2034 -2790
rect 2028 -2802 2034 -2796
rect 2028 -2808 2034 -2802
rect 2028 -2814 2034 -2808
rect 2028 -2820 2034 -2814
rect 2028 -2826 2034 -2820
rect 2028 -2832 2034 -2826
rect 2028 -2838 2034 -2832
rect 2028 -2844 2034 -2838
rect 2028 -2850 2034 -2844
rect 2028 -2856 2034 -2850
rect 2028 -2862 2034 -2856
rect 2028 -2868 2034 -2862
rect 2028 -2874 2034 -2868
rect 2028 -2880 2034 -2874
rect 2028 -2886 2034 -2880
rect 2028 -2892 2034 -2886
rect 2028 -2898 2034 -2892
rect 2028 -2904 2034 -2898
rect 2028 -2910 2034 -2904
rect 2028 -2916 2034 -2910
rect 2028 -2922 2034 -2916
rect 2028 -2928 2034 -2922
rect 2028 -2934 2034 -2928
rect 2028 -2940 2034 -2934
rect 2028 -2946 2034 -2940
rect 2028 -2952 2034 -2946
rect 2028 -2958 2034 -2952
rect 2028 -2964 2034 -2958
rect 2028 -2970 2034 -2964
rect 2028 -2976 2034 -2970
rect 2028 -2982 2034 -2976
rect 2028 -2988 2034 -2982
rect 2028 -2994 2034 -2988
rect 2028 -3000 2034 -2994
rect 2028 -3006 2034 -3000
rect 2028 -3012 2034 -3006
rect 2028 -3018 2034 -3012
rect 2028 -3024 2034 -3018
rect 2028 -3030 2034 -3024
rect 2028 -3036 2034 -3030
rect 2028 -3042 2034 -3036
rect 2028 -3048 2034 -3042
rect 2028 -3054 2034 -3048
rect 2028 -3060 2034 -3054
rect 2028 -3066 2034 -3060
rect 2028 -3072 2034 -3066
rect 2028 -3078 2034 -3072
rect 2028 -3084 2034 -3078
rect 2028 -3090 2034 -3084
rect 2028 -3096 2034 -3090
rect 2028 -3150 2034 -3144
rect 2028 -3156 2034 -3150
rect 2028 -3162 2034 -3156
rect 2028 -3168 2034 -3162
rect 2028 -3174 2034 -3168
rect 2028 -3180 2034 -3174
rect 2028 -3186 2034 -3180
rect 2028 -3192 2034 -3186
rect 2034 -408 2040 -402
rect 2034 -414 2040 -408
rect 2034 -420 2040 -414
rect 2034 -426 2040 -420
rect 2034 -432 2040 -426
rect 2034 -438 2040 -432
rect 2034 -444 2040 -438
rect 2034 -450 2040 -444
rect 2034 -456 2040 -450
rect 2034 -462 2040 -456
rect 2034 -468 2040 -462
rect 2034 -474 2040 -468
rect 2034 -480 2040 -474
rect 2034 -486 2040 -480
rect 2034 -492 2040 -486
rect 2034 -498 2040 -492
rect 2034 -504 2040 -498
rect 2034 -510 2040 -504
rect 2034 -516 2040 -510
rect 2034 -522 2040 -516
rect 2034 -528 2040 -522
rect 2034 -534 2040 -528
rect 2034 -540 2040 -534
rect 2034 -546 2040 -540
rect 2034 -552 2040 -546
rect 2034 -558 2040 -552
rect 2034 -564 2040 -558
rect 2034 -570 2040 -564
rect 2034 -576 2040 -570
rect 2034 -582 2040 -576
rect 2034 -588 2040 -582
rect 2034 -594 2040 -588
rect 2034 -600 2040 -594
rect 2034 -606 2040 -600
rect 2034 -612 2040 -606
rect 2034 -618 2040 -612
rect 2034 -624 2040 -618
rect 2034 -630 2040 -624
rect 2034 -636 2040 -630
rect 2034 -642 2040 -636
rect 2034 -648 2040 -642
rect 2034 -654 2040 -648
rect 2034 -660 2040 -654
rect 2034 -666 2040 -660
rect 2034 -672 2040 -666
rect 2034 -678 2040 -672
rect 2034 -684 2040 -678
rect 2034 -690 2040 -684
rect 2034 -696 2040 -690
rect 2034 -702 2040 -696
rect 2034 -708 2040 -702
rect 2034 -714 2040 -708
rect 2034 -720 2040 -714
rect 2034 -726 2040 -720
rect 2034 -732 2040 -726
rect 2034 -738 2040 -732
rect 2034 -744 2040 -738
rect 2034 -750 2040 -744
rect 2034 -756 2040 -750
rect 2034 -762 2040 -756
rect 2034 -768 2040 -762
rect 2034 -774 2040 -768
rect 2034 -780 2040 -774
rect 2034 -786 2040 -780
rect 2034 -792 2040 -786
rect 2034 -798 2040 -792
rect 2034 -804 2040 -798
rect 2034 -810 2040 -804
rect 2034 -816 2040 -810
rect 2034 -822 2040 -816
rect 2034 -828 2040 -822
rect 2034 -834 2040 -828
rect 2034 -840 2040 -834
rect 2034 -846 2040 -840
rect 2034 -852 2040 -846
rect 2034 -858 2040 -852
rect 2034 -864 2040 -858
rect 2034 -870 2040 -864
rect 2034 -876 2040 -870
rect 2034 -882 2040 -876
rect 2034 -888 2040 -882
rect 2034 -894 2040 -888
rect 2034 -900 2040 -894
rect 2034 -906 2040 -900
rect 2034 -912 2040 -906
rect 2034 -918 2040 -912
rect 2034 -924 2040 -918
rect 2034 -930 2040 -924
rect 2034 -936 2040 -930
rect 2034 -942 2040 -936
rect 2034 -948 2040 -942
rect 2034 -954 2040 -948
rect 2034 -960 2040 -954
rect 2034 -966 2040 -960
rect 2034 -972 2040 -966
rect 2034 -978 2040 -972
rect 2034 -984 2040 -978
rect 2034 -990 2040 -984
rect 2034 -996 2040 -990
rect 2034 -1002 2040 -996
rect 2034 -1008 2040 -1002
rect 2034 -1014 2040 -1008
rect 2034 -1020 2040 -1014
rect 2034 -1026 2040 -1020
rect 2034 -1032 2040 -1026
rect 2034 -1038 2040 -1032
rect 2034 -1044 2040 -1038
rect 2034 -1050 2040 -1044
rect 2034 -1056 2040 -1050
rect 2034 -1062 2040 -1056
rect 2034 -1068 2040 -1062
rect 2034 -1074 2040 -1068
rect 2034 -1080 2040 -1074
rect 2034 -1086 2040 -1080
rect 2034 -1092 2040 -1086
rect 2034 -1098 2040 -1092
rect 2034 -1104 2040 -1098
rect 2034 -1110 2040 -1104
rect 2034 -1116 2040 -1110
rect 2034 -1122 2040 -1116
rect 2034 -1128 2040 -1122
rect 2034 -1134 2040 -1128
rect 2034 -1140 2040 -1134
rect 2034 -1146 2040 -1140
rect 2034 -1152 2040 -1146
rect 2034 -1158 2040 -1152
rect 2034 -1164 2040 -1158
rect 2034 -1170 2040 -1164
rect 2034 -1176 2040 -1170
rect 2034 -1182 2040 -1176
rect 2034 -1188 2040 -1182
rect 2034 -1194 2040 -1188
rect 2034 -1200 2040 -1194
rect 2034 -1206 2040 -1200
rect 2034 -1212 2040 -1206
rect 2034 -1218 2040 -1212
rect 2034 -1224 2040 -1218
rect 2034 -1230 2040 -1224
rect 2034 -1236 2040 -1230
rect 2034 -1242 2040 -1236
rect 2034 -1248 2040 -1242
rect 2034 -1254 2040 -1248
rect 2034 -1260 2040 -1254
rect 2034 -1266 2040 -1260
rect 2034 -1272 2040 -1266
rect 2034 -1278 2040 -1272
rect 2034 -1284 2040 -1278
rect 2034 -1290 2040 -1284
rect 2034 -1296 2040 -1290
rect 2034 -1302 2040 -1296
rect 2034 -1308 2040 -1302
rect 2034 -1314 2040 -1308
rect 2034 -1320 2040 -1314
rect 2034 -1326 2040 -1320
rect 2034 -1332 2040 -1326
rect 2034 -1338 2040 -1332
rect 2034 -1344 2040 -1338
rect 2034 -1350 2040 -1344
rect 2034 -1356 2040 -1350
rect 2034 -1362 2040 -1356
rect 2034 -1368 2040 -1362
rect 2034 -1374 2040 -1368
rect 2034 -1380 2040 -1374
rect 2034 -1386 2040 -1380
rect 2034 -1392 2040 -1386
rect 2034 -1398 2040 -1392
rect 2034 -1404 2040 -1398
rect 2034 -1410 2040 -1404
rect 2034 -1416 2040 -1410
rect 2034 -1422 2040 -1416
rect 2034 -1428 2040 -1422
rect 2034 -1434 2040 -1428
rect 2034 -1440 2040 -1434
rect 2034 -1446 2040 -1440
rect 2034 -1452 2040 -1446
rect 2034 -1458 2040 -1452
rect 2034 -1464 2040 -1458
rect 2034 -1470 2040 -1464
rect 2034 -1476 2040 -1470
rect 2034 -1482 2040 -1476
rect 2034 -1488 2040 -1482
rect 2034 -1494 2040 -1488
rect 2034 -1500 2040 -1494
rect 2034 -1506 2040 -1500
rect 2034 -1512 2040 -1506
rect 2034 -1518 2040 -1512
rect 2034 -1524 2040 -1518
rect 2034 -1530 2040 -1524
rect 2034 -1536 2040 -1530
rect 2034 -1542 2040 -1536
rect 2034 -1548 2040 -1542
rect 2034 -1554 2040 -1548
rect 2034 -1560 2040 -1554
rect 2034 -1566 2040 -1560
rect 2034 -1572 2040 -1566
rect 2034 -1578 2040 -1572
rect 2034 -1584 2040 -1578
rect 2034 -1590 2040 -1584
rect 2034 -1596 2040 -1590
rect 2034 -1602 2040 -1596
rect 2034 -1608 2040 -1602
rect 2034 -1704 2040 -1698
rect 2034 -1710 2040 -1704
rect 2034 -1716 2040 -1710
rect 2034 -1722 2040 -1716
rect 2034 -1728 2040 -1722
rect 2034 -1734 2040 -1728
rect 2034 -1740 2040 -1734
rect 2034 -1746 2040 -1740
rect 2034 -1752 2040 -1746
rect 2034 -1758 2040 -1752
rect 2034 -1764 2040 -1758
rect 2034 -1770 2040 -1764
rect 2034 -1776 2040 -1770
rect 2034 -1782 2040 -1776
rect 2034 -1788 2040 -1782
rect 2034 -1794 2040 -1788
rect 2034 -1800 2040 -1794
rect 2034 -1806 2040 -1800
rect 2034 -1812 2040 -1806
rect 2034 -1818 2040 -1812
rect 2034 -1824 2040 -1818
rect 2034 -1830 2040 -1824
rect 2034 -1836 2040 -1830
rect 2034 -1842 2040 -1836
rect 2034 -1848 2040 -1842
rect 2034 -1854 2040 -1848
rect 2034 -1860 2040 -1854
rect 2034 -1866 2040 -1860
rect 2034 -1872 2040 -1866
rect 2034 -1878 2040 -1872
rect 2034 -1884 2040 -1878
rect 2034 -1890 2040 -1884
rect 2034 -1896 2040 -1890
rect 2034 -1902 2040 -1896
rect 2034 -1908 2040 -1902
rect 2034 -1914 2040 -1908
rect 2034 -1920 2040 -1914
rect 2034 -1926 2040 -1920
rect 2034 -1932 2040 -1926
rect 2034 -1938 2040 -1932
rect 2034 -1944 2040 -1938
rect 2034 -1950 2040 -1944
rect 2034 -1956 2040 -1950
rect 2034 -1962 2040 -1956
rect 2034 -1968 2040 -1962
rect 2034 -1974 2040 -1968
rect 2034 -1980 2040 -1974
rect 2034 -1986 2040 -1980
rect 2034 -1992 2040 -1986
rect 2034 -1998 2040 -1992
rect 2034 -2004 2040 -1998
rect 2034 -2010 2040 -2004
rect 2034 -2016 2040 -2010
rect 2034 -2022 2040 -2016
rect 2034 -2028 2040 -2022
rect 2034 -2034 2040 -2028
rect 2034 -2040 2040 -2034
rect 2034 -2046 2040 -2040
rect 2034 -2052 2040 -2046
rect 2034 -2058 2040 -2052
rect 2034 -2064 2040 -2058
rect 2034 -2070 2040 -2064
rect 2034 -2076 2040 -2070
rect 2034 -2082 2040 -2076
rect 2034 -2088 2040 -2082
rect 2034 -2094 2040 -2088
rect 2034 -2100 2040 -2094
rect 2034 -2106 2040 -2100
rect 2034 -2112 2040 -2106
rect 2034 -2118 2040 -2112
rect 2034 -2124 2040 -2118
rect 2034 -2130 2040 -2124
rect 2034 -2136 2040 -2130
rect 2034 -2142 2040 -2136
rect 2034 -2148 2040 -2142
rect 2034 -2154 2040 -2148
rect 2034 -2160 2040 -2154
rect 2034 -2166 2040 -2160
rect 2034 -2172 2040 -2166
rect 2034 -2178 2040 -2172
rect 2034 -2184 2040 -2178
rect 2034 -2190 2040 -2184
rect 2034 -2196 2040 -2190
rect 2034 -2202 2040 -2196
rect 2034 -2208 2040 -2202
rect 2034 -2214 2040 -2208
rect 2034 -2220 2040 -2214
rect 2034 -2226 2040 -2220
rect 2034 -2232 2040 -2226
rect 2034 -2238 2040 -2232
rect 2034 -2244 2040 -2238
rect 2034 -2250 2040 -2244
rect 2034 -2256 2040 -2250
rect 2034 -2262 2040 -2256
rect 2034 -2268 2040 -2262
rect 2034 -2274 2040 -2268
rect 2034 -2280 2040 -2274
rect 2034 -2286 2040 -2280
rect 2034 -2292 2040 -2286
rect 2034 -2298 2040 -2292
rect 2034 -2304 2040 -2298
rect 2034 -2310 2040 -2304
rect 2034 -2316 2040 -2310
rect 2034 -2322 2040 -2316
rect 2034 -2328 2040 -2322
rect 2034 -2334 2040 -2328
rect 2034 -2340 2040 -2334
rect 2034 -2346 2040 -2340
rect 2034 -2352 2040 -2346
rect 2034 -2358 2040 -2352
rect 2034 -2364 2040 -2358
rect 2034 -2370 2040 -2364
rect 2034 -2376 2040 -2370
rect 2034 -2382 2040 -2376
rect 2034 -2388 2040 -2382
rect 2034 -2394 2040 -2388
rect 2034 -2400 2040 -2394
rect 2034 -2406 2040 -2400
rect 2034 -2412 2040 -2406
rect 2034 -2418 2040 -2412
rect 2034 -2424 2040 -2418
rect 2034 -2430 2040 -2424
rect 2034 -2436 2040 -2430
rect 2034 -2442 2040 -2436
rect 2034 -2448 2040 -2442
rect 2034 -2454 2040 -2448
rect 2034 -2460 2040 -2454
rect 2034 -2466 2040 -2460
rect 2034 -2472 2040 -2466
rect 2034 -2478 2040 -2472
rect 2034 -2484 2040 -2478
rect 2034 -2490 2040 -2484
rect 2034 -2496 2040 -2490
rect 2034 -2502 2040 -2496
rect 2034 -2508 2040 -2502
rect 2034 -2598 2040 -2592
rect 2034 -2604 2040 -2598
rect 2034 -2610 2040 -2604
rect 2034 -2616 2040 -2610
rect 2034 -2622 2040 -2616
rect 2034 -2628 2040 -2622
rect 2034 -2634 2040 -2628
rect 2034 -2640 2040 -2634
rect 2034 -2646 2040 -2640
rect 2034 -2652 2040 -2646
rect 2034 -2658 2040 -2652
rect 2034 -2664 2040 -2658
rect 2034 -2670 2040 -2664
rect 2034 -2676 2040 -2670
rect 2034 -2682 2040 -2676
rect 2034 -2688 2040 -2682
rect 2034 -2694 2040 -2688
rect 2034 -2700 2040 -2694
rect 2034 -2706 2040 -2700
rect 2034 -2712 2040 -2706
rect 2034 -2718 2040 -2712
rect 2034 -2724 2040 -2718
rect 2034 -2730 2040 -2724
rect 2034 -2736 2040 -2730
rect 2034 -2742 2040 -2736
rect 2034 -2748 2040 -2742
rect 2034 -2754 2040 -2748
rect 2034 -2760 2040 -2754
rect 2034 -2766 2040 -2760
rect 2034 -2772 2040 -2766
rect 2034 -2778 2040 -2772
rect 2034 -2784 2040 -2778
rect 2034 -2790 2040 -2784
rect 2034 -2796 2040 -2790
rect 2034 -2802 2040 -2796
rect 2034 -2808 2040 -2802
rect 2034 -2814 2040 -2808
rect 2034 -2820 2040 -2814
rect 2034 -2826 2040 -2820
rect 2034 -2832 2040 -2826
rect 2034 -2838 2040 -2832
rect 2034 -2844 2040 -2838
rect 2034 -2850 2040 -2844
rect 2034 -2856 2040 -2850
rect 2034 -2862 2040 -2856
rect 2034 -2868 2040 -2862
rect 2034 -2874 2040 -2868
rect 2034 -2880 2040 -2874
rect 2034 -2886 2040 -2880
rect 2034 -2892 2040 -2886
rect 2034 -2898 2040 -2892
rect 2034 -2904 2040 -2898
rect 2034 -2910 2040 -2904
rect 2034 -2916 2040 -2910
rect 2034 -2922 2040 -2916
rect 2034 -2928 2040 -2922
rect 2034 -2934 2040 -2928
rect 2034 -2940 2040 -2934
rect 2034 -2946 2040 -2940
rect 2034 -2952 2040 -2946
rect 2034 -2958 2040 -2952
rect 2034 -2964 2040 -2958
rect 2034 -2970 2040 -2964
rect 2034 -2976 2040 -2970
rect 2034 -2982 2040 -2976
rect 2034 -2988 2040 -2982
rect 2034 -2994 2040 -2988
rect 2034 -3000 2040 -2994
rect 2034 -3006 2040 -3000
rect 2034 -3012 2040 -3006
rect 2034 -3018 2040 -3012
rect 2034 -3024 2040 -3018
rect 2034 -3030 2040 -3024
rect 2034 -3036 2040 -3030
rect 2034 -3042 2040 -3036
rect 2034 -3048 2040 -3042
rect 2034 -3054 2040 -3048
rect 2034 -3060 2040 -3054
rect 2034 -3066 2040 -3060
rect 2034 -3072 2040 -3066
rect 2034 -3078 2040 -3072
rect 2034 -3084 2040 -3078
rect 2034 -3090 2040 -3084
rect 2034 -3144 2040 -3138
rect 2034 -3150 2040 -3144
rect 2034 -3156 2040 -3150
rect 2034 -3162 2040 -3156
rect 2034 -3168 2040 -3162
rect 2034 -3174 2040 -3168
rect 2034 -3180 2040 -3174
rect 2034 -3186 2040 -3180
rect 2040 -402 2046 -396
rect 2040 -408 2046 -402
rect 2040 -414 2046 -408
rect 2040 -420 2046 -414
rect 2040 -426 2046 -420
rect 2040 -432 2046 -426
rect 2040 -438 2046 -432
rect 2040 -444 2046 -438
rect 2040 -450 2046 -444
rect 2040 -456 2046 -450
rect 2040 -462 2046 -456
rect 2040 -468 2046 -462
rect 2040 -474 2046 -468
rect 2040 -480 2046 -474
rect 2040 -486 2046 -480
rect 2040 -492 2046 -486
rect 2040 -498 2046 -492
rect 2040 -504 2046 -498
rect 2040 -510 2046 -504
rect 2040 -516 2046 -510
rect 2040 -522 2046 -516
rect 2040 -528 2046 -522
rect 2040 -534 2046 -528
rect 2040 -540 2046 -534
rect 2040 -546 2046 -540
rect 2040 -552 2046 -546
rect 2040 -558 2046 -552
rect 2040 -564 2046 -558
rect 2040 -570 2046 -564
rect 2040 -576 2046 -570
rect 2040 -582 2046 -576
rect 2040 -588 2046 -582
rect 2040 -594 2046 -588
rect 2040 -600 2046 -594
rect 2040 -606 2046 -600
rect 2040 -612 2046 -606
rect 2040 -618 2046 -612
rect 2040 -624 2046 -618
rect 2040 -630 2046 -624
rect 2040 -636 2046 -630
rect 2040 -642 2046 -636
rect 2040 -648 2046 -642
rect 2040 -654 2046 -648
rect 2040 -660 2046 -654
rect 2040 -666 2046 -660
rect 2040 -672 2046 -666
rect 2040 -678 2046 -672
rect 2040 -684 2046 -678
rect 2040 -690 2046 -684
rect 2040 -696 2046 -690
rect 2040 -702 2046 -696
rect 2040 -708 2046 -702
rect 2040 -714 2046 -708
rect 2040 -720 2046 -714
rect 2040 -726 2046 -720
rect 2040 -732 2046 -726
rect 2040 -738 2046 -732
rect 2040 -744 2046 -738
rect 2040 -750 2046 -744
rect 2040 -756 2046 -750
rect 2040 -762 2046 -756
rect 2040 -768 2046 -762
rect 2040 -774 2046 -768
rect 2040 -780 2046 -774
rect 2040 -786 2046 -780
rect 2040 -792 2046 -786
rect 2040 -798 2046 -792
rect 2040 -804 2046 -798
rect 2040 -810 2046 -804
rect 2040 -816 2046 -810
rect 2040 -822 2046 -816
rect 2040 -828 2046 -822
rect 2040 -834 2046 -828
rect 2040 -840 2046 -834
rect 2040 -846 2046 -840
rect 2040 -852 2046 -846
rect 2040 -858 2046 -852
rect 2040 -864 2046 -858
rect 2040 -870 2046 -864
rect 2040 -876 2046 -870
rect 2040 -882 2046 -876
rect 2040 -888 2046 -882
rect 2040 -894 2046 -888
rect 2040 -900 2046 -894
rect 2040 -906 2046 -900
rect 2040 -912 2046 -906
rect 2040 -918 2046 -912
rect 2040 -924 2046 -918
rect 2040 -930 2046 -924
rect 2040 -936 2046 -930
rect 2040 -942 2046 -936
rect 2040 -948 2046 -942
rect 2040 -954 2046 -948
rect 2040 -960 2046 -954
rect 2040 -966 2046 -960
rect 2040 -972 2046 -966
rect 2040 -978 2046 -972
rect 2040 -984 2046 -978
rect 2040 -990 2046 -984
rect 2040 -996 2046 -990
rect 2040 -1002 2046 -996
rect 2040 -1008 2046 -1002
rect 2040 -1014 2046 -1008
rect 2040 -1020 2046 -1014
rect 2040 -1026 2046 -1020
rect 2040 -1032 2046 -1026
rect 2040 -1038 2046 -1032
rect 2040 -1044 2046 -1038
rect 2040 -1050 2046 -1044
rect 2040 -1056 2046 -1050
rect 2040 -1062 2046 -1056
rect 2040 -1068 2046 -1062
rect 2040 -1074 2046 -1068
rect 2040 -1080 2046 -1074
rect 2040 -1086 2046 -1080
rect 2040 -1092 2046 -1086
rect 2040 -1098 2046 -1092
rect 2040 -1104 2046 -1098
rect 2040 -1110 2046 -1104
rect 2040 -1116 2046 -1110
rect 2040 -1122 2046 -1116
rect 2040 -1128 2046 -1122
rect 2040 -1134 2046 -1128
rect 2040 -1140 2046 -1134
rect 2040 -1146 2046 -1140
rect 2040 -1152 2046 -1146
rect 2040 -1158 2046 -1152
rect 2040 -1164 2046 -1158
rect 2040 -1170 2046 -1164
rect 2040 -1176 2046 -1170
rect 2040 -1182 2046 -1176
rect 2040 -1188 2046 -1182
rect 2040 -1194 2046 -1188
rect 2040 -1200 2046 -1194
rect 2040 -1206 2046 -1200
rect 2040 -1212 2046 -1206
rect 2040 -1218 2046 -1212
rect 2040 -1224 2046 -1218
rect 2040 -1230 2046 -1224
rect 2040 -1236 2046 -1230
rect 2040 -1242 2046 -1236
rect 2040 -1248 2046 -1242
rect 2040 -1254 2046 -1248
rect 2040 -1260 2046 -1254
rect 2040 -1266 2046 -1260
rect 2040 -1272 2046 -1266
rect 2040 -1278 2046 -1272
rect 2040 -1284 2046 -1278
rect 2040 -1290 2046 -1284
rect 2040 -1296 2046 -1290
rect 2040 -1302 2046 -1296
rect 2040 -1308 2046 -1302
rect 2040 -1314 2046 -1308
rect 2040 -1320 2046 -1314
rect 2040 -1326 2046 -1320
rect 2040 -1332 2046 -1326
rect 2040 -1338 2046 -1332
rect 2040 -1344 2046 -1338
rect 2040 -1350 2046 -1344
rect 2040 -1356 2046 -1350
rect 2040 -1362 2046 -1356
rect 2040 -1368 2046 -1362
rect 2040 -1374 2046 -1368
rect 2040 -1380 2046 -1374
rect 2040 -1386 2046 -1380
rect 2040 -1392 2046 -1386
rect 2040 -1398 2046 -1392
rect 2040 -1404 2046 -1398
rect 2040 -1410 2046 -1404
rect 2040 -1416 2046 -1410
rect 2040 -1422 2046 -1416
rect 2040 -1428 2046 -1422
rect 2040 -1434 2046 -1428
rect 2040 -1440 2046 -1434
rect 2040 -1446 2046 -1440
rect 2040 -1452 2046 -1446
rect 2040 -1458 2046 -1452
rect 2040 -1464 2046 -1458
rect 2040 -1470 2046 -1464
rect 2040 -1476 2046 -1470
rect 2040 -1482 2046 -1476
rect 2040 -1488 2046 -1482
rect 2040 -1494 2046 -1488
rect 2040 -1500 2046 -1494
rect 2040 -1506 2046 -1500
rect 2040 -1512 2046 -1506
rect 2040 -1518 2046 -1512
rect 2040 -1524 2046 -1518
rect 2040 -1530 2046 -1524
rect 2040 -1536 2046 -1530
rect 2040 -1542 2046 -1536
rect 2040 -1548 2046 -1542
rect 2040 -1554 2046 -1548
rect 2040 -1560 2046 -1554
rect 2040 -1566 2046 -1560
rect 2040 -1572 2046 -1566
rect 2040 -1578 2046 -1572
rect 2040 -1584 2046 -1578
rect 2040 -1590 2046 -1584
rect 2040 -1596 2046 -1590
rect 2040 -1602 2046 -1596
rect 2040 -1698 2046 -1692
rect 2040 -1704 2046 -1698
rect 2040 -1710 2046 -1704
rect 2040 -1716 2046 -1710
rect 2040 -1722 2046 -1716
rect 2040 -1728 2046 -1722
rect 2040 -1734 2046 -1728
rect 2040 -1740 2046 -1734
rect 2040 -1746 2046 -1740
rect 2040 -1752 2046 -1746
rect 2040 -1758 2046 -1752
rect 2040 -1764 2046 -1758
rect 2040 -1770 2046 -1764
rect 2040 -1776 2046 -1770
rect 2040 -1782 2046 -1776
rect 2040 -1788 2046 -1782
rect 2040 -1794 2046 -1788
rect 2040 -1800 2046 -1794
rect 2040 -1806 2046 -1800
rect 2040 -1812 2046 -1806
rect 2040 -1818 2046 -1812
rect 2040 -1824 2046 -1818
rect 2040 -1830 2046 -1824
rect 2040 -1836 2046 -1830
rect 2040 -1842 2046 -1836
rect 2040 -1848 2046 -1842
rect 2040 -1854 2046 -1848
rect 2040 -1860 2046 -1854
rect 2040 -1866 2046 -1860
rect 2040 -1872 2046 -1866
rect 2040 -1878 2046 -1872
rect 2040 -1884 2046 -1878
rect 2040 -1890 2046 -1884
rect 2040 -1896 2046 -1890
rect 2040 -1902 2046 -1896
rect 2040 -1908 2046 -1902
rect 2040 -1914 2046 -1908
rect 2040 -1920 2046 -1914
rect 2040 -1926 2046 -1920
rect 2040 -1932 2046 -1926
rect 2040 -1938 2046 -1932
rect 2040 -1944 2046 -1938
rect 2040 -1950 2046 -1944
rect 2040 -1956 2046 -1950
rect 2040 -1962 2046 -1956
rect 2040 -1968 2046 -1962
rect 2040 -1974 2046 -1968
rect 2040 -1980 2046 -1974
rect 2040 -1986 2046 -1980
rect 2040 -1992 2046 -1986
rect 2040 -1998 2046 -1992
rect 2040 -2004 2046 -1998
rect 2040 -2010 2046 -2004
rect 2040 -2016 2046 -2010
rect 2040 -2022 2046 -2016
rect 2040 -2028 2046 -2022
rect 2040 -2034 2046 -2028
rect 2040 -2040 2046 -2034
rect 2040 -2046 2046 -2040
rect 2040 -2052 2046 -2046
rect 2040 -2058 2046 -2052
rect 2040 -2064 2046 -2058
rect 2040 -2070 2046 -2064
rect 2040 -2076 2046 -2070
rect 2040 -2082 2046 -2076
rect 2040 -2088 2046 -2082
rect 2040 -2094 2046 -2088
rect 2040 -2100 2046 -2094
rect 2040 -2106 2046 -2100
rect 2040 -2112 2046 -2106
rect 2040 -2118 2046 -2112
rect 2040 -2124 2046 -2118
rect 2040 -2130 2046 -2124
rect 2040 -2136 2046 -2130
rect 2040 -2142 2046 -2136
rect 2040 -2148 2046 -2142
rect 2040 -2154 2046 -2148
rect 2040 -2160 2046 -2154
rect 2040 -2166 2046 -2160
rect 2040 -2172 2046 -2166
rect 2040 -2178 2046 -2172
rect 2040 -2184 2046 -2178
rect 2040 -2190 2046 -2184
rect 2040 -2196 2046 -2190
rect 2040 -2202 2046 -2196
rect 2040 -2208 2046 -2202
rect 2040 -2214 2046 -2208
rect 2040 -2220 2046 -2214
rect 2040 -2226 2046 -2220
rect 2040 -2232 2046 -2226
rect 2040 -2238 2046 -2232
rect 2040 -2244 2046 -2238
rect 2040 -2250 2046 -2244
rect 2040 -2256 2046 -2250
rect 2040 -2262 2046 -2256
rect 2040 -2268 2046 -2262
rect 2040 -2274 2046 -2268
rect 2040 -2280 2046 -2274
rect 2040 -2286 2046 -2280
rect 2040 -2292 2046 -2286
rect 2040 -2298 2046 -2292
rect 2040 -2304 2046 -2298
rect 2040 -2310 2046 -2304
rect 2040 -2316 2046 -2310
rect 2040 -2322 2046 -2316
rect 2040 -2328 2046 -2322
rect 2040 -2334 2046 -2328
rect 2040 -2340 2046 -2334
rect 2040 -2346 2046 -2340
rect 2040 -2352 2046 -2346
rect 2040 -2358 2046 -2352
rect 2040 -2364 2046 -2358
rect 2040 -2370 2046 -2364
rect 2040 -2376 2046 -2370
rect 2040 -2382 2046 -2376
rect 2040 -2388 2046 -2382
rect 2040 -2394 2046 -2388
rect 2040 -2400 2046 -2394
rect 2040 -2406 2046 -2400
rect 2040 -2412 2046 -2406
rect 2040 -2418 2046 -2412
rect 2040 -2424 2046 -2418
rect 2040 -2430 2046 -2424
rect 2040 -2436 2046 -2430
rect 2040 -2442 2046 -2436
rect 2040 -2448 2046 -2442
rect 2040 -2454 2046 -2448
rect 2040 -2460 2046 -2454
rect 2040 -2466 2046 -2460
rect 2040 -2472 2046 -2466
rect 2040 -2478 2046 -2472
rect 2040 -2484 2046 -2478
rect 2040 -2490 2046 -2484
rect 2040 -2496 2046 -2490
rect 2040 -2502 2046 -2496
rect 2040 -2508 2046 -2502
rect 2040 -2598 2046 -2592
rect 2040 -2604 2046 -2598
rect 2040 -2610 2046 -2604
rect 2040 -2616 2046 -2610
rect 2040 -2622 2046 -2616
rect 2040 -2628 2046 -2622
rect 2040 -2634 2046 -2628
rect 2040 -2640 2046 -2634
rect 2040 -2646 2046 -2640
rect 2040 -2652 2046 -2646
rect 2040 -2658 2046 -2652
rect 2040 -2664 2046 -2658
rect 2040 -2670 2046 -2664
rect 2040 -2676 2046 -2670
rect 2040 -2682 2046 -2676
rect 2040 -2688 2046 -2682
rect 2040 -2694 2046 -2688
rect 2040 -2700 2046 -2694
rect 2040 -2706 2046 -2700
rect 2040 -2712 2046 -2706
rect 2040 -2718 2046 -2712
rect 2040 -2724 2046 -2718
rect 2040 -2730 2046 -2724
rect 2040 -2736 2046 -2730
rect 2040 -2742 2046 -2736
rect 2040 -2748 2046 -2742
rect 2040 -2754 2046 -2748
rect 2040 -2760 2046 -2754
rect 2040 -2766 2046 -2760
rect 2040 -2772 2046 -2766
rect 2040 -2778 2046 -2772
rect 2040 -2784 2046 -2778
rect 2040 -2790 2046 -2784
rect 2040 -2796 2046 -2790
rect 2040 -2802 2046 -2796
rect 2040 -2808 2046 -2802
rect 2040 -2814 2046 -2808
rect 2040 -2820 2046 -2814
rect 2040 -2826 2046 -2820
rect 2040 -2832 2046 -2826
rect 2040 -2838 2046 -2832
rect 2040 -2844 2046 -2838
rect 2040 -2850 2046 -2844
rect 2040 -2856 2046 -2850
rect 2040 -2862 2046 -2856
rect 2040 -2868 2046 -2862
rect 2040 -2874 2046 -2868
rect 2040 -2880 2046 -2874
rect 2040 -2886 2046 -2880
rect 2040 -2892 2046 -2886
rect 2040 -2898 2046 -2892
rect 2040 -2904 2046 -2898
rect 2040 -2910 2046 -2904
rect 2040 -2916 2046 -2910
rect 2040 -2922 2046 -2916
rect 2040 -2928 2046 -2922
rect 2040 -2934 2046 -2928
rect 2040 -2940 2046 -2934
rect 2040 -2946 2046 -2940
rect 2040 -2952 2046 -2946
rect 2040 -2958 2046 -2952
rect 2040 -2964 2046 -2958
rect 2040 -2970 2046 -2964
rect 2040 -2976 2046 -2970
rect 2040 -2982 2046 -2976
rect 2040 -2988 2046 -2982
rect 2040 -2994 2046 -2988
rect 2040 -3000 2046 -2994
rect 2040 -3006 2046 -3000
rect 2040 -3012 2046 -3006
rect 2040 -3018 2046 -3012
rect 2040 -3024 2046 -3018
rect 2040 -3030 2046 -3024
rect 2040 -3036 2046 -3030
rect 2040 -3042 2046 -3036
rect 2040 -3048 2046 -3042
rect 2040 -3054 2046 -3048
rect 2040 -3060 2046 -3054
rect 2040 -3066 2046 -3060
rect 2040 -3072 2046 -3066
rect 2040 -3078 2046 -3072
rect 2040 -3084 2046 -3078
rect 2040 -3090 2046 -3084
rect 2040 -3144 2046 -3138
rect 2040 -3150 2046 -3144
rect 2040 -3156 2046 -3150
rect 2040 -3162 2046 -3156
rect 2040 -3168 2046 -3162
rect 2040 -3174 2046 -3168
rect 2040 -3180 2046 -3174
rect 2046 -390 2052 -384
rect 2046 -396 2052 -390
rect 2046 -402 2052 -396
rect 2046 -408 2052 -402
rect 2046 -414 2052 -408
rect 2046 -420 2052 -414
rect 2046 -426 2052 -420
rect 2046 -432 2052 -426
rect 2046 -438 2052 -432
rect 2046 -444 2052 -438
rect 2046 -450 2052 -444
rect 2046 -456 2052 -450
rect 2046 -462 2052 -456
rect 2046 -468 2052 -462
rect 2046 -474 2052 -468
rect 2046 -480 2052 -474
rect 2046 -486 2052 -480
rect 2046 -492 2052 -486
rect 2046 -498 2052 -492
rect 2046 -504 2052 -498
rect 2046 -510 2052 -504
rect 2046 -516 2052 -510
rect 2046 -522 2052 -516
rect 2046 -528 2052 -522
rect 2046 -534 2052 -528
rect 2046 -540 2052 -534
rect 2046 -546 2052 -540
rect 2046 -552 2052 -546
rect 2046 -558 2052 -552
rect 2046 -564 2052 -558
rect 2046 -570 2052 -564
rect 2046 -576 2052 -570
rect 2046 -582 2052 -576
rect 2046 -588 2052 -582
rect 2046 -594 2052 -588
rect 2046 -600 2052 -594
rect 2046 -606 2052 -600
rect 2046 -612 2052 -606
rect 2046 -618 2052 -612
rect 2046 -624 2052 -618
rect 2046 -630 2052 -624
rect 2046 -636 2052 -630
rect 2046 -642 2052 -636
rect 2046 -648 2052 -642
rect 2046 -654 2052 -648
rect 2046 -660 2052 -654
rect 2046 -666 2052 -660
rect 2046 -672 2052 -666
rect 2046 -678 2052 -672
rect 2046 -684 2052 -678
rect 2046 -690 2052 -684
rect 2046 -696 2052 -690
rect 2046 -702 2052 -696
rect 2046 -708 2052 -702
rect 2046 -714 2052 -708
rect 2046 -720 2052 -714
rect 2046 -726 2052 -720
rect 2046 -732 2052 -726
rect 2046 -738 2052 -732
rect 2046 -744 2052 -738
rect 2046 -750 2052 -744
rect 2046 -756 2052 -750
rect 2046 -762 2052 -756
rect 2046 -768 2052 -762
rect 2046 -774 2052 -768
rect 2046 -780 2052 -774
rect 2046 -786 2052 -780
rect 2046 -792 2052 -786
rect 2046 -798 2052 -792
rect 2046 -804 2052 -798
rect 2046 -810 2052 -804
rect 2046 -816 2052 -810
rect 2046 -822 2052 -816
rect 2046 -828 2052 -822
rect 2046 -834 2052 -828
rect 2046 -840 2052 -834
rect 2046 -846 2052 -840
rect 2046 -852 2052 -846
rect 2046 -858 2052 -852
rect 2046 -864 2052 -858
rect 2046 -870 2052 -864
rect 2046 -876 2052 -870
rect 2046 -882 2052 -876
rect 2046 -888 2052 -882
rect 2046 -894 2052 -888
rect 2046 -900 2052 -894
rect 2046 -906 2052 -900
rect 2046 -912 2052 -906
rect 2046 -918 2052 -912
rect 2046 -924 2052 -918
rect 2046 -930 2052 -924
rect 2046 -936 2052 -930
rect 2046 -942 2052 -936
rect 2046 -948 2052 -942
rect 2046 -954 2052 -948
rect 2046 -960 2052 -954
rect 2046 -966 2052 -960
rect 2046 -972 2052 -966
rect 2046 -978 2052 -972
rect 2046 -984 2052 -978
rect 2046 -990 2052 -984
rect 2046 -996 2052 -990
rect 2046 -1002 2052 -996
rect 2046 -1008 2052 -1002
rect 2046 -1014 2052 -1008
rect 2046 -1020 2052 -1014
rect 2046 -1026 2052 -1020
rect 2046 -1032 2052 -1026
rect 2046 -1038 2052 -1032
rect 2046 -1044 2052 -1038
rect 2046 -1050 2052 -1044
rect 2046 -1056 2052 -1050
rect 2046 -1062 2052 -1056
rect 2046 -1068 2052 -1062
rect 2046 -1074 2052 -1068
rect 2046 -1080 2052 -1074
rect 2046 -1086 2052 -1080
rect 2046 -1092 2052 -1086
rect 2046 -1098 2052 -1092
rect 2046 -1104 2052 -1098
rect 2046 -1110 2052 -1104
rect 2046 -1116 2052 -1110
rect 2046 -1122 2052 -1116
rect 2046 -1128 2052 -1122
rect 2046 -1134 2052 -1128
rect 2046 -1140 2052 -1134
rect 2046 -1146 2052 -1140
rect 2046 -1152 2052 -1146
rect 2046 -1158 2052 -1152
rect 2046 -1164 2052 -1158
rect 2046 -1170 2052 -1164
rect 2046 -1176 2052 -1170
rect 2046 -1182 2052 -1176
rect 2046 -1188 2052 -1182
rect 2046 -1194 2052 -1188
rect 2046 -1200 2052 -1194
rect 2046 -1206 2052 -1200
rect 2046 -1212 2052 -1206
rect 2046 -1218 2052 -1212
rect 2046 -1224 2052 -1218
rect 2046 -1230 2052 -1224
rect 2046 -1236 2052 -1230
rect 2046 -1242 2052 -1236
rect 2046 -1248 2052 -1242
rect 2046 -1254 2052 -1248
rect 2046 -1260 2052 -1254
rect 2046 -1266 2052 -1260
rect 2046 -1272 2052 -1266
rect 2046 -1278 2052 -1272
rect 2046 -1284 2052 -1278
rect 2046 -1290 2052 -1284
rect 2046 -1296 2052 -1290
rect 2046 -1302 2052 -1296
rect 2046 -1308 2052 -1302
rect 2046 -1314 2052 -1308
rect 2046 -1320 2052 -1314
rect 2046 -1326 2052 -1320
rect 2046 -1332 2052 -1326
rect 2046 -1338 2052 -1332
rect 2046 -1344 2052 -1338
rect 2046 -1350 2052 -1344
rect 2046 -1356 2052 -1350
rect 2046 -1362 2052 -1356
rect 2046 -1368 2052 -1362
rect 2046 -1374 2052 -1368
rect 2046 -1380 2052 -1374
rect 2046 -1386 2052 -1380
rect 2046 -1392 2052 -1386
rect 2046 -1398 2052 -1392
rect 2046 -1404 2052 -1398
rect 2046 -1410 2052 -1404
rect 2046 -1416 2052 -1410
rect 2046 -1422 2052 -1416
rect 2046 -1428 2052 -1422
rect 2046 -1434 2052 -1428
rect 2046 -1440 2052 -1434
rect 2046 -1446 2052 -1440
rect 2046 -1452 2052 -1446
rect 2046 -1458 2052 -1452
rect 2046 -1464 2052 -1458
rect 2046 -1470 2052 -1464
rect 2046 -1476 2052 -1470
rect 2046 -1482 2052 -1476
rect 2046 -1488 2052 -1482
rect 2046 -1494 2052 -1488
rect 2046 -1500 2052 -1494
rect 2046 -1506 2052 -1500
rect 2046 -1512 2052 -1506
rect 2046 -1518 2052 -1512
rect 2046 -1524 2052 -1518
rect 2046 -1530 2052 -1524
rect 2046 -1536 2052 -1530
rect 2046 -1542 2052 -1536
rect 2046 -1548 2052 -1542
rect 2046 -1554 2052 -1548
rect 2046 -1560 2052 -1554
rect 2046 -1566 2052 -1560
rect 2046 -1572 2052 -1566
rect 2046 -1578 2052 -1572
rect 2046 -1584 2052 -1578
rect 2046 -1590 2052 -1584
rect 2046 -1596 2052 -1590
rect 2046 -1692 2052 -1686
rect 2046 -1698 2052 -1692
rect 2046 -1704 2052 -1698
rect 2046 -1710 2052 -1704
rect 2046 -1716 2052 -1710
rect 2046 -1722 2052 -1716
rect 2046 -1728 2052 -1722
rect 2046 -1734 2052 -1728
rect 2046 -1740 2052 -1734
rect 2046 -1746 2052 -1740
rect 2046 -1752 2052 -1746
rect 2046 -1758 2052 -1752
rect 2046 -1764 2052 -1758
rect 2046 -1770 2052 -1764
rect 2046 -1776 2052 -1770
rect 2046 -1782 2052 -1776
rect 2046 -1788 2052 -1782
rect 2046 -1794 2052 -1788
rect 2046 -1800 2052 -1794
rect 2046 -1806 2052 -1800
rect 2046 -1812 2052 -1806
rect 2046 -1818 2052 -1812
rect 2046 -1824 2052 -1818
rect 2046 -1830 2052 -1824
rect 2046 -1836 2052 -1830
rect 2046 -1842 2052 -1836
rect 2046 -1848 2052 -1842
rect 2046 -1854 2052 -1848
rect 2046 -1860 2052 -1854
rect 2046 -1866 2052 -1860
rect 2046 -1872 2052 -1866
rect 2046 -1878 2052 -1872
rect 2046 -1884 2052 -1878
rect 2046 -1890 2052 -1884
rect 2046 -1896 2052 -1890
rect 2046 -1902 2052 -1896
rect 2046 -1908 2052 -1902
rect 2046 -1914 2052 -1908
rect 2046 -1920 2052 -1914
rect 2046 -1926 2052 -1920
rect 2046 -1932 2052 -1926
rect 2046 -1938 2052 -1932
rect 2046 -1944 2052 -1938
rect 2046 -1950 2052 -1944
rect 2046 -1956 2052 -1950
rect 2046 -1962 2052 -1956
rect 2046 -1968 2052 -1962
rect 2046 -1974 2052 -1968
rect 2046 -1980 2052 -1974
rect 2046 -1986 2052 -1980
rect 2046 -1992 2052 -1986
rect 2046 -1998 2052 -1992
rect 2046 -2004 2052 -1998
rect 2046 -2010 2052 -2004
rect 2046 -2016 2052 -2010
rect 2046 -2022 2052 -2016
rect 2046 -2028 2052 -2022
rect 2046 -2034 2052 -2028
rect 2046 -2040 2052 -2034
rect 2046 -2046 2052 -2040
rect 2046 -2052 2052 -2046
rect 2046 -2058 2052 -2052
rect 2046 -2064 2052 -2058
rect 2046 -2070 2052 -2064
rect 2046 -2076 2052 -2070
rect 2046 -2082 2052 -2076
rect 2046 -2088 2052 -2082
rect 2046 -2094 2052 -2088
rect 2046 -2100 2052 -2094
rect 2046 -2106 2052 -2100
rect 2046 -2112 2052 -2106
rect 2046 -2118 2052 -2112
rect 2046 -2124 2052 -2118
rect 2046 -2130 2052 -2124
rect 2046 -2136 2052 -2130
rect 2046 -2142 2052 -2136
rect 2046 -2148 2052 -2142
rect 2046 -2154 2052 -2148
rect 2046 -2160 2052 -2154
rect 2046 -2166 2052 -2160
rect 2046 -2172 2052 -2166
rect 2046 -2178 2052 -2172
rect 2046 -2184 2052 -2178
rect 2046 -2190 2052 -2184
rect 2046 -2196 2052 -2190
rect 2046 -2202 2052 -2196
rect 2046 -2208 2052 -2202
rect 2046 -2214 2052 -2208
rect 2046 -2220 2052 -2214
rect 2046 -2226 2052 -2220
rect 2046 -2232 2052 -2226
rect 2046 -2238 2052 -2232
rect 2046 -2244 2052 -2238
rect 2046 -2250 2052 -2244
rect 2046 -2256 2052 -2250
rect 2046 -2262 2052 -2256
rect 2046 -2268 2052 -2262
rect 2046 -2274 2052 -2268
rect 2046 -2280 2052 -2274
rect 2046 -2286 2052 -2280
rect 2046 -2292 2052 -2286
rect 2046 -2298 2052 -2292
rect 2046 -2304 2052 -2298
rect 2046 -2310 2052 -2304
rect 2046 -2316 2052 -2310
rect 2046 -2322 2052 -2316
rect 2046 -2328 2052 -2322
rect 2046 -2334 2052 -2328
rect 2046 -2340 2052 -2334
rect 2046 -2346 2052 -2340
rect 2046 -2352 2052 -2346
rect 2046 -2358 2052 -2352
rect 2046 -2364 2052 -2358
rect 2046 -2370 2052 -2364
rect 2046 -2376 2052 -2370
rect 2046 -2382 2052 -2376
rect 2046 -2388 2052 -2382
rect 2046 -2394 2052 -2388
rect 2046 -2400 2052 -2394
rect 2046 -2406 2052 -2400
rect 2046 -2412 2052 -2406
rect 2046 -2418 2052 -2412
rect 2046 -2424 2052 -2418
rect 2046 -2430 2052 -2424
rect 2046 -2436 2052 -2430
rect 2046 -2442 2052 -2436
rect 2046 -2448 2052 -2442
rect 2046 -2454 2052 -2448
rect 2046 -2460 2052 -2454
rect 2046 -2466 2052 -2460
rect 2046 -2472 2052 -2466
rect 2046 -2478 2052 -2472
rect 2046 -2484 2052 -2478
rect 2046 -2490 2052 -2484
rect 2046 -2496 2052 -2490
rect 2046 -2502 2052 -2496
rect 2046 -2592 2052 -2586
rect 2046 -2598 2052 -2592
rect 2046 -2604 2052 -2598
rect 2046 -2610 2052 -2604
rect 2046 -2616 2052 -2610
rect 2046 -2622 2052 -2616
rect 2046 -2628 2052 -2622
rect 2046 -2634 2052 -2628
rect 2046 -2640 2052 -2634
rect 2046 -2646 2052 -2640
rect 2046 -2652 2052 -2646
rect 2046 -2658 2052 -2652
rect 2046 -2664 2052 -2658
rect 2046 -2670 2052 -2664
rect 2046 -2676 2052 -2670
rect 2046 -2682 2052 -2676
rect 2046 -2688 2052 -2682
rect 2046 -2694 2052 -2688
rect 2046 -2700 2052 -2694
rect 2046 -2706 2052 -2700
rect 2046 -2712 2052 -2706
rect 2046 -2718 2052 -2712
rect 2046 -2724 2052 -2718
rect 2046 -2730 2052 -2724
rect 2046 -2736 2052 -2730
rect 2046 -2742 2052 -2736
rect 2046 -2748 2052 -2742
rect 2046 -2754 2052 -2748
rect 2046 -2760 2052 -2754
rect 2046 -2766 2052 -2760
rect 2046 -2772 2052 -2766
rect 2046 -2778 2052 -2772
rect 2046 -2784 2052 -2778
rect 2046 -2790 2052 -2784
rect 2046 -2796 2052 -2790
rect 2046 -2802 2052 -2796
rect 2046 -2808 2052 -2802
rect 2046 -2814 2052 -2808
rect 2046 -2820 2052 -2814
rect 2046 -2826 2052 -2820
rect 2046 -2832 2052 -2826
rect 2046 -2838 2052 -2832
rect 2046 -2844 2052 -2838
rect 2046 -2850 2052 -2844
rect 2046 -2856 2052 -2850
rect 2046 -2862 2052 -2856
rect 2046 -2868 2052 -2862
rect 2046 -2874 2052 -2868
rect 2046 -2880 2052 -2874
rect 2046 -2886 2052 -2880
rect 2046 -2892 2052 -2886
rect 2046 -2898 2052 -2892
rect 2046 -2904 2052 -2898
rect 2046 -2910 2052 -2904
rect 2046 -2916 2052 -2910
rect 2046 -2922 2052 -2916
rect 2046 -2928 2052 -2922
rect 2046 -2934 2052 -2928
rect 2046 -2940 2052 -2934
rect 2046 -2946 2052 -2940
rect 2046 -2952 2052 -2946
rect 2046 -2958 2052 -2952
rect 2046 -2964 2052 -2958
rect 2046 -2970 2052 -2964
rect 2046 -2976 2052 -2970
rect 2046 -2982 2052 -2976
rect 2046 -2988 2052 -2982
rect 2046 -2994 2052 -2988
rect 2046 -3000 2052 -2994
rect 2046 -3006 2052 -3000
rect 2046 -3012 2052 -3006
rect 2046 -3018 2052 -3012
rect 2046 -3024 2052 -3018
rect 2046 -3030 2052 -3024
rect 2046 -3036 2052 -3030
rect 2046 -3042 2052 -3036
rect 2046 -3048 2052 -3042
rect 2046 -3054 2052 -3048
rect 2046 -3060 2052 -3054
rect 2046 -3066 2052 -3060
rect 2046 -3072 2052 -3066
rect 2046 -3078 2052 -3072
rect 2046 -3084 2052 -3078
rect 2046 -3144 2052 -3138
rect 2046 -3150 2052 -3144
rect 2046 -3156 2052 -3150
rect 2046 -3162 2052 -3156
rect 2046 -3168 2052 -3162
rect 2046 -3174 2052 -3168
rect 2052 -384 2058 -378
rect 2052 -390 2058 -384
rect 2052 -396 2058 -390
rect 2052 -402 2058 -396
rect 2052 -408 2058 -402
rect 2052 -414 2058 -408
rect 2052 -420 2058 -414
rect 2052 -426 2058 -420
rect 2052 -432 2058 -426
rect 2052 -438 2058 -432
rect 2052 -444 2058 -438
rect 2052 -450 2058 -444
rect 2052 -456 2058 -450
rect 2052 -462 2058 -456
rect 2052 -468 2058 -462
rect 2052 -474 2058 -468
rect 2052 -480 2058 -474
rect 2052 -486 2058 -480
rect 2052 -492 2058 -486
rect 2052 -498 2058 -492
rect 2052 -504 2058 -498
rect 2052 -510 2058 -504
rect 2052 -516 2058 -510
rect 2052 -522 2058 -516
rect 2052 -528 2058 -522
rect 2052 -534 2058 -528
rect 2052 -540 2058 -534
rect 2052 -546 2058 -540
rect 2052 -552 2058 -546
rect 2052 -558 2058 -552
rect 2052 -564 2058 -558
rect 2052 -570 2058 -564
rect 2052 -576 2058 -570
rect 2052 -582 2058 -576
rect 2052 -588 2058 -582
rect 2052 -594 2058 -588
rect 2052 -600 2058 -594
rect 2052 -606 2058 -600
rect 2052 -612 2058 -606
rect 2052 -618 2058 -612
rect 2052 -624 2058 -618
rect 2052 -630 2058 -624
rect 2052 -636 2058 -630
rect 2052 -642 2058 -636
rect 2052 -648 2058 -642
rect 2052 -654 2058 -648
rect 2052 -660 2058 -654
rect 2052 -666 2058 -660
rect 2052 -672 2058 -666
rect 2052 -678 2058 -672
rect 2052 -684 2058 -678
rect 2052 -690 2058 -684
rect 2052 -696 2058 -690
rect 2052 -702 2058 -696
rect 2052 -708 2058 -702
rect 2052 -714 2058 -708
rect 2052 -720 2058 -714
rect 2052 -726 2058 -720
rect 2052 -732 2058 -726
rect 2052 -738 2058 -732
rect 2052 -744 2058 -738
rect 2052 -750 2058 -744
rect 2052 -756 2058 -750
rect 2052 -762 2058 -756
rect 2052 -768 2058 -762
rect 2052 -774 2058 -768
rect 2052 -780 2058 -774
rect 2052 -786 2058 -780
rect 2052 -792 2058 -786
rect 2052 -798 2058 -792
rect 2052 -804 2058 -798
rect 2052 -810 2058 -804
rect 2052 -816 2058 -810
rect 2052 -822 2058 -816
rect 2052 -828 2058 -822
rect 2052 -834 2058 -828
rect 2052 -840 2058 -834
rect 2052 -846 2058 -840
rect 2052 -852 2058 -846
rect 2052 -858 2058 -852
rect 2052 -864 2058 -858
rect 2052 -870 2058 -864
rect 2052 -876 2058 -870
rect 2052 -882 2058 -876
rect 2052 -888 2058 -882
rect 2052 -894 2058 -888
rect 2052 -900 2058 -894
rect 2052 -906 2058 -900
rect 2052 -912 2058 -906
rect 2052 -918 2058 -912
rect 2052 -924 2058 -918
rect 2052 -930 2058 -924
rect 2052 -936 2058 -930
rect 2052 -942 2058 -936
rect 2052 -948 2058 -942
rect 2052 -954 2058 -948
rect 2052 -960 2058 -954
rect 2052 -966 2058 -960
rect 2052 -972 2058 -966
rect 2052 -978 2058 -972
rect 2052 -984 2058 -978
rect 2052 -990 2058 -984
rect 2052 -996 2058 -990
rect 2052 -1002 2058 -996
rect 2052 -1008 2058 -1002
rect 2052 -1014 2058 -1008
rect 2052 -1020 2058 -1014
rect 2052 -1026 2058 -1020
rect 2052 -1032 2058 -1026
rect 2052 -1038 2058 -1032
rect 2052 -1044 2058 -1038
rect 2052 -1050 2058 -1044
rect 2052 -1056 2058 -1050
rect 2052 -1062 2058 -1056
rect 2052 -1068 2058 -1062
rect 2052 -1074 2058 -1068
rect 2052 -1080 2058 -1074
rect 2052 -1086 2058 -1080
rect 2052 -1092 2058 -1086
rect 2052 -1098 2058 -1092
rect 2052 -1104 2058 -1098
rect 2052 -1110 2058 -1104
rect 2052 -1116 2058 -1110
rect 2052 -1122 2058 -1116
rect 2052 -1128 2058 -1122
rect 2052 -1134 2058 -1128
rect 2052 -1140 2058 -1134
rect 2052 -1146 2058 -1140
rect 2052 -1152 2058 -1146
rect 2052 -1158 2058 -1152
rect 2052 -1164 2058 -1158
rect 2052 -1170 2058 -1164
rect 2052 -1176 2058 -1170
rect 2052 -1182 2058 -1176
rect 2052 -1188 2058 -1182
rect 2052 -1194 2058 -1188
rect 2052 -1200 2058 -1194
rect 2052 -1206 2058 -1200
rect 2052 -1212 2058 -1206
rect 2052 -1218 2058 -1212
rect 2052 -1224 2058 -1218
rect 2052 -1230 2058 -1224
rect 2052 -1236 2058 -1230
rect 2052 -1242 2058 -1236
rect 2052 -1248 2058 -1242
rect 2052 -1254 2058 -1248
rect 2052 -1260 2058 -1254
rect 2052 -1266 2058 -1260
rect 2052 -1272 2058 -1266
rect 2052 -1278 2058 -1272
rect 2052 -1284 2058 -1278
rect 2052 -1290 2058 -1284
rect 2052 -1296 2058 -1290
rect 2052 -1302 2058 -1296
rect 2052 -1308 2058 -1302
rect 2052 -1314 2058 -1308
rect 2052 -1320 2058 -1314
rect 2052 -1326 2058 -1320
rect 2052 -1332 2058 -1326
rect 2052 -1338 2058 -1332
rect 2052 -1344 2058 -1338
rect 2052 -1350 2058 -1344
rect 2052 -1356 2058 -1350
rect 2052 -1362 2058 -1356
rect 2052 -1368 2058 -1362
rect 2052 -1374 2058 -1368
rect 2052 -1380 2058 -1374
rect 2052 -1386 2058 -1380
rect 2052 -1392 2058 -1386
rect 2052 -1398 2058 -1392
rect 2052 -1404 2058 -1398
rect 2052 -1410 2058 -1404
rect 2052 -1416 2058 -1410
rect 2052 -1422 2058 -1416
rect 2052 -1428 2058 -1422
rect 2052 -1434 2058 -1428
rect 2052 -1440 2058 -1434
rect 2052 -1446 2058 -1440
rect 2052 -1452 2058 -1446
rect 2052 -1458 2058 -1452
rect 2052 -1464 2058 -1458
rect 2052 -1470 2058 -1464
rect 2052 -1476 2058 -1470
rect 2052 -1482 2058 -1476
rect 2052 -1488 2058 -1482
rect 2052 -1494 2058 -1488
rect 2052 -1500 2058 -1494
rect 2052 -1506 2058 -1500
rect 2052 -1512 2058 -1506
rect 2052 -1518 2058 -1512
rect 2052 -1524 2058 -1518
rect 2052 -1530 2058 -1524
rect 2052 -1536 2058 -1530
rect 2052 -1542 2058 -1536
rect 2052 -1548 2058 -1542
rect 2052 -1554 2058 -1548
rect 2052 -1560 2058 -1554
rect 2052 -1566 2058 -1560
rect 2052 -1572 2058 -1566
rect 2052 -1578 2058 -1572
rect 2052 -1584 2058 -1578
rect 2052 -1590 2058 -1584
rect 2052 -1686 2058 -1680
rect 2052 -1692 2058 -1686
rect 2052 -1698 2058 -1692
rect 2052 -1704 2058 -1698
rect 2052 -1710 2058 -1704
rect 2052 -1716 2058 -1710
rect 2052 -1722 2058 -1716
rect 2052 -1728 2058 -1722
rect 2052 -1734 2058 -1728
rect 2052 -1740 2058 -1734
rect 2052 -1746 2058 -1740
rect 2052 -1752 2058 -1746
rect 2052 -1758 2058 -1752
rect 2052 -1764 2058 -1758
rect 2052 -1770 2058 -1764
rect 2052 -1776 2058 -1770
rect 2052 -1782 2058 -1776
rect 2052 -1788 2058 -1782
rect 2052 -1794 2058 -1788
rect 2052 -1800 2058 -1794
rect 2052 -1806 2058 -1800
rect 2052 -1812 2058 -1806
rect 2052 -1818 2058 -1812
rect 2052 -1824 2058 -1818
rect 2052 -1830 2058 -1824
rect 2052 -1836 2058 -1830
rect 2052 -1842 2058 -1836
rect 2052 -1848 2058 -1842
rect 2052 -1854 2058 -1848
rect 2052 -1860 2058 -1854
rect 2052 -1866 2058 -1860
rect 2052 -1872 2058 -1866
rect 2052 -1878 2058 -1872
rect 2052 -1884 2058 -1878
rect 2052 -1890 2058 -1884
rect 2052 -1896 2058 -1890
rect 2052 -1902 2058 -1896
rect 2052 -1908 2058 -1902
rect 2052 -1914 2058 -1908
rect 2052 -1920 2058 -1914
rect 2052 -1926 2058 -1920
rect 2052 -1932 2058 -1926
rect 2052 -1938 2058 -1932
rect 2052 -1944 2058 -1938
rect 2052 -1950 2058 -1944
rect 2052 -1956 2058 -1950
rect 2052 -1962 2058 -1956
rect 2052 -1968 2058 -1962
rect 2052 -1974 2058 -1968
rect 2052 -1980 2058 -1974
rect 2052 -1986 2058 -1980
rect 2052 -1992 2058 -1986
rect 2052 -1998 2058 -1992
rect 2052 -2004 2058 -1998
rect 2052 -2010 2058 -2004
rect 2052 -2016 2058 -2010
rect 2052 -2022 2058 -2016
rect 2052 -2028 2058 -2022
rect 2052 -2034 2058 -2028
rect 2052 -2040 2058 -2034
rect 2052 -2046 2058 -2040
rect 2052 -2052 2058 -2046
rect 2052 -2058 2058 -2052
rect 2052 -2064 2058 -2058
rect 2052 -2070 2058 -2064
rect 2052 -2076 2058 -2070
rect 2052 -2082 2058 -2076
rect 2052 -2088 2058 -2082
rect 2052 -2094 2058 -2088
rect 2052 -2100 2058 -2094
rect 2052 -2106 2058 -2100
rect 2052 -2112 2058 -2106
rect 2052 -2118 2058 -2112
rect 2052 -2124 2058 -2118
rect 2052 -2130 2058 -2124
rect 2052 -2136 2058 -2130
rect 2052 -2142 2058 -2136
rect 2052 -2148 2058 -2142
rect 2052 -2154 2058 -2148
rect 2052 -2160 2058 -2154
rect 2052 -2166 2058 -2160
rect 2052 -2172 2058 -2166
rect 2052 -2178 2058 -2172
rect 2052 -2184 2058 -2178
rect 2052 -2190 2058 -2184
rect 2052 -2196 2058 -2190
rect 2052 -2202 2058 -2196
rect 2052 -2208 2058 -2202
rect 2052 -2214 2058 -2208
rect 2052 -2220 2058 -2214
rect 2052 -2226 2058 -2220
rect 2052 -2232 2058 -2226
rect 2052 -2238 2058 -2232
rect 2052 -2244 2058 -2238
rect 2052 -2250 2058 -2244
rect 2052 -2256 2058 -2250
rect 2052 -2262 2058 -2256
rect 2052 -2268 2058 -2262
rect 2052 -2274 2058 -2268
rect 2052 -2280 2058 -2274
rect 2052 -2286 2058 -2280
rect 2052 -2292 2058 -2286
rect 2052 -2298 2058 -2292
rect 2052 -2304 2058 -2298
rect 2052 -2310 2058 -2304
rect 2052 -2316 2058 -2310
rect 2052 -2322 2058 -2316
rect 2052 -2328 2058 -2322
rect 2052 -2334 2058 -2328
rect 2052 -2340 2058 -2334
rect 2052 -2346 2058 -2340
rect 2052 -2352 2058 -2346
rect 2052 -2358 2058 -2352
rect 2052 -2364 2058 -2358
rect 2052 -2370 2058 -2364
rect 2052 -2376 2058 -2370
rect 2052 -2382 2058 -2376
rect 2052 -2388 2058 -2382
rect 2052 -2394 2058 -2388
rect 2052 -2400 2058 -2394
rect 2052 -2406 2058 -2400
rect 2052 -2412 2058 -2406
rect 2052 -2418 2058 -2412
rect 2052 -2424 2058 -2418
rect 2052 -2430 2058 -2424
rect 2052 -2436 2058 -2430
rect 2052 -2442 2058 -2436
rect 2052 -2448 2058 -2442
rect 2052 -2454 2058 -2448
rect 2052 -2460 2058 -2454
rect 2052 -2466 2058 -2460
rect 2052 -2472 2058 -2466
rect 2052 -2478 2058 -2472
rect 2052 -2484 2058 -2478
rect 2052 -2490 2058 -2484
rect 2052 -2496 2058 -2490
rect 2052 -2502 2058 -2496
rect 2052 -2592 2058 -2586
rect 2052 -2598 2058 -2592
rect 2052 -2604 2058 -2598
rect 2052 -2610 2058 -2604
rect 2052 -2616 2058 -2610
rect 2052 -2622 2058 -2616
rect 2052 -2628 2058 -2622
rect 2052 -2634 2058 -2628
rect 2052 -2640 2058 -2634
rect 2052 -2646 2058 -2640
rect 2052 -2652 2058 -2646
rect 2052 -2658 2058 -2652
rect 2052 -2664 2058 -2658
rect 2052 -2670 2058 -2664
rect 2052 -2676 2058 -2670
rect 2052 -2682 2058 -2676
rect 2052 -2688 2058 -2682
rect 2052 -2694 2058 -2688
rect 2052 -2700 2058 -2694
rect 2052 -2706 2058 -2700
rect 2052 -2712 2058 -2706
rect 2052 -2718 2058 -2712
rect 2052 -2724 2058 -2718
rect 2052 -2730 2058 -2724
rect 2052 -2736 2058 -2730
rect 2052 -2742 2058 -2736
rect 2052 -2748 2058 -2742
rect 2052 -2754 2058 -2748
rect 2052 -2760 2058 -2754
rect 2052 -2766 2058 -2760
rect 2052 -2772 2058 -2766
rect 2052 -2778 2058 -2772
rect 2052 -2784 2058 -2778
rect 2052 -2790 2058 -2784
rect 2052 -2796 2058 -2790
rect 2052 -2802 2058 -2796
rect 2052 -2808 2058 -2802
rect 2052 -2814 2058 -2808
rect 2052 -2820 2058 -2814
rect 2052 -2826 2058 -2820
rect 2052 -2832 2058 -2826
rect 2052 -2838 2058 -2832
rect 2052 -2844 2058 -2838
rect 2052 -2850 2058 -2844
rect 2052 -2856 2058 -2850
rect 2052 -2862 2058 -2856
rect 2052 -2868 2058 -2862
rect 2052 -2874 2058 -2868
rect 2052 -2880 2058 -2874
rect 2052 -2886 2058 -2880
rect 2052 -2892 2058 -2886
rect 2052 -2898 2058 -2892
rect 2052 -2904 2058 -2898
rect 2052 -2910 2058 -2904
rect 2052 -2916 2058 -2910
rect 2052 -2922 2058 -2916
rect 2052 -2928 2058 -2922
rect 2052 -2934 2058 -2928
rect 2052 -2940 2058 -2934
rect 2052 -2946 2058 -2940
rect 2052 -2952 2058 -2946
rect 2052 -2958 2058 -2952
rect 2052 -2964 2058 -2958
rect 2052 -2970 2058 -2964
rect 2052 -2976 2058 -2970
rect 2052 -2982 2058 -2976
rect 2052 -2988 2058 -2982
rect 2052 -2994 2058 -2988
rect 2052 -3000 2058 -2994
rect 2052 -3006 2058 -3000
rect 2052 -3012 2058 -3006
rect 2052 -3018 2058 -3012
rect 2052 -3024 2058 -3018
rect 2052 -3030 2058 -3024
rect 2052 -3036 2058 -3030
rect 2052 -3042 2058 -3036
rect 2052 -3048 2058 -3042
rect 2052 -3054 2058 -3048
rect 2052 -3060 2058 -3054
rect 2052 -3066 2058 -3060
rect 2052 -3072 2058 -3066
rect 2052 -3078 2058 -3072
rect 2052 -3084 2058 -3078
rect 2052 -3138 2058 -3132
rect 2052 -3144 2058 -3138
rect 2052 -3150 2058 -3144
rect 2052 -3156 2058 -3150
rect 2052 -3162 2058 -3156
rect 2052 -3168 2058 -3162
rect 2058 -378 2064 -372
rect 2058 -384 2064 -378
rect 2058 -390 2064 -384
rect 2058 -396 2064 -390
rect 2058 -402 2064 -396
rect 2058 -408 2064 -402
rect 2058 -414 2064 -408
rect 2058 -420 2064 -414
rect 2058 -426 2064 -420
rect 2058 -432 2064 -426
rect 2058 -438 2064 -432
rect 2058 -444 2064 -438
rect 2058 -450 2064 -444
rect 2058 -456 2064 -450
rect 2058 -462 2064 -456
rect 2058 -468 2064 -462
rect 2058 -474 2064 -468
rect 2058 -480 2064 -474
rect 2058 -486 2064 -480
rect 2058 -492 2064 -486
rect 2058 -498 2064 -492
rect 2058 -504 2064 -498
rect 2058 -510 2064 -504
rect 2058 -516 2064 -510
rect 2058 -522 2064 -516
rect 2058 -528 2064 -522
rect 2058 -534 2064 -528
rect 2058 -540 2064 -534
rect 2058 -546 2064 -540
rect 2058 -552 2064 -546
rect 2058 -558 2064 -552
rect 2058 -564 2064 -558
rect 2058 -570 2064 -564
rect 2058 -576 2064 -570
rect 2058 -582 2064 -576
rect 2058 -588 2064 -582
rect 2058 -594 2064 -588
rect 2058 -600 2064 -594
rect 2058 -606 2064 -600
rect 2058 -612 2064 -606
rect 2058 -618 2064 -612
rect 2058 -624 2064 -618
rect 2058 -630 2064 -624
rect 2058 -636 2064 -630
rect 2058 -642 2064 -636
rect 2058 -648 2064 -642
rect 2058 -654 2064 -648
rect 2058 -660 2064 -654
rect 2058 -666 2064 -660
rect 2058 -672 2064 -666
rect 2058 -678 2064 -672
rect 2058 -684 2064 -678
rect 2058 -690 2064 -684
rect 2058 -696 2064 -690
rect 2058 -702 2064 -696
rect 2058 -708 2064 -702
rect 2058 -714 2064 -708
rect 2058 -720 2064 -714
rect 2058 -726 2064 -720
rect 2058 -732 2064 -726
rect 2058 -738 2064 -732
rect 2058 -744 2064 -738
rect 2058 -750 2064 -744
rect 2058 -756 2064 -750
rect 2058 -762 2064 -756
rect 2058 -768 2064 -762
rect 2058 -774 2064 -768
rect 2058 -780 2064 -774
rect 2058 -786 2064 -780
rect 2058 -792 2064 -786
rect 2058 -798 2064 -792
rect 2058 -804 2064 -798
rect 2058 -810 2064 -804
rect 2058 -816 2064 -810
rect 2058 -822 2064 -816
rect 2058 -828 2064 -822
rect 2058 -834 2064 -828
rect 2058 -840 2064 -834
rect 2058 -846 2064 -840
rect 2058 -852 2064 -846
rect 2058 -858 2064 -852
rect 2058 -864 2064 -858
rect 2058 -870 2064 -864
rect 2058 -876 2064 -870
rect 2058 -882 2064 -876
rect 2058 -888 2064 -882
rect 2058 -894 2064 -888
rect 2058 -900 2064 -894
rect 2058 -906 2064 -900
rect 2058 -912 2064 -906
rect 2058 -918 2064 -912
rect 2058 -924 2064 -918
rect 2058 -930 2064 -924
rect 2058 -936 2064 -930
rect 2058 -942 2064 -936
rect 2058 -948 2064 -942
rect 2058 -954 2064 -948
rect 2058 -960 2064 -954
rect 2058 -966 2064 -960
rect 2058 -972 2064 -966
rect 2058 -978 2064 -972
rect 2058 -984 2064 -978
rect 2058 -990 2064 -984
rect 2058 -996 2064 -990
rect 2058 -1002 2064 -996
rect 2058 -1008 2064 -1002
rect 2058 -1014 2064 -1008
rect 2058 -1020 2064 -1014
rect 2058 -1026 2064 -1020
rect 2058 -1032 2064 -1026
rect 2058 -1038 2064 -1032
rect 2058 -1044 2064 -1038
rect 2058 -1050 2064 -1044
rect 2058 -1056 2064 -1050
rect 2058 -1062 2064 -1056
rect 2058 -1068 2064 -1062
rect 2058 -1074 2064 -1068
rect 2058 -1080 2064 -1074
rect 2058 -1086 2064 -1080
rect 2058 -1092 2064 -1086
rect 2058 -1098 2064 -1092
rect 2058 -1104 2064 -1098
rect 2058 -1110 2064 -1104
rect 2058 -1116 2064 -1110
rect 2058 -1122 2064 -1116
rect 2058 -1128 2064 -1122
rect 2058 -1134 2064 -1128
rect 2058 -1140 2064 -1134
rect 2058 -1146 2064 -1140
rect 2058 -1152 2064 -1146
rect 2058 -1158 2064 -1152
rect 2058 -1164 2064 -1158
rect 2058 -1170 2064 -1164
rect 2058 -1176 2064 -1170
rect 2058 -1182 2064 -1176
rect 2058 -1188 2064 -1182
rect 2058 -1194 2064 -1188
rect 2058 -1200 2064 -1194
rect 2058 -1206 2064 -1200
rect 2058 -1212 2064 -1206
rect 2058 -1218 2064 -1212
rect 2058 -1224 2064 -1218
rect 2058 -1230 2064 -1224
rect 2058 -1236 2064 -1230
rect 2058 -1242 2064 -1236
rect 2058 -1248 2064 -1242
rect 2058 -1254 2064 -1248
rect 2058 -1260 2064 -1254
rect 2058 -1266 2064 -1260
rect 2058 -1272 2064 -1266
rect 2058 -1278 2064 -1272
rect 2058 -1284 2064 -1278
rect 2058 -1290 2064 -1284
rect 2058 -1296 2064 -1290
rect 2058 -1302 2064 -1296
rect 2058 -1308 2064 -1302
rect 2058 -1314 2064 -1308
rect 2058 -1320 2064 -1314
rect 2058 -1326 2064 -1320
rect 2058 -1332 2064 -1326
rect 2058 -1338 2064 -1332
rect 2058 -1344 2064 -1338
rect 2058 -1350 2064 -1344
rect 2058 -1356 2064 -1350
rect 2058 -1362 2064 -1356
rect 2058 -1368 2064 -1362
rect 2058 -1374 2064 -1368
rect 2058 -1380 2064 -1374
rect 2058 -1386 2064 -1380
rect 2058 -1392 2064 -1386
rect 2058 -1398 2064 -1392
rect 2058 -1404 2064 -1398
rect 2058 -1410 2064 -1404
rect 2058 -1416 2064 -1410
rect 2058 -1422 2064 -1416
rect 2058 -1428 2064 -1422
rect 2058 -1434 2064 -1428
rect 2058 -1440 2064 -1434
rect 2058 -1446 2064 -1440
rect 2058 -1452 2064 -1446
rect 2058 -1458 2064 -1452
rect 2058 -1464 2064 -1458
rect 2058 -1470 2064 -1464
rect 2058 -1476 2064 -1470
rect 2058 -1482 2064 -1476
rect 2058 -1488 2064 -1482
rect 2058 -1494 2064 -1488
rect 2058 -1500 2064 -1494
rect 2058 -1506 2064 -1500
rect 2058 -1512 2064 -1506
rect 2058 -1518 2064 -1512
rect 2058 -1524 2064 -1518
rect 2058 -1530 2064 -1524
rect 2058 -1536 2064 -1530
rect 2058 -1542 2064 -1536
rect 2058 -1548 2064 -1542
rect 2058 -1554 2064 -1548
rect 2058 -1560 2064 -1554
rect 2058 -1566 2064 -1560
rect 2058 -1572 2064 -1566
rect 2058 -1578 2064 -1572
rect 2058 -1680 2064 -1674
rect 2058 -1686 2064 -1680
rect 2058 -1692 2064 -1686
rect 2058 -1698 2064 -1692
rect 2058 -1704 2064 -1698
rect 2058 -1710 2064 -1704
rect 2058 -1716 2064 -1710
rect 2058 -1722 2064 -1716
rect 2058 -1728 2064 -1722
rect 2058 -1734 2064 -1728
rect 2058 -1740 2064 -1734
rect 2058 -1746 2064 -1740
rect 2058 -1752 2064 -1746
rect 2058 -1758 2064 -1752
rect 2058 -1764 2064 -1758
rect 2058 -1770 2064 -1764
rect 2058 -1776 2064 -1770
rect 2058 -1782 2064 -1776
rect 2058 -1788 2064 -1782
rect 2058 -1794 2064 -1788
rect 2058 -1800 2064 -1794
rect 2058 -1806 2064 -1800
rect 2058 -1812 2064 -1806
rect 2058 -1818 2064 -1812
rect 2058 -1824 2064 -1818
rect 2058 -1830 2064 -1824
rect 2058 -1836 2064 -1830
rect 2058 -1842 2064 -1836
rect 2058 -1848 2064 -1842
rect 2058 -1854 2064 -1848
rect 2058 -1860 2064 -1854
rect 2058 -1866 2064 -1860
rect 2058 -1872 2064 -1866
rect 2058 -1878 2064 -1872
rect 2058 -1884 2064 -1878
rect 2058 -1890 2064 -1884
rect 2058 -1896 2064 -1890
rect 2058 -1902 2064 -1896
rect 2058 -1908 2064 -1902
rect 2058 -1914 2064 -1908
rect 2058 -1920 2064 -1914
rect 2058 -1926 2064 -1920
rect 2058 -1932 2064 -1926
rect 2058 -1938 2064 -1932
rect 2058 -1944 2064 -1938
rect 2058 -1950 2064 -1944
rect 2058 -1956 2064 -1950
rect 2058 -1962 2064 -1956
rect 2058 -1968 2064 -1962
rect 2058 -1974 2064 -1968
rect 2058 -1980 2064 -1974
rect 2058 -1986 2064 -1980
rect 2058 -1992 2064 -1986
rect 2058 -1998 2064 -1992
rect 2058 -2004 2064 -1998
rect 2058 -2010 2064 -2004
rect 2058 -2016 2064 -2010
rect 2058 -2022 2064 -2016
rect 2058 -2028 2064 -2022
rect 2058 -2034 2064 -2028
rect 2058 -2040 2064 -2034
rect 2058 -2046 2064 -2040
rect 2058 -2052 2064 -2046
rect 2058 -2058 2064 -2052
rect 2058 -2064 2064 -2058
rect 2058 -2070 2064 -2064
rect 2058 -2076 2064 -2070
rect 2058 -2082 2064 -2076
rect 2058 -2088 2064 -2082
rect 2058 -2094 2064 -2088
rect 2058 -2100 2064 -2094
rect 2058 -2106 2064 -2100
rect 2058 -2112 2064 -2106
rect 2058 -2118 2064 -2112
rect 2058 -2124 2064 -2118
rect 2058 -2130 2064 -2124
rect 2058 -2136 2064 -2130
rect 2058 -2142 2064 -2136
rect 2058 -2148 2064 -2142
rect 2058 -2154 2064 -2148
rect 2058 -2160 2064 -2154
rect 2058 -2166 2064 -2160
rect 2058 -2172 2064 -2166
rect 2058 -2178 2064 -2172
rect 2058 -2184 2064 -2178
rect 2058 -2190 2064 -2184
rect 2058 -2196 2064 -2190
rect 2058 -2202 2064 -2196
rect 2058 -2208 2064 -2202
rect 2058 -2214 2064 -2208
rect 2058 -2220 2064 -2214
rect 2058 -2226 2064 -2220
rect 2058 -2232 2064 -2226
rect 2058 -2238 2064 -2232
rect 2058 -2244 2064 -2238
rect 2058 -2250 2064 -2244
rect 2058 -2256 2064 -2250
rect 2058 -2262 2064 -2256
rect 2058 -2268 2064 -2262
rect 2058 -2274 2064 -2268
rect 2058 -2280 2064 -2274
rect 2058 -2286 2064 -2280
rect 2058 -2292 2064 -2286
rect 2058 -2298 2064 -2292
rect 2058 -2304 2064 -2298
rect 2058 -2310 2064 -2304
rect 2058 -2316 2064 -2310
rect 2058 -2322 2064 -2316
rect 2058 -2328 2064 -2322
rect 2058 -2334 2064 -2328
rect 2058 -2340 2064 -2334
rect 2058 -2346 2064 -2340
rect 2058 -2352 2064 -2346
rect 2058 -2358 2064 -2352
rect 2058 -2364 2064 -2358
rect 2058 -2370 2064 -2364
rect 2058 -2376 2064 -2370
rect 2058 -2382 2064 -2376
rect 2058 -2388 2064 -2382
rect 2058 -2394 2064 -2388
rect 2058 -2400 2064 -2394
rect 2058 -2406 2064 -2400
rect 2058 -2412 2064 -2406
rect 2058 -2418 2064 -2412
rect 2058 -2424 2064 -2418
rect 2058 -2430 2064 -2424
rect 2058 -2436 2064 -2430
rect 2058 -2442 2064 -2436
rect 2058 -2448 2064 -2442
rect 2058 -2454 2064 -2448
rect 2058 -2460 2064 -2454
rect 2058 -2466 2064 -2460
rect 2058 -2472 2064 -2466
rect 2058 -2478 2064 -2472
rect 2058 -2484 2064 -2478
rect 2058 -2490 2064 -2484
rect 2058 -2496 2064 -2490
rect 2058 -2586 2064 -2580
rect 2058 -2592 2064 -2586
rect 2058 -2598 2064 -2592
rect 2058 -2604 2064 -2598
rect 2058 -2610 2064 -2604
rect 2058 -2616 2064 -2610
rect 2058 -2622 2064 -2616
rect 2058 -2628 2064 -2622
rect 2058 -2634 2064 -2628
rect 2058 -2640 2064 -2634
rect 2058 -2646 2064 -2640
rect 2058 -2652 2064 -2646
rect 2058 -2658 2064 -2652
rect 2058 -2664 2064 -2658
rect 2058 -2670 2064 -2664
rect 2058 -2676 2064 -2670
rect 2058 -2682 2064 -2676
rect 2058 -2688 2064 -2682
rect 2058 -2694 2064 -2688
rect 2058 -2700 2064 -2694
rect 2058 -2706 2064 -2700
rect 2058 -2712 2064 -2706
rect 2058 -2718 2064 -2712
rect 2058 -2724 2064 -2718
rect 2058 -2730 2064 -2724
rect 2058 -2736 2064 -2730
rect 2058 -2742 2064 -2736
rect 2058 -2748 2064 -2742
rect 2058 -2754 2064 -2748
rect 2058 -2760 2064 -2754
rect 2058 -2766 2064 -2760
rect 2058 -2772 2064 -2766
rect 2058 -2778 2064 -2772
rect 2058 -2784 2064 -2778
rect 2058 -2790 2064 -2784
rect 2058 -2796 2064 -2790
rect 2058 -2802 2064 -2796
rect 2058 -2808 2064 -2802
rect 2058 -2814 2064 -2808
rect 2058 -2820 2064 -2814
rect 2058 -2826 2064 -2820
rect 2058 -2832 2064 -2826
rect 2058 -2838 2064 -2832
rect 2058 -2844 2064 -2838
rect 2058 -2850 2064 -2844
rect 2058 -2856 2064 -2850
rect 2058 -2862 2064 -2856
rect 2058 -2868 2064 -2862
rect 2058 -2874 2064 -2868
rect 2058 -2880 2064 -2874
rect 2058 -2886 2064 -2880
rect 2058 -2892 2064 -2886
rect 2058 -2898 2064 -2892
rect 2058 -2904 2064 -2898
rect 2058 -2910 2064 -2904
rect 2058 -2916 2064 -2910
rect 2058 -2922 2064 -2916
rect 2058 -2928 2064 -2922
rect 2058 -2934 2064 -2928
rect 2058 -2940 2064 -2934
rect 2058 -2946 2064 -2940
rect 2058 -2952 2064 -2946
rect 2058 -2958 2064 -2952
rect 2058 -2964 2064 -2958
rect 2058 -2970 2064 -2964
rect 2058 -2976 2064 -2970
rect 2058 -2982 2064 -2976
rect 2058 -2988 2064 -2982
rect 2058 -2994 2064 -2988
rect 2058 -3000 2064 -2994
rect 2058 -3006 2064 -3000
rect 2058 -3012 2064 -3006
rect 2058 -3018 2064 -3012
rect 2058 -3024 2064 -3018
rect 2058 -3030 2064 -3024
rect 2058 -3036 2064 -3030
rect 2058 -3042 2064 -3036
rect 2058 -3048 2064 -3042
rect 2058 -3054 2064 -3048
rect 2058 -3060 2064 -3054
rect 2058 -3066 2064 -3060
rect 2058 -3072 2064 -3066
rect 2058 -3078 2064 -3072
rect 2058 -3084 2064 -3078
rect 2058 -3138 2064 -3132
rect 2058 -3144 2064 -3138
rect 2058 -3150 2064 -3144
rect 2058 -3156 2064 -3150
rect 2058 -3162 2064 -3156
rect 2058 -3168 2064 -3162
rect 2064 -366 2070 -360
rect 2064 -372 2070 -366
rect 2064 -378 2070 -372
rect 2064 -384 2070 -378
rect 2064 -390 2070 -384
rect 2064 -396 2070 -390
rect 2064 -402 2070 -396
rect 2064 -408 2070 -402
rect 2064 -414 2070 -408
rect 2064 -420 2070 -414
rect 2064 -426 2070 -420
rect 2064 -432 2070 -426
rect 2064 -438 2070 -432
rect 2064 -444 2070 -438
rect 2064 -450 2070 -444
rect 2064 -456 2070 -450
rect 2064 -462 2070 -456
rect 2064 -468 2070 -462
rect 2064 -474 2070 -468
rect 2064 -480 2070 -474
rect 2064 -486 2070 -480
rect 2064 -492 2070 -486
rect 2064 -498 2070 -492
rect 2064 -504 2070 -498
rect 2064 -510 2070 -504
rect 2064 -516 2070 -510
rect 2064 -522 2070 -516
rect 2064 -528 2070 -522
rect 2064 -534 2070 -528
rect 2064 -540 2070 -534
rect 2064 -546 2070 -540
rect 2064 -552 2070 -546
rect 2064 -558 2070 -552
rect 2064 -564 2070 -558
rect 2064 -570 2070 -564
rect 2064 -576 2070 -570
rect 2064 -582 2070 -576
rect 2064 -588 2070 -582
rect 2064 -594 2070 -588
rect 2064 -600 2070 -594
rect 2064 -606 2070 -600
rect 2064 -612 2070 -606
rect 2064 -618 2070 -612
rect 2064 -624 2070 -618
rect 2064 -630 2070 -624
rect 2064 -636 2070 -630
rect 2064 -642 2070 -636
rect 2064 -648 2070 -642
rect 2064 -654 2070 -648
rect 2064 -660 2070 -654
rect 2064 -666 2070 -660
rect 2064 -672 2070 -666
rect 2064 -678 2070 -672
rect 2064 -684 2070 -678
rect 2064 -690 2070 -684
rect 2064 -696 2070 -690
rect 2064 -702 2070 -696
rect 2064 -708 2070 -702
rect 2064 -714 2070 -708
rect 2064 -720 2070 -714
rect 2064 -726 2070 -720
rect 2064 -732 2070 -726
rect 2064 -738 2070 -732
rect 2064 -744 2070 -738
rect 2064 -750 2070 -744
rect 2064 -756 2070 -750
rect 2064 -762 2070 -756
rect 2064 -768 2070 -762
rect 2064 -774 2070 -768
rect 2064 -780 2070 -774
rect 2064 -786 2070 -780
rect 2064 -792 2070 -786
rect 2064 -798 2070 -792
rect 2064 -804 2070 -798
rect 2064 -810 2070 -804
rect 2064 -816 2070 -810
rect 2064 -822 2070 -816
rect 2064 -828 2070 -822
rect 2064 -834 2070 -828
rect 2064 -840 2070 -834
rect 2064 -846 2070 -840
rect 2064 -852 2070 -846
rect 2064 -858 2070 -852
rect 2064 -864 2070 -858
rect 2064 -870 2070 -864
rect 2064 -876 2070 -870
rect 2064 -882 2070 -876
rect 2064 -888 2070 -882
rect 2064 -894 2070 -888
rect 2064 -900 2070 -894
rect 2064 -906 2070 -900
rect 2064 -912 2070 -906
rect 2064 -918 2070 -912
rect 2064 -924 2070 -918
rect 2064 -930 2070 -924
rect 2064 -936 2070 -930
rect 2064 -942 2070 -936
rect 2064 -948 2070 -942
rect 2064 -954 2070 -948
rect 2064 -960 2070 -954
rect 2064 -966 2070 -960
rect 2064 -972 2070 -966
rect 2064 -978 2070 -972
rect 2064 -984 2070 -978
rect 2064 -990 2070 -984
rect 2064 -996 2070 -990
rect 2064 -1002 2070 -996
rect 2064 -1008 2070 -1002
rect 2064 -1014 2070 -1008
rect 2064 -1020 2070 -1014
rect 2064 -1026 2070 -1020
rect 2064 -1032 2070 -1026
rect 2064 -1038 2070 -1032
rect 2064 -1044 2070 -1038
rect 2064 -1050 2070 -1044
rect 2064 -1056 2070 -1050
rect 2064 -1062 2070 -1056
rect 2064 -1068 2070 -1062
rect 2064 -1074 2070 -1068
rect 2064 -1080 2070 -1074
rect 2064 -1086 2070 -1080
rect 2064 -1092 2070 -1086
rect 2064 -1098 2070 -1092
rect 2064 -1104 2070 -1098
rect 2064 -1110 2070 -1104
rect 2064 -1116 2070 -1110
rect 2064 -1122 2070 -1116
rect 2064 -1128 2070 -1122
rect 2064 -1134 2070 -1128
rect 2064 -1140 2070 -1134
rect 2064 -1146 2070 -1140
rect 2064 -1152 2070 -1146
rect 2064 -1158 2070 -1152
rect 2064 -1164 2070 -1158
rect 2064 -1170 2070 -1164
rect 2064 -1176 2070 -1170
rect 2064 -1182 2070 -1176
rect 2064 -1188 2070 -1182
rect 2064 -1194 2070 -1188
rect 2064 -1200 2070 -1194
rect 2064 -1206 2070 -1200
rect 2064 -1212 2070 -1206
rect 2064 -1218 2070 -1212
rect 2064 -1224 2070 -1218
rect 2064 -1230 2070 -1224
rect 2064 -1236 2070 -1230
rect 2064 -1242 2070 -1236
rect 2064 -1248 2070 -1242
rect 2064 -1254 2070 -1248
rect 2064 -1260 2070 -1254
rect 2064 -1266 2070 -1260
rect 2064 -1272 2070 -1266
rect 2064 -1278 2070 -1272
rect 2064 -1284 2070 -1278
rect 2064 -1290 2070 -1284
rect 2064 -1296 2070 -1290
rect 2064 -1302 2070 -1296
rect 2064 -1308 2070 -1302
rect 2064 -1314 2070 -1308
rect 2064 -1320 2070 -1314
rect 2064 -1326 2070 -1320
rect 2064 -1332 2070 -1326
rect 2064 -1338 2070 -1332
rect 2064 -1344 2070 -1338
rect 2064 -1350 2070 -1344
rect 2064 -1356 2070 -1350
rect 2064 -1362 2070 -1356
rect 2064 -1368 2070 -1362
rect 2064 -1374 2070 -1368
rect 2064 -1380 2070 -1374
rect 2064 -1386 2070 -1380
rect 2064 -1392 2070 -1386
rect 2064 -1398 2070 -1392
rect 2064 -1404 2070 -1398
rect 2064 -1410 2070 -1404
rect 2064 -1416 2070 -1410
rect 2064 -1422 2070 -1416
rect 2064 -1428 2070 -1422
rect 2064 -1434 2070 -1428
rect 2064 -1440 2070 -1434
rect 2064 -1446 2070 -1440
rect 2064 -1452 2070 -1446
rect 2064 -1458 2070 -1452
rect 2064 -1464 2070 -1458
rect 2064 -1470 2070 -1464
rect 2064 -1476 2070 -1470
rect 2064 -1482 2070 -1476
rect 2064 -1488 2070 -1482
rect 2064 -1494 2070 -1488
rect 2064 -1500 2070 -1494
rect 2064 -1506 2070 -1500
rect 2064 -1512 2070 -1506
rect 2064 -1518 2070 -1512
rect 2064 -1524 2070 -1518
rect 2064 -1530 2070 -1524
rect 2064 -1536 2070 -1530
rect 2064 -1542 2070 -1536
rect 2064 -1548 2070 -1542
rect 2064 -1554 2070 -1548
rect 2064 -1560 2070 -1554
rect 2064 -1566 2070 -1560
rect 2064 -1674 2070 -1668
rect 2064 -1680 2070 -1674
rect 2064 -1686 2070 -1680
rect 2064 -1692 2070 -1686
rect 2064 -1698 2070 -1692
rect 2064 -1704 2070 -1698
rect 2064 -1710 2070 -1704
rect 2064 -1716 2070 -1710
rect 2064 -1722 2070 -1716
rect 2064 -1728 2070 -1722
rect 2064 -1734 2070 -1728
rect 2064 -1740 2070 -1734
rect 2064 -1746 2070 -1740
rect 2064 -1752 2070 -1746
rect 2064 -1758 2070 -1752
rect 2064 -1764 2070 -1758
rect 2064 -1770 2070 -1764
rect 2064 -1776 2070 -1770
rect 2064 -1782 2070 -1776
rect 2064 -1788 2070 -1782
rect 2064 -1794 2070 -1788
rect 2064 -1800 2070 -1794
rect 2064 -1806 2070 -1800
rect 2064 -1812 2070 -1806
rect 2064 -1818 2070 -1812
rect 2064 -1824 2070 -1818
rect 2064 -1830 2070 -1824
rect 2064 -1836 2070 -1830
rect 2064 -1842 2070 -1836
rect 2064 -1848 2070 -1842
rect 2064 -1854 2070 -1848
rect 2064 -1860 2070 -1854
rect 2064 -1866 2070 -1860
rect 2064 -1872 2070 -1866
rect 2064 -1878 2070 -1872
rect 2064 -1884 2070 -1878
rect 2064 -1890 2070 -1884
rect 2064 -1896 2070 -1890
rect 2064 -1902 2070 -1896
rect 2064 -1908 2070 -1902
rect 2064 -1914 2070 -1908
rect 2064 -1920 2070 -1914
rect 2064 -1926 2070 -1920
rect 2064 -1932 2070 -1926
rect 2064 -1938 2070 -1932
rect 2064 -1944 2070 -1938
rect 2064 -1950 2070 -1944
rect 2064 -1956 2070 -1950
rect 2064 -1962 2070 -1956
rect 2064 -1968 2070 -1962
rect 2064 -1974 2070 -1968
rect 2064 -1980 2070 -1974
rect 2064 -1986 2070 -1980
rect 2064 -1992 2070 -1986
rect 2064 -1998 2070 -1992
rect 2064 -2004 2070 -1998
rect 2064 -2010 2070 -2004
rect 2064 -2016 2070 -2010
rect 2064 -2022 2070 -2016
rect 2064 -2028 2070 -2022
rect 2064 -2034 2070 -2028
rect 2064 -2040 2070 -2034
rect 2064 -2046 2070 -2040
rect 2064 -2052 2070 -2046
rect 2064 -2058 2070 -2052
rect 2064 -2064 2070 -2058
rect 2064 -2070 2070 -2064
rect 2064 -2076 2070 -2070
rect 2064 -2082 2070 -2076
rect 2064 -2088 2070 -2082
rect 2064 -2094 2070 -2088
rect 2064 -2100 2070 -2094
rect 2064 -2106 2070 -2100
rect 2064 -2112 2070 -2106
rect 2064 -2118 2070 -2112
rect 2064 -2124 2070 -2118
rect 2064 -2130 2070 -2124
rect 2064 -2136 2070 -2130
rect 2064 -2142 2070 -2136
rect 2064 -2148 2070 -2142
rect 2064 -2154 2070 -2148
rect 2064 -2160 2070 -2154
rect 2064 -2166 2070 -2160
rect 2064 -2172 2070 -2166
rect 2064 -2178 2070 -2172
rect 2064 -2184 2070 -2178
rect 2064 -2190 2070 -2184
rect 2064 -2196 2070 -2190
rect 2064 -2202 2070 -2196
rect 2064 -2208 2070 -2202
rect 2064 -2214 2070 -2208
rect 2064 -2220 2070 -2214
rect 2064 -2226 2070 -2220
rect 2064 -2232 2070 -2226
rect 2064 -2238 2070 -2232
rect 2064 -2244 2070 -2238
rect 2064 -2250 2070 -2244
rect 2064 -2256 2070 -2250
rect 2064 -2262 2070 -2256
rect 2064 -2268 2070 -2262
rect 2064 -2274 2070 -2268
rect 2064 -2280 2070 -2274
rect 2064 -2286 2070 -2280
rect 2064 -2292 2070 -2286
rect 2064 -2298 2070 -2292
rect 2064 -2304 2070 -2298
rect 2064 -2310 2070 -2304
rect 2064 -2316 2070 -2310
rect 2064 -2322 2070 -2316
rect 2064 -2328 2070 -2322
rect 2064 -2334 2070 -2328
rect 2064 -2340 2070 -2334
rect 2064 -2346 2070 -2340
rect 2064 -2352 2070 -2346
rect 2064 -2358 2070 -2352
rect 2064 -2364 2070 -2358
rect 2064 -2370 2070 -2364
rect 2064 -2376 2070 -2370
rect 2064 -2382 2070 -2376
rect 2064 -2388 2070 -2382
rect 2064 -2394 2070 -2388
rect 2064 -2400 2070 -2394
rect 2064 -2406 2070 -2400
rect 2064 -2412 2070 -2406
rect 2064 -2418 2070 -2412
rect 2064 -2424 2070 -2418
rect 2064 -2430 2070 -2424
rect 2064 -2436 2070 -2430
rect 2064 -2442 2070 -2436
rect 2064 -2448 2070 -2442
rect 2064 -2454 2070 -2448
rect 2064 -2460 2070 -2454
rect 2064 -2466 2070 -2460
rect 2064 -2472 2070 -2466
rect 2064 -2478 2070 -2472
rect 2064 -2484 2070 -2478
rect 2064 -2490 2070 -2484
rect 2064 -2496 2070 -2490
rect 2064 -2586 2070 -2580
rect 2064 -2592 2070 -2586
rect 2064 -2598 2070 -2592
rect 2064 -2604 2070 -2598
rect 2064 -2610 2070 -2604
rect 2064 -2616 2070 -2610
rect 2064 -2622 2070 -2616
rect 2064 -2628 2070 -2622
rect 2064 -2634 2070 -2628
rect 2064 -2640 2070 -2634
rect 2064 -2646 2070 -2640
rect 2064 -2652 2070 -2646
rect 2064 -2658 2070 -2652
rect 2064 -2664 2070 -2658
rect 2064 -2670 2070 -2664
rect 2064 -2676 2070 -2670
rect 2064 -2682 2070 -2676
rect 2064 -2688 2070 -2682
rect 2064 -2694 2070 -2688
rect 2064 -2700 2070 -2694
rect 2064 -2706 2070 -2700
rect 2064 -2712 2070 -2706
rect 2064 -2718 2070 -2712
rect 2064 -2724 2070 -2718
rect 2064 -2730 2070 -2724
rect 2064 -2736 2070 -2730
rect 2064 -2742 2070 -2736
rect 2064 -2748 2070 -2742
rect 2064 -2754 2070 -2748
rect 2064 -2760 2070 -2754
rect 2064 -2766 2070 -2760
rect 2064 -2772 2070 -2766
rect 2064 -2778 2070 -2772
rect 2064 -2784 2070 -2778
rect 2064 -2790 2070 -2784
rect 2064 -2796 2070 -2790
rect 2064 -2802 2070 -2796
rect 2064 -2808 2070 -2802
rect 2064 -2814 2070 -2808
rect 2064 -2820 2070 -2814
rect 2064 -2826 2070 -2820
rect 2064 -2832 2070 -2826
rect 2064 -2838 2070 -2832
rect 2064 -2844 2070 -2838
rect 2064 -2850 2070 -2844
rect 2064 -2856 2070 -2850
rect 2064 -2862 2070 -2856
rect 2064 -2868 2070 -2862
rect 2064 -2874 2070 -2868
rect 2064 -2880 2070 -2874
rect 2064 -2886 2070 -2880
rect 2064 -2892 2070 -2886
rect 2064 -2898 2070 -2892
rect 2064 -2904 2070 -2898
rect 2064 -2910 2070 -2904
rect 2064 -2916 2070 -2910
rect 2064 -2922 2070 -2916
rect 2064 -2928 2070 -2922
rect 2064 -2934 2070 -2928
rect 2064 -2940 2070 -2934
rect 2064 -2946 2070 -2940
rect 2064 -2952 2070 -2946
rect 2064 -2958 2070 -2952
rect 2064 -2964 2070 -2958
rect 2064 -2970 2070 -2964
rect 2064 -2976 2070 -2970
rect 2064 -2982 2070 -2976
rect 2064 -2988 2070 -2982
rect 2064 -2994 2070 -2988
rect 2064 -3000 2070 -2994
rect 2064 -3006 2070 -3000
rect 2064 -3012 2070 -3006
rect 2064 -3018 2070 -3012
rect 2064 -3024 2070 -3018
rect 2064 -3030 2070 -3024
rect 2064 -3036 2070 -3030
rect 2064 -3042 2070 -3036
rect 2064 -3048 2070 -3042
rect 2064 -3054 2070 -3048
rect 2064 -3060 2070 -3054
rect 2064 -3066 2070 -3060
rect 2064 -3072 2070 -3066
rect 2064 -3078 2070 -3072
rect 2064 -3138 2070 -3132
rect 2064 -3144 2070 -3138
rect 2064 -3150 2070 -3144
rect 2064 -3156 2070 -3150
rect 2064 -3162 2070 -3156
rect 2070 -360 2076 -354
rect 2070 -366 2076 -360
rect 2070 -372 2076 -366
rect 2070 -378 2076 -372
rect 2070 -384 2076 -378
rect 2070 -390 2076 -384
rect 2070 -396 2076 -390
rect 2070 -402 2076 -396
rect 2070 -408 2076 -402
rect 2070 -414 2076 -408
rect 2070 -420 2076 -414
rect 2070 -426 2076 -420
rect 2070 -432 2076 -426
rect 2070 -438 2076 -432
rect 2070 -444 2076 -438
rect 2070 -450 2076 -444
rect 2070 -456 2076 -450
rect 2070 -462 2076 -456
rect 2070 -468 2076 -462
rect 2070 -474 2076 -468
rect 2070 -480 2076 -474
rect 2070 -486 2076 -480
rect 2070 -492 2076 -486
rect 2070 -498 2076 -492
rect 2070 -504 2076 -498
rect 2070 -510 2076 -504
rect 2070 -516 2076 -510
rect 2070 -522 2076 -516
rect 2070 -528 2076 -522
rect 2070 -534 2076 -528
rect 2070 -540 2076 -534
rect 2070 -546 2076 -540
rect 2070 -552 2076 -546
rect 2070 -558 2076 -552
rect 2070 -564 2076 -558
rect 2070 -570 2076 -564
rect 2070 -576 2076 -570
rect 2070 -582 2076 -576
rect 2070 -588 2076 -582
rect 2070 -594 2076 -588
rect 2070 -600 2076 -594
rect 2070 -606 2076 -600
rect 2070 -612 2076 -606
rect 2070 -618 2076 -612
rect 2070 -624 2076 -618
rect 2070 -630 2076 -624
rect 2070 -636 2076 -630
rect 2070 -642 2076 -636
rect 2070 -648 2076 -642
rect 2070 -654 2076 -648
rect 2070 -660 2076 -654
rect 2070 -666 2076 -660
rect 2070 -672 2076 -666
rect 2070 -678 2076 -672
rect 2070 -684 2076 -678
rect 2070 -690 2076 -684
rect 2070 -696 2076 -690
rect 2070 -702 2076 -696
rect 2070 -708 2076 -702
rect 2070 -714 2076 -708
rect 2070 -720 2076 -714
rect 2070 -726 2076 -720
rect 2070 -732 2076 -726
rect 2070 -738 2076 -732
rect 2070 -744 2076 -738
rect 2070 -750 2076 -744
rect 2070 -756 2076 -750
rect 2070 -762 2076 -756
rect 2070 -768 2076 -762
rect 2070 -774 2076 -768
rect 2070 -780 2076 -774
rect 2070 -786 2076 -780
rect 2070 -792 2076 -786
rect 2070 -798 2076 -792
rect 2070 -804 2076 -798
rect 2070 -810 2076 -804
rect 2070 -816 2076 -810
rect 2070 -822 2076 -816
rect 2070 -828 2076 -822
rect 2070 -834 2076 -828
rect 2070 -840 2076 -834
rect 2070 -846 2076 -840
rect 2070 -852 2076 -846
rect 2070 -858 2076 -852
rect 2070 -864 2076 -858
rect 2070 -870 2076 -864
rect 2070 -876 2076 -870
rect 2070 -882 2076 -876
rect 2070 -888 2076 -882
rect 2070 -894 2076 -888
rect 2070 -900 2076 -894
rect 2070 -906 2076 -900
rect 2070 -912 2076 -906
rect 2070 -918 2076 -912
rect 2070 -924 2076 -918
rect 2070 -930 2076 -924
rect 2070 -936 2076 -930
rect 2070 -942 2076 -936
rect 2070 -948 2076 -942
rect 2070 -954 2076 -948
rect 2070 -960 2076 -954
rect 2070 -966 2076 -960
rect 2070 -972 2076 -966
rect 2070 -978 2076 -972
rect 2070 -984 2076 -978
rect 2070 -990 2076 -984
rect 2070 -996 2076 -990
rect 2070 -1002 2076 -996
rect 2070 -1008 2076 -1002
rect 2070 -1014 2076 -1008
rect 2070 -1020 2076 -1014
rect 2070 -1026 2076 -1020
rect 2070 -1032 2076 -1026
rect 2070 -1038 2076 -1032
rect 2070 -1044 2076 -1038
rect 2070 -1050 2076 -1044
rect 2070 -1056 2076 -1050
rect 2070 -1062 2076 -1056
rect 2070 -1068 2076 -1062
rect 2070 -1074 2076 -1068
rect 2070 -1080 2076 -1074
rect 2070 -1086 2076 -1080
rect 2070 -1092 2076 -1086
rect 2070 -1098 2076 -1092
rect 2070 -1104 2076 -1098
rect 2070 -1110 2076 -1104
rect 2070 -1116 2076 -1110
rect 2070 -1122 2076 -1116
rect 2070 -1128 2076 -1122
rect 2070 -1134 2076 -1128
rect 2070 -1140 2076 -1134
rect 2070 -1146 2076 -1140
rect 2070 -1152 2076 -1146
rect 2070 -1158 2076 -1152
rect 2070 -1164 2076 -1158
rect 2070 -1170 2076 -1164
rect 2070 -1176 2076 -1170
rect 2070 -1182 2076 -1176
rect 2070 -1188 2076 -1182
rect 2070 -1194 2076 -1188
rect 2070 -1200 2076 -1194
rect 2070 -1206 2076 -1200
rect 2070 -1212 2076 -1206
rect 2070 -1218 2076 -1212
rect 2070 -1224 2076 -1218
rect 2070 -1230 2076 -1224
rect 2070 -1236 2076 -1230
rect 2070 -1242 2076 -1236
rect 2070 -1248 2076 -1242
rect 2070 -1254 2076 -1248
rect 2070 -1260 2076 -1254
rect 2070 -1266 2076 -1260
rect 2070 -1272 2076 -1266
rect 2070 -1278 2076 -1272
rect 2070 -1284 2076 -1278
rect 2070 -1290 2076 -1284
rect 2070 -1296 2076 -1290
rect 2070 -1302 2076 -1296
rect 2070 -1308 2076 -1302
rect 2070 -1314 2076 -1308
rect 2070 -1320 2076 -1314
rect 2070 -1326 2076 -1320
rect 2070 -1332 2076 -1326
rect 2070 -1338 2076 -1332
rect 2070 -1344 2076 -1338
rect 2070 -1350 2076 -1344
rect 2070 -1356 2076 -1350
rect 2070 -1362 2076 -1356
rect 2070 -1368 2076 -1362
rect 2070 -1374 2076 -1368
rect 2070 -1380 2076 -1374
rect 2070 -1386 2076 -1380
rect 2070 -1392 2076 -1386
rect 2070 -1398 2076 -1392
rect 2070 -1404 2076 -1398
rect 2070 -1410 2076 -1404
rect 2070 -1416 2076 -1410
rect 2070 -1422 2076 -1416
rect 2070 -1428 2076 -1422
rect 2070 -1434 2076 -1428
rect 2070 -1440 2076 -1434
rect 2070 -1446 2076 -1440
rect 2070 -1452 2076 -1446
rect 2070 -1458 2076 -1452
rect 2070 -1464 2076 -1458
rect 2070 -1470 2076 -1464
rect 2070 -1476 2076 -1470
rect 2070 -1482 2076 -1476
rect 2070 -1488 2076 -1482
rect 2070 -1494 2076 -1488
rect 2070 -1500 2076 -1494
rect 2070 -1506 2076 -1500
rect 2070 -1512 2076 -1506
rect 2070 -1518 2076 -1512
rect 2070 -1524 2076 -1518
rect 2070 -1530 2076 -1524
rect 2070 -1536 2076 -1530
rect 2070 -1542 2076 -1536
rect 2070 -1548 2076 -1542
rect 2070 -1554 2076 -1548
rect 2070 -1668 2076 -1662
rect 2070 -1674 2076 -1668
rect 2070 -1680 2076 -1674
rect 2070 -1686 2076 -1680
rect 2070 -1692 2076 -1686
rect 2070 -1698 2076 -1692
rect 2070 -1704 2076 -1698
rect 2070 -1710 2076 -1704
rect 2070 -1716 2076 -1710
rect 2070 -1722 2076 -1716
rect 2070 -1728 2076 -1722
rect 2070 -1734 2076 -1728
rect 2070 -1740 2076 -1734
rect 2070 -1746 2076 -1740
rect 2070 -1752 2076 -1746
rect 2070 -1758 2076 -1752
rect 2070 -1764 2076 -1758
rect 2070 -1770 2076 -1764
rect 2070 -1776 2076 -1770
rect 2070 -1782 2076 -1776
rect 2070 -1788 2076 -1782
rect 2070 -1794 2076 -1788
rect 2070 -1800 2076 -1794
rect 2070 -1806 2076 -1800
rect 2070 -1812 2076 -1806
rect 2070 -1818 2076 -1812
rect 2070 -1824 2076 -1818
rect 2070 -1830 2076 -1824
rect 2070 -1836 2076 -1830
rect 2070 -1842 2076 -1836
rect 2070 -1848 2076 -1842
rect 2070 -1854 2076 -1848
rect 2070 -1860 2076 -1854
rect 2070 -1866 2076 -1860
rect 2070 -1872 2076 -1866
rect 2070 -1878 2076 -1872
rect 2070 -1884 2076 -1878
rect 2070 -1890 2076 -1884
rect 2070 -1896 2076 -1890
rect 2070 -1902 2076 -1896
rect 2070 -1908 2076 -1902
rect 2070 -1914 2076 -1908
rect 2070 -1920 2076 -1914
rect 2070 -1926 2076 -1920
rect 2070 -1932 2076 -1926
rect 2070 -1938 2076 -1932
rect 2070 -1944 2076 -1938
rect 2070 -1950 2076 -1944
rect 2070 -1956 2076 -1950
rect 2070 -1962 2076 -1956
rect 2070 -1968 2076 -1962
rect 2070 -1974 2076 -1968
rect 2070 -1980 2076 -1974
rect 2070 -1986 2076 -1980
rect 2070 -1992 2076 -1986
rect 2070 -1998 2076 -1992
rect 2070 -2004 2076 -1998
rect 2070 -2010 2076 -2004
rect 2070 -2016 2076 -2010
rect 2070 -2022 2076 -2016
rect 2070 -2028 2076 -2022
rect 2070 -2034 2076 -2028
rect 2070 -2040 2076 -2034
rect 2070 -2046 2076 -2040
rect 2070 -2052 2076 -2046
rect 2070 -2058 2076 -2052
rect 2070 -2064 2076 -2058
rect 2070 -2070 2076 -2064
rect 2070 -2076 2076 -2070
rect 2070 -2082 2076 -2076
rect 2070 -2088 2076 -2082
rect 2070 -2094 2076 -2088
rect 2070 -2100 2076 -2094
rect 2070 -2106 2076 -2100
rect 2070 -2112 2076 -2106
rect 2070 -2118 2076 -2112
rect 2070 -2124 2076 -2118
rect 2070 -2130 2076 -2124
rect 2070 -2136 2076 -2130
rect 2070 -2142 2076 -2136
rect 2070 -2148 2076 -2142
rect 2070 -2154 2076 -2148
rect 2070 -2160 2076 -2154
rect 2070 -2166 2076 -2160
rect 2070 -2172 2076 -2166
rect 2070 -2178 2076 -2172
rect 2070 -2184 2076 -2178
rect 2070 -2190 2076 -2184
rect 2070 -2196 2076 -2190
rect 2070 -2202 2076 -2196
rect 2070 -2208 2076 -2202
rect 2070 -2214 2076 -2208
rect 2070 -2220 2076 -2214
rect 2070 -2226 2076 -2220
rect 2070 -2232 2076 -2226
rect 2070 -2238 2076 -2232
rect 2070 -2244 2076 -2238
rect 2070 -2250 2076 -2244
rect 2070 -2256 2076 -2250
rect 2070 -2262 2076 -2256
rect 2070 -2268 2076 -2262
rect 2070 -2274 2076 -2268
rect 2070 -2280 2076 -2274
rect 2070 -2286 2076 -2280
rect 2070 -2292 2076 -2286
rect 2070 -2298 2076 -2292
rect 2070 -2304 2076 -2298
rect 2070 -2310 2076 -2304
rect 2070 -2316 2076 -2310
rect 2070 -2322 2076 -2316
rect 2070 -2328 2076 -2322
rect 2070 -2334 2076 -2328
rect 2070 -2340 2076 -2334
rect 2070 -2346 2076 -2340
rect 2070 -2352 2076 -2346
rect 2070 -2358 2076 -2352
rect 2070 -2364 2076 -2358
rect 2070 -2370 2076 -2364
rect 2070 -2376 2076 -2370
rect 2070 -2382 2076 -2376
rect 2070 -2388 2076 -2382
rect 2070 -2394 2076 -2388
rect 2070 -2400 2076 -2394
rect 2070 -2406 2076 -2400
rect 2070 -2412 2076 -2406
rect 2070 -2418 2076 -2412
rect 2070 -2424 2076 -2418
rect 2070 -2430 2076 -2424
rect 2070 -2436 2076 -2430
rect 2070 -2442 2076 -2436
rect 2070 -2448 2076 -2442
rect 2070 -2454 2076 -2448
rect 2070 -2460 2076 -2454
rect 2070 -2466 2076 -2460
rect 2070 -2472 2076 -2466
rect 2070 -2478 2076 -2472
rect 2070 -2484 2076 -2478
rect 2070 -2490 2076 -2484
rect 2070 -2586 2076 -2580
rect 2070 -2592 2076 -2586
rect 2070 -2598 2076 -2592
rect 2070 -2604 2076 -2598
rect 2070 -2610 2076 -2604
rect 2070 -2616 2076 -2610
rect 2070 -2622 2076 -2616
rect 2070 -2628 2076 -2622
rect 2070 -2634 2076 -2628
rect 2070 -2640 2076 -2634
rect 2070 -2646 2076 -2640
rect 2070 -2652 2076 -2646
rect 2070 -2658 2076 -2652
rect 2070 -2664 2076 -2658
rect 2070 -2670 2076 -2664
rect 2070 -2676 2076 -2670
rect 2070 -2682 2076 -2676
rect 2070 -2688 2076 -2682
rect 2070 -2694 2076 -2688
rect 2070 -2700 2076 -2694
rect 2070 -2706 2076 -2700
rect 2070 -2712 2076 -2706
rect 2070 -2718 2076 -2712
rect 2070 -2724 2076 -2718
rect 2070 -2730 2076 -2724
rect 2070 -2736 2076 -2730
rect 2070 -2742 2076 -2736
rect 2070 -2748 2076 -2742
rect 2070 -2754 2076 -2748
rect 2070 -2760 2076 -2754
rect 2070 -2766 2076 -2760
rect 2070 -2772 2076 -2766
rect 2070 -2778 2076 -2772
rect 2070 -2784 2076 -2778
rect 2070 -2790 2076 -2784
rect 2070 -2796 2076 -2790
rect 2070 -2802 2076 -2796
rect 2070 -2808 2076 -2802
rect 2070 -2814 2076 -2808
rect 2070 -2820 2076 -2814
rect 2070 -2826 2076 -2820
rect 2070 -2832 2076 -2826
rect 2070 -2838 2076 -2832
rect 2070 -2844 2076 -2838
rect 2070 -2850 2076 -2844
rect 2070 -2856 2076 -2850
rect 2070 -2862 2076 -2856
rect 2070 -2868 2076 -2862
rect 2070 -2874 2076 -2868
rect 2070 -2880 2076 -2874
rect 2070 -2886 2076 -2880
rect 2070 -2892 2076 -2886
rect 2070 -2898 2076 -2892
rect 2070 -2904 2076 -2898
rect 2070 -2910 2076 -2904
rect 2070 -2916 2076 -2910
rect 2070 -2922 2076 -2916
rect 2070 -2928 2076 -2922
rect 2070 -2934 2076 -2928
rect 2070 -2940 2076 -2934
rect 2070 -2946 2076 -2940
rect 2070 -2952 2076 -2946
rect 2070 -2958 2076 -2952
rect 2070 -2964 2076 -2958
rect 2070 -2970 2076 -2964
rect 2070 -2976 2076 -2970
rect 2070 -2982 2076 -2976
rect 2070 -2988 2076 -2982
rect 2070 -2994 2076 -2988
rect 2070 -3000 2076 -2994
rect 2070 -3006 2076 -3000
rect 2070 -3012 2076 -3006
rect 2070 -3018 2076 -3012
rect 2070 -3024 2076 -3018
rect 2070 -3030 2076 -3024
rect 2070 -3036 2076 -3030
rect 2070 -3042 2076 -3036
rect 2070 -3048 2076 -3042
rect 2070 -3054 2076 -3048
rect 2070 -3060 2076 -3054
rect 2070 -3066 2076 -3060
rect 2070 -3072 2076 -3066
rect 2070 -3078 2076 -3072
rect 2070 -3132 2076 -3126
rect 2070 -3138 2076 -3132
rect 2070 -3144 2076 -3138
rect 2070 -3150 2076 -3144
rect 2070 -3156 2076 -3150
rect 2076 -354 2082 -348
rect 2076 -360 2082 -354
rect 2076 -366 2082 -360
rect 2076 -372 2082 -366
rect 2076 -378 2082 -372
rect 2076 -384 2082 -378
rect 2076 -390 2082 -384
rect 2076 -396 2082 -390
rect 2076 -402 2082 -396
rect 2076 -408 2082 -402
rect 2076 -414 2082 -408
rect 2076 -420 2082 -414
rect 2076 -426 2082 -420
rect 2076 -432 2082 -426
rect 2076 -438 2082 -432
rect 2076 -444 2082 -438
rect 2076 -450 2082 -444
rect 2076 -456 2082 -450
rect 2076 -462 2082 -456
rect 2076 -468 2082 -462
rect 2076 -474 2082 -468
rect 2076 -480 2082 -474
rect 2076 -486 2082 -480
rect 2076 -492 2082 -486
rect 2076 -498 2082 -492
rect 2076 -504 2082 -498
rect 2076 -510 2082 -504
rect 2076 -516 2082 -510
rect 2076 -522 2082 -516
rect 2076 -528 2082 -522
rect 2076 -534 2082 -528
rect 2076 -540 2082 -534
rect 2076 -546 2082 -540
rect 2076 -552 2082 -546
rect 2076 -558 2082 -552
rect 2076 -564 2082 -558
rect 2076 -570 2082 -564
rect 2076 -576 2082 -570
rect 2076 -582 2082 -576
rect 2076 -588 2082 -582
rect 2076 -594 2082 -588
rect 2076 -600 2082 -594
rect 2076 -606 2082 -600
rect 2076 -612 2082 -606
rect 2076 -618 2082 -612
rect 2076 -624 2082 -618
rect 2076 -630 2082 -624
rect 2076 -636 2082 -630
rect 2076 -642 2082 -636
rect 2076 -648 2082 -642
rect 2076 -654 2082 -648
rect 2076 -660 2082 -654
rect 2076 -666 2082 -660
rect 2076 -672 2082 -666
rect 2076 -678 2082 -672
rect 2076 -684 2082 -678
rect 2076 -690 2082 -684
rect 2076 -696 2082 -690
rect 2076 -702 2082 -696
rect 2076 -708 2082 -702
rect 2076 -714 2082 -708
rect 2076 -720 2082 -714
rect 2076 -726 2082 -720
rect 2076 -732 2082 -726
rect 2076 -738 2082 -732
rect 2076 -744 2082 -738
rect 2076 -750 2082 -744
rect 2076 -756 2082 -750
rect 2076 -762 2082 -756
rect 2076 -768 2082 -762
rect 2076 -774 2082 -768
rect 2076 -780 2082 -774
rect 2076 -786 2082 -780
rect 2076 -792 2082 -786
rect 2076 -798 2082 -792
rect 2076 -804 2082 -798
rect 2076 -810 2082 -804
rect 2076 -816 2082 -810
rect 2076 -822 2082 -816
rect 2076 -828 2082 -822
rect 2076 -834 2082 -828
rect 2076 -840 2082 -834
rect 2076 -846 2082 -840
rect 2076 -852 2082 -846
rect 2076 -858 2082 -852
rect 2076 -864 2082 -858
rect 2076 -870 2082 -864
rect 2076 -876 2082 -870
rect 2076 -882 2082 -876
rect 2076 -888 2082 -882
rect 2076 -894 2082 -888
rect 2076 -900 2082 -894
rect 2076 -906 2082 -900
rect 2076 -912 2082 -906
rect 2076 -918 2082 -912
rect 2076 -924 2082 -918
rect 2076 -930 2082 -924
rect 2076 -936 2082 -930
rect 2076 -942 2082 -936
rect 2076 -948 2082 -942
rect 2076 -954 2082 -948
rect 2076 -960 2082 -954
rect 2076 -966 2082 -960
rect 2076 -972 2082 -966
rect 2076 -978 2082 -972
rect 2076 -984 2082 -978
rect 2076 -990 2082 -984
rect 2076 -996 2082 -990
rect 2076 -1002 2082 -996
rect 2076 -1008 2082 -1002
rect 2076 -1014 2082 -1008
rect 2076 -1020 2082 -1014
rect 2076 -1026 2082 -1020
rect 2076 -1032 2082 -1026
rect 2076 -1038 2082 -1032
rect 2076 -1044 2082 -1038
rect 2076 -1050 2082 -1044
rect 2076 -1056 2082 -1050
rect 2076 -1062 2082 -1056
rect 2076 -1068 2082 -1062
rect 2076 -1074 2082 -1068
rect 2076 -1080 2082 -1074
rect 2076 -1086 2082 -1080
rect 2076 -1092 2082 -1086
rect 2076 -1098 2082 -1092
rect 2076 -1104 2082 -1098
rect 2076 -1110 2082 -1104
rect 2076 -1116 2082 -1110
rect 2076 -1122 2082 -1116
rect 2076 -1128 2082 -1122
rect 2076 -1134 2082 -1128
rect 2076 -1140 2082 -1134
rect 2076 -1146 2082 -1140
rect 2076 -1152 2082 -1146
rect 2076 -1158 2082 -1152
rect 2076 -1164 2082 -1158
rect 2076 -1170 2082 -1164
rect 2076 -1176 2082 -1170
rect 2076 -1182 2082 -1176
rect 2076 -1188 2082 -1182
rect 2076 -1194 2082 -1188
rect 2076 -1200 2082 -1194
rect 2076 -1206 2082 -1200
rect 2076 -1212 2082 -1206
rect 2076 -1218 2082 -1212
rect 2076 -1224 2082 -1218
rect 2076 -1230 2082 -1224
rect 2076 -1236 2082 -1230
rect 2076 -1242 2082 -1236
rect 2076 -1248 2082 -1242
rect 2076 -1254 2082 -1248
rect 2076 -1260 2082 -1254
rect 2076 -1266 2082 -1260
rect 2076 -1272 2082 -1266
rect 2076 -1278 2082 -1272
rect 2076 -1284 2082 -1278
rect 2076 -1290 2082 -1284
rect 2076 -1296 2082 -1290
rect 2076 -1302 2082 -1296
rect 2076 -1308 2082 -1302
rect 2076 -1314 2082 -1308
rect 2076 -1320 2082 -1314
rect 2076 -1326 2082 -1320
rect 2076 -1332 2082 -1326
rect 2076 -1338 2082 -1332
rect 2076 -1344 2082 -1338
rect 2076 -1350 2082 -1344
rect 2076 -1356 2082 -1350
rect 2076 -1362 2082 -1356
rect 2076 -1368 2082 -1362
rect 2076 -1374 2082 -1368
rect 2076 -1380 2082 -1374
rect 2076 -1386 2082 -1380
rect 2076 -1392 2082 -1386
rect 2076 -1398 2082 -1392
rect 2076 -1404 2082 -1398
rect 2076 -1410 2082 -1404
rect 2076 -1416 2082 -1410
rect 2076 -1422 2082 -1416
rect 2076 -1428 2082 -1422
rect 2076 -1434 2082 -1428
rect 2076 -1440 2082 -1434
rect 2076 -1446 2082 -1440
rect 2076 -1452 2082 -1446
rect 2076 -1458 2082 -1452
rect 2076 -1464 2082 -1458
rect 2076 -1470 2082 -1464
rect 2076 -1476 2082 -1470
rect 2076 -1482 2082 -1476
rect 2076 -1488 2082 -1482
rect 2076 -1494 2082 -1488
rect 2076 -1500 2082 -1494
rect 2076 -1506 2082 -1500
rect 2076 -1512 2082 -1506
rect 2076 -1518 2082 -1512
rect 2076 -1524 2082 -1518
rect 2076 -1530 2082 -1524
rect 2076 -1536 2082 -1530
rect 2076 -1662 2082 -1656
rect 2076 -1668 2082 -1662
rect 2076 -1674 2082 -1668
rect 2076 -1680 2082 -1674
rect 2076 -1686 2082 -1680
rect 2076 -1692 2082 -1686
rect 2076 -1698 2082 -1692
rect 2076 -1704 2082 -1698
rect 2076 -1710 2082 -1704
rect 2076 -1716 2082 -1710
rect 2076 -1722 2082 -1716
rect 2076 -1728 2082 -1722
rect 2076 -1734 2082 -1728
rect 2076 -1740 2082 -1734
rect 2076 -1746 2082 -1740
rect 2076 -1752 2082 -1746
rect 2076 -1758 2082 -1752
rect 2076 -1764 2082 -1758
rect 2076 -1770 2082 -1764
rect 2076 -1776 2082 -1770
rect 2076 -1782 2082 -1776
rect 2076 -1788 2082 -1782
rect 2076 -1794 2082 -1788
rect 2076 -1800 2082 -1794
rect 2076 -1806 2082 -1800
rect 2076 -1812 2082 -1806
rect 2076 -1818 2082 -1812
rect 2076 -1824 2082 -1818
rect 2076 -1830 2082 -1824
rect 2076 -1836 2082 -1830
rect 2076 -1842 2082 -1836
rect 2076 -1848 2082 -1842
rect 2076 -1854 2082 -1848
rect 2076 -1860 2082 -1854
rect 2076 -1866 2082 -1860
rect 2076 -1872 2082 -1866
rect 2076 -1878 2082 -1872
rect 2076 -1884 2082 -1878
rect 2076 -1890 2082 -1884
rect 2076 -1896 2082 -1890
rect 2076 -1902 2082 -1896
rect 2076 -1908 2082 -1902
rect 2076 -1914 2082 -1908
rect 2076 -1920 2082 -1914
rect 2076 -1926 2082 -1920
rect 2076 -1932 2082 -1926
rect 2076 -1938 2082 -1932
rect 2076 -1944 2082 -1938
rect 2076 -1950 2082 -1944
rect 2076 -1956 2082 -1950
rect 2076 -1962 2082 -1956
rect 2076 -1968 2082 -1962
rect 2076 -1974 2082 -1968
rect 2076 -1980 2082 -1974
rect 2076 -1986 2082 -1980
rect 2076 -1992 2082 -1986
rect 2076 -1998 2082 -1992
rect 2076 -2004 2082 -1998
rect 2076 -2010 2082 -2004
rect 2076 -2016 2082 -2010
rect 2076 -2022 2082 -2016
rect 2076 -2028 2082 -2022
rect 2076 -2034 2082 -2028
rect 2076 -2040 2082 -2034
rect 2076 -2046 2082 -2040
rect 2076 -2052 2082 -2046
rect 2076 -2058 2082 -2052
rect 2076 -2064 2082 -2058
rect 2076 -2070 2082 -2064
rect 2076 -2076 2082 -2070
rect 2076 -2082 2082 -2076
rect 2076 -2088 2082 -2082
rect 2076 -2094 2082 -2088
rect 2076 -2100 2082 -2094
rect 2076 -2106 2082 -2100
rect 2076 -2112 2082 -2106
rect 2076 -2118 2082 -2112
rect 2076 -2124 2082 -2118
rect 2076 -2130 2082 -2124
rect 2076 -2136 2082 -2130
rect 2076 -2142 2082 -2136
rect 2076 -2148 2082 -2142
rect 2076 -2154 2082 -2148
rect 2076 -2160 2082 -2154
rect 2076 -2166 2082 -2160
rect 2076 -2172 2082 -2166
rect 2076 -2178 2082 -2172
rect 2076 -2184 2082 -2178
rect 2076 -2190 2082 -2184
rect 2076 -2196 2082 -2190
rect 2076 -2202 2082 -2196
rect 2076 -2208 2082 -2202
rect 2076 -2214 2082 -2208
rect 2076 -2220 2082 -2214
rect 2076 -2226 2082 -2220
rect 2076 -2232 2082 -2226
rect 2076 -2238 2082 -2232
rect 2076 -2244 2082 -2238
rect 2076 -2250 2082 -2244
rect 2076 -2256 2082 -2250
rect 2076 -2262 2082 -2256
rect 2076 -2268 2082 -2262
rect 2076 -2274 2082 -2268
rect 2076 -2280 2082 -2274
rect 2076 -2286 2082 -2280
rect 2076 -2292 2082 -2286
rect 2076 -2298 2082 -2292
rect 2076 -2304 2082 -2298
rect 2076 -2310 2082 -2304
rect 2076 -2316 2082 -2310
rect 2076 -2322 2082 -2316
rect 2076 -2328 2082 -2322
rect 2076 -2334 2082 -2328
rect 2076 -2340 2082 -2334
rect 2076 -2346 2082 -2340
rect 2076 -2352 2082 -2346
rect 2076 -2358 2082 -2352
rect 2076 -2364 2082 -2358
rect 2076 -2370 2082 -2364
rect 2076 -2376 2082 -2370
rect 2076 -2382 2082 -2376
rect 2076 -2388 2082 -2382
rect 2076 -2394 2082 -2388
rect 2076 -2400 2082 -2394
rect 2076 -2406 2082 -2400
rect 2076 -2412 2082 -2406
rect 2076 -2418 2082 -2412
rect 2076 -2424 2082 -2418
rect 2076 -2430 2082 -2424
rect 2076 -2436 2082 -2430
rect 2076 -2442 2082 -2436
rect 2076 -2448 2082 -2442
rect 2076 -2454 2082 -2448
rect 2076 -2460 2082 -2454
rect 2076 -2466 2082 -2460
rect 2076 -2472 2082 -2466
rect 2076 -2478 2082 -2472
rect 2076 -2484 2082 -2478
rect 2076 -2490 2082 -2484
rect 2076 -2580 2082 -2574
rect 2076 -2586 2082 -2580
rect 2076 -2592 2082 -2586
rect 2076 -2598 2082 -2592
rect 2076 -2604 2082 -2598
rect 2076 -2610 2082 -2604
rect 2076 -2616 2082 -2610
rect 2076 -2622 2082 -2616
rect 2076 -2628 2082 -2622
rect 2076 -2634 2082 -2628
rect 2076 -2640 2082 -2634
rect 2076 -2646 2082 -2640
rect 2076 -2652 2082 -2646
rect 2076 -2658 2082 -2652
rect 2076 -2664 2082 -2658
rect 2076 -2670 2082 -2664
rect 2076 -2676 2082 -2670
rect 2076 -2682 2082 -2676
rect 2076 -2688 2082 -2682
rect 2076 -2694 2082 -2688
rect 2076 -2700 2082 -2694
rect 2076 -2706 2082 -2700
rect 2076 -2712 2082 -2706
rect 2076 -2718 2082 -2712
rect 2076 -2724 2082 -2718
rect 2076 -2730 2082 -2724
rect 2076 -2736 2082 -2730
rect 2076 -2742 2082 -2736
rect 2076 -2748 2082 -2742
rect 2076 -2754 2082 -2748
rect 2076 -2760 2082 -2754
rect 2076 -2766 2082 -2760
rect 2076 -2772 2082 -2766
rect 2076 -2778 2082 -2772
rect 2076 -2784 2082 -2778
rect 2076 -2790 2082 -2784
rect 2076 -2796 2082 -2790
rect 2076 -2802 2082 -2796
rect 2076 -2808 2082 -2802
rect 2076 -2814 2082 -2808
rect 2076 -2820 2082 -2814
rect 2076 -2826 2082 -2820
rect 2076 -2832 2082 -2826
rect 2076 -2838 2082 -2832
rect 2076 -2844 2082 -2838
rect 2076 -2850 2082 -2844
rect 2076 -2856 2082 -2850
rect 2076 -2862 2082 -2856
rect 2076 -2868 2082 -2862
rect 2076 -2874 2082 -2868
rect 2076 -2880 2082 -2874
rect 2076 -2886 2082 -2880
rect 2076 -2892 2082 -2886
rect 2076 -2898 2082 -2892
rect 2076 -2904 2082 -2898
rect 2076 -2910 2082 -2904
rect 2076 -2916 2082 -2910
rect 2076 -2922 2082 -2916
rect 2076 -2928 2082 -2922
rect 2076 -2934 2082 -2928
rect 2076 -2940 2082 -2934
rect 2076 -2946 2082 -2940
rect 2076 -2952 2082 -2946
rect 2076 -2958 2082 -2952
rect 2076 -2964 2082 -2958
rect 2076 -2970 2082 -2964
rect 2076 -2976 2082 -2970
rect 2076 -2982 2082 -2976
rect 2076 -2988 2082 -2982
rect 2076 -2994 2082 -2988
rect 2076 -3000 2082 -2994
rect 2076 -3006 2082 -3000
rect 2076 -3012 2082 -3006
rect 2076 -3018 2082 -3012
rect 2076 -3024 2082 -3018
rect 2076 -3030 2082 -3024
rect 2076 -3036 2082 -3030
rect 2076 -3042 2082 -3036
rect 2076 -3048 2082 -3042
rect 2076 -3054 2082 -3048
rect 2076 -3060 2082 -3054
rect 2076 -3066 2082 -3060
rect 2076 -3072 2082 -3066
rect 2076 -3132 2082 -3126
rect 2076 -3138 2082 -3132
rect 2076 -3144 2082 -3138
rect 2076 -3150 2082 -3144
rect 2082 -348 2088 -342
rect 2082 -354 2088 -348
rect 2082 -360 2088 -354
rect 2082 -366 2088 -360
rect 2082 -372 2088 -366
rect 2082 -378 2088 -372
rect 2082 -384 2088 -378
rect 2082 -390 2088 -384
rect 2082 -396 2088 -390
rect 2082 -402 2088 -396
rect 2082 -408 2088 -402
rect 2082 -414 2088 -408
rect 2082 -420 2088 -414
rect 2082 -426 2088 -420
rect 2082 -432 2088 -426
rect 2082 -438 2088 -432
rect 2082 -444 2088 -438
rect 2082 -450 2088 -444
rect 2082 -456 2088 -450
rect 2082 -462 2088 -456
rect 2082 -468 2088 -462
rect 2082 -474 2088 -468
rect 2082 -480 2088 -474
rect 2082 -486 2088 -480
rect 2082 -492 2088 -486
rect 2082 -498 2088 -492
rect 2082 -504 2088 -498
rect 2082 -510 2088 -504
rect 2082 -516 2088 -510
rect 2082 -522 2088 -516
rect 2082 -528 2088 -522
rect 2082 -534 2088 -528
rect 2082 -540 2088 -534
rect 2082 -546 2088 -540
rect 2082 -552 2088 -546
rect 2082 -558 2088 -552
rect 2082 -564 2088 -558
rect 2082 -570 2088 -564
rect 2082 -576 2088 -570
rect 2082 -582 2088 -576
rect 2082 -588 2088 -582
rect 2082 -594 2088 -588
rect 2082 -600 2088 -594
rect 2082 -606 2088 -600
rect 2082 -612 2088 -606
rect 2082 -618 2088 -612
rect 2082 -624 2088 -618
rect 2082 -630 2088 -624
rect 2082 -636 2088 -630
rect 2082 -642 2088 -636
rect 2082 -648 2088 -642
rect 2082 -654 2088 -648
rect 2082 -660 2088 -654
rect 2082 -666 2088 -660
rect 2082 -672 2088 -666
rect 2082 -678 2088 -672
rect 2082 -684 2088 -678
rect 2082 -690 2088 -684
rect 2082 -696 2088 -690
rect 2082 -702 2088 -696
rect 2082 -708 2088 -702
rect 2082 -714 2088 -708
rect 2082 -720 2088 -714
rect 2082 -726 2088 -720
rect 2082 -732 2088 -726
rect 2082 -738 2088 -732
rect 2082 -744 2088 -738
rect 2082 -750 2088 -744
rect 2082 -756 2088 -750
rect 2082 -762 2088 -756
rect 2082 -768 2088 -762
rect 2082 -774 2088 -768
rect 2082 -780 2088 -774
rect 2082 -786 2088 -780
rect 2082 -792 2088 -786
rect 2082 -798 2088 -792
rect 2082 -804 2088 -798
rect 2082 -810 2088 -804
rect 2082 -816 2088 -810
rect 2082 -822 2088 -816
rect 2082 -828 2088 -822
rect 2082 -834 2088 -828
rect 2082 -840 2088 -834
rect 2082 -846 2088 -840
rect 2082 -852 2088 -846
rect 2082 -858 2088 -852
rect 2082 -864 2088 -858
rect 2082 -870 2088 -864
rect 2082 -876 2088 -870
rect 2082 -882 2088 -876
rect 2082 -888 2088 -882
rect 2082 -894 2088 -888
rect 2082 -900 2088 -894
rect 2082 -906 2088 -900
rect 2082 -912 2088 -906
rect 2082 -918 2088 -912
rect 2082 -924 2088 -918
rect 2082 -930 2088 -924
rect 2082 -936 2088 -930
rect 2082 -942 2088 -936
rect 2082 -948 2088 -942
rect 2082 -954 2088 -948
rect 2082 -960 2088 -954
rect 2082 -966 2088 -960
rect 2082 -972 2088 -966
rect 2082 -978 2088 -972
rect 2082 -984 2088 -978
rect 2082 -990 2088 -984
rect 2082 -996 2088 -990
rect 2082 -1002 2088 -996
rect 2082 -1008 2088 -1002
rect 2082 -1014 2088 -1008
rect 2082 -1020 2088 -1014
rect 2082 -1026 2088 -1020
rect 2082 -1032 2088 -1026
rect 2082 -1038 2088 -1032
rect 2082 -1044 2088 -1038
rect 2082 -1050 2088 -1044
rect 2082 -1056 2088 -1050
rect 2082 -1062 2088 -1056
rect 2082 -1068 2088 -1062
rect 2082 -1074 2088 -1068
rect 2082 -1080 2088 -1074
rect 2082 -1086 2088 -1080
rect 2082 -1092 2088 -1086
rect 2082 -1098 2088 -1092
rect 2082 -1104 2088 -1098
rect 2082 -1110 2088 -1104
rect 2082 -1116 2088 -1110
rect 2082 -1122 2088 -1116
rect 2082 -1128 2088 -1122
rect 2082 -1134 2088 -1128
rect 2082 -1140 2088 -1134
rect 2082 -1146 2088 -1140
rect 2082 -1152 2088 -1146
rect 2082 -1158 2088 -1152
rect 2082 -1164 2088 -1158
rect 2082 -1170 2088 -1164
rect 2082 -1176 2088 -1170
rect 2082 -1182 2088 -1176
rect 2082 -1188 2088 -1182
rect 2082 -1194 2088 -1188
rect 2082 -1200 2088 -1194
rect 2082 -1206 2088 -1200
rect 2082 -1212 2088 -1206
rect 2082 -1218 2088 -1212
rect 2082 -1224 2088 -1218
rect 2082 -1230 2088 -1224
rect 2082 -1236 2088 -1230
rect 2082 -1242 2088 -1236
rect 2082 -1248 2088 -1242
rect 2082 -1254 2088 -1248
rect 2082 -1260 2088 -1254
rect 2082 -1266 2088 -1260
rect 2082 -1272 2088 -1266
rect 2082 -1278 2088 -1272
rect 2082 -1284 2088 -1278
rect 2082 -1290 2088 -1284
rect 2082 -1296 2088 -1290
rect 2082 -1302 2088 -1296
rect 2082 -1308 2088 -1302
rect 2082 -1314 2088 -1308
rect 2082 -1320 2088 -1314
rect 2082 -1326 2088 -1320
rect 2082 -1332 2088 -1326
rect 2082 -1338 2088 -1332
rect 2082 -1344 2088 -1338
rect 2082 -1350 2088 -1344
rect 2082 -1356 2088 -1350
rect 2082 -1362 2088 -1356
rect 2082 -1368 2088 -1362
rect 2082 -1374 2088 -1368
rect 2082 -1380 2088 -1374
rect 2082 -1386 2088 -1380
rect 2082 -1392 2088 -1386
rect 2082 -1398 2088 -1392
rect 2082 -1404 2088 -1398
rect 2082 -1410 2088 -1404
rect 2082 -1416 2088 -1410
rect 2082 -1422 2088 -1416
rect 2082 -1428 2088 -1422
rect 2082 -1434 2088 -1428
rect 2082 -1440 2088 -1434
rect 2082 -1446 2088 -1440
rect 2082 -1452 2088 -1446
rect 2082 -1458 2088 -1452
rect 2082 -1464 2088 -1458
rect 2082 -1470 2088 -1464
rect 2082 -1476 2088 -1470
rect 2082 -1482 2088 -1476
rect 2082 -1488 2088 -1482
rect 2082 -1494 2088 -1488
rect 2082 -1500 2088 -1494
rect 2082 -1506 2088 -1500
rect 2082 -1512 2088 -1506
rect 2082 -1518 2088 -1512
rect 2082 -1524 2088 -1518
rect 2082 -1656 2088 -1650
rect 2082 -1662 2088 -1656
rect 2082 -1668 2088 -1662
rect 2082 -1674 2088 -1668
rect 2082 -1680 2088 -1674
rect 2082 -1686 2088 -1680
rect 2082 -1692 2088 -1686
rect 2082 -1698 2088 -1692
rect 2082 -1704 2088 -1698
rect 2082 -1710 2088 -1704
rect 2082 -1716 2088 -1710
rect 2082 -1722 2088 -1716
rect 2082 -1728 2088 -1722
rect 2082 -1734 2088 -1728
rect 2082 -1740 2088 -1734
rect 2082 -1746 2088 -1740
rect 2082 -1752 2088 -1746
rect 2082 -1758 2088 -1752
rect 2082 -1764 2088 -1758
rect 2082 -1770 2088 -1764
rect 2082 -1776 2088 -1770
rect 2082 -1782 2088 -1776
rect 2082 -1788 2088 -1782
rect 2082 -1794 2088 -1788
rect 2082 -1800 2088 -1794
rect 2082 -1806 2088 -1800
rect 2082 -1812 2088 -1806
rect 2082 -1818 2088 -1812
rect 2082 -1824 2088 -1818
rect 2082 -1830 2088 -1824
rect 2082 -1836 2088 -1830
rect 2082 -1842 2088 -1836
rect 2082 -1848 2088 -1842
rect 2082 -1854 2088 -1848
rect 2082 -1860 2088 -1854
rect 2082 -1866 2088 -1860
rect 2082 -1872 2088 -1866
rect 2082 -1878 2088 -1872
rect 2082 -1884 2088 -1878
rect 2082 -1890 2088 -1884
rect 2082 -1896 2088 -1890
rect 2082 -1902 2088 -1896
rect 2082 -1908 2088 -1902
rect 2082 -1914 2088 -1908
rect 2082 -1920 2088 -1914
rect 2082 -1926 2088 -1920
rect 2082 -1932 2088 -1926
rect 2082 -1938 2088 -1932
rect 2082 -1944 2088 -1938
rect 2082 -1950 2088 -1944
rect 2082 -1956 2088 -1950
rect 2082 -1962 2088 -1956
rect 2082 -1968 2088 -1962
rect 2082 -1974 2088 -1968
rect 2082 -1980 2088 -1974
rect 2082 -1986 2088 -1980
rect 2082 -1992 2088 -1986
rect 2082 -1998 2088 -1992
rect 2082 -2004 2088 -1998
rect 2082 -2010 2088 -2004
rect 2082 -2016 2088 -2010
rect 2082 -2022 2088 -2016
rect 2082 -2028 2088 -2022
rect 2082 -2034 2088 -2028
rect 2082 -2040 2088 -2034
rect 2082 -2046 2088 -2040
rect 2082 -2052 2088 -2046
rect 2082 -2058 2088 -2052
rect 2082 -2064 2088 -2058
rect 2082 -2070 2088 -2064
rect 2082 -2076 2088 -2070
rect 2082 -2082 2088 -2076
rect 2082 -2088 2088 -2082
rect 2082 -2094 2088 -2088
rect 2082 -2100 2088 -2094
rect 2082 -2106 2088 -2100
rect 2082 -2112 2088 -2106
rect 2082 -2118 2088 -2112
rect 2082 -2124 2088 -2118
rect 2082 -2130 2088 -2124
rect 2082 -2136 2088 -2130
rect 2082 -2142 2088 -2136
rect 2082 -2148 2088 -2142
rect 2082 -2154 2088 -2148
rect 2082 -2160 2088 -2154
rect 2082 -2166 2088 -2160
rect 2082 -2172 2088 -2166
rect 2082 -2178 2088 -2172
rect 2082 -2184 2088 -2178
rect 2082 -2190 2088 -2184
rect 2082 -2196 2088 -2190
rect 2082 -2202 2088 -2196
rect 2082 -2208 2088 -2202
rect 2082 -2214 2088 -2208
rect 2082 -2220 2088 -2214
rect 2082 -2226 2088 -2220
rect 2082 -2232 2088 -2226
rect 2082 -2238 2088 -2232
rect 2082 -2244 2088 -2238
rect 2082 -2250 2088 -2244
rect 2082 -2256 2088 -2250
rect 2082 -2262 2088 -2256
rect 2082 -2268 2088 -2262
rect 2082 -2274 2088 -2268
rect 2082 -2280 2088 -2274
rect 2082 -2286 2088 -2280
rect 2082 -2292 2088 -2286
rect 2082 -2298 2088 -2292
rect 2082 -2304 2088 -2298
rect 2082 -2310 2088 -2304
rect 2082 -2316 2088 -2310
rect 2082 -2322 2088 -2316
rect 2082 -2328 2088 -2322
rect 2082 -2334 2088 -2328
rect 2082 -2340 2088 -2334
rect 2082 -2346 2088 -2340
rect 2082 -2352 2088 -2346
rect 2082 -2358 2088 -2352
rect 2082 -2364 2088 -2358
rect 2082 -2370 2088 -2364
rect 2082 -2376 2088 -2370
rect 2082 -2382 2088 -2376
rect 2082 -2388 2088 -2382
rect 2082 -2394 2088 -2388
rect 2082 -2400 2088 -2394
rect 2082 -2406 2088 -2400
rect 2082 -2412 2088 -2406
rect 2082 -2418 2088 -2412
rect 2082 -2424 2088 -2418
rect 2082 -2430 2088 -2424
rect 2082 -2436 2088 -2430
rect 2082 -2442 2088 -2436
rect 2082 -2448 2088 -2442
rect 2082 -2454 2088 -2448
rect 2082 -2460 2088 -2454
rect 2082 -2466 2088 -2460
rect 2082 -2472 2088 -2466
rect 2082 -2478 2088 -2472
rect 2082 -2484 2088 -2478
rect 2082 -2580 2088 -2574
rect 2082 -2586 2088 -2580
rect 2082 -2592 2088 -2586
rect 2082 -2598 2088 -2592
rect 2082 -2604 2088 -2598
rect 2082 -2610 2088 -2604
rect 2082 -2616 2088 -2610
rect 2082 -2622 2088 -2616
rect 2082 -2628 2088 -2622
rect 2082 -2634 2088 -2628
rect 2082 -2640 2088 -2634
rect 2082 -2646 2088 -2640
rect 2082 -2652 2088 -2646
rect 2082 -2658 2088 -2652
rect 2082 -2664 2088 -2658
rect 2082 -2670 2088 -2664
rect 2082 -2676 2088 -2670
rect 2082 -2682 2088 -2676
rect 2082 -2688 2088 -2682
rect 2082 -2694 2088 -2688
rect 2082 -2700 2088 -2694
rect 2082 -2706 2088 -2700
rect 2082 -2712 2088 -2706
rect 2082 -2718 2088 -2712
rect 2082 -2724 2088 -2718
rect 2082 -2730 2088 -2724
rect 2082 -2736 2088 -2730
rect 2082 -2742 2088 -2736
rect 2082 -2748 2088 -2742
rect 2082 -2754 2088 -2748
rect 2082 -2760 2088 -2754
rect 2082 -2766 2088 -2760
rect 2082 -2772 2088 -2766
rect 2082 -2778 2088 -2772
rect 2082 -2784 2088 -2778
rect 2082 -2790 2088 -2784
rect 2082 -2796 2088 -2790
rect 2082 -2802 2088 -2796
rect 2082 -2808 2088 -2802
rect 2082 -2814 2088 -2808
rect 2082 -2820 2088 -2814
rect 2082 -2826 2088 -2820
rect 2082 -2832 2088 -2826
rect 2082 -2838 2088 -2832
rect 2082 -2844 2088 -2838
rect 2082 -2850 2088 -2844
rect 2082 -2856 2088 -2850
rect 2082 -2862 2088 -2856
rect 2082 -2868 2088 -2862
rect 2082 -2874 2088 -2868
rect 2082 -2880 2088 -2874
rect 2082 -2886 2088 -2880
rect 2082 -2892 2088 -2886
rect 2082 -2898 2088 -2892
rect 2082 -2904 2088 -2898
rect 2082 -2910 2088 -2904
rect 2082 -2916 2088 -2910
rect 2082 -2922 2088 -2916
rect 2082 -2928 2088 -2922
rect 2082 -2934 2088 -2928
rect 2082 -2940 2088 -2934
rect 2082 -2946 2088 -2940
rect 2082 -2952 2088 -2946
rect 2082 -2958 2088 -2952
rect 2082 -2964 2088 -2958
rect 2082 -2970 2088 -2964
rect 2082 -2976 2088 -2970
rect 2082 -2982 2088 -2976
rect 2082 -2988 2088 -2982
rect 2082 -2994 2088 -2988
rect 2082 -3000 2088 -2994
rect 2082 -3006 2088 -3000
rect 2082 -3012 2088 -3006
rect 2082 -3018 2088 -3012
rect 2082 -3024 2088 -3018
rect 2082 -3030 2088 -3024
rect 2082 -3036 2088 -3030
rect 2082 -3042 2088 -3036
rect 2082 -3048 2088 -3042
rect 2082 -3054 2088 -3048
rect 2082 -3060 2088 -3054
rect 2082 -3066 2088 -3060
rect 2082 -3072 2088 -3066
rect 2082 -3126 2088 -3120
rect 2082 -3132 2088 -3126
rect 2082 -3138 2088 -3132
rect 2082 -3144 2088 -3138
rect 2088 -336 2094 -330
rect 2088 -342 2094 -336
rect 2088 -348 2094 -342
rect 2088 -354 2094 -348
rect 2088 -360 2094 -354
rect 2088 -366 2094 -360
rect 2088 -372 2094 -366
rect 2088 -378 2094 -372
rect 2088 -384 2094 -378
rect 2088 -390 2094 -384
rect 2088 -396 2094 -390
rect 2088 -402 2094 -396
rect 2088 -408 2094 -402
rect 2088 -414 2094 -408
rect 2088 -420 2094 -414
rect 2088 -426 2094 -420
rect 2088 -432 2094 -426
rect 2088 -438 2094 -432
rect 2088 -444 2094 -438
rect 2088 -450 2094 -444
rect 2088 -456 2094 -450
rect 2088 -462 2094 -456
rect 2088 -468 2094 -462
rect 2088 -474 2094 -468
rect 2088 -480 2094 -474
rect 2088 -486 2094 -480
rect 2088 -492 2094 -486
rect 2088 -498 2094 -492
rect 2088 -504 2094 -498
rect 2088 -510 2094 -504
rect 2088 -516 2094 -510
rect 2088 -522 2094 -516
rect 2088 -528 2094 -522
rect 2088 -534 2094 -528
rect 2088 -540 2094 -534
rect 2088 -546 2094 -540
rect 2088 -552 2094 -546
rect 2088 -558 2094 -552
rect 2088 -564 2094 -558
rect 2088 -570 2094 -564
rect 2088 -576 2094 -570
rect 2088 -582 2094 -576
rect 2088 -588 2094 -582
rect 2088 -594 2094 -588
rect 2088 -600 2094 -594
rect 2088 -606 2094 -600
rect 2088 -612 2094 -606
rect 2088 -618 2094 -612
rect 2088 -624 2094 -618
rect 2088 -630 2094 -624
rect 2088 -636 2094 -630
rect 2088 -642 2094 -636
rect 2088 -648 2094 -642
rect 2088 -654 2094 -648
rect 2088 -660 2094 -654
rect 2088 -666 2094 -660
rect 2088 -672 2094 -666
rect 2088 -678 2094 -672
rect 2088 -684 2094 -678
rect 2088 -690 2094 -684
rect 2088 -696 2094 -690
rect 2088 -702 2094 -696
rect 2088 -708 2094 -702
rect 2088 -714 2094 -708
rect 2088 -720 2094 -714
rect 2088 -726 2094 -720
rect 2088 -732 2094 -726
rect 2088 -738 2094 -732
rect 2088 -744 2094 -738
rect 2088 -750 2094 -744
rect 2088 -756 2094 -750
rect 2088 -762 2094 -756
rect 2088 -768 2094 -762
rect 2088 -774 2094 -768
rect 2088 -780 2094 -774
rect 2088 -786 2094 -780
rect 2088 -792 2094 -786
rect 2088 -798 2094 -792
rect 2088 -804 2094 -798
rect 2088 -810 2094 -804
rect 2088 -816 2094 -810
rect 2088 -822 2094 -816
rect 2088 -828 2094 -822
rect 2088 -834 2094 -828
rect 2088 -840 2094 -834
rect 2088 -846 2094 -840
rect 2088 -852 2094 -846
rect 2088 -858 2094 -852
rect 2088 -864 2094 -858
rect 2088 -870 2094 -864
rect 2088 -876 2094 -870
rect 2088 -882 2094 -876
rect 2088 -888 2094 -882
rect 2088 -894 2094 -888
rect 2088 -900 2094 -894
rect 2088 -906 2094 -900
rect 2088 -912 2094 -906
rect 2088 -918 2094 -912
rect 2088 -924 2094 -918
rect 2088 -930 2094 -924
rect 2088 -936 2094 -930
rect 2088 -942 2094 -936
rect 2088 -948 2094 -942
rect 2088 -954 2094 -948
rect 2088 -960 2094 -954
rect 2088 -966 2094 -960
rect 2088 -972 2094 -966
rect 2088 -978 2094 -972
rect 2088 -984 2094 -978
rect 2088 -990 2094 -984
rect 2088 -996 2094 -990
rect 2088 -1002 2094 -996
rect 2088 -1008 2094 -1002
rect 2088 -1014 2094 -1008
rect 2088 -1020 2094 -1014
rect 2088 -1026 2094 -1020
rect 2088 -1032 2094 -1026
rect 2088 -1038 2094 -1032
rect 2088 -1044 2094 -1038
rect 2088 -1050 2094 -1044
rect 2088 -1056 2094 -1050
rect 2088 -1062 2094 -1056
rect 2088 -1068 2094 -1062
rect 2088 -1074 2094 -1068
rect 2088 -1080 2094 -1074
rect 2088 -1086 2094 -1080
rect 2088 -1092 2094 -1086
rect 2088 -1098 2094 -1092
rect 2088 -1104 2094 -1098
rect 2088 -1110 2094 -1104
rect 2088 -1116 2094 -1110
rect 2088 -1122 2094 -1116
rect 2088 -1128 2094 -1122
rect 2088 -1134 2094 -1128
rect 2088 -1140 2094 -1134
rect 2088 -1146 2094 -1140
rect 2088 -1152 2094 -1146
rect 2088 -1158 2094 -1152
rect 2088 -1164 2094 -1158
rect 2088 -1170 2094 -1164
rect 2088 -1176 2094 -1170
rect 2088 -1182 2094 -1176
rect 2088 -1188 2094 -1182
rect 2088 -1194 2094 -1188
rect 2088 -1200 2094 -1194
rect 2088 -1206 2094 -1200
rect 2088 -1212 2094 -1206
rect 2088 -1218 2094 -1212
rect 2088 -1224 2094 -1218
rect 2088 -1230 2094 -1224
rect 2088 -1236 2094 -1230
rect 2088 -1242 2094 -1236
rect 2088 -1248 2094 -1242
rect 2088 -1254 2094 -1248
rect 2088 -1260 2094 -1254
rect 2088 -1266 2094 -1260
rect 2088 -1272 2094 -1266
rect 2088 -1278 2094 -1272
rect 2088 -1284 2094 -1278
rect 2088 -1290 2094 -1284
rect 2088 -1296 2094 -1290
rect 2088 -1302 2094 -1296
rect 2088 -1308 2094 -1302
rect 2088 -1314 2094 -1308
rect 2088 -1320 2094 -1314
rect 2088 -1326 2094 -1320
rect 2088 -1332 2094 -1326
rect 2088 -1338 2094 -1332
rect 2088 -1344 2094 -1338
rect 2088 -1350 2094 -1344
rect 2088 -1356 2094 -1350
rect 2088 -1362 2094 -1356
rect 2088 -1368 2094 -1362
rect 2088 -1374 2094 -1368
rect 2088 -1380 2094 -1374
rect 2088 -1386 2094 -1380
rect 2088 -1392 2094 -1386
rect 2088 -1398 2094 -1392
rect 2088 -1404 2094 -1398
rect 2088 -1410 2094 -1404
rect 2088 -1416 2094 -1410
rect 2088 -1422 2094 -1416
rect 2088 -1428 2094 -1422
rect 2088 -1434 2094 -1428
rect 2088 -1440 2094 -1434
rect 2088 -1446 2094 -1440
rect 2088 -1452 2094 -1446
rect 2088 -1458 2094 -1452
rect 2088 -1464 2094 -1458
rect 2088 -1470 2094 -1464
rect 2088 -1476 2094 -1470
rect 2088 -1482 2094 -1476
rect 2088 -1488 2094 -1482
rect 2088 -1494 2094 -1488
rect 2088 -1500 2094 -1494
rect 2088 -1506 2094 -1500
rect 2088 -1512 2094 -1506
rect 2088 -1650 2094 -1644
rect 2088 -1656 2094 -1650
rect 2088 -1662 2094 -1656
rect 2088 -1668 2094 -1662
rect 2088 -1674 2094 -1668
rect 2088 -1680 2094 -1674
rect 2088 -1686 2094 -1680
rect 2088 -1692 2094 -1686
rect 2088 -1698 2094 -1692
rect 2088 -1704 2094 -1698
rect 2088 -1710 2094 -1704
rect 2088 -1716 2094 -1710
rect 2088 -1722 2094 -1716
rect 2088 -1728 2094 -1722
rect 2088 -1734 2094 -1728
rect 2088 -1740 2094 -1734
rect 2088 -1746 2094 -1740
rect 2088 -1752 2094 -1746
rect 2088 -1758 2094 -1752
rect 2088 -1764 2094 -1758
rect 2088 -1770 2094 -1764
rect 2088 -1776 2094 -1770
rect 2088 -1782 2094 -1776
rect 2088 -1788 2094 -1782
rect 2088 -1794 2094 -1788
rect 2088 -1800 2094 -1794
rect 2088 -1806 2094 -1800
rect 2088 -1812 2094 -1806
rect 2088 -1818 2094 -1812
rect 2088 -1824 2094 -1818
rect 2088 -1830 2094 -1824
rect 2088 -1836 2094 -1830
rect 2088 -1842 2094 -1836
rect 2088 -1848 2094 -1842
rect 2088 -1854 2094 -1848
rect 2088 -1860 2094 -1854
rect 2088 -1866 2094 -1860
rect 2088 -1872 2094 -1866
rect 2088 -1878 2094 -1872
rect 2088 -1884 2094 -1878
rect 2088 -1890 2094 -1884
rect 2088 -1896 2094 -1890
rect 2088 -1902 2094 -1896
rect 2088 -1908 2094 -1902
rect 2088 -1914 2094 -1908
rect 2088 -1920 2094 -1914
rect 2088 -1926 2094 -1920
rect 2088 -1932 2094 -1926
rect 2088 -1938 2094 -1932
rect 2088 -1944 2094 -1938
rect 2088 -1950 2094 -1944
rect 2088 -1956 2094 -1950
rect 2088 -1962 2094 -1956
rect 2088 -1968 2094 -1962
rect 2088 -1974 2094 -1968
rect 2088 -1980 2094 -1974
rect 2088 -1986 2094 -1980
rect 2088 -1992 2094 -1986
rect 2088 -1998 2094 -1992
rect 2088 -2004 2094 -1998
rect 2088 -2010 2094 -2004
rect 2088 -2016 2094 -2010
rect 2088 -2022 2094 -2016
rect 2088 -2028 2094 -2022
rect 2088 -2034 2094 -2028
rect 2088 -2040 2094 -2034
rect 2088 -2046 2094 -2040
rect 2088 -2052 2094 -2046
rect 2088 -2058 2094 -2052
rect 2088 -2064 2094 -2058
rect 2088 -2070 2094 -2064
rect 2088 -2076 2094 -2070
rect 2088 -2082 2094 -2076
rect 2088 -2088 2094 -2082
rect 2088 -2094 2094 -2088
rect 2088 -2100 2094 -2094
rect 2088 -2106 2094 -2100
rect 2088 -2112 2094 -2106
rect 2088 -2118 2094 -2112
rect 2088 -2124 2094 -2118
rect 2088 -2130 2094 -2124
rect 2088 -2136 2094 -2130
rect 2088 -2142 2094 -2136
rect 2088 -2148 2094 -2142
rect 2088 -2154 2094 -2148
rect 2088 -2160 2094 -2154
rect 2088 -2166 2094 -2160
rect 2088 -2172 2094 -2166
rect 2088 -2178 2094 -2172
rect 2088 -2184 2094 -2178
rect 2088 -2190 2094 -2184
rect 2088 -2196 2094 -2190
rect 2088 -2202 2094 -2196
rect 2088 -2208 2094 -2202
rect 2088 -2214 2094 -2208
rect 2088 -2220 2094 -2214
rect 2088 -2226 2094 -2220
rect 2088 -2232 2094 -2226
rect 2088 -2238 2094 -2232
rect 2088 -2244 2094 -2238
rect 2088 -2250 2094 -2244
rect 2088 -2256 2094 -2250
rect 2088 -2262 2094 -2256
rect 2088 -2268 2094 -2262
rect 2088 -2274 2094 -2268
rect 2088 -2280 2094 -2274
rect 2088 -2286 2094 -2280
rect 2088 -2292 2094 -2286
rect 2088 -2298 2094 -2292
rect 2088 -2304 2094 -2298
rect 2088 -2310 2094 -2304
rect 2088 -2316 2094 -2310
rect 2088 -2322 2094 -2316
rect 2088 -2328 2094 -2322
rect 2088 -2334 2094 -2328
rect 2088 -2340 2094 -2334
rect 2088 -2346 2094 -2340
rect 2088 -2352 2094 -2346
rect 2088 -2358 2094 -2352
rect 2088 -2364 2094 -2358
rect 2088 -2370 2094 -2364
rect 2088 -2376 2094 -2370
rect 2088 -2382 2094 -2376
rect 2088 -2388 2094 -2382
rect 2088 -2394 2094 -2388
rect 2088 -2400 2094 -2394
rect 2088 -2406 2094 -2400
rect 2088 -2412 2094 -2406
rect 2088 -2418 2094 -2412
rect 2088 -2424 2094 -2418
rect 2088 -2430 2094 -2424
rect 2088 -2436 2094 -2430
rect 2088 -2442 2094 -2436
rect 2088 -2448 2094 -2442
rect 2088 -2454 2094 -2448
rect 2088 -2460 2094 -2454
rect 2088 -2466 2094 -2460
rect 2088 -2472 2094 -2466
rect 2088 -2478 2094 -2472
rect 2088 -2580 2094 -2574
rect 2088 -2586 2094 -2580
rect 2088 -2592 2094 -2586
rect 2088 -2598 2094 -2592
rect 2088 -2604 2094 -2598
rect 2088 -2610 2094 -2604
rect 2088 -2616 2094 -2610
rect 2088 -2622 2094 -2616
rect 2088 -2628 2094 -2622
rect 2088 -2634 2094 -2628
rect 2088 -2640 2094 -2634
rect 2088 -2646 2094 -2640
rect 2088 -2652 2094 -2646
rect 2088 -2658 2094 -2652
rect 2088 -2664 2094 -2658
rect 2088 -2670 2094 -2664
rect 2088 -2676 2094 -2670
rect 2088 -2682 2094 -2676
rect 2088 -2688 2094 -2682
rect 2088 -2694 2094 -2688
rect 2088 -2700 2094 -2694
rect 2088 -2706 2094 -2700
rect 2088 -2712 2094 -2706
rect 2088 -2718 2094 -2712
rect 2088 -2724 2094 -2718
rect 2088 -2730 2094 -2724
rect 2088 -2736 2094 -2730
rect 2088 -2742 2094 -2736
rect 2088 -2748 2094 -2742
rect 2088 -2754 2094 -2748
rect 2088 -2760 2094 -2754
rect 2088 -2766 2094 -2760
rect 2088 -2772 2094 -2766
rect 2088 -2778 2094 -2772
rect 2088 -2784 2094 -2778
rect 2088 -2790 2094 -2784
rect 2088 -2796 2094 -2790
rect 2088 -2802 2094 -2796
rect 2088 -2808 2094 -2802
rect 2088 -2814 2094 -2808
rect 2088 -2820 2094 -2814
rect 2088 -2826 2094 -2820
rect 2088 -2832 2094 -2826
rect 2088 -2838 2094 -2832
rect 2088 -2844 2094 -2838
rect 2088 -2850 2094 -2844
rect 2088 -2856 2094 -2850
rect 2088 -2862 2094 -2856
rect 2088 -2868 2094 -2862
rect 2088 -2874 2094 -2868
rect 2088 -2880 2094 -2874
rect 2088 -2886 2094 -2880
rect 2088 -2892 2094 -2886
rect 2088 -2898 2094 -2892
rect 2088 -2904 2094 -2898
rect 2088 -2910 2094 -2904
rect 2088 -2916 2094 -2910
rect 2088 -2922 2094 -2916
rect 2088 -2928 2094 -2922
rect 2088 -2934 2094 -2928
rect 2088 -2940 2094 -2934
rect 2088 -2946 2094 -2940
rect 2088 -2952 2094 -2946
rect 2088 -2958 2094 -2952
rect 2088 -2964 2094 -2958
rect 2088 -2970 2094 -2964
rect 2088 -2976 2094 -2970
rect 2088 -2982 2094 -2976
rect 2088 -2988 2094 -2982
rect 2088 -2994 2094 -2988
rect 2088 -3000 2094 -2994
rect 2088 -3006 2094 -3000
rect 2088 -3012 2094 -3006
rect 2088 -3018 2094 -3012
rect 2088 -3024 2094 -3018
rect 2088 -3030 2094 -3024
rect 2088 -3036 2094 -3030
rect 2088 -3042 2094 -3036
rect 2088 -3048 2094 -3042
rect 2088 -3054 2094 -3048
rect 2088 -3060 2094 -3054
rect 2088 -3066 2094 -3060
rect 2088 -3072 2094 -3066
rect 2088 -3126 2094 -3120
rect 2088 -3132 2094 -3126
rect 2088 -3138 2094 -3132
rect 2094 -330 2100 -324
rect 2094 -336 2100 -330
rect 2094 -342 2100 -336
rect 2094 -348 2100 -342
rect 2094 -354 2100 -348
rect 2094 -360 2100 -354
rect 2094 -366 2100 -360
rect 2094 -372 2100 -366
rect 2094 -378 2100 -372
rect 2094 -384 2100 -378
rect 2094 -390 2100 -384
rect 2094 -396 2100 -390
rect 2094 -402 2100 -396
rect 2094 -408 2100 -402
rect 2094 -414 2100 -408
rect 2094 -420 2100 -414
rect 2094 -426 2100 -420
rect 2094 -432 2100 -426
rect 2094 -438 2100 -432
rect 2094 -444 2100 -438
rect 2094 -450 2100 -444
rect 2094 -456 2100 -450
rect 2094 -462 2100 -456
rect 2094 -468 2100 -462
rect 2094 -474 2100 -468
rect 2094 -480 2100 -474
rect 2094 -486 2100 -480
rect 2094 -492 2100 -486
rect 2094 -498 2100 -492
rect 2094 -504 2100 -498
rect 2094 -510 2100 -504
rect 2094 -516 2100 -510
rect 2094 -522 2100 -516
rect 2094 -528 2100 -522
rect 2094 -534 2100 -528
rect 2094 -540 2100 -534
rect 2094 -546 2100 -540
rect 2094 -552 2100 -546
rect 2094 -558 2100 -552
rect 2094 -564 2100 -558
rect 2094 -570 2100 -564
rect 2094 -576 2100 -570
rect 2094 -582 2100 -576
rect 2094 -588 2100 -582
rect 2094 -594 2100 -588
rect 2094 -600 2100 -594
rect 2094 -606 2100 -600
rect 2094 -612 2100 -606
rect 2094 -618 2100 -612
rect 2094 -624 2100 -618
rect 2094 -630 2100 -624
rect 2094 -636 2100 -630
rect 2094 -642 2100 -636
rect 2094 -648 2100 -642
rect 2094 -654 2100 -648
rect 2094 -660 2100 -654
rect 2094 -666 2100 -660
rect 2094 -672 2100 -666
rect 2094 -678 2100 -672
rect 2094 -684 2100 -678
rect 2094 -690 2100 -684
rect 2094 -696 2100 -690
rect 2094 -702 2100 -696
rect 2094 -708 2100 -702
rect 2094 -714 2100 -708
rect 2094 -720 2100 -714
rect 2094 -726 2100 -720
rect 2094 -732 2100 -726
rect 2094 -738 2100 -732
rect 2094 -744 2100 -738
rect 2094 -750 2100 -744
rect 2094 -756 2100 -750
rect 2094 -762 2100 -756
rect 2094 -768 2100 -762
rect 2094 -774 2100 -768
rect 2094 -780 2100 -774
rect 2094 -786 2100 -780
rect 2094 -792 2100 -786
rect 2094 -798 2100 -792
rect 2094 -804 2100 -798
rect 2094 -810 2100 -804
rect 2094 -816 2100 -810
rect 2094 -822 2100 -816
rect 2094 -828 2100 -822
rect 2094 -834 2100 -828
rect 2094 -840 2100 -834
rect 2094 -846 2100 -840
rect 2094 -852 2100 -846
rect 2094 -858 2100 -852
rect 2094 -864 2100 -858
rect 2094 -870 2100 -864
rect 2094 -876 2100 -870
rect 2094 -882 2100 -876
rect 2094 -888 2100 -882
rect 2094 -894 2100 -888
rect 2094 -900 2100 -894
rect 2094 -906 2100 -900
rect 2094 -912 2100 -906
rect 2094 -918 2100 -912
rect 2094 -924 2100 -918
rect 2094 -930 2100 -924
rect 2094 -936 2100 -930
rect 2094 -942 2100 -936
rect 2094 -948 2100 -942
rect 2094 -954 2100 -948
rect 2094 -960 2100 -954
rect 2094 -966 2100 -960
rect 2094 -972 2100 -966
rect 2094 -978 2100 -972
rect 2094 -984 2100 -978
rect 2094 -990 2100 -984
rect 2094 -996 2100 -990
rect 2094 -1002 2100 -996
rect 2094 -1008 2100 -1002
rect 2094 -1014 2100 -1008
rect 2094 -1020 2100 -1014
rect 2094 -1026 2100 -1020
rect 2094 -1032 2100 -1026
rect 2094 -1038 2100 -1032
rect 2094 -1044 2100 -1038
rect 2094 -1050 2100 -1044
rect 2094 -1056 2100 -1050
rect 2094 -1062 2100 -1056
rect 2094 -1068 2100 -1062
rect 2094 -1074 2100 -1068
rect 2094 -1080 2100 -1074
rect 2094 -1086 2100 -1080
rect 2094 -1092 2100 -1086
rect 2094 -1098 2100 -1092
rect 2094 -1104 2100 -1098
rect 2094 -1110 2100 -1104
rect 2094 -1116 2100 -1110
rect 2094 -1122 2100 -1116
rect 2094 -1128 2100 -1122
rect 2094 -1134 2100 -1128
rect 2094 -1140 2100 -1134
rect 2094 -1146 2100 -1140
rect 2094 -1152 2100 -1146
rect 2094 -1158 2100 -1152
rect 2094 -1164 2100 -1158
rect 2094 -1170 2100 -1164
rect 2094 -1176 2100 -1170
rect 2094 -1182 2100 -1176
rect 2094 -1188 2100 -1182
rect 2094 -1194 2100 -1188
rect 2094 -1200 2100 -1194
rect 2094 -1206 2100 -1200
rect 2094 -1212 2100 -1206
rect 2094 -1218 2100 -1212
rect 2094 -1224 2100 -1218
rect 2094 -1230 2100 -1224
rect 2094 -1236 2100 -1230
rect 2094 -1242 2100 -1236
rect 2094 -1248 2100 -1242
rect 2094 -1254 2100 -1248
rect 2094 -1260 2100 -1254
rect 2094 -1266 2100 -1260
rect 2094 -1272 2100 -1266
rect 2094 -1278 2100 -1272
rect 2094 -1284 2100 -1278
rect 2094 -1290 2100 -1284
rect 2094 -1296 2100 -1290
rect 2094 -1302 2100 -1296
rect 2094 -1308 2100 -1302
rect 2094 -1314 2100 -1308
rect 2094 -1320 2100 -1314
rect 2094 -1326 2100 -1320
rect 2094 -1332 2100 -1326
rect 2094 -1338 2100 -1332
rect 2094 -1344 2100 -1338
rect 2094 -1350 2100 -1344
rect 2094 -1356 2100 -1350
rect 2094 -1362 2100 -1356
rect 2094 -1368 2100 -1362
rect 2094 -1374 2100 -1368
rect 2094 -1380 2100 -1374
rect 2094 -1386 2100 -1380
rect 2094 -1392 2100 -1386
rect 2094 -1398 2100 -1392
rect 2094 -1404 2100 -1398
rect 2094 -1410 2100 -1404
rect 2094 -1416 2100 -1410
rect 2094 -1422 2100 -1416
rect 2094 -1428 2100 -1422
rect 2094 -1434 2100 -1428
rect 2094 -1440 2100 -1434
rect 2094 -1446 2100 -1440
rect 2094 -1452 2100 -1446
rect 2094 -1458 2100 -1452
rect 2094 -1464 2100 -1458
rect 2094 -1470 2100 -1464
rect 2094 -1476 2100 -1470
rect 2094 -1482 2100 -1476
rect 2094 -1488 2100 -1482
rect 2094 -1494 2100 -1488
rect 2094 -1644 2100 -1638
rect 2094 -1650 2100 -1644
rect 2094 -1656 2100 -1650
rect 2094 -1662 2100 -1656
rect 2094 -1668 2100 -1662
rect 2094 -1674 2100 -1668
rect 2094 -1680 2100 -1674
rect 2094 -1686 2100 -1680
rect 2094 -1692 2100 -1686
rect 2094 -1698 2100 -1692
rect 2094 -1704 2100 -1698
rect 2094 -1710 2100 -1704
rect 2094 -1716 2100 -1710
rect 2094 -1722 2100 -1716
rect 2094 -1728 2100 -1722
rect 2094 -1734 2100 -1728
rect 2094 -1740 2100 -1734
rect 2094 -1746 2100 -1740
rect 2094 -1752 2100 -1746
rect 2094 -1758 2100 -1752
rect 2094 -1764 2100 -1758
rect 2094 -1770 2100 -1764
rect 2094 -1776 2100 -1770
rect 2094 -1782 2100 -1776
rect 2094 -1788 2100 -1782
rect 2094 -1794 2100 -1788
rect 2094 -1800 2100 -1794
rect 2094 -1806 2100 -1800
rect 2094 -1812 2100 -1806
rect 2094 -1818 2100 -1812
rect 2094 -1824 2100 -1818
rect 2094 -1830 2100 -1824
rect 2094 -1836 2100 -1830
rect 2094 -1842 2100 -1836
rect 2094 -1848 2100 -1842
rect 2094 -1854 2100 -1848
rect 2094 -1860 2100 -1854
rect 2094 -1866 2100 -1860
rect 2094 -1872 2100 -1866
rect 2094 -1878 2100 -1872
rect 2094 -1884 2100 -1878
rect 2094 -1890 2100 -1884
rect 2094 -1896 2100 -1890
rect 2094 -1902 2100 -1896
rect 2094 -1908 2100 -1902
rect 2094 -1914 2100 -1908
rect 2094 -1920 2100 -1914
rect 2094 -1926 2100 -1920
rect 2094 -1932 2100 -1926
rect 2094 -1938 2100 -1932
rect 2094 -1944 2100 -1938
rect 2094 -1950 2100 -1944
rect 2094 -1956 2100 -1950
rect 2094 -1962 2100 -1956
rect 2094 -1968 2100 -1962
rect 2094 -1974 2100 -1968
rect 2094 -1980 2100 -1974
rect 2094 -1986 2100 -1980
rect 2094 -1992 2100 -1986
rect 2094 -1998 2100 -1992
rect 2094 -2004 2100 -1998
rect 2094 -2010 2100 -2004
rect 2094 -2016 2100 -2010
rect 2094 -2022 2100 -2016
rect 2094 -2028 2100 -2022
rect 2094 -2034 2100 -2028
rect 2094 -2040 2100 -2034
rect 2094 -2046 2100 -2040
rect 2094 -2052 2100 -2046
rect 2094 -2058 2100 -2052
rect 2094 -2064 2100 -2058
rect 2094 -2070 2100 -2064
rect 2094 -2076 2100 -2070
rect 2094 -2082 2100 -2076
rect 2094 -2088 2100 -2082
rect 2094 -2094 2100 -2088
rect 2094 -2100 2100 -2094
rect 2094 -2106 2100 -2100
rect 2094 -2112 2100 -2106
rect 2094 -2118 2100 -2112
rect 2094 -2124 2100 -2118
rect 2094 -2130 2100 -2124
rect 2094 -2136 2100 -2130
rect 2094 -2142 2100 -2136
rect 2094 -2148 2100 -2142
rect 2094 -2154 2100 -2148
rect 2094 -2160 2100 -2154
rect 2094 -2166 2100 -2160
rect 2094 -2172 2100 -2166
rect 2094 -2178 2100 -2172
rect 2094 -2184 2100 -2178
rect 2094 -2190 2100 -2184
rect 2094 -2196 2100 -2190
rect 2094 -2202 2100 -2196
rect 2094 -2208 2100 -2202
rect 2094 -2214 2100 -2208
rect 2094 -2220 2100 -2214
rect 2094 -2226 2100 -2220
rect 2094 -2232 2100 -2226
rect 2094 -2238 2100 -2232
rect 2094 -2244 2100 -2238
rect 2094 -2250 2100 -2244
rect 2094 -2256 2100 -2250
rect 2094 -2262 2100 -2256
rect 2094 -2268 2100 -2262
rect 2094 -2274 2100 -2268
rect 2094 -2280 2100 -2274
rect 2094 -2286 2100 -2280
rect 2094 -2292 2100 -2286
rect 2094 -2298 2100 -2292
rect 2094 -2304 2100 -2298
rect 2094 -2310 2100 -2304
rect 2094 -2316 2100 -2310
rect 2094 -2322 2100 -2316
rect 2094 -2328 2100 -2322
rect 2094 -2334 2100 -2328
rect 2094 -2340 2100 -2334
rect 2094 -2346 2100 -2340
rect 2094 -2352 2100 -2346
rect 2094 -2358 2100 -2352
rect 2094 -2364 2100 -2358
rect 2094 -2370 2100 -2364
rect 2094 -2376 2100 -2370
rect 2094 -2382 2100 -2376
rect 2094 -2388 2100 -2382
rect 2094 -2394 2100 -2388
rect 2094 -2400 2100 -2394
rect 2094 -2406 2100 -2400
rect 2094 -2412 2100 -2406
rect 2094 -2418 2100 -2412
rect 2094 -2424 2100 -2418
rect 2094 -2430 2100 -2424
rect 2094 -2436 2100 -2430
rect 2094 -2442 2100 -2436
rect 2094 -2448 2100 -2442
rect 2094 -2454 2100 -2448
rect 2094 -2460 2100 -2454
rect 2094 -2466 2100 -2460
rect 2094 -2472 2100 -2466
rect 2094 -2574 2100 -2568
rect 2094 -2580 2100 -2574
rect 2094 -2586 2100 -2580
rect 2094 -2592 2100 -2586
rect 2094 -2598 2100 -2592
rect 2094 -2604 2100 -2598
rect 2094 -2610 2100 -2604
rect 2094 -2616 2100 -2610
rect 2094 -2622 2100 -2616
rect 2094 -2628 2100 -2622
rect 2094 -2634 2100 -2628
rect 2094 -2640 2100 -2634
rect 2094 -2646 2100 -2640
rect 2094 -2652 2100 -2646
rect 2094 -2658 2100 -2652
rect 2094 -2664 2100 -2658
rect 2094 -2670 2100 -2664
rect 2094 -2676 2100 -2670
rect 2094 -2682 2100 -2676
rect 2094 -2688 2100 -2682
rect 2094 -2694 2100 -2688
rect 2094 -2700 2100 -2694
rect 2094 -2706 2100 -2700
rect 2094 -2712 2100 -2706
rect 2094 -2718 2100 -2712
rect 2094 -2724 2100 -2718
rect 2094 -2730 2100 -2724
rect 2094 -2736 2100 -2730
rect 2094 -2742 2100 -2736
rect 2094 -2748 2100 -2742
rect 2094 -2754 2100 -2748
rect 2094 -2760 2100 -2754
rect 2094 -2766 2100 -2760
rect 2094 -2772 2100 -2766
rect 2094 -2778 2100 -2772
rect 2094 -2784 2100 -2778
rect 2094 -2790 2100 -2784
rect 2094 -2796 2100 -2790
rect 2094 -2802 2100 -2796
rect 2094 -2808 2100 -2802
rect 2094 -2814 2100 -2808
rect 2094 -2820 2100 -2814
rect 2094 -2826 2100 -2820
rect 2094 -2832 2100 -2826
rect 2094 -2838 2100 -2832
rect 2094 -2844 2100 -2838
rect 2094 -2850 2100 -2844
rect 2094 -2856 2100 -2850
rect 2094 -2862 2100 -2856
rect 2094 -2868 2100 -2862
rect 2094 -2874 2100 -2868
rect 2094 -2880 2100 -2874
rect 2094 -2886 2100 -2880
rect 2094 -2892 2100 -2886
rect 2094 -2898 2100 -2892
rect 2094 -2904 2100 -2898
rect 2094 -2910 2100 -2904
rect 2094 -2916 2100 -2910
rect 2094 -2922 2100 -2916
rect 2094 -2928 2100 -2922
rect 2094 -2934 2100 -2928
rect 2094 -2940 2100 -2934
rect 2094 -2946 2100 -2940
rect 2094 -2952 2100 -2946
rect 2094 -2958 2100 -2952
rect 2094 -2964 2100 -2958
rect 2094 -2970 2100 -2964
rect 2094 -2976 2100 -2970
rect 2094 -2982 2100 -2976
rect 2094 -2988 2100 -2982
rect 2094 -2994 2100 -2988
rect 2094 -3000 2100 -2994
rect 2094 -3006 2100 -3000
rect 2094 -3012 2100 -3006
rect 2094 -3018 2100 -3012
rect 2094 -3024 2100 -3018
rect 2094 -3030 2100 -3024
rect 2094 -3036 2100 -3030
rect 2094 -3042 2100 -3036
rect 2094 -3048 2100 -3042
rect 2094 -3054 2100 -3048
rect 2094 -3060 2100 -3054
rect 2094 -3066 2100 -3060
rect 2094 -3126 2100 -3120
rect 2094 -3132 2100 -3126
rect 2100 -324 2106 -318
rect 2100 -330 2106 -324
rect 2100 -336 2106 -330
rect 2100 -342 2106 -336
rect 2100 -348 2106 -342
rect 2100 -354 2106 -348
rect 2100 -360 2106 -354
rect 2100 -366 2106 -360
rect 2100 -372 2106 -366
rect 2100 -378 2106 -372
rect 2100 -384 2106 -378
rect 2100 -390 2106 -384
rect 2100 -396 2106 -390
rect 2100 -402 2106 -396
rect 2100 -408 2106 -402
rect 2100 -414 2106 -408
rect 2100 -420 2106 -414
rect 2100 -426 2106 -420
rect 2100 -432 2106 -426
rect 2100 -438 2106 -432
rect 2100 -444 2106 -438
rect 2100 -450 2106 -444
rect 2100 -456 2106 -450
rect 2100 -462 2106 -456
rect 2100 -468 2106 -462
rect 2100 -474 2106 -468
rect 2100 -480 2106 -474
rect 2100 -486 2106 -480
rect 2100 -492 2106 -486
rect 2100 -498 2106 -492
rect 2100 -504 2106 -498
rect 2100 -510 2106 -504
rect 2100 -516 2106 -510
rect 2100 -522 2106 -516
rect 2100 -528 2106 -522
rect 2100 -534 2106 -528
rect 2100 -540 2106 -534
rect 2100 -546 2106 -540
rect 2100 -552 2106 -546
rect 2100 -558 2106 -552
rect 2100 -564 2106 -558
rect 2100 -570 2106 -564
rect 2100 -576 2106 -570
rect 2100 -582 2106 -576
rect 2100 -588 2106 -582
rect 2100 -594 2106 -588
rect 2100 -600 2106 -594
rect 2100 -606 2106 -600
rect 2100 -612 2106 -606
rect 2100 -618 2106 -612
rect 2100 -624 2106 -618
rect 2100 -630 2106 -624
rect 2100 -636 2106 -630
rect 2100 -642 2106 -636
rect 2100 -648 2106 -642
rect 2100 -654 2106 -648
rect 2100 -660 2106 -654
rect 2100 -666 2106 -660
rect 2100 -672 2106 -666
rect 2100 -678 2106 -672
rect 2100 -684 2106 -678
rect 2100 -690 2106 -684
rect 2100 -696 2106 -690
rect 2100 -702 2106 -696
rect 2100 -708 2106 -702
rect 2100 -714 2106 -708
rect 2100 -720 2106 -714
rect 2100 -726 2106 -720
rect 2100 -732 2106 -726
rect 2100 -738 2106 -732
rect 2100 -744 2106 -738
rect 2100 -750 2106 -744
rect 2100 -756 2106 -750
rect 2100 -762 2106 -756
rect 2100 -768 2106 -762
rect 2100 -774 2106 -768
rect 2100 -780 2106 -774
rect 2100 -786 2106 -780
rect 2100 -792 2106 -786
rect 2100 -798 2106 -792
rect 2100 -804 2106 -798
rect 2100 -810 2106 -804
rect 2100 -816 2106 -810
rect 2100 -822 2106 -816
rect 2100 -828 2106 -822
rect 2100 -834 2106 -828
rect 2100 -840 2106 -834
rect 2100 -846 2106 -840
rect 2100 -852 2106 -846
rect 2100 -858 2106 -852
rect 2100 -864 2106 -858
rect 2100 -870 2106 -864
rect 2100 -876 2106 -870
rect 2100 -882 2106 -876
rect 2100 -888 2106 -882
rect 2100 -894 2106 -888
rect 2100 -900 2106 -894
rect 2100 -906 2106 -900
rect 2100 -912 2106 -906
rect 2100 -918 2106 -912
rect 2100 -924 2106 -918
rect 2100 -930 2106 -924
rect 2100 -936 2106 -930
rect 2100 -942 2106 -936
rect 2100 -948 2106 -942
rect 2100 -954 2106 -948
rect 2100 -960 2106 -954
rect 2100 -966 2106 -960
rect 2100 -972 2106 -966
rect 2100 -978 2106 -972
rect 2100 -984 2106 -978
rect 2100 -990 2106 -984
rect 2100 -996 2106 -990
rect 2100 -1002 2106 -996
rect 2100 -1008 2106 -1002
rect 2100 -1014 2106 -1008
rect 2100 -1020 2106 -1014
rect 2100 -1026 2106 -1020
rect 2100 -1032 2106 -1026
rect 2100 -1038 2106 -1032
rect 2100 -1044 2106 -1038
rect 2100 -1050 2106 -1044
rect 2100 -1056 2106 -1050
rect 2100 -1062 2106 -1056
rect 2100 -1068 2106 -1062
rect 2100 -1074 2106 -1068
rect 2100 -1080 2106 -1074
rect 2100 -1086 2106 -1080
rect 2100 -1092 2106 -1086
rect 2100 -1098 2106 -1092
rect 2100 -1104 2106 -1098
rect 2100 -1110 2106 -1104
rect 2100 -1116 2106 -1110
rect 2100 -1122 2106 -1116
rect 2100 -1128 2106 -1122
rect 2100 -1134 2106 -1128
rect 2100 -1140 2106 -1134
rect 2100 -1146 2106 -1140
rect 2100 -1152 2106 -1146
rect 2100 -1158 2106 -1152
rect 2100 -1164 2106 -1158
rect 2100 -1170 2106 -1164
rect 2100 -1176 2106 -1170
rect 2100 -1182 2106 -1176
rect 2100 -1188 2106 -1182
rect 2100 -1194 2106 -1188
rect 2100 -1200 2106 -1194
rect 2100 -1206 2106 -1200
rect 2100 -1212 2106 -1206
rect 2100 -1218 2106 -1212
rect 2100 -1224 2106 -1218
rect 2100 -1230 2106 -1224
rect 2100 -1236 2106 -1230
rect 2100 -1242 2106 -1236
rect 2100 -1248 2106 -1242
rect 2100 -1254 2106 -1248
rect 2100 -1260 2106 -1254
rect 2100 -1266 2106 -1260
rect 2100 -1272 2106 -1266
rect 2100 -1278 2106 -1272
rect 2100 -1284 2106 -1278
rect 2100 -1290 2106 -1284
rect 2100 -1296 2106 -1290
rect 2100 -1302 2106 -1296
rect 2100 -1308 2106 -1302
rect 2100 -1314 2106 -1308
rect 2100 -1320 2106 -1314
rect 2100 -1326 2106 -1320
rect 2100 -1332 2106 -1326
rect 2100 -1338 2106 -1332
rect 2100 -1344 2106 -1338
rect 2100 -1350 2106 -1344
rect 2100 -1356 2106 -1350
rect 2100 -1362 2106 -1356
rect 2100 -1368 2106 -1362
rect 2100 -1374 2106 -1368
rect 2100 -1380 2106 -1374
rect 2100 -1386 2106 -1380
rect 2100 -1392 2106 -1386
rect 2100 -1398 2106 -1392
rect 2100 -1404 2106 -1398
rect 2100 -1410 2106 -1404
rect 2100 -1416 2106 -1410
rect 2100 -1422 2106 -1416
rect 2100 -1428 2106 -1422
rect 2100 -1434 2106 -1428
rect 2100 -1440 2106 -1434
rect 2100 -1446 2106 -1440
rect 2100 -1452 2106 -1446
rect 2100 -1458 2106 -1452
rect 2100 -1464 2106 -1458
rect 2100 -1470 2106 -1464
rect 2100 -1476 2106 -1470
rect 2100 -1482 2106 -1476
rect 2100 -1644 2106 -1638
rect 2100 -1650 2106 -1644
rect 2100 -1656 2106 -1650
rect 2100 -1662 2106 -1656
rect 2100 -1668 2106 -1662
rect 2100 -1674 2106 -1668
rect 2100 -1680 2106 -1674
rect 2100 -1686 2106 -1680
rect 2100 -1692 2106 -1686
rect 2100 -1698 2106 -1692
rect 2100 -1704 2106 -1698
rect 2100 -1710 2106 -1704
rect 2100 -1716 2106 -1710
rect 2100 -1722 2106 -1716
rect 2100 -1728 2106 -1722
rect 2100 -1734 2106 -1728
rect 2100 -1740 2106 -1734
rect 2100 -1746 2106 -1740
rect 2100 -1752 2106 -1746
rect 2100 -1758 2106 -1752
rect 2100 -1764 2106 -1758
rect 2100 -1770 2106 -1764
rect 2100 -1776 2106 -1770
rect 2100 -1782 2106 -1776
rect 2100 -1788 2106 -1782
rect 2100 -1794 2106 -1788
rect 2100 -1800 2106 -1794
rect 2100 -1806 2106 -1800
rect 2100 -1812 2106 -1806
rect 2100 -1818 2106 -1812
rect 2100 -1824 2106 -1818
rect 2100 -1830 2106 -1824
rect 2100 -1836 2106 -1830
rect 2100 -1842 2106 -1836
rect 2100 -1848 2106 -1842
rect 2100 -1854 2106 -1848
rect 2100 -1860 2106 -1854
rect 2100 -1866 2106 -1860
rect 2100 -1872 2106 -1866
rect 2100 -1878 2106 -1872
rect 2100 -1884 2106 -1878
rect 2100 -1890 2106 -1884
rect 2100 -1896 2106 -1890
rect 2100 -1902 2106 -1896
rect 2100 -1908 2106 -1902
rect 2100 -1914 2106 -1908
rect 2100 -1920 2106 -1914
rect 2100 -1926 2106 -1920
rect 2100 -1932 2106 -1926
rect 2100 -1938 2106 -1932
rect 2100 -1944 2106 -1938
rect 2100 -1950 2106 -1944
rect 2100 -1956 2106 -1950
rect 2100 -1962 2106 -1956
rect 2100 -1968 2106 -1962
rect 2100 -1974 2106 -1968
rect 2100 -1980 2106 -1974
rect 2100 -1986 2106 -1980
rect 2100 -1992 2106 -1986
rect 2100 -1998 2106 -1992
rect 2100 -2004 2106 -1998
rect 2100 -2010 2106 -2004
rect 2100 -2016 2106 -2010
rect 2100 -2022 2106 -2016
rect 2100 -2028 2106 -2022
rect 2100 -2034 2106 -2028
rect 2100 -2040 2106 -2034
rect 2100 -2046 2106 -2040
rect 2100 -2052 2106 -2046
rect 2100 -2058 2106 -2052
rect 2100 -2064 2106 -2058
rect 2100 -2070 2106 -2064
rect 2100 -2076 2106 -2070
rect 2100 -2082 2106 -2076
rect 2100 -2088 2106 -2082
rect 2100 -2094 2106 -2088
rect 2100 -2100 2106 -2094
rect 2100 -2106 2106 -2100
rect 2100 -2112 2106 -2106
rect 2100 -2118 2106 -2112
rect 2100 -2124 2106 -2118
rect 2100 -2130 2106 -2124
rect 2100 -2136 2106 -2130
rect 2100 -2142 2106 -2136
rect 2100 -2148 2106 -2142
rect 2100 -2154 2106 -2148
rect 2100 -2160 2106 -2154
rect 2100 -2166 2106 -2160
rect 2100 -2172 2106 -2166
rect 2100 -2178 2106 -2172
rect 2100 -2184 2106 -2178
rect 2100 -2190 2106 -2184
rect 2100 -2196 2106 -2190
rect 2100 -2202 2106 -2196
rect 2100 -2208 2106 -2202
rect 2100 -2214 2106 -2208
rect 2100 -2220 2106 -2214
rect 2100 -2226 2106 -2220
rect 2100 -2232 2106 -2226
rect 2100 -2238 2106 -2232
rect 2100 -2244 2106 -2238
rect 2100 -2250 2106 -2244
rect 2100 -2256 2106 -2250
rect 2100 -2262 2106 -2256
rect 2100 -2268 2106 -2262
rect 2100 -2274 2106 -2268
rect 2100 -2280 2106 -2274
rect 2100 -2286 2106 -2280
rect 2100 -2292 2106 -2286
rect 2100 -2298 2106 -2292
rect 2100 -2304 2106 -2298
rect 2100 -2310 2106 -2304
rect 2100 -2316 2106 -2310
rect 2100 -2322 2106 -2316
rect 2100 -2328 2106 -2322
rect 2100 -2334 2106 -2328
rect 2100 -2340 2106 -2334
rect 2100 -2346 2106 -2340
rect 2100 -2352 2106 -2346
rect 2100 -2358 2106 -2352
rect 2100 -2364 2106 -2358
rect 2100 -2370 2106 -2364
rect 2100 -2376 2106 -2370
rect 2100 -2382 2106 -2376
rect 2100 -2388 2106 -2382
rect 2100 -2394 2106 -2388
rect 2100 -2400 2106 -2394
rect 2100 -2406 2106 -2400
rect 2100 -2412 2106 -2406
rect 2100 -2418 2106 -2412
rect 2100 -2424 2106 -2418
rect 2100 -2430 2106 -2424
rect 2100 -2436 2106 -2430
rect 2100 -2442 2106 -2436
rect 2100 -2448 2106 -2442
rect 2100 -2454 2106 -2448
rect 2100 -2460 2106 -2454
rect 2100 -2466 2106 -2460
rect 2100 -2574 2106 -2568
rect 2100 -2580 2106 -2574
rect 2100 -2586 2106 -2580
rect 2100 -2592 2106 -2586
rect 2100 -2598 2106 -2592
rect 2100 -2604 2106 -2598
rect 2100 -2610 2106 -2604
rect 2100 -2616 2106 -2610
rect 2100 -2622 2106 -2616
rect 2100 -2628 2106 -2622
rect 2100 -2634 2106 -2628
rect 2100 -2640 2106 -2634
rect 2100 -2646 2106 -2640
rect 2100 -2652 2106 -2646
rect 2100 -2658 2106 -2652
rect 2100 -2664 2106 -2658
rect 2100 -2670 2106 -2664
rect 2100 -2676 2106 -2670
rect 2100 -2682 2106 -2676
rect 2100 -2688 2106 -2682
rect 2100 -2694 2106 -2688
rect 2100 -2700 2106 -2694
rect 2100 -2706 2106 -2700
rect 2100 -2712 2106 -2706
rect 2100 -2718 2106 -2712
rect 2100 -2724 2106 -2718
rect 2100 -2730 2106 -2724
rect 2100 -2736 2106 -2730
rect 2100 -2742 2106 -2736
rect 2100 -2748 2106 -2742
rect 2100 -2754 2106 -2748
rect 2100 -2760 2106 -2754
rect 2100 -2766 2106 -2760
rect 2100 -2772 2106 -2766
rect 2100 -2778 2106 -2772
rect 2100 -2784 2106 -2778
rect 2100 -2790 2106 -2784
rect 2100 -2796 2106 -2790
rect 2100 -2802 2106 -2796
rect 2100 -2808 2106 -2802
rect 2100 -2814 2106 -2808
rect 2100 -2820 2106 -2814
rect 2100 -2826 2106 -2820
rect 2100 -2832 2106 -2826
rect 2100 -2838 2106 -2832
rect 2100 -2844 2106 -2838
rect 2100 -2850 2106 -2844
rect 2100 -2856 2106 -2850
rect 2100 -2862 2106 -2856
rect 2100 -2868 2106 -2862
rect 2100 -2874 2106 -2868
rect 2100 -2880 2106 -2874
rect 2100 -2886 2106 -2880
rect 2100 -2892 2106 -2886
rect 2100 -2898 2106 -2892
rect 2100 -2904 2106 -2898
rect 2100 -2910 2106 -2904
rect 2100 -2916 2106 -2910
rect 2100 -2922 2106 -2916
rect 2100 -2928 2106 -2922
rect 2100 -2934 2106 -2928
rect 2100 -2940 2106 -2934
rect 2100 -2946 2106 -2940
rect 2100 -2952 2106 -2946
rect 2100 -2958 2106 -2952
rect 2100 -2964 2106 -2958
rect 2100 -2970 2106 -2964
rect 2100 -2976 2106 -2970
rect 2100 -2982 2106 -2976
rect 2100 -2988 2106 -2982
rect 2100 -2994 2106 -2988
rect 2100 -3000 2106 -2994
rect 2100 -3006 2106 -3000
rect 2100 -3012 2106 -3006
rect 2100 -3018 2106 -3012
rect 2100 -3024 2106 -3018
rect 2100 -3030 2106 -3024
rect 2100 -3036 2106 -3030
rect 2100 -3042 2106 -3036
rect 2100 -3048 2106 -3042
rect 2100 -3054 2106 -3048
rect 2100 -3060 2106 -3054
rect 2100 -3066 2106 -3060
rect 2100 -3120 2106 -3114
rect 2100 -3126 2106 -3120
rect 2106 -318 2112 -312
rect 2106 -324 2112 -318
rect 2106 -330 2112 -324
rect 2106 -336 2112 -330
rect 2106 -342 2112 -336
rect 2106 -348 2112 -342
rect 2106 -354 2112 -348
rect 2106 -360 2112 -354
rect 2106 -366 2112 -360
rect 2106 -372 2112 -366
rect 2106 -378 2112 -372
rect 2106 -384 2112 -378
rect 2106 -390 2112 -384
rect 2106 -396 2112 -390
rect 2106 -402 2112 -396
rect 2106 -408 2112 -402
rect 2106 -414 2112 -408
rect 2106 -420 2112 -414
rect 2106 -426 2112 -420
rect 2106 -432 2112 -426
rect 2106 -438 2112 -432
rect 2106 -444 2112 -438
rect 2106 -450 2112 -444
rect 2106 -456 2112 -450
rect 2106 -462 2112 -456
rect 2106 -468 2112 -462
rect 2106 -474 2112 -468
rect 2106 -480 2112 -474
rect 2106 -486 2112 -480
rect 2106 -492 2112 -486
rect 2106 -498 2112 -492
rect 2106 -504 2112 -498
rect 2106 -510 2112 -504
rect 2106 -516 2112 -510
rect 2106 -522 2112 -516
rect 2106 -528 2112 -522
rect 2106 -534 2112 -528
rect 2106 -540 2112 -534
rect 2106 -546 2112 -540
rect 2106 -552 2112 -546
rect 2106 -558 2112 -552
rect 2106 -564 2112 -558
rect 2106 -570 2112 -564
rect 2106 -576 2112 -570
rect 2106 -582 2112 -576
rect 2106 -588 2112 -582
rect 2106 -594 2112 -588
rect 2106 -600 2112 -594
rect 2106 -606 2112 -600
rect 2106 -612 2112 -606
rect 2106 -618 2112 -612
rect 2106 -624 2112 -618
rect 2106 -630 2112 -624
rect 2106 -636 2112 -630
rect 2106 -642 2112 -636
rect 2106 -648 2112 -642
rect 2106 -654 2112 -648
rect 2106 -660 2112 -654
rect 2106 -666 2112 -660
rect 2106 -672 2112 -666
rect 2106 -678 2112 -672
rect 2106 -684 2112 -678
rect 2106 -690 2112 -684
rect 2106 -696 2112 -690
rect 2106 -702 2112 -696
rect 2106 -708 2112 -702
rect 2106 -714 2112 -708
rect 2106 -720 2112 -714
rect 2106 -726 2112 -720
rect 2106 -732 2112 -726
rect 2106 -738 2112 -732
rect 2106 -744 2112 -738
rect 2106 -750 2112 -744
rect 2106 -756 2112 -750
rect 2106 -762 2112 -756
rect 2106 -768 2112 -762
rect 2106 -774 2112 -768
rect 2106 -780 2112 -774
rect 2106 -786 2112 -780
rect 2106 -792 2112 -786
rect 2106 -798 2112 -792
rect 2106 -804 2112 -798
rect 2106 -810 2112 -804
rect 2106 -816 2112 -810
rect 2106 -822 2112 -816
rect 2106 -828 2112 -822
rect 2106 -834 2112 -828
rect 2106 -840 2112 -834
rect 2106 -846 2112 -840
rect 2106 -852 2112 -846
rect 2106 -858 2112 -852
rect 2106 -864 2112 -858
rect 2106 -870 2112 -864
rect 2106 -876 2112 -870
rect 2106 -882 2112 -876
rect 2106 -888 2112 -882
rect 2106 -894 2112 -888
rect 2106 -900 2112 -894
rect 2106 -906 2112 -900
rect 2106 -912 2112 -906
rect 2106 -918 2112 -912
rect 2106 -924 2112 -918
rect 2106 -930 2112 -924
rect 2106 -936 2112 -930
rect 2106 -942 2112 -936
rect 2106 -948 2112 -942
rect 2106 -954 2112 -948
rect 2106 -960 2112 -954
rect 2106 -966 2112 -960
rect 2106 -972 2112 -966
rect 2106 -978 2112 -972
rect 2106 -984 2112 -978
rect 2106 -990 2112 -984
rect 2106 -996 2112 -990
rect 2106 -1002 2112 -996
rect 2106 -1008 2112 -1002
rect 2106 -1014 2112 -1008
rect 2106 -1020 2112 -1014
rect 2106 -1026 2112 -1020
rect 2106 -1032 2112 -1026
rect 2106 -1038 2112 -1032
rect 2106 -1044 2112 -1038
rect 2106 -1050 2112 -1044
rect 2106 -1056 2112 -1050
rect 2106 -1062 2112 -1056
rect 2106 -1068 2112 -1062
rect 2106 -1074 2112 -1068
rect 2106 -1080 2112 -1074
rect 2106 -1086 2112 -1080
rect 2106 -1092 2112 -1086
rect 2106 -1098 2112 -1092
rect 2106 -1104 2112 -1098
rect 2106 -1110 2112 -1104
rect 2106 -1116 2112 -1110
rect 2106 -1122 2112 -1116
rect 2106 -1128 2112 -1122
rect 2106 -1134 2112 -1128
rect 2106 -1140 2112 -1134
rect 2106 -1146 2112 -1140
rect 2106 -1152 2112 -1146
rect 2106 -1158 2112 -1152
rect 2106 -1164 2112 -1158
rect 2106 -1170 2112 -1164
rect 2106 -1176 2112 -1170
rect 2106 -1182 2112 -1176
rect 2106 -1188 2112 -1182
rect 2106 -1194 2112 -1188
rect 2106 -1200 2112 -1194
rect 2106 -1206 2112 -1200
rect 2106 -1212 2112 -1206
rect 2106 -1218 2112 -1212
rect 2106 -1224 2112 -1218
rect 2106 -1230 2112 -1224
rect 2106 -1236 2112 -1230
rect 2106 -1242 2112 -1236
rect 2106 -1248 2112 -1242
rect 2106 -1254 2112 -1248
rect 2106 -1260 2112 -1254
rect 2106 -1266 2112 -1260
rect 2106 -1272 2112 -1266
rect 2106 -1278 2112 -1272
rect 2106 -1284 2112 -1278
rect 2106 -1290 2112 -1284
rect 2106 -1296 2112 -1290
rect 2106 -1302 2112 -1296
rect 2106 -1308 2112 -1302
rect 2106 -1314 2112 -1308
rect 2106 -1320 2112 -1314
rect 2106 -1326 2112 -1320
rect 2106 -1332 2112 -1326
rect 2106 -1338 2112 -1332
rect 2106 -1344 2112 -1338
rect 2106 -1350 2112 -1344
rect 2106 -1356 2112 -1350
rect 2106 -1362 2112 -1356
rect 2106 -1368 2112 -1362
rect 2106 -1374 2112 -1368
rect 2106 -1380 2112 -1374
rect 2106 -1386 2112 -1380
rect 2106 -1392 2112 -1386
rect 2106 -1398 2112 -1392
rect 2106 -1404 2112 -1398
rect 2106 -1410 2112 -1404
rect 2106 -1416 2112 -1410
rect 2106 -1422 2112 -1416
rect 2106 -1428 2112 -1422
rect 2106 -1434 2112 -1428
rect 2106 -1440 2112 -1434
rect 2106 -1446 2112 -1440
rect 2106 -1452 2112 -1446
rect 2106 -1458 2112 -1452
rect 2106 -1464 2112 -1458
rect 2106 -1470 2112 -1464
rect 2106 -1638 2112 -1632
rect 2106 -1644 2112 -1638
rect 2106 -1650 2112 -1644
rect 2106 -1656 2112 -1650
rect 2106 -1662 2112 -1656
rect 2106 -1668 2112 -1662
rect 2106 -1674 2112 -1668
rect 2106 -1680 2112 -1674
rect 2106 -1686 2112 -1680
rect 2106 -1692 2112 -1686
rect 2106 -1698 2112 -1692
rect 2106 -1704 2112 -1698
rect 2106 -1710 2112 -1704
rect 2106 -1716 2112 -1710
rect 2106 -1722 2112 -1716
rect 2106 -1728 2112 -1722
rect 2106 -1734 2112 -1728
rect 2106 -1740 2112 -1734
rect 2106 -1746 2112 -1740
rect 2106 -1752 2112 -1746
rect 2106 -1758 2112 -1752
rect 2106 -1764 2112 -1758
rect 2106 -1770 2112 -1764
rect 2106 -1776 2112 -1770
rect 2106 -1782 2112 -1776
rect 2106 -1788 2112 -1782
rect 2106 -1794 2112 -1788
rect 2106 -1800 2112 -1794
rect 2106 -1806 2112 -1800
rect 2106 -1812 2112 -1806
rect 2106 -1818 2112 -1812
rect 2106 -1824 2112 -1818
rect 2106 -1830 2112 -1824
rect 2106 -1836 2112 -1830
rect 2106 -1842 2112 -1836
rect 2106 -1848 2112 -1842
rect 2106 -1854 2112 -1848
rect 2106 -1860 2112 -1854
rect 2106 -1866 2112 -1860
rect 2106 -1872 2112 -1866
rect 2106 -1878 2112 -1872
rect 2106 -1884 2112 -1878
rect 2106 -1890 2112 -1884
rect 2106 -1896 2112 -1890
rect 2106 -1902 2112 -1896
rect 2106 -1908 2112 -1902
rect 2106 -1914 2112 -1908
rect 2106 -1920 2112 -1914
rect 2106 -1926 2112 -1920
rect 2106 -1932 2112 -1926
rect 2106 -1938 2112 -1932
rect 2106 -1944 2112 -1938
rect 2106 -1950 2112 -1944
rect 2106 -1956 2112 -1950
rect 2106 -1962 2112 -1956
rect 2106 -1968 2112 -1962
rect 2106 -1974 2112 -1968
rect 2106 -1980 2112 -1974
rect 2106 -1986 2112 -1980
rect 2106 -1992 2112 -1986
rect 2106 -1998 2112 -1992
rect 2106 -2004 2112 -1998
rect 2106 -2010 2112 -2004
rect 2106 -2016 2112 -2010
rect 2106 -2022 2112 -2016
rect 2106 -2028 2112 -2022
rect 2106 -2034 2112 -2028
rect 2106 -2040 2112 -2034
rect 2106 -2046 2112 -2040
rect 2106 -2052 2112 -2046
rect 2106 -2058 2112 -2052
rect 2106 -2064 2112 -2058
rect 2106 -2070 2112 -2064
rect 2106 -2076 2112 -2070
rect 2106 -2082 2112 -2076
rect 2106 -2088 2112 -2082
rect 2106 -2094 2112 -2088
rect 2106 -2100 2112 -2094
rect 2106 -2106 2112 -2100
rect 2106 -2112 2112 -2106
rect 2106 -2118 2112 -2112
rect 2106 -2124 2112 -2118
rect 2106 -2130 2112 -2124
rect 2106 -2136 2112 -2130
rect 2106 -2142 2112 -2136
rect 2106 -2148 2112 -2142
rect 2106 -2154 2112 -2148
rect 2106 -2160 2112 -2154
rect 2106 -2166 2112 -2160
rect 2106 -2172 2112 -2166
rect 2106 -2178 2112 -2172
rect 2106 -2184 2112 -2178
rect 2106 -2190 2112 -2184
rect 2106 -2196 2112 -2190
rect 2106 -2202 2112 -2196
rect 2106 -2208 2112 -2202
rect 2106 -2214 2112 -2208
rect 2106 -2220 2112 -2214
rect 2106 -2226 2112 -2220
rect 2106 -2232 2112 -2226
rect 2106 -2238 2112 -2232
rect 2106 -2244 2112 -2238
rect 2106 -2250 2112 -2244
rect 2106 -2256 2112 -2250
rect 2106 -2262 2112 -2256
rect 2106 -2268 2112 -2262
rect 2106 -2274 2112 -2268
rect 2106 -2280 2112 -2274
rect 2106 -2286 2112 -2280
rect 2106 -2292 2112 -2286
rect 2106 -2298 2112 -2292
rect 2106 -2304 2112 -2298
rect 2106 -2310 2112 -2304
rect 2106 -2316 2112 -2310
rect 2106 -2322 2112 -2316
rect 2106 -2328 2112 -2322
rect 2106 -2334 2112 -2328
rect 2106 -2340 2112 -2334
rect 2106 -2346 2112 -2340
rect 2106 -2352 2112 -2346
rect 2106 -2358 2112 -2352
rect 2106 -2364 2112 -2358
rect 2106 -2370 2112 -2364
rect 2106 -2376 2112 -2370
rect 2106 -2382 2112 -2376
rect 2106 -2388 2112 -2382
rect 2106 -2394 2112 -2388
rect 2106 -2400 2112 -2394
rect 2106 -2406 2112 -2400
rect 2106 -2412 2112 -2406
rect 2106 -2418 2112 -2412
rect 2106 -2424 2112 -2418
rect 2106 -2430 2112 -2424
rect 2106 -2436 2112 -2430
rect 2106 -2442 2112 -2436
rect 2106 -2448 2112 -2442
rect 2106 -2454 2112 -2448
rect 2106 -2460 2112 -2454
rect 2106 -2568 2112 -2562
rect 2106 -2574 2112 -2568
rect 2106 -2580 2112 -2574
rect 2106 -2586 2112 -2580
rect 2106 -2592 2112 -2586
rect 2106 -2598 2112 -2592
rect 2106 -2604 2112 -2598
rect 2106 -2610 2112 -2604
rect 2106 -2616 2112 -2610
rect 2106 -2622 2112 -2616
rect 2106 -2628 2112 -2622
rect 2106 -2634 2112 -2628
rect 2106 -2640 2112 -2634
rect 2106 -2646 2112 -2640
rect 2106 -2652 2112 -2646
rect 2106 -2658 2112 -2652
rect 2106 -2664 2112 -2658
rect 2106 -2670 2112 -2664
rect 2106 -2676 2112 -2670
rect 2106 -2682 2112 -2676
rect 2106 -2688 2112 -2682
rect 2106 -2694 2112 -2688
rect 2106 -2700 2112 -2694
rect 2106 -2706 2112 -2700
rect 2106 -2712 2112 -2706
rect 2106 -2718 2112 -2712
rect 2106 -2724 2112 -2718
rect 2106 -2730 2112 -2724
rect 2106 -2736 2112 -2730
rect 2106 -2742 2112 -2736
rect 2106 -2748 2112 -2742
rect 2106 -2754 2112 -2748
rect 2106 -2760 2112 -2754
rect 2106 -2766 2112 -2760
rect 2106 -2772 2112 -2766
rect 2106 -2778 2112 -2772
rect 2106 -2784 2112 -2778
rect 2106 -2790 2112 -2784
rect 2106 -2796 2112 -2790
rect 2106 -2802 2112 -2796
rect 2106 -2808 2112 -2802
rect 2106 -2814 2112 -2808
rect 2106 -2820 2112 -2814
rect 2106 -2826 2112 -2820
rect 2106 -2832 2112 -2826
rect 2106 -2838 2112 -2832
rect 2106 -2844 2112 -2838
rect 2106 -2850 2112 -2844
rect 2106 -2856 2112 -2850
rect 2106 -2862 2112 -2856
rect 2106 -2868 2112 -2862
rect 2106 -2874 2112 -2868
rect 2106 -2880 2112 -2874
rect 2106 -2886 2112 -2880
rect 2106 -2892 2112 -2886
rect 2106 -2898 2112 -2892
rect 2106 -2904 2112 -2898
rect 2106 -2910 2112 -2904
rect 2106 -2916 2112 -2910
rect 2106 -2922 2112 -2916
rect 2106 -2928 2112 -2922
rect 2106 -2934 2112 -2928
rect 2106 -2940 2112 -2934
rect 2106 -2946 2112 -2940
rect 2106 -2952 2112 -2946
rect 2106 -2958 2112 -2952
rect 2106 -2964 2112 -2958
rect 2106 -2970 2112 -2964
rect 2106 -2976 2112 -2970
rect 2106 -2982 2112 -2976
rect 2106 -2988 2112 -2982
rect 2106 -2994 2112 -2988
rect 2106 -3000 2112 -2994
rect 2106 -3006 2112 -3000
rect 2106 -3012 2112 -3006
rect 2106 -3018 2112 -3012
rect 2106 -3024 2112 -3018
rect 2106 -3030 2112 -3024
rect 2106 -3036 2112 -3030
rect 2106 -3042 2112 -3036
rect 2106 -3048 2112 -3042
rect 2106 -3054 2112 -3048
rect 2106 -3060 2112 -3054
rect 2106 -3120 2112 -3114
rect 2112 -306 2118 -300
rect 2112 -312 2118 -306
rect 2112 -318 2118 -312
rect 2112 -324 2118 -318
rect 2112 -330 2118 -324
rect 2112 -336 2118 -330
rect 2112 -342 2118 -336
rect 2112 -348 2118 -342
rect 2112 -354 2118 -348
rect 2112 -360 2118 -354
rect 2112 -366 2118 -360
rect 2112 -372 2118 -366
rect 2112 -378 2118 -372
rect 2112 -384 2118 -378
rect 2112 -390 2118 -384
rect 2112 -396 2118 -390
rect 2112 -402 2118 -396
rect 2112 -408 2118 -402
rect 2112 -414 2118 -408
rect 2112 -420 2118 -414
rect 2112 -426 2118 -420
rect 2112 -432 2118 -426
rect 2112 -438 2118 -432
rect 2112 -444 2118 -438
rect 2112 -450 2118 -444
rect 2112 -456 2118 -450
rect 2112 -462 2118 -456
rect 2112 -468 2118 -462
rect 2112 -474 2118 -468
rect 2112 -480 2118 -474
rect 2112 -486 2118 -480
rect 2112 -492 2118 -486
rect 2112 -498 2118 -492
rect 2112 -504 2118 -498
rect 2112 -510 2118 -504
rect 2112 -516 2118 -510
rect 2112 -522 2118 -516
rect 2112 -528 2118 -522
rect 2112 -534 2118 -528
rect 2112 -540 2118 -534
rect 2112 -546 2118 -540
rect 2112 -552 2118 -546
rect 2112 -558 2118 -552
rect 2112 -564 2118 -558
rect 2112 -570 2118 -564
rect 2112 -576 2118 -570
rect 2112 -582 2118 -576
rect 2112 -588 2118 -582
rect 2112 -594 2118 -588
rect 2112 -600 2118 -594
rect 2112 -606 2118 -600
rect 2112 -612 2118 -606
rect 2112 -618 2118 -612
rect 2112 -624 2118 -618
rect 2112 -630 2118 -624
rect 2112 -636 2118 -630
rect 2112 -642 2118 -636
rect 2112 -648 2118 -642
rect 2112 -654 2118 -648
rect 2112 -660 2118 -654
rect 2112 -666 2118 -660
rect 2112 -672 2118 -666
rect 2112 -678 2118 -672
rect 2112 -684 2118 -678
rect 2112 -690 2118 -684
rect 2112 -696 2118 -690
rect 2112 -702 2118 -696
rect 2112 -708 2118 -702
rect 2112 -714 2118 -708
rect 2112 -720 2118 -714
rect 2112 -726 2118 -720
rect 2112 -732 2118 -726
rect 2112 -738 2118 -732
rect 2112 -744 2118 -738
rect 2112 -750 2118 -744
rect 2112 -756 2118 -750
rect 2112 -762 2118 -756
rect 2112 -768 2118 -762
rect 2112 -774 2118 -768
rect 2112 -780 2118 -774
rect 2112 -786 2118 -780
rect 2112 -792 2118 -786
rect 2112 -798 2118 -792
rect 2112 -804 2118 -798
rect 2112 -810 2118 -804
rect 2112 -816 2118 -810
rect 2112 -822 2118 -816
rect 2112 -828 2118 -822
rect 2112 -834 2118 -828
rect 2112 -840 2118 -834
rect 2112 -846 2118 -840
rect 2112 -852 2118 -846
rect 2112 -858 2118 -852
rect 2112 -864 2118 -858
rect 2112 -870 2118 -864
rect 2112 -876 2118 -870
rect 2112 -882 2118 -876
rect 2112 -888 2118 -882
rect 2112 -894 2118 -888
rect 2112 -900 2118 -894
rect 2112 -906 2118 -900
rect 2112 -912 2118 -906
rect 2112 -918 2118 -912
rect 2112 -924 2118 -918
rect 2112 -930 2118 -924
rect 2112 -936 2118 -930
rect 2112 -942 2118 -936
rect 2112 -948 2118 -942
rect 2112 -954 2118 -948
rect 2112 -960 2118 -954
rect 2112 -966 2118 -960
rect 2112 -972 2118 -966
rect 2112 -978 2118 -972
rect 2112 -984 2118 -978
rect 2112 -990 2118 -984
rect 2112 -996 2118 -990
rect 2112 -1002 2118 -996
rect 2112 -1008 2118 -1002
rect 2112 -1014 2118 -1008
rect 2112 -1020 2118 -1014
rect 2112 -1026 2118 -1020
rect 2112 -1032 2118 -1026
rect 2112 -1038 2118 -1032
rect 2112 -1044 2118 -1038
rect 2112 -1050 2118 -1044
rect 2112 -1056 2118 -1050
rect 2112 -1062 2118 -1056
rect 2112 -1068 2118 -1062
rect 2112 -1074 2118 -1068
rect 2112 -1080 2118 -1074
rect 2112 -1086 2118 -1080
rect 2112 -1092 2118 -1086
rect 2112 -1098 2118 -1092
rect 2112 -1104 2118 -1098
rect 2112 -1110 2118 -1104
rect 2112 -1116 2118 -1110
rect 2112 -1122 2118 -1116
rect 2112 -1128 2118 -1122
rect 2112 -1134 2118 -1128
rect 2112 -1140 2118 -1134
rect 2112 -1146 2118 -1140
rect 2112 -1152 2118 -1146
rect 2112 -1158 2118 -1152
rect 2112 -1164 2118 -1158
rect 2112 -1170 2118 -1164
rect 2112 -1176 2118 -1170
rect 2112 -1182 2118 -1176
rect 2112 -1188 2118 -1182
rect 2112 -1194 2118 -1188
rect 2112 -1200 2118 -1194
rect 2112 -1206 2118 -1200
rect 2112 -1212 2118 -1206
rect 2112 -1218 2118 -1212
rect 2112 -1224 2118 -1218
rect 2112 -1230 2118 -1224
rect 2112 -1236 2118 -1230
rect 2112 -1242 2118 -1236
rect 2112 -1248 2118 -1242
rect 2112 -1254 2118 -1248
rect 2112 -1260 2118 -1254
rect 2112 -1266 2118 -1260
rect 2112 -1272 2118 -1266
rect 2112 -1278 2118 -1272
rect 2112 -1284 2118 -1278
rect 2112 -1290 2118 -1284
rect 2112 -1296 2118 -1290
rect 2112 -1302 2118 -1296
rect 2112 -1308 2118 -1302
rect 2112 -1314 2118 -1308
rect 2112 -1320 2118 -1314
rect 2112 -1326 2118 -1320
rect 2112 -1332 2118 -1326
rect 2112 -1338 2118 -1332
rect 2112 -1344 2118 -1338
rect 2112 -1350 2118 -1344
rect 2112 -1356 2118 -1350
rect 2112 -1362 2118 -1356
rect 2112 -1368 2118 -1362
rect 2112 -1374 2118 -1368
rect 2112 -1380 2118 -1374
rect 2112 -1386 2118 -1380
rect 2112 -1392 2118 -1386
rect 2112 -1398 2118 -1392
rect 2112 -1404 2118 -1398
rect 2112 -1410 2118 -1404
rect 2112 -1416 2118 -1410
rect 2112 -1422 2118 -1416
rect 2112 -1428 2118 -1422
rect 2112 -1434 2118 -1428
rect 2112 -1440 2118 -1434
rect 2112 -1446 2118 -1440
rect 2112 -1452 2118 -1446
rect 2112 -1632 2118 -1626
rect 2112 -1638 2118 -1632
rect 2112 -1644 2118 -1638
rect 2112 -1650 2118 -1644
rect 2112 -1656 2118 -1650
rect 2112 -1662 2118 -1656
rect 2112 -1668 2118 -1662
rect 2112 -1674 2118 -1668
rect 2112 -1680 2118 -1674
rect 2112 -1686 2118 -1680
rect 2112 -1692 2118 -1686
rect 2112 -1698 2118 -1692
rect 2112 -1704 2118 -1698
rect 2112 -1710 2118 -1704
rect 2112 -1716 2118 -1710
rect 2112 -1722 2118 -1716
rect 2112 -1728 2118 -1722
rect 2112 -1734 2118 -1728
rect 2112 -1740 2118 -1734
rect 2112 -1746 2118 -1740
rect 2112 -1752 2118 -1746
rect 2112 -1758 2118 -1752
rect 2112 -1764 2118 -1758
rect 2112 -1770 2118 -1764
rect 2112 -1776 2118 -1770
rect 2112 -1782 2118 -1776
rect 2112 -1788 2118 -1782
rect 2112 -1794 2118 -1788
rect 2112 -1800 2118 -1794
rect 2112 -1806 2118 -1800
rect 2112 -1812 2118 -1806
rect 2112 -1818 2118 -1812
rect 2112 -1824 2118 -1818
rect 2112 -1830 2118 -1824
rect 2112 -1836 2118 -1830
rect 2112 -1842 2118 -1836
rect 2112 -1848 2118 -1842
rect 2112 -1854 2118 -1848
rect 2112 -1860 2118 -1854
rect 2112 -1866 2118 -1860
rect 2112 -1872 2118 -1866
rect 2112 -1878 2118 -1872
rect 2112 -1884 2118 -1878
rect 2112 -1890 2118 -1884
rect 2112 -1896 2118 -1890
rect 2112 -1902 2118 -1896
rect 2112 -1908 2118 -1902
rect 2112 -1914 2118 -1908
rect 2112 -1920 2118 -1914
rect 2112 -1926 2118 -1920
rect 2112 -1932 2118 -1926
rect 2112 -1938 2118 -1932
rect 2112 -1944 2118 -1938
rect 2112 -1950 2118 -1944
rect 2112 -1956 2118 -1950
rect 2112 -1962 2118 -1956
rect 2112 -1968 2118 -1962
rect 2112 -1974 2118 -1968
rect 2112 -1980 2118 -1974
rect 2112 -1986 2118 -1980
rect 2112 -1992 2118 -1986
rect 2112 -1998 2118 -1992
rect 2112 -2004 2118 -1998
rect 2112 -2010 2118 -2004
rect 2112 -2016 2118 -2010
rect 2112 -2022 2118 -2016
rect 2112 -2028 2118 -2022
rect 2112 -2034 2118 -2028
rect 2112 -2040 2118 -2034
rect 2112 -2046 2118 -2040
rect 2112 -2052 2118 -2046
rect 2112 -2058 2118 -2052
rect 2112 -2064 2118 -2058
rect 2112 -2070 2118 -2064
rect 2112 -2076 2118 -2070
rect 2112 -2082 2118 -2076
rect 2112 -2088 2118 -2082
rect 2112 -2094 2118 -2088
rect 2112 -2100 2118 -2094
rect 2112 -2106 2118 -2100
rect 2112 -2112 2118 -2106
rect 2112 -2118 2118 -2112
rect 2112 -2124 2118 -2118
rect 2112 -2130 2118 -2124
rect 2112 -2136 2118 -2130
rect 2112 -2142 2118 -2136
rect 2112 -2148 2118 -2142
rect 2112 -2154 2118 -2148
rect 2112 -2160 2118 -2154
rect 2112 -2166 2118 -2160
rect 2112 -2172 2118 -2166
rect 2112 -2178 2118 -2172
rect 2112 -2184 2118 -2178
rect 2112 -2190 2118 -2184
rect 2112 -2196 2118 -2190
rect 2112 -2202 2118 -2196
rect 2112 -2208 2118 -2202
rect 2112 -2214 2118 -2208
rect 2112 -2220 2118 -2214
rect 2112 -2226 2118 -2220
rect 2112 -2232 2118 -2226
rect 2112 -2238 2118 -2232
rect 2112 -2244 2118 -2238
rect 2112 -2250 2118 -2244
rect 2112 -2256 2118 -2250
rect 2112 -2262 2118 -2256
rect 2112 -2268 2118 -2262
rect 2112 -2274 2118 -2268
rect 2112 -2280 2118 -2274
rect 2112 -2286 2118 -2280
rect 2112 -2292 2118 -2286
rect 2112 -2298 2118 -2292
rect 2112 -2304 2118 -2298
rect 2112 -2310 2118 -2304
rect 2112 -2316 2118 -2310
rect 2112 -2322 2118 -2316
rect 2112 -2328 2118 -2322
rect 2112 -2334 2118 -2328
rect 2112 -2340 2118 -2334
rect 2112 -2346 2118 -2340
rect 2112 -2352 2118 -2346
rect 2112 -2358 2118 -2352
rect 2112 -2364 2118 -2358
rect 2112 -2370 2118 -2364
rect 2112 -2376 2118 -2370
rect 2112 -2382 2118 -2376
rect 2112 -2388 2118 -2382
rect 2112 -2394 2118 -2388
rect 2112 -2400 2118 -2394
rect 2112 -2406 2118 -2400
rect 2112 -2412 2118 -2406
rect 2112 -2418 2118 -2412
rect 2112 -2424 2118 -2418
rect 2112 -2430 2118 -2424
rect 2112 -2436 2118 -2430
rect 2112 -2442 2118 -2436
rect 2112 -2448 2118 -2442
rect 2112 -2568 2118 -2562
rect 2112 -2574 2118 -2568
rect 2112 -2580 2118 -2574
rect 2112 -2586 2118 -2580
rect 2112 -2592 2118 -2586
rect 2112 -2598 2118 -2592
rect 2112 -2604 2118 -2598
rect 2112 -2610 2118 -2604
rect 2112 -2616 2118 -2610
rect 2112 -2622 2118 -2616
rect 2112 -2628 2118 -2622
rect 2112 -2634 2118 -2628
rect 2112 -2640 2118 -2634
rect 2112 -2646 2118 -2640
rect 2112 -2652 2118 -2646
rect 2112 -2658 2118 -2652
rect 2112 -2664 2118 -2658
rect 2112 -2670 2118 -2664
rect 2112 -2676 2118 -2670
rect 2112 -2682 2118 -2676
rect 2112 -2688 2118 -2682
rect 2112 -2694 2118 -2688
rect 2112 -2700 2118 -2694
rect 2112 -2706 2118 -2700
rect 2112 -2712 2118 -2706
rect 2112 -2718 2118 -2712
rect 2112 -2724 2118 -2718
rect 2112 -2730 2118 -2724
rect 2112 -2736 2118 -2730
rect 2112 -2742 2118 -2736
rect 2112 -2748 2118 -2742
rect 2112 -2754 2118 -2748
rect 2112 -2760 2118 -2754
rect 2112 -2766 2118 -2760
rect 2112 -2772 2118 -2766
rect 2112 -2778 2118 -2772
rect 2112 -2784 2118 -2778
rect 2112 -2790 2118 -2784
rect 2112 -2796 2118 -2790
rect 2112 -2802 2118 -2796
rect 2112 -2808 2118 -2802
rect 2112 -2814 2118 -2808
rect 2112 -2820 2118 -2814
rect 2112 -2826 2118 -2820
rect 2112 -2832 2118 -2826
rect 2112 -2838 2118 -2832
rect 2112 -2844 2118 -2838
rect 2112 -2850 2118 -2844
rect 2112 -2856 2118 -2850
rect 2112 -2862 2118 -2856
rect 2112 -2868 2118 -2862
rect 2112 -2874 2118 -2868
rect 2112 -2880 2118 -2874
rect 2112 -2886 2118 -2880
rect 2112 -2892 2118 -2886
rect 2112 -2898 2118 -2892
rect 2112 -2904 2118 -2898
rect 2112 -2910 2118 -2904
rect 2112 -2916 2118 -2910
rect 2112 -2922 2118 -2916
rect 2112 -2928 2118 -2922
rect 2112 -2934 2118 -2928
rect 2112 -2940 2118 -2934
rect 2112 -2946 2118 -2940
rect 2112 -2952 2118 -2946
rect 2112 -2958 2118 -2952
rect 2112 -2964 2118 -2958
rect 2112 -2970 2118 -2964
rect 2112 -2976 2118 -2970
rect 2112 -2982 2118 -2976
rect 2112 -2988 2118 -2982
rect 2112 -2994 2118 -2988
rect 2112 -3000 2118 -2994
rect 2112 -3006 2118 -3000
rect 2112 -3012 2118 -3006
rect 2112 -3018 2118 -3012
rect 2112 -3024 2118 -3018
rect 2112 -3030 2118 -3024
rect 2112 -3036 2118 -3030
rect 2112 -3042 2118 -3036
rect 2112 -3048 2118 -3042
rect 2112 -3054 2118 -3048
rect 2112 -3060 2118 -3054
rect 2118 -300 2124 -294
rect 2118 -306 2124 -300
rect 2118 -312 2124 -306
rect 2118 -318 2124 -312
rect 2118 -324 2124 -318
rect 2118 -330 2124 -324
rect 2118 -336 2124 -330
rect 2118 -342 2124 -336
rect 2118 -348 2124 -342
rect 2118 -354 2124 -348
rect 2118 -360 2124 -354
rect 2118 -366 2124 -360
rect 2118 -372 2124 -366
rect 2118 -378 2124 -372
rect 2118 -384 2124 -378
rect 2118 -390 2124 -384
rect 2118 -396 2124 -390
rect 2118 -402 2124 -396
rect 2118 -408 2124 -402
rect 2118 -414 2124 -408
rect 2118 -420 2124 -414
rect 2118 -426 2124 -420
rect 2118 -432 2124 -426
rect 2118 -438 2124 -432
rect 2118 -444 2124 -438
rect 2118 -450 2124 -444
rect 2118 -456 2124 -450
rect 2118 -462 2124 -456
rect 2118 -468 2124 -462
rect 2118 -474 2124 -468
rect 2118 -480 2124 -474
rect 2118 -486 2124 -480
rect 2118 -492 2124 -486
rect 2118 -498 2124 -492
rect 2118 -504 2124 -498
rect 2118 -510 2124 -504
rect 2118 -516 2124 -510
rect 2118 -522 2124 -516
rect 2118 -528 2124 -522
rect 2118 -534 2124 -528
rect 2118 -540 2124 -534
rect 2118 -546 2124 -540
rect 2118 -552 2124 -546
rect 2118 -558 2124 -552
rect 2118 -564 2124 -558
rect 2118 -570 2124 -564
rect 2118 -576 2124 -570
rect 2118 -582 2124 -576
rect 2118 -588 2124 -582
rect 2118 -594 2124 -588
rect 2118 -600 2124 -594
rect 2118 -606 2124 -600
rect 2118 -612 2124 -606
rect 2118 -618 2124 -612
rect 2118 -624 2124 -618
rect 2118 -630 2124 -624
rect 2118 -636 2124 -630
rect 2118 -642 2124 -636
rect 2118 -648 2124 -642
rect 2118 -654 2124 -648
rect 2118 -660 2124 -654
rect 2118 -666 2124 -660
rect 2118 -672 2124 -666
rect 2118 -678 2124 -672
rect 2118 -684 2124 -678
rect 2118 -690 2124 -684
rect 2118 -696 2124 -690
rect 2118 -702 2124 -696
rect 2118 -708 2124 -702
rect 2118 -714 2124 -708
rect 2118 -720 2124 -714
rect 2118 -726 2124 -720
rect 2118 -732 2124 -726
rect 2118 -738 2124 -732
rect 2118 -744 2124 -738
rect 2118 -750 2124 -744
rect 2118 -756 2124 -750
rect 2118 -762 2124 -756
rect 2118 -768 2124 -762
rect 2118 -774 2124 -768
rect 2118 -780 2124 -774
rect 2118 -786 2124 -780
rect 2118 -792 2124 -786
rect 2118 -798 2124 -792
rect 2118 -804 2124 -798
rect 2118 -810 2124 -804
rect 2118 -816 2124 -810
rect 2118 -822 2124 -816
rect 2118 -828 2124 -822
rect 2118 -834 2124 -828
rect 2118 -840 2124 -834
rect 2118 -846 2124 -840
rect 2118 -852 2124 -846
rect 2118 -858 2124 -852
rect 2118 -864 2124 -858
rect 2118 -870 2124 -864
rect 2118 -876 2124 -870
rect 2118 -882 2124 -876
rect 2118 -888 2124 -882
rect 2118 -894 2124 -888
rect 2118 -900 2124 -894
rect 2118 -906 2124 -900
rect 2118 -912 2124 -906
rect 2118 -918 2124 -912
rect 2118 -924 2124 -918
rect 2118 -930 2124 -924
rect 2118 -936 2124 -930
rect 2118 -942 2124 -936
rect 2118 -948 2124 -942
rect 2118 -954 2124 -948
rect 2118 -960 2124 -954
rect 2118 -966 2124 -960
rect 2118 -972 2124 -966
rect 2118 -978 2124 -972
rect 2118 -984 2124 -978
rect 2118 -990 2124 -984
rect 2118 -996 2124 -990
rect 2118 -1002 2124 -996
rect 2118 -1008 2124 -1002
rect 2118 -1014 2124 -1008
rect 2118 -1020 2124 -1014
rect 2118 -1026 2124 -1020
rect 2118 -1032 2124 -1026
rect 2118 -1038 2124 -1032
rect 2118 -1044 2124 -1038
rect 2118 -1050 2124 -1044
rect 2118 -1056 2124 -1050
rect 2118 -1062 2124 -1056
rect 2118 -1068 2124 -1062
rect 2118 -1074 2124 -1068
rect 2118 -1080 2124 -1074
rect 2118 -1086 2124 -1080
rect 2118 -1092 2124 -1086
rect 2118 -1098 2124 -1092
rect 2118 -1104 2124 -1098
rect 2118 -1110 2124 -1104
rect 2118 -1116 2124 -1110
rect 2118 -1122 2124 -1116
rect 2118 -1128 2124 -1122
rect 2118 -1134 2124 -1128
rect 2118 -1140 2124 -1134
rect 2118 -1146 2124 -1140
rect 2118 -1152 2124 -1146
rect 2118 -1158 2124 -1152
rect 2118 -1164 2124 -1158
rect 2118 -1170 2124 -1164
rect 2118 -1176 2124 -1170
rect 2118 -1182 2124 -1176
rect 2118 -1188 2124 -1182
rect 2118 -1194 2124 -1188
rect 2118 -1200 2124 -1194
rect 2118 -1206 2124 -1200
rect 2118 -1212 2124 -1206
rect 2118 -1218 2124 -1212
rect 2118 -1224 2124 -1218
rect 2118 -1230 2124 -1224
rect 2118 -1236 2124 -1230
rect 2118 -1242 2124 -1236
rect 2118 -1248 2124 -1242
rect 2118 -1254 2124 -1248
rect 2118 -1260 2124 -1254
rect 2118 -1266 2124 -1260
rect 2118 -1272 2124 -1266
rect 2118 -1278 2124 -1272
rect 2118 -1284 2124 -1278
rect 2118 -1290 2124 -1284
rect 2118 -1296 2124 -1290
rect 2118 -1302 2124 -1296
rect 2118 -1308 2124 -1302
rect 2118 -1314 2124 -1308
rect 2118 -1320 2124 -1314
rect 2118 -1326 2124 -1320
rect 2118 -1332 2124 -1326
rect 2118 -1338 2124 -1332
rect 2118 -1344 2124 -1338
rect 2118 -1350 2124 -1344
rect 2118 -1356 2124 -1350
rect 2118 -1362 2124 -1356
rect 2118 -1368 2124 -1362
rect 2118 -1374 2124 -1368
rect 2118 -1380 2124 -1374
rect 2118 -1386 2124 -1380
rect 2118 -1392 2124 -1386
rect 2118 -1398 2124 -1392
rect 2118 -1404 2124 -1398
rect 2118 -1410 2124 -1404
rect 2118 -1416 2124 -1410
rect 2118 -1422 2124 -1416
rect 2118 -1428 2124 -1422
rect 2118 -1434 2124 -1428
rect 2118 -1440 2124 -1434
rect 2118 -1626 2124 -1620
rect 2118 -1632 2124 -1626
rect 2118 -1638 2124 -1632
rect 2118 -1644 2124 -1638
rect 2118 -1650 2124 -1644
rect 2118 -1656 2124 -1650
rect 2118 -1662 2124 -1656
rect 2118 -1668 2124 -1662
rect 2118 -1674 2124 -1668
rect 2118 -1680 2124 -1674
rect 2118 -1686 2124 -1680
rect 2118 -1692 2124 -1686
rect 2118 -1698 2124 -1692
rect 2118 -1704 2124 -1698
rect 2118 -1710 2124 -1704
rect 2118 -1716 2124 -1710
rect 2118 -1722 2124 -1716
rect 2118 -1728 2124 -1722
rect 2118 -1734 2124 -1728
rect 2118 -1740 2124 -1734
rect 2118 -1746 2124 -1740
rect 2118 -1752 2124 -1746
rect 2118 -1758 2124 -1752
rect 2118 -1764 2124 -1758
rect 2118 -1770 2124 -1764
rect 2118 -1776 2124 -1770
rect 2118 -1782 2124 -1776
rect 2118 -1788 2124 -1782
rect 2118 -1794 2124 -1788
rect 2118 -1800 2124 -1794
rect 2118 -1806 2124 -1800
rect 2118 -1812 2124 -1806
rect 2118 -1818 2124 -1812
rect 2118 -1824 2124 -1818
rect 2118 -1830 2124 -1824
rect 2118 -1836 2124 -1830
rect 2118 -1842 2124 -1836
rect 2118 -1848 2124 -1842
rect 2118 -1854 2124 -1848
rect 2118 -1860 2124 -1854
rect 2118 -1866 2124 -1860
rect 2118 -1872 2124 -1866
rect 2118 -1878 2124 -1872
rect 2118 -1884 2124 -1878
rect 2118 -1890 2124 -1884
rect 2118 -1896 2124 -1890
rect 2118 -1902 2124 -1896
rect 2118 -1908 2124 -1902
rect 2118 -1914 2124 -1908
rect 2118 -1920 2124 -1914
rect 2118 -1926 2124 -1920
rect 2118 -1932 2124 -1926
rect 2118 -1938 2124 -1932
rect 2118 -1944 2124 -1938
rect 2118 -1950 2124 -1944
rect 2118 -1956 2124 -1950
rect 2118 -1962 2124 -1956
rect 2118 -1968 2124 -1962
rect 2118 -1974 2124 -1968
rect 2118 -1980 2124 -1974
rect 2118 -1986 2124 -1980
rect 2118 -1992 2124 -1986
rect 2118 -1998 2124 -1992
rect 2118 -2004 2124 -1998
rect 2118 -2010 2124 -2004
rect 2118 -2016 2124 -2010
rect 2118 -2022 2124 -2016
rect 2118 -2028 2124 -2022
rect 2118 -2034 2124 -2028
rect 2118 -2040 2124 -2034
rect 2118 -2046 2124 -2040
rect 2118 -2052 2124 -2046
rect 2118 -2058 2124 -2052
rect 2118 -2064 2124 -2058
rect 2118 -2070 2124 -2064
rect 2118 -2076 2124 -2070
rect 2118 -2082 2124 -2076
rect 2118 -2088 2124 -2082
rect 2118 -2094 2124 -2088
rect 2118 -2100 2124 -2094
rect 2118 -2106 2124 -2100
rect 2118 -2112 2124 -2106
rect 2118 -2118 2124 -2112
rect 2118 -2124 2124 -2118
rect 2118 -2130 2124 -2124
rect 2118 -2136 2124 -2130
rect 2118 -2142 2124 -2136
rect 2118 -2148 2124 -2142
rect 2118 -2154 2124 -2148
rect 2118 -2160 2124 -2154
rect 2118 -2166 2124 -2160
rect 2118 -2172 2124 -2166
rect 2118 -2178 2124 -2172
rect 2118 -2184 2124 -2178
rect 2118 -2190 2124 -2184
rect 2118 -2196 2124 -2190
rect 2118 -2202 2124 -2196
rect 2118 -2208 2124 -2202
rect 2118 -2214 2124 -2208
rect 2118 -2220 2124 -2214
rect 2118 -2226 2124 -2220
rect 2118 -2232 2124 -2226
rect 2118 -2238 2124 -2232
rect 2118 -2244 2124 -2238
rect 2118 -2250 2124 -2244
rect 2118 -2256 2124 -2250
rect 2118 -2262 2124 -2256
rect 2118 -2268 2124 -2262
rect 2118 -2274 2124 -2268
rect 2118 -2280 2124 -2274
rect 2118 -2286 2124 -2280
rect 2118 -2292 2124 -2286
rect 2118 -2298 2124 -2292
rect 2118 -2304 2124 -2298
rect 2118 -2310 2124 -2304
rect 2118 -2316 2124 -2310
rect 2118 -2322 2124 -2316
rect 2118 -2328 2124 -2322
rect 2118 -2334 2124 -2328
rect 2118 -2340 2124 -2334
rect 2118 -2346 2124 -2340
rect 2118 -2352 2124 -2346
rect 2118 -2358 2124 -2352
rect 2118 -2364 2124 -2358
rect 2118 -2370 2124 -2364
rect 2118 -2376 2124 -2370
rect 2118 -2382 2124 -2376
rect 2118 -2388 2124 -2382
rect 2118 -2394 2124 -2388
rect 2118 -2400 2124 -2394
rect 2118 -2406 2124 -2400
rect 2118 -2412 2124 -2406
rect 2118 -2418 2124 -2412
rect 2118 -2424 2124 -2418
rect 2118 -2430 2124 -2424
rect 2118 -2436 2124 -2430
rect 2118 -2442 2124 -2436
rect 2118 -2568 2124 -2562
rect 2118 -2574 2124 -2568
rect 2118 -2580 2124 -2574
rect 2118 -2586 2124 -2580
rect 2118 -2592 2124 -2586
rect 2118 -2598 2124 -2592
rect 2118 -2604 2124 -2598
rect 2118 -2610 2124 -2604
rect 2118 -2616 2124 -2610
rect 2118 -2622 2124 -2616
rect 2118 -2628 2124 -2622
rect 2118 -2634 2124 -2628
rect 2118 -2640 2124 -2634
rect 2118 -2646 2124 -2640
rect 2118 -2652 2124 -2646
rect 2118 -2658 2124 -2652
rect 2118 -2664 2124 -2658
rect 2118 -2670 2124 -2664
rect 2118 -2676 2124 -2670
rect 2118 -2682 2124 -2676
rect 2118 -2688 2124 -2682
rect 2118 -2694 2124 -2688
rect 2118 -2700 2124 -2694
rect 2118 -2706 2124 -2700
rect 2118 -2712 2124 -2706
rect 2118 -2718 2124 -2712
rect 2118 -2724 2124 -2718
rect 2118 -2730 2124 -2724
rect 2118 -2736 2124 -2730
rect 2118 -2742 2124 -2736
rect 2118 -2748 2124 -2742
rect 2118 -2754 2124 -2748
rect 2118 -2760 2124 -2754
rect 2118 -2766 2124 -2760
rect 2118 -2772 2124 -2766
rect 2118 -2778 2124 -2772
rect 2118 -2784 2124 -2778
rect 2118 -2790 2124 -2784
rect 2118 -2796 2124 -2790
rect 2118 -2802 2124 -2796
rect 2118 -2808 2124 -2802
rect 2118 -2814 2124 -2808
rect 2118 -2820 2124 -2814
rect 2118 -2826 2124 -2820
rect 2118 -2832 2124 -2826
rect 2118 -2838 2124 -2832
rect 2118 -2844 2124 -2838
rect 2118 -2850 2124 -2844
rect 2118 -2856 2124 -2850
rect 2118 -2862 2124 -2856
rect 2118 -2868 2124 -2862
rect 2118 -2874 2124 -2868
rect 2118 -2880 2124 -2874
rect 2118 -2886 2124 -2880
rect 2118 -2892 2124 -2886
rect 2118 -2898 2124 -2892
rect 2118 -2904 2124 -2898
rect 2118 -2910 2124 -2904
rect 2118 -2916 2124 -2910
rect 2118 -2922 2124 -2916
rect 2118 -2928 2124 -2922
rect 2118 -2934 2124 -2928
rect 2118 -2940 2124 -2934
rect 2118 -2946 2124 -2940
rect 2118 -2952 2124 -2946
rect 2118 -2958 2124 -2952
rect 2118 -2964 2124 -2958
rect 2118 -2970 2124 -2964
rect 2118 -2976 2124 -2970
rect 2118 -2982 2124 -2976
rect 2118 -2988 2124 -2982
rect 2118 -2994 2124 -2988
rect 2118 -3000 2124 -2994
rect 2118 -3006 2124 -3000
rect 2118 -3012 2124 -3006
rect 2118 -3018 2124 -3012
rect 2118 -3024 2124 -3018
rect 2118 -3030 2124 -3024
rect 2118 -3036 2124 -3030
rect 2118 -3042 2124 -3036
rect 2118 -3048 2124 -3042
rect 2118 -3054 2124 -3048
rect 2124 -294 2130 -288
rect 2124 -300 2130 -294
rect 2124 -306 2130 -300
rect 2124 -312 2130 -306
rect 2124 -318 2130 -312
rect 2124 -324 2130 -318
rect 2124 -330 2130 -324
rect 2124 -336 2130 -330
rect 2124 -342 2130 -336
rect 2124 -348 2130 -342
rect 2124 -354 2130 -348
rect 2124 -360 2130 -354
rect 2124 -366 2130 -360
rect 2124 -372 2130 -366
rect 2124 -378 2130 -372
rect 2124 -384 2130 -378
rect 2124 -390 2130 -384
rect 2124 -396 2130 -390
rect 2124 -402 2130 -396
rect 2124 -408 2130 -402
rect 2124 -414 2130 -408
rect 2124 -420 2130 -414
rect 2124 -426 2130 -420
rect 2124 -432 2130 -426
rect 2124 -438 2130 -432
rect 2124 -444 2130 -438
rect 2124 -450 2130 -444
rect 2124 -456 2130 -450
rect 2124 -462 2130 -456
rect 2124 -468 2130 -462
rect 2124 -474 2130 -468
rect 2124 -480 2130 -474
rect 2124 -486 2130 -480
rect 2124 -492 2130 -486
rect 2124 -498 2130 -492
rect 2124 -504 2130 -498
rect 2124 -510 2130 -504
rect 2124 -516 2130 -510
rect 2124 -522 2130 -516
rect 2124 -528 2130 -522
rect 2124 -534 2130 -528
rect 2124 -540 2130 -534
rect 2124 -546 2130 -540
rect 2124 -552 2130 -546
rect 2124 -558 2130 -552
rect 2124 -564 2130 -558
rect 2124 -570 2130 -564
rect 2124 -576 2130 -570
rect 2124 -582 2130 -576
rect 2124 -588 2130 -582
rect 2124 -594 2130 -588
rect 2124 -600 2130 -594
rect 2124 -606 2130 -600
rect 2124 -612 2130 -606
rect 2124 -618 2130 -612
rect 2124 -624 2130 -618
rect 2124 -630 2130 -624
rect 2124 -636 2130 -630
rect 2124 -642 2130 -636
rect 2124 -648 2130 -642
rect 2124 -654 2130 -648
rect 2124 -660 2130 -654
rect 2124 -666 2130 -660
rect 2124 -672 2130 -666
rect 2124 -678 2130 -672
rect 2124 -684 2130 -678
rect 2124 -690 2130 -684
rect 2124 -696 2130 -690
rect 2124 -702 2130 -696
rect 2124 -708 2130 -702
rect 2124 -714 2130 -708
rect 2124 -720 2130 -714
rect 2124 -726 2130 -720
rect 2124 -732 2130 -726
rect 2124 -738 2130 -732
rect 2124 -744 2130 -738
rect 2124 -750 2130 -744
rect 2124 -756 2130 -750
rect 2124 -762 2130 -756
rect 2124 -768 2130 -762
rect 2124 -774 2130 -768
rect 2124 -780 2130 -774
rect 2124 -786 2130 -780
rect 2124 -792 2130 -786
rect 2124 -798 2130 -792
rect 2124 -804 2130 -798
rect 2124 -810 2130 -804
rect 2124 -816 2130 -810
rect 2124 -822 2130 -816
rect 2124 -828 2130 -822
rect 2124 -834 2130 -828
rect 2124 -840 2130 -834
rect 2124 -846 2130 -840
rect 2124 -852 2130 -846
rect 2124 -858 2130 -852
rect 2124 -864 2130 -858
rect 2124 -870 2130 -864
rect 2124 -876 2130 -870
rect 2124 -882 2130 -876
rect 2124 -888 2130 -882
rect 2124 -894 2130 -888
rect 2124 -900 2130 -894
rect 2124 -906 2130 -900
rect 2124 -912 2130 -906
rect 2124 -918 2130 -912
rect 2124 -924 2130 -918
rect 2124 -930 2130 -924
rect 2124 -936 2130 -930
rect 2124 -942 2130 -936
rect 2124 -948 2130 -942
rect 2124 -954 2130 -948
rect 2124 -960 2130 -954
rect 2124 -966 2130 -960
rect 2124 -972 2130 -966
rect 2124 -978 2130 -972
rect 2124 -984 2130 -978
rect 2124 -990 2130 -984
rect 2124 -996 2130 -990
rect 2124 -1002 2130 -996
rect 2124 -1008 2130 -1002
rect 2124 -1014 2130 -1008
rect 2124 -1020 2130 -1014
rect 2124 -1026 2130 -1020
rect 2124 -1032 2130 -1026
rect 2124 -1038 2130 -1032
rect 2124 -1044 2130 -1038
rect 2124 -1050 2130 -1044
rect 2124 -1056 2130 -1050
rect 2124 -1062 2130 -1056
rect 2124 -1068 2130 -1062
rect 2124 -1074 2130 -1068
rect 2124 -1080 2130 -1074
rect 2124 -1086 2130 -1080
rect 2124 -1092 2130 -1086
rect 2124 -1098 2130 -1092
rect 2124 -1104 2130 -1098
rect 2124 -1110 2130 -1104
rect 2124 -1116 2130 -1110
rect 2124 -1122 2130 -1116
rect 2124 -1128 2130 -1122
rect 2124 -1134 2130 -1128
rect 2124 -1140 2130 -1134
rect 2124 -1146 2130 -1140
rect 2124 -1152 2130 -1146
rect 2124 -1158 2130 -1152
rect 2124 -1164 2130 -1158
rect 2124 -1170 2130 -1164
rect 2124 -1176 2130 -1170
rect 2124 -1182 2130 -1176
rect 2124 -1188 2130 -1182
rect 2124 -1194 2130 -1188
rect 2124 -1200 2130 -1194
rect 2124 -1206 2130 -1200
rect 2124 -1212 2130 -1206
rect 2124 -1218 2130 -1212
rect 2124 -1224 2130 -1218
rect 2124 -1230 2130 -1224
rect 2124 -1236 2130 -1230
rect 2124 -1242 2130 -1236
rect 2124 -1248 2130 -1242
rect 2124 -1254 2130 -1248
rect 2124 -1260 2130 -1254
rect 2124 -1266 2130 -1260
rect 2124 -1272 2130 -1266
rect 2124 -1278 2130 -1272
rect 2124 -1284 2130 -1278
rect 2124 -1290 2130 -1284
rect 2124 -1296 2130 -1290
rect 2124 -1302 2130 -1296
rect 2124 -1308 2130 -1302
rect 2124 -1314 2130 -1308
rect 2124 -1320 2130 -1314
rect 2124 -1326 2130 -1320
rect 2124 -1332 2130 -1326
rect 2124 -1338 2130 -1332
rect 2124 -1344 2130 -1338
rect 2124 -1350 2130 -1344
rect 2124 -1356 2130 -1350
rect 2124 -1362 2130 -1356
rect 2124 -1368 2130 -1362
rect 2124 -1374 2130 -1368
rect 2124 -1380 2130 -1374
rect 2124 -1386 2130 -1380
rect 2124 -1392 2130 -1386
rect 2124 -1398 2130 -1392
rect 2124 -1404 2130 -1398
rect 2124 -1410 2130 -1404
rect 2124 -1416 2130 -1410
rect 2124 -1422 2130 -1416
rect 2124 -1428 2130 -1422
rect 2124 -1620 2130 -1614
rect 2124 -1626 2130 -1620
rect 2124 -1632 2130 -1626
rect 2124 -1638 2130 -1632
rect 2124 -1644 2130 -1638
rect 2124 -1650 2130 -1644
rect 2124 -1656 2130 -1650
rect 2124 -1662 2130 -1656
rect 2124 -1668 2130 -1662
rect 2124 -1674 2130 -1668
rect 2124 -1680 2130 -1674
rect 2124 -1686 2130 -1680
rect 2124 -1692 2130 -1686
rect 2124 -1698 2130 -1692
rect 2124 -1704 2130 -1698
rect 2124 -1710 2130 -1704
rect 2124 -1716 2130 -1710
rect 2124 -1722 2130 -1716
rect 2124 -1728 2130 -1722
rect 2124 -1734 2130 -1728
rect 2124 -1740 2130 -1734
rect 2124 -1746 2130 -1740
rect 2124 -1752 2130 -1746
rect 2124 -1758 2130 -1752
rect 2124 -1764 2130 -1758
rect 2124 -1770 2130 -1764
rect 2124 -1776 2130 -1770
rect 2124 -1782 2130 -1776
rect 2124 -1788 2130 -1782
rect 2124 -1794 2130 -1788
rect 2124 -1800 2130 -1794
rect 2124 -1806 2130 -1800
rect 2124 -1812 2130 -1806
rect 2124 -1818 2130 -1812
rect 2124 -1824 2130 -1818
rect 2124 -1830 2130 -1824
rect 2124 -1836 2130 -1830
rect 2124 -1842 2130 -1836
rect 2124 -1848 2130 -1842
rect 2124 -1854 2130 -1848
rect 2124 -1860 2130 -1854
rect 2124 -1866 2130 -1860
rect 2124 -1872 2130 -1866
rect 2124 -1878 2130 -1872
rect 2124 -1884 2130 -1878
rect 2124 -1890 2130 -1884
rect 2124 -1896 2130 -1890
rect 2124 -1902 2130 -1896
rect 2124 -1908 2130 -1902
rect 2124 -1914 2130 -1908
rect 2124 -1920 2130 -1914
rect 2124 -1926 2130 -1920
rect 2124 -1932 2130 -1926
rect 2124 -1938 2130 -1932
rect 2124 -1944 2130 -1938
rect 2124 -1950 2130 -1944
rect 2124 -1956 2130 -1950
rect 2124 -1962 2130 -1956
rect 2124 -1968 2130 -1962
rect 2124 -1974 2130 -1968
rect 2124 -1980 2130 -1974
rect 2124 -1986 2130 -1980
rect 2124 -1992 2130 -1986
rect 2124 -1998 2130 -1992
rect 2124 -2004 2130 -1998
rect 2124 -2010 2130 -2004
rect 2124 -2016 2130 -2010
rect 2124 -2022 2130 -2016
rect 2124 -2028 2130 -2022
rect 2124 -2034 2130 -2028
rect 2124 -2040 2130 -2034
rect 2124 -2046 2130 -2040
rect 2124 -2052 2130 -2046
rect 2124 -2058 2130 -2052
rect 2124 -2064 2130 -2058
rect 2124 -2070 2130 -2064
rect 2124 -2076 2130 -2070
rect 2124 -2082 2130 -2076
rect 2124 -2088 2130 -2082
rect 2124 -2094 2130 -2088
rect 2124 -2100 2130 -2094
rect 2124 -2106 2130 -2100
rect 2124 -2112 2130 -2106
rect 2124 -2118 2130 -2112
rect 2124 -2124 2130 -2118
rect 2124 -2130 2130 -2124
rect 2124 -2136 2130 -2130
rect 2124 -2142 2130 -2136
rect 2124 -2148 2130 -2142
rect 2124 -2154 2130 -2148
rect 2124 -2160 2130 -2154
rect 2124 -2166 2130 -2160
rect 2124 -2172 2130 -2166
rect 2124 -2178 2130 -2172
rect 2124 -2184 2130 -2178
rect 2124 -2190 2130 -2184
rect 2124 -2196 2130 -2190
rect 2124 -2202 2130 -2196
rect 2124 -2208 2130 -2202
rect 2124 -2214 2130 -2208
rect 2124 -2220 2130 -2214
rect 2124 -2226 2130 -2220
rect 2124 -2232 2130 -2226
rect 2124 -2238 2130 -2232
rect 2124 -2244 2130 -2238
rect 2124 -2250 2130 -2244
rect 2124 -2256 2130 -2250
rect 2124 -2262 2130 -2256
rect 2124 -2268 2130 -2262
rect 2124 -2274 2130 -2268
rect 2124 -2280 2130 -2274
rect 2124 -2286 2130 -2280
rect 2124 -2292 2130 -2286
rect 2124 -2298 2130 -2292
rect 2124 -2304 2130 -2298
rect 2124 -2310 2130 -2304
rect 2124 -2316 2130 -2310
rect 2124 -2322 2130 -2316
rect 2124 -2328 2130 -2322
rect 2124 -2334 2130 -2328
rect 2124 -2340 2130 -2334
rect 2124 -2346 2130 -2340
rect 2124 -2352 2130 -2346
rect 2124 -2358 2130 -2352
rect 2124 -2364 2130 -2358
rect 2124 -2370 2130 -2364
rect 2124 -2376 2130 -2370
rect 2124 -2382 2130 -2376
rect 2124 -2388 2130 -2382
rect 2124 -2394 2130 -2388
rect 2124 -2400 2130 -2394
rect 2124 -2406 2130 -2400
rect 2124 -2412 2130 -2406
rect 2124 -2418 2130 -2412
rect 2124 -2424 2130 -2418
rect 2124 -2430 2130 -2424
rect 2124 -2436 2130 -2430
rect 2124 -2562 2130 -2556
rect 2124 -2568 2130 -2562
rect 2124 -2574 2130 -2568
rect 2124 -2580 2130 -2574
rect 2124 -2586 2130 -2580
rect 2124 -2592 2130 -2586
rect 2124 -2598 2130 -2592
rect 2124 -2604 2130 -2598
rect 2124 -2610 2130 -2604
rect 2124 -2616 2130 -2610
rect 2124 -2622 2130 -2616
rect 2124 -2628 2130 -2622
rect 2124 -2634 2130 -2628
rect 2124 -2640 2130 -2634
rect 2124 -2646 2130 -2640
rect 2124 -2652 2130 -2646
rect 2124 -2658 2130 -2652
rect 2124 -2664 2130 -2658
rect 2124 -2670 2130 -2664
rect 2124 -2676 2130 -2670
rect 2124 -2682 2130 -2676
rect 2124 -2688 2130 -2682
rect 2124 -2694 2130 -2688
rect 2124 -2700 2130 -2694
rect 2124 -2706 2130 -2700
rect 2124 -2712 2130 -2706
rect 2124 -2718 2130 -2712
rect 2124 -2724 2130 -2718
rect 2124 -2730 2130 -2724
rect 2124 -2736 2130 -2730
rect 2124 -2742 2130 -2736
rect 2124 -2748 2130 -2742
rect 2124 -2754 2130 -2748
rect 2124 -2760 2130 -2754
rect 2124 -2766 2130 -2760
rect 2124 -2772 2130 -2766
rect 2124 -2778 2130 -2772
rect 2124 -2784 2130 -2778
rect 2124 -2790 2130 -2784
rect 2124 -2796 2130 -2790
rect 2124 -2802 2130 -2796
rect 2124 -2808 2130 -2802
rect 2124 -2814 2130 -2808
rect 2124 -2820 2130 -2814
rect 2124 -2826 2130 -2820
rect 2124 -2832 2130 -2826
rect 2124 -2838 2130 -2832
rect 2124 -2844 2130 -2838
rect 2124 -2850 2130 -2844
rect 2124 -2856 2130 -2850
rect 2124 -2862 2130 -2856
rect 2124 -2868 2130 -2862
rect 2124 -2874 2130 -2868
rect 2124 -2880 2130 -2874
rect 2124 -2886 2130 -2880
rect 2124 -2892 2130 -2886
rect 2124 -2898 2130 -2892
rect 2124 -2904 2130 -2898
rect 2124 -2910 2130 -2904
rect 2124 -2916 2130 -2910
rect 2124 -2922 2130 -2916
rect 2124 -2928 2130 -2922
rect 2124 -2934 2130 -2928
rect 2124 -2940 2130 -2934
rect 2124 -2946 2130 -2940
rect 2124 -2952 2130 -2946
rect 2124 -2958 2130 -2952
rect 2124 -2964 2130 -2958
rect 2124 -2970 2130 -2964
rect 2124 -2976 2130 -2970
rect 2124 -2982 2130 -2976
rect 2124 -2988 2130 -2982
rect 2124 -2994 2130 -2988
rect 2124 -3000 2130 -2994
rect 2124 -3006 2130 -3000
rect 2124 -3012 2130 -3006
rect 2124 -3018 2130 -3012
rect 2124 -3024 2130 -3018
rect 2124 -3030 2130 -3024
rect 2124 -3036 2130 -3030
rect 2124 -3042 2130 -3036
rect 2124 -3048 2130 -3042
rect 2124 -3054 2130 -3048
rect 2130 -288 2136 -282
rect 2130 -294 2136 -288
rect 2130 -300 2136 -294
rect 2130 -306 2136 -300
rect 2130 -312 2136 -306
rect 2130 -318 2136 -312
rect 2130 -324 2136 -318
rect 2130 -330 2136 -324
rect 2130 -336 2136 -330
rect 2130 -342 2136 -336
rect 2130 -348 2136 -342
rect 2130 -354 2136 -348
rect 2130 -360 2136 -354
rect 2130 -366 2136 -360
rect 2130 -372 2136 -366
rect 2130 -378 2136 -372
rect 2130 -384 2136 -378
rect 2130 -390 2136 -384
rect 2130 -396 2136 -390
rect 2130 -402 2136 -396
rect 2130 -408 2136 -402
rect 2130 -414 2136 -408
rect 2130 -420 2136 -414
rect 2130 -426 2136 -420
rect 2130 -432 2136 -426
rect 2130 -438 2136 -432
rect 2130 -444 2136 -438
rect 2130 -450 2136 -444
rect 2130 -456 2136 -450
rect 2130 -462 2136 -456
rect 2130 -468 2136 -462
rect 2130 -474 2136 -468
rect 2130 -480 2136 -474
rect 2130 -486 2136 -480
rect 2130 -492 2136 -486
rect 2130 -498 2136 -492
rect 2130 -504 2136 -498
rect 2130 -510 2136 -504
rect 2130 -516 2136 -510
rect 2130 -522 2136 -516
rect 2130 -528 2136 -522
rect 2130 -534 2136 -528
rect 2130 -540 2136 -534
rect 2130 -546 2136 -540
rect 2130 -552 2136 -546
rect 2130 -558 2136 -552
rect 2130 -564 2136 -558
rect 2130 -570 2136 -564
rect 2130 -576 2136 -570
rect 2130 -582 2136 -576
rect 2130 -588 2136 -582
rect 2130 -594 2136 -588
rect 2130 -600 2136 -594
rect 2130 -606 2136 -600
rect 2130 -612 2136 -606
rect 2130 -618 2136 -612
rect 2130 -624 2136 -618
rect 2130 -630 2136 -624
rect 2130 -636 2136 -630
rect 2130 -642 2136 -636
rect 2130 -648 2136 -642
rect 2130 -654 2136 -648
rect 2130 -660 2136 -654
rect 2130 -666 2136 -660
rect 2130 -672 2136 -666
rect 2130 -678 2136 -672
rect 2130 -684 2136 -678
rect 2130 -690 2136 -684
rect 2130 -696 2136 -690
rect 2130 -702 2136 -696
rect 2130 -708 2136 -702
rect 2130 -714 2136 -708
rect 2130 -720 2136 -714
rect 2130 -726 2136 -720
rect 2130 -732 2136 -726
rect 2130 -738 2136 -732
rect 2130 -744 2136 -738
rect 2130 -750 2136 -744
rect 2130 -756 2136 -750
rect 2130 -762 2136 -756
rect 2130 -768 2136 -762
rect 2130 -774 2136 -768
rect 2130 -780 2136 -774
rect 2130 -786 2136 -780
rect 2130 -792 2136 -786
rect 2130 -798 2136 -792
rect 2130 -804 2136 -798
rect 2130 -810 2136 -804
rect 2130 -816 2136 -810
rect 2130 -822 2136 -816
rect 2130 -828 2136 -822
rect 2130 -834 2136 -828
rect 2130 -840 2136 -834
rect 2130 -846 2136 -840
rect 2130 -852 2136 -846
rect 2130 -858 2136 -852
rect 2130 -864 2136 -858
rect 2130 -870 2136 -864
rect 2130 -876 2136 -870
rect 2130 -882 2136 -876
rect 2130 -888 2136 -882
rect 2130 -894 2136 -888
rect 2130 -900 2136 -894
rect 2130 -906 2136 -900
rect 2130 -912 2136 -906
rect 2130 -918 2136 -912
rect 2130 -924 2136 -918
rect 2130 -930 2136 -924
rect 2130 -936 2136 -930
rect 2130 -942 2136 -936
rect 2130 -948 2136 -942
rect 2130 -954 2136 -948
rect 2130 -960 2136 -954
rect 2130 -966 2136 -960
rect 2130 -972 2136 -966
rect 2130 -978 2136 -972
rect 2130 -984 2136 -978
rect 2130 -990 2136 -984
rect 2130 -996 2136 -990
rect 2130 -1002 2136 -996
rect 2130 -1008 2136 -1002
rect 2130 -1014 2136 -1008
rect 2130 -1020 2136 -1014
rect 2130 -1026 2136 -1020
rect 2130 -1032 2136 -1026
rect 2130 -1038 2136 -1032
rect 2130 -1044 2136 -1038
rect 2130 -1050 2136 -1044
rect 2130 -1056 2136 -1050
rect 2130 -1062 2136 -1056
rect 2130 -1068 2136 -1062
rect 2130 -1074 2136 -1068
rect 2130 -1080 2136 -1074
rect 2130 -1086 2136 -1080
rect 2130 -1092 2136 -1086
rect 2130 -1098 2136 -1092
rect 2130 -1104 2136 -1098
rect 2130 -1110 2136 -1104
rect 2130 -1116 2136 -1110
rect 2130 -1122 2136 -1116
rect 2130 -1128 2136 -1122
rect 2130 -1134 2136 -1128
rect 2130 -1140 2136 -1134
rect 2130 -1146 2136 -1140
rect 2130 -1152 2136 -1146
rect 2130 -1158 2136 -1152
rect 2130 -1164 2136 -1158
rect 2130 -1170 2136 -1164
rect 2130 -1176 2136 -1170
rect 2130 -1182 2136 -1176
rect 2130 -1188 2136 -1182
rect 2130 -1194 2136 -1188
rect 2130 -1200 2136 -1194
rect 2130 -1206 2136 -1200
rect 2130 -1212 2136 -1206
rect 2130 -1218 2136 -1212
rect 2130 -1224 2136 -1218
rect 2130 -1230 2136 -1224
rect 2130 -1236 2136 -1230
rect 2130 -1242 2136 -1236
rect 2130 -1248 2136 -1242
rect 2130 -1254 2136 -1248
rect 2130 -1260 2136 -1254
rect 2130 -1266 2136 -1260
rect 2130 -1272 2136 -1266
rect 2130 -1278 2136 -1272
rect 2130 -1284 2136 -1278
rect 2130 -1290 2136 -1284
rect 2130 -1296 2136 -1290
rect 2130 -1302 2136 -1296
rect 2130 -1308 2136 -1302
rect 2130 -1314 2136 -1308
rect 2130 -1320 2136 -1314
rect 2130 -1326 2136 -1320
rect 2130 -1332 2136 -1326
rect 2130 -1338 2136 -1332
rect 2130 -1344 2136 -1338
rect 2130 -1350 2136 -1344
rect 2130 -1356 2136 -1350
rect 2130 -1362 2136 -1356
rect 2130 -1368 2136 -1362
rect 2130 -1374 2136 -1368
rect 2130 -1380 2136 -1374
rect 2130 -1386 2136 -1380
rect 2130 -1392 2136 -1386
rect 2130 -1398 2136 -1392
rect 2130 -1404 2136 -1398
rect 2130 -1410 2136 -1404
rect 2130 -1614 2136 -1608
rect 2130 -1620 2136 -1614
rect 2130 -1626 2136 -1620
rect 2130 -1632 2136 -1626
rect 2130 -1638 2136 -1632
rect 2130 -1644 2136 -1638
rect 2130 -1650 2136 -1644
rect 2130 -1656 2136 -1650
rect 2130 -1662 2136 -1656
rect 2130 -1668 2136 -1662
rect 2130 -1674 2136 -1668
rect 2130 -1680 2136 -1674
rect 2130 -1686 2136 -1680
rect 2130 -1692 2136 -1686
rect 2130 -1698 2136 -1692
rect 2130 -1704 2136 -1698
rect 2130 -1710 2136 -1704
rect 2130 -1716 2136 -1710
rect 2130 -1722 2136 -1716
rect 2130 -1728 2136 -1722
rect 2130 -1734 2136 -1728
rect 2130 -1740 2136 -1734
rect 2130 -1746 2136 -1740
rect 2130 -1752 2136 -1746
rect 2130 -1758 2136 -1752
rect 2130 -1764 2136 -1758
rect 2130 -1770 2136 -1764
rect 2130 -1776 2136 -1770
rect 2130 -1782 2136 -1776
rect 2130 -1788 2136 -1782
rect 2130 -1794 2136 -1788
rect 2130 -1800 2136 -1794
rect 2130 -1806 2136 -1800
rect 2130 -1812 2136 -1806
rect 2130 -1818 2136 -1812
rect 2130 -1824 2136 -1818
rect 2130 -1830 2136 -1824
rect 2130 -1836 2136 -1830
rect 2130 -1842 2136 -1836
rect 2130 -1848 2136 -1842
rect 2130 -1854 2136 -1848
rect 2130 -1860 2136 -1854
rect 2130 -1866 2136 -1860
rect 2130 -1872 2136 -1866
rect 2130 -1878 2136 -1872
rect 2130 -1884 2136 -1878
rect 2130 -1890 2136 -1884
rect 2130 -1896 2136 -1890
rect 2130 -1902 2136 -1896
rect 2130 -1908 2136 -1902
rect 2130 -1914 2136 -1908
rect 2130 -1920 2136 -1914
rect 2130 -1926 2136 -1920
rect 2130 -1932 2136 -1926
rect 2130 -1938 2136 -1932
rect 2130 -1944 2136 -1938
rect 2130 -1950 2136 -1944
rect 2130 -1956 2136 -1950
rect 2130 -1962 2136 -1956
rect 2130 -1968 2136 -1962
rect 2130 -1974 2136 -1968
rect 2130 -1980 2136 -1974
rect 2130 -1986 2136 -1980
rect 2130 -1992 2136 -1986
rect 2130 -1998 2136 -1992
rect 2130 -2004 2136 -1998
rect 2130 -2010 2136 -2004
rect 2130 -2016 2136 -2010
rect 2130 -2022 2136 -2016
rect 2130 -2028 2136 -2022
rect 2130 -2034 2136 -2028
rect 2130 -2040 2136 -2034
rect 2130 -2046 2136 -2040
rect 2130 -2052 2136 -2046
rect 2130 -2058 2136 -2052
rect 2130 -2064 2136 -2058
rect 2130 -2070 2136 -2064
rect 2130 -2076 2136 -2070
rect 2130 -2082 2136 -2076
rect 2130 -2088 2136 -2082
rect 2130 -2094 2136 -2088
rect 2130 -2100 2136 -2094
rect 2130 -2106 2136 -2100
rect 2130 -2112 2136 -2106
rect 2130 -2118 2136 -2112
rect 2130 -2124 2136 -2118
rect 2130 -2130 2136 -2124
rect 2130 -2136 2136 -2130
rect 2130 -2142 2136 -2136
rect 2130 -2148 2136 -2142
rect 2130 -2154 2136 -2148
rect 2130 -2160 2136 -2154
rect 2130 -2166 2136 -2160
rect 2130 -2172 2136 -2166
rect 2130 -2178 2136 -2172
rect 2130 -2184 2136 -2178
rect 2130 -2190 2136 -2184
rect 2130 -2196 2136 -2190
rect 2130 -2202 2136 -2196
rect 2130 -2208 2136 -2202
rect 2130 -2214 2136 -2208
rect 2130 -2220 2136 -2214
rect 2130 -2226 2136 -2220
rect 2130 -2232 2136 -2226
rect 2130 -2238 2136 -2232
rect 2130 -2244 2136 -2238
rect 2130 -2250 2136 -2244
rect 2130 -2256 2136 -2250
rect 2130 -2262 2136 -2256
rect 2130 -2268 2136 -2262
rect 2130 -2274 2136 -2268
rect 2130 -2280 2136 -2274
rect 2130 -2286 2136 -2280
rect 2130 -2292 2136 -2286
rect 2130 -2298 2136 -2292
rect 2130 -2304 2136 -2298
rect 2130 -2310 2136 -2304
rect 2130 -2316 2136 -2310
rect 2130 -2322 2136 -2316
rect 2130 -2328 2136 -2322
rect 2130 -2334 2136 -2328
rect 2130 -2340 2136 -2334
rect 2130 -2346 2136 -2340
rect 2130 -2352 2136 -2346
rect 2130 -2358 2136 -2352
rect 2130 -2364 2136 -2358
rect 2130 -2370 2136 -2364
rect 2130 -2376 2136 -2370
rect 2130 -2382 2136 -2376
rect 2130 -2388 2136 -2382
rect 2130 -2394 2136 -2388
rect 2130 -2400 2136 -2394
rect 2130 -2406 2136 -2400
rect 2130 -2412 2136 -2406
rect 2130 -2418 2136 -2412
rect 2130 -2424 2136 -2418
rect 2130 -2430 2136 -2424
rect 2130 -2562 2136 -2556
rect 2130 -2568 2136 -2562
rect 2130 -2574 2136 -2568
rect 2130 -2580 2136 -2574
rect 2130 -2586 2136 -2580
rect 2130 -2592 2136 -2586
rect 2130 -2598 2136 -2592
rect 2130 -2604 2136 -2598
rect 2130 -2610 2136 -2604
rect 2130 -2616 2136 -2610
rect 2130 -2622 2136 -2616
rect 2130 -2628 2136 -2622
rect 2130 -2634 2136 -2628
rect 2130 -2640 2136 -2634
rect 2130 -2646 2136 -2640
rect 2130 -2652 2136 -2646
rect 2130 -2658 2136 -2652
rect 2130 -2664 2136 -2658
rect 2130 -2670 2136 -2664
rect 2130 -2676 2136 -2670
rect 2130 -2682 2136 -2676
rect 2130 -2688 2136 -2682
rect 2130 -2694 2136 -2688
rect 2130 -2700 2136 -2694
rect 2130 -2706 2136 -2700
rect 2130 -2712 2136 -2706
rect 2130 -2718 2136 -2712
rect 2130 -2724 2136 -2718
rect 2130 -2730 2136 -2724
rect 2130 -2736 2136 -2730
rect 2130 -2742 2136 -2736
rect 2130 -2748 2136 -2742
rect 2130 -2754 2136 -2748
rect 2130 -2760 2136 -2754
rect 2130 -2766 2136 -2760
rect 2130 -2772 2136 -2766
rect 2130 -2778 2136 -2772
rect 2130 -2784 2136 -2778
rect 2130 -2790 2136 -2784
rect 2130 -2796 2136 -2790
rect 2130 -2802 2136 -2796
rect 2130 -2808 2136 -2802
rect 2130 -2814 2136 -2808
rect 2130 -2820 2136 -2814
rect 2130 -2826 2136 -2820
rect 2130 -2832 2136 -2826
rect 2130 -2838 2136 -2832
rect 2130 -2844 2136 -2838
rect 2130 -2850 2136 -2844
rect 2130 -2856 2136 -2850
rect 2130 -2862 2136 -2856
rect 2130 -2868 2136 -2862
rect 2130 -2874 2136 -2868
rect 2130 -2880 2136 -2874
rect 2130 -2886 2136 -2880
rect 2130 -2892 2136 -2886
rect 2130 -2898 2136 -2892
rect 2130 -2904 2136 -2898
rect 2130 -2910 2136 -2904
rect 2130 -2916 2136 -2910
rect 2130 -2922 2136 -2916
rect 2130 -2928 2136 -2922
rect 2130 -2934 2136 -2928
rect 2130 -2940 2136 -2934
rect 2130 -2946 2136 -2940
rect 2130 -2952 2136 -2946
rect 2130 -2958 2136 -2952
rect 2130 -2964 2136 -2958
rect 2130 -2970 2136 -2964
rect 2130 -2976 2136 -2970
rect 2130 -2982 2136 -2976
rect 2130 -2988 2136 -2982
rect 2130 -2994 2136 -2988
rect 2130 -3000 2136 -2994
rect 2130 -3006 2136 -3000
rect 2130 -3012 2136 -3006
rect 2130 -3018 2136 -3012
rect 2130 -3024 2136 -3018
rect 2130 -3030 2136 -3024
rect 2130 -3036 2136 -3030
rect 2130 -3042 2136 -3036
rect 2130 -3048 2136 -3042
rect 2136 -276 2142 -270
rect 2136 -282 2142 -276
rect 2136 -288 2142 -282
rect 2136 -294 2142 -288
rect 2136 -300 2142 -294
rect 2136 -306 2142 -300
rect 2136 -312 2142 -306
rect 2136 -318 2142 -312
rect 2136 -324 2142 -318
rect 2136 -330 2142 -324
rect 2136 -336 2142 -330
rect 2136 -342 2142 -336
rect 2136 -348 2142 -342
rect 2136 -354 2142 -348
rect 2136 -360 2142 -354
rect 2136 -366 2142 -360
rect 2136 -372 2142 -366
rect 2136 -378 2142 -372
rect 2136 -384 2142 -378
rect 2136 -390 2142 -384
rect 2136 -396 2142 -390
rect 2136 -402 2142 -396
rect 2136 -408 2142 -402
rect 2136 -414 2142 -408
rect 2136 -420 2142 -414
rect 2136 -426 2142 -420
rect 2136 -432 2142 -426
rect 2136 -438 2142 -432
rect 2136 -444 2142 -438
rect 2136 -450 2142 -444
rect 2136 -456 2142 -450
rect 2136 -462 2142 -456
rect 2136 -468 2142 -462
rect 2136 -474 2142 -468
rect 2136 -480 2142 -474
rect 2136 -486 2142 -480
rect 2136 -492 2142 -486
rect 2136 -498 2142 -492
rect 2136 -504 2142 -498
rect 2136 -510 2142 -504
rect 2136 -516 2142 -510
rect 2136 -522 2142 -516
rect 2136 -528 2142 -522
rect 2136 -534 2142 -528
rect 2136 -540 2142 -534
rect 2136 -546 2142 -540
rect 2136 -552 2142 -546
rect 2136 -558 2142 -552
rect 2136 -564 2142 -558
rect 2136 -570 2142 -564
rect 2136 -576 2142 -570
rect 2136 -582 2142 -576
rect 2136 -588 2142 -582
rect 2136 -594 2142 -588
rect 2136 -600 2142 -594
rect 2136 -606 2142 -600
rect 2136 -612 2142 -606
rect 2136 -618 2142 -612
rect 2136 -624 2142 -618
rect 2136 -630 2142 -624
rect 2136 -636 2142 -630
rect 2136 -642 2142 -636
rect 2136 -648 2142 -642
rect 2136 -654 2142 -648
rect 2136 -660 2142 -654
rect 2136 -666 2142 -660
rect 2136 -672 2142 -666
rect 2136 -678 2142 -672
rect 2136 -684 2142 -678
rect 2136 -690 2142 -684
rect 2136 -696 2142 -690
rect 2136 -702 2142 -696
rect 2136 -708 2142 -702
rect 2136 -714 2142 -708
rect 2136 -720 2142 -714
rect 2136 -726 2142 -720
rect 2136 -732 2142 -726
rect 2136 -738 2142 -732
rect 2136 -744 2142 -738
rect 2136 -750 2142 -744
rect 2136 -756 2142 -750
rect 2136 -762 2142 -756
rect 2136 -768 2142 -762
rect 2136 -774 2142 -768
rect 2136 -780 2142 -774
rect 2136 -786 2142 -780
rect 2136 -792 2142 -786
rect 2136 -798 2142 -792
rect 2136 -804 2142 -798
rect 2136 -810 2142 -804
rect 2136 -816 2142 -810
rect 2136 -822 2142 -816
rect 2136 -828 2142 -822
rect 2136 -834 2142 -828
rect 2136 -840 2142 -834
rect 2136 -846 2142 -840
rect 2136 -852 2142 -846
rect 2136 -858 2142 -852
rect 2136 -864 2142 -858
rect 2136 -870 2142 -864
rect 2136 -876 2142 -870
rect 2136 -882 2142 -876
rect 2136 -888 2142 -882
rect 2136 -894 2142 -888
rect 2136 -900 2142 -894
rect 2136 -906 2142 -900
rect 2136 -912 2142 -906
rect 2136 -918 2142 -912
rect 2136 -924 2142 -918
rect 2136 -930 2142 -924
rect 2136 -936 2142 -930
rect 2136 -942 2142 -936
rect 2136 -948 2142 -942
rect 2136 -954 2142 -948
rect 2136 -960 2142 -954
rect 2136 -966 2142 -960
rect 2136 -972 2142 -966
rect 2136 -978 2142 -972
rect 2136 -984 2142 -978
rect 2136 -990 2142 -984
rect 2136 -996 2142 -990
rect 2136 -1002 2142 -996
rect 2136 -1008 2142 -1002
rect 2136 -1014 2142 -1008
rect 2136 -1020 2142 -1014
rect 2136 -1026 2142 -1020
rect 2136 -1032 2142 -1026
rect 2136 -1038 2142 -1032
rect 2136 -1044 2142 -1038
rect 2136 -1050 2142 -1044
rect 2136 -1056 2142 -1050
rect 2136 -1062 2142 -1056
rect 2136 -1068 2142 -1062
rect 2136 -1074 2142 -1068
rect 2136 -1080 2142 -1074
rect 2136 -1086 2142 -1080
rect 2136 -1092 2142 -1086
rect 2136 -1098 2142 -1092
rect 2136 -1104 2142 -1098
rect 2136 -1110 2142 -1104
rect 2136 -1116 2142 -1110
rect 2136 -1122 2142 -1116
rect 2136 -1128 2142 -1122
rect 2136 -1134 2142 -1128
rect 2136 -1140 2142 -1134
rect 2136 -1146 2142 -1140
rect 2136 -1152 2142 -1146
rect 2136 -1158 2142 -1152
rect 2136 -1164 2142 -1158
rect 2136 -1170 2142 -1164
rect 2136 -1176 2142 -1170
rect 2136 -1182 2142 -1176
rect 2136 -1188 2142 -1182
rect 2136 -1194 2142 -1188
rect 2136 -1200 2142 -1194
rect 2136 -1206 2142 -1200
rect 2136 -1212 2142 -1206
rect 2136 -1218 2142 -1212
rect 2136 -1224 2142 -1218
rect 2136 -1230 2142 -1224
rect 2136 -1236 2142 -1230
rect 2136 -1242 2142 -1236
rect 2136 -1248 2142 -1242
rect 2136 -1254 2142 -1248
rect 2136 -1260 2142 -1254
rect 2136 -1266 2142 -1260
rect 2136 -1272 2142 -1266
rect 2136 -1278 2142 -1272
rect 2136 -1284 2142 -1278
rect 2136 -1290 2142 -1284
rect 2136 -1296 2142 -1290
rect 2136 -1302 2142 -1296
rect 2136 -1308 2142 -1302
rect 2136 -1314 2142 -1308
rect 2136 -1320 2142 -1314
rect 2136 -1326 2142 -1320
rect 2136 -1332 2142 -1326
rect 2136 -1338 2142 -1332
rect 2136 -1344 2142 -1338
rect 2136 -1350 2142 -1344
rect 2136 -1356 2142 -1350
rect 2136 -1362 2142 -1356
rect 2136 -1368 2142 -1362
rect 2136 -1374 2142 -1368
rect 2136 -1380 2142 -1374
rect 2136 -1386 2142 -1380
rect 2136 -1392 2142 -1386
rect 2136 -1398 2142 -1392
rect 2136 -1608 2142 -1602
rect 2136 -1614 2142 -1608
rect 2136 -1620 2142 -1614
rect 2136 -1626 2142 -1620
rect 2136 -1632 2142 -1626
rect 2136 -1638 2142 -1632
rect 2136 -1644 2142 -1638
rect 2136 -1650 2142 -1644
rect 2136 -1656 2142 -1650
rect 2136 -1662 2142 -1656
rect 2136 -1668 2142 -1662
rect 2136 -1674 2142 -1668
rect 2136 -1680 2142 -1674
rect 2136 -1686 2142 -1680
rect 2136 -1692 2142 -1686
rect 2136 -1698 2142 -1692
rect 2136 -1704 2142 -1698
rect 2136 -1710 2142 -1704
rect 2136 -1716 2142 -1710
rect 2136 -1722 2142 -1716
rect 2136 -1728 2142 -1722
rect 2136 -1734 2142 -1728
rect 2136 -1740 2142 -1734
rect 2136 -1746 2142 -1740
rect 2136 -1752 2142 -1746
rect 2136 -1758 2142 -1752
rect 2136 -1764 2142 -1758
rect 2136 -1770 2142 -1764
rect 2136 -1776 2142 -1770
rect 2136 -1782 2142 -1776
rect 2136 -1788 2142 -1782
rect 2136 -1794 2142 -1788
rect 2136 -1800 2142 -1794
rect 2136 -1806 2142 -1800
rect 2136 -1812 2142 -1806
rect 2136 -1818 2142 -1812
rect 2136 -1824 2142 -1818
rect 2136 -1830 2142 -1824
rect 2136 -1836 2142 -1830
rect 2136 -1842 2142 -1836
rect 2136 -1848 2142 -1842
rect 2136 -1854 2142 -1848
rect 2136 -1860 2142 -1854
rect 2136 -1866 2142 -1860
rect 2136 -1872 2142 -1866
rect 2136 -1878 2142 -1872
rect 2136 -1884 2142 -1878
rect 2136 -1890 2142 -1884
rect 2136 -1896 2142 -1890
rect 2136 -1902 2142 -1896
rect 2136 -1908 2142 -1902
rect 2136 -1914 2142 -1908
rect 2136 -1920 2142 -1914
rect 2136 -1926 2142 -1920
rect 2136 -1932 2142 -1926
rect 2136 -1938 2142 -1932
rect 2136 -1944 2142 -1938
rect 2136 -1950 2142 -1944
rect 2136 -1956 2142 -1950
rect 2136 -1962 2142 -1956
rect 2136 -1968 2142 -1962
rect 2136 -1974 2142 -1968
rect 2136 -1980 2142 -1974
rect 2136 -1986 2142 -1980
rect 2136 -1992 2142 -1986
rect 2136 -1998 2142 -1992
rect 2136 -2004 2142 -1998
rect 2136 -2010 2142 -2004
rect 2136 -2016 2142 -2010
rect 2136 -2022 2142 -2016
rect 2136 -2028 2142 -2022
rect 2136 -2034 2142 -2028
rect 2136 -2040 2142 -2034
rect 2136 -2046 2142 -2040
rect 2136 -2052 2142 -2046
rect 2136 -2058 2142 -2052
rect 2136 -2064 2142 -2058
rect 2136 -2070 2142 -2064
rect 2136 -2076 2142 -2070
rect 2136 -2082 2142 -2076
rect 2136 -2088 2142 -2082
rect 2136 -2094 2142 -2088
rect 2136 -2100 2142 -2094
rect 2136 -2106 2142 -2100
rect 2136 -2112 2142 -2106
rect 2136 -2118 2142 -2112
rect 2136 -2124 2142 -2118
rect 2136 -2130 2142 -2124
rect 2136 -2136 2142 -2130
rect 2136 -2142 2142 -2136
rect 2136 -2148 2142 -2142
rect 2136 -2154 2142 -2148
rect 2136 -2160 2142 -2154
rect 2136 -2166 2142 -2160
rect 2136 -2172 2142 -2166
rect 2136 -2178 2142 -2172
rect 2136 -2184 2142 -2178
rect 2136 -2190 2142 -2184
rect 2136 -2196 2142 -2190
rect 2136 -2202 2142 -2196
rect 2136 -2208 2142 -2202
rect 2136 -2214 2142 -2208
rect 2136 -2220 2142 -2214
rect 2136 -2226 2142 -2220
rect 2136 -2232 2142 -2226
rect 2136 -2238 2142 -2232
rect 2136 -2244 2142 -2238
rect 2136 -2250 2142 -2244
rect 2136 -2256 2142 -2250
rect 2136 -2262 2142 -2256
rect 2136 -2268 2142 -2262
rect 2136 -2274 2142 -2268
rect 2136 -2280 2142 -2274
rect 2136 -2286 2142 -2280
rect 2136 -2292 2142 -2286
rect 2136 -2298 2142 -2292
rect 2136 -2304 2142 -2298
rect 2136 -2310 2142 -2304
rect 2136 -2316 2142 -2310
rect 2136 -2322 2142 -2316
rect 2136 -2328 2142 -2322
rect 2136 -2334 2142 -2328
rect 2136 -2340 2142 -2334
rect 2136 -2346 2142 -2340
rect 2136 -2352 2142 -2346
rect 2136 -2358 2142 -2352
rect 2136 -2364 2142 -2358
rect 2136 -2370 2142 -2364
rect 2136 -2376 2142 -2370
rect 2136 -2382 2142 -2376
rect 2136 -2388 2142 -2382
rect 2136 -2394 2142 -2388
rect 2136 -2400 2142 -2394
rect 2136 -2406 2142 -2400
rect 2136 -2412 2142 -2406
rect 2136 -2418 2142 -2412
rect 2136 -2424 2142 -2418
rect 2136 -2562 2142 -2556
rect 2136 -2568 2142 -2562
rect 2136 -2574 2142 -2568
rect 2136 -2580 2142 -2574
rect 2136 -2586 2142 -2580
rect 2136 -2592 2142 -2586
rect 2136 -2598 2142 -2592
rect 2136 -2604 2142 -2598
rect 2136 -2610 2142 -2604
rect 2136 -2616 2142 -2610
rect 2136 -2622 2142 -2616
rect 2136 -2628 2142 -2622
rect 2136 -2634 2142 -2628
rect 2136 -2640 2142 -2634
rect 2136 -2646 2142 -2640
rect 2136 -2652 2142 -2646
rect 2136 -2658 2142 -2652
rect 2136 -2664 2142 -2658
rect 2136 -2670 2142 -2664
rect 2136 -2676 2142 -2670
rect 2136 -2682 2142 -2676
rect 2136 -2688 2142 -2682
rect 2136 -2694 2142 -2688
rect 2136 -2700 2142 -2694
rect 2136 -2706 2142 -2700
rect 2136 -2712 2142 -2706
rect 2136 -2718 2142 -2712
rect 2136 -2724 2142 -2718
rect 2136 -2730 2142 -2724
rect 2136 -2736 2142 -2730
rect 2136 -2742 2142 -2736
rect 2136 -2748 2142 -2742
rect 2136 -2754 2142 -2748
rect 2136 -2760 2142 -2754
rect 2136 -2766 2142 -2760
rect 2136 -2772 2142 -2766
rect 2136 -2778 2142 -2772
rect 2136 -2784 2142 -2778
rect 2136 -2790 2142 -2784
rect 2136 -2796 2142 -2790
rect 2136 -2802 2142 -2796
rect 2136 -2808 2142 -2802
rect 2136 -2814 2142 -2808
rect 2136 -2820 2142 -2814
rect 2136 -2826 2142 -2820
rect 2136 -2832 2142 -2826
rect 2136 -2838 2142 -2832
rect 2136 -2844 2142 -2838
rect 2136 -2850 2142 -2844
rect 2136 -2856 2142 -2850
rect 2136 -2862 2142 -2856
rect 2136 -2868 2142 -2862
rect 2136 -2874 2142 -2868
rect 2136 -2880 2142 -2874
rect 2136 -2886 2142 -2880
rect 2136 -2892 2142 -2886
rect 2136 -2898 2142 -2892
rect 2136 -2904 2142 -2898
rect 2136 -2910 2142 -2904
rect 2136 -2916 2142 -2910
rect 2136 -2922 2142 -2916
rect 2136 -2928 2142 -2922
rect 2136 -2934 2142 -2928
rect 2136 -2940 2142 -2934
rect 2136 -2946 2142 -2940
rect 2136 -2952 2142 -2946
rect 2136 -2958 2142 -2952
rect 2136 -2964 2142 -2958
rect 2136 -2970 2142 -2964
rect 2136 -2976 2142 -2970
rect 2136 -2982 2142 -2976
rect 2136 -2988 2142 -2982
rect 2136 -2994 2142 -2988
rect 2136 -3000 2142 -2994
rect 2136 -3006 2142 -3000
rect 2136 -3012 2142 -3006
rect 2136 -3018 2142 -3012
rect 2136 -3024 2142 -3018
rect 2136 -3030 2142 -3024
rect 2136 -3036 2142 -3030
rect 2136 -3042 2142 -3036
rect 2136 -3048 2142 -3042
rect 2142 -270 2148 -264
rect 2142 -276 2148 -270
rect 2142 -282 2148 -276
rect 2142 -288 2148 -282
rect 2142 -294 2148 -288
rect 2142 -300 2148 -294
rect 2142 -306 2148 -300
rect 2142 -312 2148 -306
rect 2142 -318 2148 -312
rect 2142 -324 2148 -318
rect 2142 -330 2148 -324
rect 2142 -336 2148 -330
rect 2142 -342 2148 -336
rect 2142 -348 2148 -342
rect 2142 -354 2148 -348
rect 2142 -360 2148 -354
rect 2142 -366 2148 -360
rect 2142 -372 2148 -366
rect 2142 -378 2148 -372
rect 2142 -384 2148 -378
rect 2142 -390 2148 -384
rect 2142 -396 2148 -390
rect 2142 -402 2148 -396
rect 2142 -408 2148 -402
rect 2142 -414 2148 -408
rect 2142 -420 2148 -414
rect 2142 -426 2148 -420
rect 2142 -432 2148 -426
rect 2142 -438 2148 -432
rect 2142 -444 2148 -438
rect 2142 -450 2148 -444
rect 2142 -456 2148 -450
rect 2142 -462 2148 -456
rect 2142 -468 2148 -462
rect 2142 -474 2148 -468
rect 2142 -480 2148 -474
rect 2142 -486 2148 -480
rect 2142 -492 2148 -486
rect 2142 -498 2148 -492
rect 2142 -504 2148 -498
rect 2142 -510 2148 -504
rect 2142 -516 2148 -510
rect 2142 -522 2148 -516
rect 2142 -528 2148 -522
rect 2142 -534 2148 -528
rect 2142 -540 2148 -534
rect 2142 -546 2148 -540
rect 2142 -552 2148 -546
rect 2142 -558 2148 -552
rect 2142 -564 2148 -558
rect 2142 -570 2148 -564
rect 2142 -576 2148 -570
rect 2142 -582 2148 -576
rect 2142 -588 2148 -582
rect 2142 -594 2148 -588
rect 2142 -600 2148 -594
rect 2142 -606 2148 -600
rect 2142 -612 2148 -606
rect 2142 -618 2148 -612
rect 2142 -624 2148 -618
rect 2142 -630 2148 -624
rect 2142 -636 2148 -630
rect 2142 -642 2148 -636
rect 2142 -648 2148 -642
rect 2142 -654 2148 -648
rect 2142 -660 2148 -654
rect 2142 -666 2148 -660
rect 2142 -672 2148 -666
rect 2142 -678 2148 -672
rect 2142 -684 2148 -678
rect 2142 -690 2148 -684
rect 2142 -696 2148 -690
rect 2142 -702 2148 -696
rect 2142 -708 2148 -702
rect 2142 -714 2148 -708
rect 2142 -720 2148 -714
rect 2142 -726 2148 -720
rect 2142 -732 2148 -726
rect 2142 -738 2148 -732
rect 2142 -744 2148 -738
rect 2142 -750 2148 -744
rect 2142 -756 2148 -750
rect 2142 -762 2148 -756
rect 2142 -768 2148 -762
rect 2142 -774 2148 -768
rect 2142 -780 2148 -774
rect 2142 -786 2148 -780
rect 2142 -792 2148 -786
rect 2142 -798 2148 -792
rect 2142 -804 2148 -798
rect 2142 -810 2148 -804
rect 2142 -816 2148 -810
rect 2142 -822 2148 -816
rect 2142 -828 2148 -822
rect 2142 -834 2148 -828
rect 2142 -840 2148 -834
rect 2142 -846 2148 -840
rect 2142 -852 2148 -846
rect 2142 -858 2148 -852
rect 2142 -864 2148 -858
rect 2142 -870 2148 -864
rect 2142 -876 2148 -870
rect 2142 -882 2148 -876
rect 2142 -888 2148 -882
rect 2142 -894 2148 -888
rect 2142 -900 2148 -894
rect 2142 -906 2148 -900
rect 2142 -912 2148 -906
rect 2142 -918 2148 -912
rect 2142 -924 2148 -918
rect 2142 -930 2148 -924
rect 2142 -936 2148 -930
rect 2142 -942 2148 -936
rect 2142 -948 2148 -942
rect 2142 -954 2148 -948
rect 2142 -960 2148 -954
rect 2142 -966 2148 -960
rect 2142 -972 2148 -966
rect 2142 -978 2148 -972
rect 2142 -984 2148 -978
rect 2142 -990 2148 -984
rect 2142 -996 2148 -990
rect 2142 -1002 2148 -996
rect 2142 -1008 2148 -1002
rect 2142 -1014 2148 -1008
rect 2142 -1020 2148 -1014
rect 2142 -1026 2148 -1020
rect 2142 -1032 2148 -1026
rect 2142 -1038 2148 -1032
rect 2142 -1044 2148 -1038
rect 2142 -1050 2148 -1044
rect 2142 -1056 2148 -1050
rect 2142 -1062 2148 -1056
rect 2142 -1068 2148 -1062
rect 2142 -1074 2148 -1068
rect 2142 -1080 2148 -1074
rect 2142 -1086 2148 -1080
rect 2142 -1092 2148 -1086
rect 2142 -1098 2148 -1092
rect 2142 -1104 2148 -1098
rect 2142 -1110 2148 -1104
rect 2142 -1116 2148 -1110
rect 2142 -1122 2148 -1116
rect 2142 -1128 2148 -1122
rect 2142 -1134 2148 -1128
rect 2142 -1140 2148 -1134
rect 2142 -1146 2148 -1140
rect 2142 -1152 2148 -1146
rect 2142 -1158 2148 -1152
rect 2142 -1164 2148 -1158
rect 2142 -1170 2148 -1164
rect 2142 -1176 2148 -1170
rect 2142 -1182 2148 -1176
rect 2142 -1188 2148 -1182
rect 2142 -1194 2148 -1188
rect 2142 -1200 2148 -1194
rect 2142 -1206 2148 -1200
rect 2142 -1212 2148 -1206
rect 2142 -1218 2148 -1212
rect 2142 -1224 2148 -1218
rect 2142 -1230 2148 -1224
rect 2142 -1236 2148 -1230
rect 2142 -1242 2148 -1236
rect 2142 -1248 2148 -1242
rect 2142 -1254 2148 -1248
rect 2142 -1260 2148 -1254
rect 2142 -1266 2148 -1260
rect 2142 -1272 2148 -1266
rect 2142 -1278 2148 -1272
rect 2142 -1284 2148 -1278
rect 2142 -1290 2148 -1284
rect 2142 -1296 2148 -1290
rect 2142 -1302 2148 -1296
rect 2142 -1308 2148 -1302
rect 2142 -1314 2148 -1308
rect 2142 -1320 2148 -1314
rect 2142 -1326 2148 -1320
rect 2142 -1332 2148 -1326
rect 2142 -1338 2148 -1332
rect 2142 -1344 2148 -1338
rect 2142 -1350 2148 -1344
rect 2142 -1356 2148 -1350
rect 2142 -1362 2148 -1356
rect 2142 -1368 2148 -1362
rect 2142 -1374 2148 -1368
rect 2142 -1380 2148 -1374
rect 2142 -1386 2148 -1380
rect 2142 -1602 2148 -1596
rect 2142 -1608 2148 -1602
rect 2142 -1614 2148 -1608
rect 2142 -1620 2148 -1614
rect 2142 -1626 2148 -1620
rect 2142 -1632 2148 -1626
rect 2142 -1638 2148 -1632
rect 2142 -1644 2148 -1638
rect 2142 -1650 2148 -1644
rect 2142 -1656 2148 -1650
rect 2142 -1662 2148 -1656
rect 2142 -1668 2148 -1662
rect 2142 -1674 2148 -1668
rect 2142 -1680 2148 -1674
rect 2142 -1686 2148 -1680
rect 2142 -1692 2148 -1686
rect 2142 -1698 2148 -1692
rect 2142 -1704 2148 -1698
rect 2142 -1710 2148 -1704
rect 2142 -1716 2148 -1710
rect 2142 -1722 2148 -1716
rect 2142 -1728 2148 -1722
rect 2142 -1734 2148 -1728
rect 2142 -1740 2148 -1734
rect 2142 -1746 2148 -1740
rect 2142 -1752 2148 -1746
rect 2142 -1758 2148 -1752
rect 2142 -1764 2148 -1758
rect 2142 -1770 2148 -1764
rect 2142 -1776 2148 -1770
rect 2142 -1782 2148 -1776
rect 2142 -1788 2148 -1782
rect 2142 -1794 2148 -1788
rect 2142 -1800 2148 -1794
rect 2142 -1806 2148 -1800
rect 2142 -1812 2148 -1806
rect 2142 -1818 2148 -1812
rect 2142 -1824 2148 -1818
rect 2142 -1830 2148 -1824
rect 2142 -1836 2148 -1830
rect 2142 -1842 2148 -1836
rect 2142 -1848 2148 -1842
rect 2142 -1854 2148 -1848
rect 2142 -1860 2148 -1854
rect 2142 -1866 2148 -1860
rect 2142 -1872 2148 -1866
rect 2142 -1878 2148 -1872
rect 2142 -1884 2148 -1878
rect 2142 -1890 2148 -1884
rect 2142 -1896 2148 -1890
rect 2142 -1902 2148 -1896
rect 2142 -1908 2148 -1902
rect 2142 -1914 2148 -1908
rect 2142 -1920 2148 -1914
rect 2142 -1926 2148 -1920
rect 2142 -1932 2148 -1926
rect 2142 -1938 2148 -1932
rect 2142 -1944 2148 -1938
rect 2142 -1950 2148 -1944
rect 2142 -1956 2148 -1950
rect 2142 -1962 2148 -1956
rect 2142 -1968 2148 -1962
rect 2142 -1974 2148 -1968
rect 2142 -1980 2148 -1974
rect 2142 -1986 2148 -1980
rect 2142 -1992 2148 -1986
rect 2142 -1998 2148 -1992
rect 2142 -2004 2148 -1998
rect 2142 -2010 2148 -2004
rect 2142 -2016 2148 -2010
rect 2142 -2022 2148 -2016
rect 2142 -2028 2148 -2022
rect 2142 -2034 2148 -2028
rect 2142 -2040 2148 -2034
rect 2142 -2046 2148 -2040
rect 2142 -2052 2148 -2046
rect 2142 -2058 2148 -2052
rect 2142 -2064 2148 -2058
rect 2142 -2070 2148 -2064
rect 2142 -2076 2148 -2070
rect 2142 -2082 2148 -2076
rect 2142 -2088 2148 -2082
rect 2142 -2094 2148 -2088
rect 2142 -2100 2148 -2094
rect 2142 -2106 2148 -2100
rect 2142 -2112 2148 -2106
rect 2142 -2118 2148 -2112
rect 2142 -2124 2148 -2118
rect 2142 -2130 2148 -2124
rect 2142 -2136 2148 -2130
rect 2142 -2142 2148 -2136
rect 2142 -2148 2148 -2142
rect 2142 -2154 2148 -2148
rect 2142 -2160 2148 -2154
rect 2142 -2166 2148 -2160
rect 2142 -2172 2148 -2166
rect 2142 -2178 2148 -2172
rect 2142 -2184 2148 -2178
rect 2142 -2190 2148 -2184
rect 2142 -2196 2148 -2190
rect 2142 -2202 2148 -2196
rect 2142 -2208 2148 -2202
rect 2142 -2214 2148 -2208
rect 2142 -2220 2148 -2214
rect 2142 -2226 2148 -2220
rect 2142 -2232 2148 -2226
rect 2142 -2238 2148 -2232
rect 2142 -2244 2148 -2238
rect 2142 -2250 2148 -2244
rect 2142 -2256 2148 -2250
rect 2142 -2262 2148 -2256
rect 2142 -2268 2148 -2262
rect 2142 -2274 2148 -2268
rect 2142 -2280 2148 -2274
rect 2142 -2286 2148 -2280
rect 2142 -2292 2148 -2286
rect 2142 -2298 2148 -2292
rect 2142 -2304 2148 -2298
rect 2142 -2310 2148 -2304
rect 2142 -2316 2148 -2310
rect 2142 -2322 2148 -2316
rect 2142 -2328 2148 -2322
rect 2142 -2334 2148 -2328
rect 2142 -2340 2148 -2334
rect 2142 -2346 2148 -2340
rect 2142 -2352 2148 -2346
rect 2142 -2358 2148 -2352
rect 2142 -2364 2148 -2358
rect 2142 -2370 2148 -2364
rect 2142 -2376 2148 -2370
rect 2142 -2382 2148 -2376
rect 2142 -2388 2148 -2382
rect 2142 -2394 2148 -2388
rect 2142 -2400 2148 -2394
rect 2142 -2406 2148 -2400
rect 2142 -2412 2148 -2406
rect 2142 -2556 2148 -2550
rect 2142 -2562 2148 -2556
rect 2142 -2568 2148 -2562
rect 2142 -2574 2148 -2568
rect 2142 -2580 2148 -2574
rect 2142 -2586 2148 -2580
rect 2142 -2592 2148 -2586
rect 2142 -2598 2148 -2592
rect 2142 -2604 2148 -2598
rect 2142 -2610 2148 -2604
rect 2142 -2616 2148 -2610
rect 2142 -2622 2148 -2616
rect 2142 -2628 2148 -2622
rect 2142 -2634 2148 -2628
rect 2142 -2640 2148 -2634
rect 2142 -2646 2148 -2640
rect 2142 -2652 2148 -2646
rect 2142 -2658 2148 -2652
rect 2142 -2664 2148 -2658
rect 2142 -2670 2148 -2664
rect 2142 -2676 2148 -2670
rect 2142 -2682 2148 -2676
rect 2142 -2688 2148 -2682
rect 2142 -2694 2148 -2688
rect 2142 -2700 2148 -2694
rect 2142 -2706 2148 -2700
rect 2142 -2712 2148 -2706
rect 2142 -2718 2148 -2712
rect 2142 -2724 2148 -2718
rect 2142 -2730 2148 -2724
rect 2142 -2736 2148 -2730
rect 2142 -2742 2148 -2736
rect 2142 -2748 2148 -2742
rect 2142 -2754 2148 -2748
rect 2142 -2760 2148 -2754
rect 2142 -2766 2148 -2760
rect 2142 -2772 2148 -2766
rect 2142 -2778 2148 -2772
rect 2142 -2784 2148 -2778
rect 2142 -2790 2148 -2784
rect 2142 -2796 2148 -2790
rect 2142 -2802 2148 -2796
rect 2142 -2808 2148 -2802
rect 2142 -2814 2148 -2808
rect 2142 -2820 2148 -2814
rect 2142 -2826 2148 -2820
rect 2142 -2832 2148 -2826
rect 2142 -2838 2148 -2832
rect 2142 -2844 2148 -2838
rect 2142 -2850 2148 -2844
rect 2142 -2856 2148 -2850
rect 2142 -2862 2148 -2856
rect 2142 -2868 2148 -2862
rect 2142 -2874 2148 -2868
rect 2142 -2880 2148 -2874
rect 2142 -2886 2148 -2880
rect 2142 -2892 2148 -2886
rect 2142 -2898 2148 -2892
rect 2142 -2904 2148 -2898
rect 2142 -2910 2148 -2904
rect 2142 -2916 2148 -2910
rect 2142 -2922 2148 -2916
rect 2142 -2928 2148 -2922
rect 2142 -2934 2148 -2928
rect 2142 -2940 2148 -2934
rect 2142 -2946 2148 -2940
rect 2142 -2952 2148 -2946
rect 2142 -2958 2148 -2952
rect 2142 -2964 2148 -2958
rect 2142 -2970 2148 -2964
rect 2142 -2976 2148 -2970
rect 2142 -2982 2148 -2976
rect 2142 -2988 2148 -2982
rect 2142 -2994 2148 -2988
rect 2142 -3000 2148 -2994
rect 2142 -3006 2148 -3000
rect 2142 -3012 2148 -3006
rect 2142 -3018 2148 -3012
rect 2142 -3024 2148 -3018
rect 2142 -3030 2148 -3024
rect 2142 -3036 2148 -3030
rect 2142 -3042 2148 -3036
rect 2148 -264 2154 -258
rect 2148 -270 2154 -264
rect 2148 -276 2154 -270
rect 2148 -282 2154 -276
rect 2148 -288 2154 -282
rect 2148 -294 2154 -288
rect 2148 -300 2154 -294
rect 2148 -306 2154 -300
rect 2148 -312 2154 -306
rect 2148 -318 2154 -312
rect 2148 -324 2154 -318
rect 2148 -330 2154 -324
rect 2148 -336 2154 -330
rect 2148 -342 2154 -336
rect 2148 -348 2154 -342
rect 2148 -354 2154 -348
rect 2148 -360 2154 -354
rect 2148 -366 2154 -360
rect 2148 -372 2154 -366
rect 2148 -378 2154 -372
rect 2148 -384 2154 -378
rect 2148 -390 2154 -384
rect 2148 -396 2154 -390
rect 2148 -402 2154 -396
rect 2148 -408 2154 -402
rect 2148 -414 2154 -408
rect 2148 -420 2154 -414
rect 2148 -426 2154 -420
rect 2148 -432 2154 -426
rect 2148 -438 2154 -432
rect 2148 -444 2154 -438
rect 2148 -450 2154 -444
rect 2148 -456 2154 -450
rect 2148 -462 2154 -456
rect 2148 -468 2154 -462
rect 2148 -474 2154 -468
rect 2148 -480 2154 -474
rect 2148 -486 2154 -480
rect 2148 -492 2154 -486
rect 2148 -498 2154 -492
rect 2148 -504 2154 -498
rect 2148 -510 2154 -504
rect 2148 -516 2154 -510
rect 2148 -522 2154 -516
rect 2148 -528 2154 -522
rect 2148 -534 2154 -528
rect 2148 -540 2154 -534
rect 2148 -546 2154 -540
rect 2148 -552 2154 -546
rect 2148 -558 2154 -552
rect 2148 -564 2154 -558
rect 2148 -570 2154 -564
rect 2148 -576 2154 -570
rect 2148 -582 2154 -576
rect 2148 -588 2154 -582
rect 2148 -594 2154 -588
rect 2148 -600 2154 -594
rect 2148 -606 2154 -600
rect 2148 -612 2154 -606
rect 2148 -618 2154 -612
rect 2148 -624 2154 -618
rect 2148 -630 2154 -624
rect 2148 -636 2154 -630
rect 2148 -642 2154 -636
rect 2148 -648 2154 -642
rect 2148 -654 2154 -648
rect 2148 -660 2154 -654
rect 2148 -666 2154 -660
rect 2148 -672 2154 -666
rect 2148 -678 2154 -672
rect 2148 -684 2154 -678
rect 2148 -690 2154 -684
rect 2148 -696 2154 -690
rect 2148 -702 2154 -696
rect 2148 -708 2154 -702
rect 2148 -714 2154 -708
rect 2148 -720 2154 -714
rect 2148 -726 2154 -720
rect 2148 -732 2154 -726
rect 2148 -738 2154 -732
rect 2148 -744 2154 -738
rect 2148 -750 2154 -744
rect 2148 -756 2154 -750
rect 2148 -762 2154 -756
rect 2148 -768 2154 -762
rect 2148 -774 2154 -768
rect 2148 -780 2154 -774
rect 2148 -786 2154 -780
rect 2148 -792 2154 -786
rect 2148 -798 2154 -792
rect 2148 -804 2154 -798
rect 2148 -810 2154 -804
rect 2148 -816 2154 -810
rect 2148 -822 2154 -816
rect 2148 -828 2154 -822
rect 2148 -834 2154 -828
rect 2148 -840 2154 -834
rect 2148 -846 2154 -840
rect 2148 -852 2154 -846
rect 2148 -858 2154 -852
rect 2148 -864 2154 -858
rect 2148 -870 2154 -864
rect 2148 -876 2154 -870
rect 2148 -882 2154 -876
rect 2148 -888 2154 -882
rect 2148 -894 2154 -888
rect 2148 -900 2154 -894
rect 2148 -906 2154 -900
rect 2148 -912 2154 -906
rect 2148 -918 2154 -912
rect 2148 -924 2154 -918
rect 2148 -930 2154 -924
rect 2148 -936 2154 -930
rect 2148 -942 2154 -936
rect 2148 -948 2154 -942
rect 2148 -954 2154 -948
rect 2148 -960 2154 -954
rect 2148 -966 2154 -960
rect 2148 -972 2154 -966
rect 2148 -978 2154 -972
rect 2148 -984 2154 -978
rect 2148 -990 2154 -984
rect 2148 -996 2154 -990
rect 2148 -1002 2154 -996
rect 2148 -1008 2154 -1002
rect 2148 -1014 2154 -1008
rect 2148 -1020 2154 -1014
rect 2148 -1026 2154 -1020
rect 2148 -1032 2154 -1026
rect 2148 -1038 2154 -1032
rect 2148 -1044 2154 -1038
rect 2148 -1050 2154 -1044
rect 2148 -1056 2154 -1050
rect 2148 -1062 2154 -1056
rect 2148 -1068 2154 -1062
rect 2148 -1074 2154 -1068
rect 2148 -1080 2154 -1074
rect 2148 -1086 2154 -1080
rect 2148 -1092 2154 -1086
rect 2148 -1098 2154 -1092
rect 2148 -1104 2154 -1098
rect 2148 -1110 2154 -1104
rect 2148 -1116 2154 -1110
rect 2148 -1122 2154 -1116
rect 2148 -1128 2154 -1122
rect 2148 -1134 2154 -1128
rect 2148 -1140 2154 -1134
rect 2148 -1146 2154 -1140
rect 2148 -1152 2154 -1146
rect 2148 -1158 2154 -1152
rect 2148 -1164 2154 -1158
rect 2148 -1170 2154 -1164
rect 2148 -1176 2154 -1170
rect 2148 -1182 2154 -1176
rect 2148 -1188 2154 -1182
rect 2148 -1194 2154 -1188
rect 2148 -1200 2154 -1194
rect 2148 -1206 2154 -1200
rect 2148 -1212 2154 -1206
rect 2148 -1218 2154 -1212
rect 2148 -1224 2154 -1218
rect 2148 -1230 2154 -1224
rect 2148 -1236 2154 -1230
rect 2148 -1242 2154 -1236
rect 2148 -1248 2154 -1242
rect 2148 -1254 2154 -1248
rect 2148 -1260 2154 -1254
rect 2148 -1266 2154 -1260
rect 2148 -1272 2154 -1266
rect 2148 -1278 2154 -1272
rect 2148 -1284 2154 -1278
rect 2148 -1290 2154 -1284
rect 2148 -1296 2154 -1290
rect 2148 -1302 2154 -1296
rect 2148 -1308 2154 -1302
rect 2148 -1314 2154 -1308
rect 2148 -1320 2154 -1314
rect 2148 -1326 2154 -1320
rect 2148 -1332 2154 -1326
rect 2148 -1338 2154 -1332
rect 2148 -1344 2154 -1338
rect 2148 -1350 2154 -1344
rect 2148 -1356 2154 -1350
rect 2148 -1362 2154 -1356
rect 2148 -1368 2154 -1362
rect 2148 -1596 2154 -1590
rect 2148 -1602 2154 -1596
rect 2148 -1608 2154 -1602
rect 2148 -1614 2154 -1608
rect 2148 -1620 2154 -1614
rect 2148 -1626 2154 -1620
rect 2148 -1632 2154 -1626
rect 2148 -1638 2154 -1632
rect 2148 -1644 2154 -1638
rect 2148 -1650 2154 -1644
rect 2148 -1656 2154 -1650
rect 2148 -1662 2154 -1656
rect 2148 -1668 2154 -1662
rect 2148 -1674 2154 -1668
rect 2148 -1680 2154 -1674
rect 2148 -1686 2154 -1680
rect 2148 -1692 2154 -1686
rect 2148 -1698 2154 -1692
rect 2148 -1704 2154 -1698
rect 2148 -1710 2154 -1704
rect 2148 -1716 2154 -1710
rect 2148 -1722 2154 -1716
rect 2148 -1728 2154 -1722
rect 2148 -1734 2154 -1728
rect 2148 -1740 2154 -1734
rect 2148 -1746 2154 -1740
rect 2148 -1752 2154 -1746
rect 2148 -1758 2154 -1752
rect 2148 -1764 2154 -1758
rect 2148 -1770 2154 -1764
rect 2148 -1776 2154 -1770
rect 2148 -1782 2154 -1776
rect 2148 -1788 2154 -1782
rect 2148 -1794 2154 -1788
rect 2148 -1800 2154 -1794
rect 2148 -1806 2154 -1800
rect 2148 -1812 2154 -1806
rect 2148 -1818 2154 -1812
rect 2148 -1824 2154 -1818
rect 2148 -1830 2154 -1824
rect 2148 -1836 2154 -1830
rect 2148 -1842 2154 -1836
rect 2148 -1848 2154 -1842
rect 2148 -1854 2154 -1848
rect 2148 -1860 2154 -1854
rect 2148 -1866 2154 -1860
rect 2148 -1872 2154 -1866
rect 2148 -1878 2154 -1872
rect 2148 -1884 2154 -1878
rect 2148 -1890 2154 -1884
rect 2148 -1896 2154 -1890
rect 2148 -1902 2154 -1896
rect 2148 -1908 2154 -1902
rect 2148 -1914 2154 -1908
rect 2148 -1920 2154 -1914
rect 2148 -1926 2154 -1920
rect 2148 -1932 2154 -1926
rect 2148 -1938 2154 -1932
rect 2148 -1944 2154 -1938
rect 2148 -1950 2154 -1944
rect 2148 -1956 2154 -1950
rect 2148 -1962 2154 -1956
rect 2148 -1968 2154 -1962
rect 2148 -1974 2154 -1968
rect 2148 -1980 2154 -1974
rect 2148 -1986 2154 -1980
rect 2148 -1992 2154 -1986
rect 2148 -1998 2154 -1992
rect 2148 -2004 2154 -1998
rect 2148 -2010 2154 -2004
rect 2148 -2016 2154 -2010
rect 2148 -2022 2154 -2016
rect 2148 -2028 2154 -2022
rect 2148 -2034 2154 -2028
rect 2148 -2040 2154 -2034
rect 2148 -2046 2154 -2040
rect 2148 -2052 2154 -2046
rect 2148 -2058 2154 -2052
rect 2148 -2064 2154 -2058
rect 2148 -2070 2154 -2064
rect 2148 -2076 2154 -2070
rect 2148 -2082 2154 -2076
rect 2148 -2088 2154 -2082
rect 2148 -2094 2154 -2088
rect 2148 -2100 2154 -2094
rect 2148 -2106 2154 -2100
rect 2148 -2112 2154 -2106
rect 2148 -2118 2154 -2112
rect 2148 -2124 2154 -2118
rect 2148 -2130 2154 -2124
rect 2148 -2136 2154 -2130
rect 2148 -2142 2154 -2136
rect 2148 -2148 2154 -2142
rect 2148 -2154 2154 -2148
rect 2148 -2160 2154 -2154
rect 2148 -2166 2154 -2160
rect 2148 -2172 2154 -2166
rect 2148 -2178 2154 -2172
rect 2148 -2184 2154 -2178
rect 2148 -2190 2154 -2184
rect 2148 -2196 2154 -2190
rect 2148 -2202 2154 -2196
rect 2148 -2208 2154 -2202
rect 2148 -2214 2154 -2208
rect 2148 -2220 2154 -2214
rect 2148 -2226 2154 -2220
rect 2148 -2232 2154 -2226
rect 2148 -2238 2154 -2232
rect 2148 -2244 2154 -2238
rect 2148 -2250 2154 -2244
rect 2148 -2256 2154 -2250
rect 2148 -2262 2154 -2256
rect 2148 -2268 2154 -2262
rect 2148 -2274 2154 -2268
rect 2148 -2280 2154 -2274
rect 2148 -2286 2154 -2280
rect 2148 -2292 2154 -2286
rect 2148 -2298 2154 -2292
rect 2148 -2304 2154 -2298
rect 2148 -2310 2154 -2304
rect 2148 -2316 2154 -2310
rect 2148 -2322 2154 -2316
rect 2148 -2328 2154 -2322
rect 2148 -2334 2154 -2328
rect 2148 -2340 2154 -2334
rect 2148 -2346 2154 -2340
rect 2148 -2352 2154 -2346
rect 2148 -2358 2154 -2352
rect 2148 -2364 2154 -2358
rect 2148 -2370 2154 -2364
rect 2148 -2376 2154 -2370
rect 2148 -2382 2154 -2376
rect 2148 -2388 2154 -2382
rect 2148 -2394 2154 -2388
rect 2148 -2400 2154 -2394
rect 2148 -2406 2154 -2400
rect 2148 -2556 2154 -2550
rect 2148 -2562 2154 -2556
rect 2148 -2568 2154 -2562
rect 2148 -2574 2154 -2568
rect 2148 -2580 2154 -2574
rect 2148 -2586 2154 -2580
rect 2148 -2592 2154 -2586
rect 2148 -2598 2154 -2592
rect 2148 -2604 2154 -2598
rect 2148 -2610 2154 -2604
rect 2148 -2616 2154 -2610
rect 2148 -2622 2154 -2616
rect 2148 -2628 2154 -2622
rect 2148 -2634 2154 -2628
rect 2148 -2640 2154 -2634
rect 2148 -2646 2154 -2640
rect 2148 -2652 2154 -2646
rect 2148 -2658 2154 -2652
rect 2148 -2664 2154 -2658
rect 2148 -2670 2154 -2664
rect 2148 -2676 2154 -2670
rect 2148 -2682 2154 -2676
rect 2148 -2688 2154 -2682
rect 2148 -2694 2154 -2688
rect 2148 -2700 2154 -2694
rect 2148 -2706 2154 -2700
rect 2148 -2712 2154 -2706
rect 2148 -2718 2154 -2712
rect 2148 -2724 2154 -2718
rect 2148 -2730 2154 -2724
rect 2148 -2736 2154 -2730
rect 2148 -2742 2154 -2736
rect 2148 -2748 2154 -2742
rect 2148 -2754 2154 -2748
rect 2148 -2760 2154 -2754
rect 2148 -2766 2154 -2760
rect 2148 -2772 2154 -2766
rect 2148 -2778 2154 -2772
rect 2148 -2784 2154 -2778
rect 2148 -2790 2154 -2784
rect 2148 -2796 2154 -2790
rect 2148 -2802 2154 -2796
rect 2148 -2808 2154 -2802
rect 2148 -2814 2154 -2808
rect 2148 -2820 2154 -2814
rect 2148 -2826 2154 -2820
rect 2148 -2832 2154 -2826
rect 2148 -2838 2154 -2832
rect 2148 -2844 2154 -2838
rect 2148 -2850 2154 -2844
rect 2148 -2856 2154 -2850
rect 2148 -2862 2154 -2856
rect 2148 -2868 2154 -2862
rect 2148 -2874 2154 -2868
rect 2148 -2880 2154 -2874
rect 2148 -2886 2154 -2880
rect 2148 -2892 2154 -2886
rect 2148 -2898 2154 -2892
rect 2148 -2904 2154 -2898
rect 2148 -2910 2154 -2904
rect 2148 -2916 2154 -2910
rect 2148 -2922 2154 -2916
rect 2148 -2928 2154 -2922
rect 2148 -2934 2154 -2928
rect 2148 -2940 2154 -2934
rect 2148 -2946 2154 -2940
rect 2148 -2952 2154 -2946
rect 2148 -2958 2154 -2952
rect 2148 -2964 2154 -2958
rect 2148 -2970 2154 -2964
rect 2148 -2976 2154 -2970
rect 2148 -2982 2154 -2976
rect 2148 -2988 2154 -2982
rect 2148 -2994 2154 -2988
rect 2148 -3000 2154 -2994
rect 2148 -3006 2154 -3000
rect 2148 -3012 2154 -3006
rect 2148 -3018 2154 -3012
rect 2148 -3024 2154 -3018
rect 2148 -3030 2154 -3024
rect 2148 -3036 2154 -3030
rect 2154 -258 2160 -252
rect 2154 -264 2160 -258
rect 2154 -270 2160 -264
rect 2154 -276 2160 -270
rect 2154 -282 2160 -276
rect 2154 -288 2160 -282
rect 2154 -294 2160 -288
rect 2154 -300 2160 -294
rect 2154 -306 2160 -300
rect 2154 -312 2160 -306
rect 2154 -318 2160 -312
rect 2154 -324 2160 -318
rect 2154 -330 2160 -324
rect 2154 -336 2160 -330
rect 2154 -342 2160 -336
rect 2154 -348 2160 -342
rect 2154 -354 2160 -348
rect 2154 -360 2160 -354
rect 2154 -366 2160 -360
rect 2154 -372 2160 -366
rect 2154 -378 2160 -372
rect 2154 -384 2160 -378
rect 2154 -390 2160 -384
rect 2154 -396 2160 -390
rect 2154 -402 2160 -396
rect 2154 -408 2160 -402
rect 2154 -414 2160 -408
rect 2154 -420 2160 -414
rect 2154 -426 2160 -420
rect 2154 -432 2160 -426
rect 2154 -438 2160 -432
rect 2154 -444 2160 -438
rect 2154 -450 2160 -444
rect 2154 -456 2160 -450
rect 2154 -462 2160 -456
rect 2154 -468 2160 -462
rect 2154 -474 2160 -468
rect 2154 -480 2160 -474
rect 2154 -486 2160 -480
rect 2154 -492 2160 -486
rect 2154 -498 2160 -492
rect 2154 -504 2160 -498
rect 2154 -510 2160 -504
rect 2154 -516 2160 -510
rect 2154 -522 2160 -516
rect 2154 -528 2160 -522
rect 2154 -534 2160 -528
rect 2154 -540 2160 -534
rect 2154 -546 2160 -540
rect 2154 -552 2160 -546
rect 2154 -558 2160 -552
rect 2154 -564 2160 -558
rect 2154 -570 2160 -564
rect 2154 -576 2160 -570
rect 2154 -582 2160 -576
rect 2154 -588 2160 -582
rect 2154 -594 2160 -588
rect 2154 -600 2160 -594
rect 2154 -606 2160 -600
rect 2154 -612 2160 -606
rect 2154 -618 2160 -612
rect 2154 -624 2160 -618
rect 2154 -630 2160 -624
rect 2154 -636 2160 -630
rect 2154 -642 2160 -636
rect 2154 -648 2160 -642
rect 2154 -654 2160 -648
rect 2154 -660 2160 -654
rect 2154 -666 2160 -660
rect 2154 -672 2160 -666
rect 2154 -678 2160 -672
rect 2154 -684 2160 -678
rect 2154 -690 2160 -684
rect 2154 -696 2160 -690
rect 2154 -702 2160 -696
rect 2154 -708 2160 -702
rect 2154 -714 2160 -708
rect 2154 -720 2160 -714
rect 2154 -726 2160 -720
rect 2154 -732 2160 -726
rect 2154 -738 2160 -732
rect 2154 -744 2160 -738
rect 2154 -750 2160 -744
rect 2154 -756 2160 -750
rect 2154 -762 2160 -756
rect 2154 -768 2160 -762
rect 2154 -774 2160 -768
rect 2154 -780 2160 -774
rect 2154 -786 2160 -780
rect 2154 -792 2160 -786
rect 2154 -798 2160 -792
rect 2154 -804 2160 -798
rect 2154 -810 2160 -804
rect 2154 -816 2160 -810
rect 2154 -822 2160 -816
rect 2154 -828 2160 -822
rect 2154 -834 2160 -828
rect 2154 -840 2160 -834
rect 2154 -846 2160 -840
rect 2154 -852 2160 -846
rect 2154 -858 2160 -852
rect 2154 -864 2160 -858
rect 2154 -870 2160 -864
rect 2154 -876 2160 -870
rect 2154 -882 2160 -876
rect 2154 -888 2160 -882
rect 2154 -894 2160 -888
rect 2154 -900 2160 -894
rect 2154 -906 2160 -900
rect 2154 -912 2160 -906
rect 2154 -918 2160 -912
rect 2154 -924 2160 -918
rect 2154 -930 2160 -924
rect 2154 -936 2160 -930
rect 2154 -942 2160 -936
rect 2154 -948 2160 -942
rect 2154 -954 2160 -948
rect 2154 -960 2160 -954
rect 2154 -966 2160 -960
rect 2154 -972 2160 -966
rect 2154 -978 2160 -972
rect 2154 -984 2160 -978
rect 2154 -990 2160 -984
rect 2154 -996 2160 -990
rect 2154 -1002 2160 -996
rect 2154 -1008 2160 -1002
rect 2154 -1014 2160 -1008
rect 2154 -1020 2160 -1014
rect 2154 -1026 2160 -1020
rect 2154 -1032 2160 -1026
rect 2154 -1038 2160 -1032
rect 2154 -1044 2160 -1038
rect 2154 -1050 2160 -1044
rect 2154 -1056 2160 -1050
rect 2154 -1062 2160 -1056
rect 2154 -1068 2160 -1062
rect 2154 -1074 2160 -1068
rect 2154 -1080 2160 -1074
rect 2154 -1086 2160 -1080
rect 2154 -1092 2160 -1086
rect 2154 -1098 2160 -1092
rect 2154 -1104 2160 -1098
rect 2154 -1110 2160 -1104
rect 2154 -1116 2160 -1110
rect 2154 -1122 2160 -1116
rect 2154 -1128 2160 -1122
rect 2154 -1134 2160 -1128
rect 2154 -1140 2160 -1134
rect 2154 -1146 2160 -1140
rect 2154 -1152 2160 -1146
rect 2154 -1158 2160 -1152
rect 2154 -1164 2160 -1158
rect 2154 -1170 2160 -1164
rect 2154 -1176 2160 -1170
rect 2154 -1182 2160 -1176
rect 2154 -1188 2160 -1182
rect 2154 -1194 2160 -1188
rect 2154 -1200 2160 -1194
rect 2154 -1206 2160 -1200
rect 2154 -1212 2160 -1206
rect 2154 -1218 2160 -1212
rect 2154 -1224 2160 -1218
rect 2154 -1230 2160 -1224
rect 2154 -1236 2160 -1230
rect 2154 -1242 2160 -1236
rect 2154 -1248 2160 -1242
rect 2154 -1254 2160 -1248
rect 2154 -1260 2160 -1254
rect 2154 -1266 2160 -1260
rect 2154 -1272 2160 -1266
rect 2154 -1278 2160 -1272
rect 2154 -1284 2160 -1278
rect 2154 -1290 2160 -1284
rect 2154 -1296 2160 -1290
rect 2154 -1302 2160 -1296
rect 2154 -1308 2160 -1302
rect 2154 -1314 2160 -1308
rect 2154 -1320 2160 -1314
rect 2154 -1326 2160 -1320
rect 2154 -1332 2160 -1326
rect 2154 -1338 2160 -1332
rect 2154 -1344 2160 -1338
rect 2154 -1350 2160 -1344
rect 2154 -1356 2160 -1350
rect 2154 -1596 2160 -1590
rect 2154 -1602 2160 -1596
rect 2154 -1608 2160 -1602
rect 2154 -1614 2160 -1608
rect 2154 -1620 2160 -1614
rect 2154 -1626 2160 -1620
rect 2154 -1632 2160 -1626
rect 2154 -1638 2160 -1632
rect 2154 -1644 2160 -1638
rect 2154 -1650 2160 -1644
rect 2154 -1656 2160 -1650
rect 2154 -1662 2160 -1656
rect 2154 -1668 2160 -1662
rect 2154 -1674 2160 -1668
rect 2154 -1680 2160 -1674
rect 2154 -1686 2160 -1680
rect 2154 -1692 2160 -1686
rect 2154 -1698 2160 -1692
rect 2154 -1704 2160 -1698
rect 2154 -1710 2160 -1704
rect 2154 -1716 2160 -1710
rect 2154 -1722 2160 -1716
rect 2154 -1728 2160 -1722
rect 2154 -1734 2160 -1728
rect 2154 -1740 2160 -1734
rect 2154 -1746 2160 -1740
rect 2154 -1752 2160 -1746
rect 2154 -1758 2160 -1752
rect 2154 -1764 2160 -1758
rect 2154 -1770 2160 -1764
rect 2154 -1776 2160 -1770
rect 2154 -1782 2160 -1776
rect 2154 -1788 2160 -1782
rect 2154 -1794 2160 -1788
rect 2154 -1800 2160 -1794
rect 2154 -1806 2160 -1800
rect 2154 -1812 2160 -1806
rect 2154 -1818 2160 -1812
rect 2154 -1824 2160 -1818
rect 2154 -1830 2160 -1824
rect 2154 -1836 2160 -1830
rect 2154 -1842 2160 -1836
rect 2154 -1848 2160 -1842
rect 2154 -1854 2160 -1848
rect 2154 -1860 2160 -1854
rect 2154 -1866 2160 -1860
rect 2154 -1872 2160 -1866
rect 2154 -1878 2160 -1872
rect 2154 -1884 2160 -1878
rect 2154 -1890 2160 -1884
rect 2154 -1896 2160 -1890
rect 2154 -1902 2160 -1896
rect 2154 -1908 2160 -1902
rect 2154 -1914 2160 -1908
rect 2154 -1920 2160 -1914
rect 2154 -1926 2160 -1920
rect 2154 -1932 2160 -1926
rect 2154 -1938 2160 -1932
rect 2154 -1944 2160 -1938
rect 2154 -1950 2160 -1944
rect 2154 -1956 2160 -1950
rect 2154 -1962 2160 -1956
rect 2154 -1968 2160 -1962
rect 2154 -1974 2160 -1968
rect 2154 -1980 2160 -1974
rect 2154 -1986 2160 -1980
rect 2154 -1992 2160 -1986
rect 2154 -1998 2160 -1992
rect 2154 -2004 2160 -1998
rect 2154 -2010 2160 -2004
rect 2154 -2016 2160 -2010
rect 2154 -2022 2160 -2016
rect 2154 -2028 2160 -2022
rect 2154 -2034 2160 -2028
rect 2154 -2040 2160 -2034
rect 2154 -2046 2160 -2040
rect 2154 -2052 2160 -2046
rect 2154 -2058 2160 -2052
rect 2154 -2064 2160 -2058
rect 2154 -2070 2160 -2064
rect 2154 -2076 2160 -2070
rect 2154 -2082 2160 -2076
rect 2154 -2088 2160 -2082
rect 2154 -2094 2160 -2088
rect 2154 -2100 2160 -2094
rect 2154 -2106 2160 -2100
rect 2154 -2112 2160 -2106
rect 2154 -2118 2160 -2112
rect 2154 -2124 2160 -2118
rect 2154 -2130 2160 -2124
rect 2154 -2136 2160 -2130
rect 2154 -2142 2160 -2136
rect 2154 -2148 2160 -2142
rect 2154 -2154 2160 -2148
rect 2154 -2160 2160 -2154
rect 2154 -2166 2160 -2160
rect 2154 -2172 2160 -2166
rect 2154 -2178 2160 -2172
rect 2154 -2184 2160 -2178
rect 2154 -2190 2160 -2184
rect 2154 -2196 2160 -2190
rect 2154 -2202 2160 -2196
rect 2154 -2208 2160 -2202
rect 2154 -2214 2160 -2208
rect 2154 -2220 2160 -2214
rect 2154 -2226 2160 -2220
rect 2154 -2232 2160 -2226
rect 2154 -2238 2160 -2232
rect 2154 -2244 2160 -2238
rect 2154 -2250 2160 -2244
rect 2154 -2256 2160 -2250
rect 2154 -2262 2160 -2256
rect 2154 -2268 2160 -2262
rect 2154 -2274 2160 -2268
rect 2154 -2280 2160 -2274
rect 2154 -2286 2160 -2280
rect 2154 -2292 2160 -2286
rect 2154 -2298 2160 -2292
rect 2154 -2304 2160 -2298
rect 2154 -2310 2160 -2304
rect 2154 -2316 2160 -2310
rect 2154 -2322 2160 -2316
rect 2154 -2328 2160 -2322
rect 2154 -2334 2160 -2328
rect 2154 -2340 2160 -2334
rect 2154 -2346 2160 -2340
rect 2154 -2352 2160 -2346
rect 2154 -2358 2160 -2352
rect 2154 -2364 2160 -2358
rect 2154 -2370 2160 -2364
rect 2154 -2376 2160 -2370
rect 2154 -2382 2160 -2376
rect 2154 -2388 2160 -2382
rect 2154 -2394 2160 -2388
rect 2154 -2400 2160 -2394
rect 2154 -2556 2160 -2550
rect 2154 -2562 2160 -2556
rect 2154 -2568 2160 -2562
rect 2154 -2574 2160 -2568
rect 2154 -2580 2160 -2574
rect 2154 -2586 2160 -2580
rect 2154 -2592 2160 -2586
rect 2154 -2598 2160 -2592
rect 2154 -2604 2160 -2598
rect 2154 -2610 2160 -2604
rect 2154 -2616 2160 -2610
rect 2154 -2622 2160 -2616
rect 2154 -2628 2160 -2622
rect 2154 -2634 2160 -2628
rect 2154 -2640 2160 -2634
rect 2154 -2646 2160 -2640
rect 2154 -2652 2160 -2646
rect 2154 -2658 2160 -2652
rect 2154 -2664 2160 -2658
rect 2154 -2670 2160 -2664
rect 2154 -2676 2160 -2670
rect 2154 -2682 2160 -2676
rect 2154 -2688 2160 -2682
rect 2154 -2694 2160 -2688
rect 2154 -2700 2160 -2694
rect 2154 -2706 2160 -2700
rect 2154 -2712 2160 -2706
rect 2154 -2718 2160 -2712
rect 2154 -2724 2160 -2718
rect 2154 -2730 2160 -2724
rect 2154 -2736 2160 -2730
rect 2154 -2742 2160 -2736
rect 2154 -2748 2160 -2742
rect 2154 -2754 2160 -2748
rect 2154 -2760 2160 -2754
rect 2154 -2766 2160 -2760
rect 2154 -2772 2160 -2766
rect 2154 -2778 2160 -2772
rect 2154 -2784 2160 -2778
rect 2154 -2790 2160 -2784
rect 2154 -2796 2160 -2790
rect 2154 -2802 2160 -2796
rect 2154 -2808 2160 -2802
rect 2154 -2814 2160 -2808
rect 2154 -2820 2160 -2814
rect 2154 -2826 2160 -2820
rect 2154 -2832 2160 -2826
rect 2154 -2838 2160 -2832
rect 2154 -2844 2160 -2838
rect 2154 -2850 2160 -2844
rect 2154 -2856 2160 -2850
rect 2154 -2862 2160 -2856
rect 2154 -2868 2160 -2862
rect 2154 -2874 2160 -2868
rect 2154 -2880 2160 -2874
rect 2154 -2886 2160 -2880
rect 2154 -2892 2160 -2886
rect 2154 -2898 2160 -2892
rect 2154 -2904 2160 -2898
rect 2154 -2910 2160 -2904
rect 2154 -2916 2160 -2910
rect 2154 -2922 2160 -2916
rect 2154 -2928 2160 -2922
rect 2154 -2934 2160 -2928
rect 2154 -2940 2160 -2934
rect 2154 -2946 2160 -2940
rect 2154 -2952 2160 -2946
rect 2154 -2958 2160 -2952
rect 2154 -2964 2160 -2958
rect 2154 -2970 2160 -2964
rect 2154 -2976 2160 -2970
rect 2154 -2982 2160 -2976
rect 2154 -2988 2160 -2982
rect 2154 -2994 2160 -2988
rect 2154 -3000 2160 -2994
rect 2154 -3006 2160 -3000
rect 2154 -3012 2160 -3006
rect 2154 -3018 2160 -3012
rect 2154 -3024 2160 -3018
rect 2154 -3030 2160 -3024
rect 2154 -3036 2160 -3030
rect 2160 -246 2166 -240
rect 2160 -252 2166 -246
rect 2160 -258 2166 -252
rect 2160 -264 2166 -258
rect 2160 -270 2166 -264
rect 2160 -276 2166 -270
rect 2160 -282 2166 -276
rect 2160 -288 2166 -282
rect 2160 -294 2166 -288
rect 2160 -300 2166 -294
rect 2160 -306 2166 -300
rect 2160 -312 2166 -306
rect 2160 -318 2166 -312
rect 2160 -324 2166 -318
rect 2160 -330 2166 -324
rect 2160 -336 2166 -330
rect 2160 -342 2166 -336
rect 2160 -348 2166 -342
rect 2160 -354 2166 -348
rect 2160 -360 2166 -354
rect 2160 -366 2166 -360
rect 2160 -372 2166 -366
rect 2160 -378 2166 -372
rect 2160 -384 2166 -378
rect 2160 -390 2166 -384
rect 2160 -396 2166 -390
rect 2160 -402 2166 -396
rect 2160 -408 2166 -402
rect 2160 -414 2166 -408
rect 2160 -420 2166 -414
rect 2160 -426 2166 -420
rect 2160 -432 2166 -426
rect 2160 -438 2166 -432
rect 2160 -444 2166 -438
rect 2160 -450 2166 -444
rect 2160 -456 2166 -450
rect 2160 -462 2166 -456
rect 2160 -468 2166 -462
rect 2160 -474 2166 -468
rect 2160 -480 2166 -474
rect 2160 -486 2166 -480
rect 2160 -492 2166 -486
rect 2160 -498 2166 -492
rect 2160 -504 2166 -498
rect 2160 -510 2166 -504
rect 2160 -516 2166 -510
rect 2160 -522 2166 -516
rect 2160 -528 2166 -522
rect 2160 -534 2166 -528
rect 2160 -540 2166 -534
rect 2160 -546 2166 -540
rect 2160 -552 2166 -546
rect 2160 -558 2166 -552
rect 2160 -564 2166 -558
rect 2160 -570 2166 -564
rect 2160 -576 2166 -570
rect 2160 -582 2166 -576
rect 2160 -588 2166 -582
rect 2160 -594 2166 -588
rect 2160 -600 2166 -594
rect 2160 -606 2166 -600
rect 2160 -612 2166 -606
rect 2160 -618 2166 -612
rect 2160 -624 2166 -618
rect 2160 -630 2166 -624
rect 2160 -636 2166 -630
rect 2160 -642 2166 -636
rect 2160 -648 2166 -642
rect 2160 -654 2166 -648
rect 2160 -660 2166 -654
rect 2160 -666 2166 -660
rect 2160 -672 2166 -666
rect 2160 -678 2166 -672
rect 2160 -684 2166 -678
rect 2160 -690 2166 -684
rect 2160 -696 2166 -690
rect 2160 -702 2166 -696
rect 2160 -708 2166 -702
rect 2160 -714 2166 -708
rect 2160 -720 2166 -714
rect 2160 -726 2166 -720
rect 2160 -732 2166 -726
rect 2160 -738 2166 -732
rect 2160 -744 2166 -738
rect 2160 -750 2166 -744
rect 2160 -756 2166 -750
rect 2160 -762 2166 -756
rect 2160 -768 2166 -762
rect 2160 -774 2166 -768
rect 2160 -780 2166 -774
rect 2160 -786 2166 -780
rect 2160 -792 2166 -786
rect 2160 -798 2166 -792
rect 2160 -804 2166 -798
rect 2160 -810 2166 -804
rect 2160 -816 2166 -810
rect 2160 -822 2166 -816
rect 2160 -828 2166 -822
rect 2160 -834 2166 -828
rect 2160 -840 2166 -834
rect 2160 -846 2166 -840
rect 2160 -852 2166 -846
rect 2160 -858 2166 -852
rect 2160 -864 2166 -858
rect 2160 -870 2166 -864
rect 2160 -876 2166 -870
rect 2160 -882 2166 -876
rect 2160 -888 2166 -882
rect 2160 -894 2166 -888
rect 2160 -900 2166 -894
rect 2160 -906 2166 -900
rect 2160 -912 2166 -906
rect 2160 -918 2166 -912
rect 2160 -924 2166 -918
rect 2160 -930 2166 -924
rect 2160 -936 2166 -930
rect 2160 -942 2166 -936
rect 2160 -948 2166 -942
rect 2160 -954 2166 -948
rect 2160 -960 2166 -954
rect 2160 -966 2166 -960
rect 2160 -972 2166 -966
rect 2160 -978 2166 -972
rect 2160 -984 2166 -978
rect 2160 -990 2166 -984
rect 2160 -996 2166 -990
rect 2160 -1002 2166 -996
rect 2160 -1008 2166 -1002
rect 2160 -1014 2166 -1008
rect 2160 -1020 2166 -1014
rect 2160 -1026 2166 -1020
rect 2160 -1032 2166 -1026
rect 2160 -1038 2166 -1032
rect 2160 -1044 2166 -1038
rect 2160 -1050 2166 -1044
rect 2160 -1056 2166 -1050
rect 2160 -1062 2166 -1056
rect 2160 -1068 2166 -1062
rect 2160 -1074 2166 -1068
rect 2160 -1080 2166 -1074
rect 2160 -1086 2166 -1080
rect 2160 -1092 2166 -1086
rect 2160 -1098 2166 -1092
rect 2160 -1104 2166 -1098
rect 2160 -1110 2166 -1104
rect 2160 -1116 2166 -1110
rect 2160 -1122 2166 -1116
rect 2160 -1128 2166 -1122
rect 2160 -1134 2166 -1128
rect 2160 -1140 2166 -1134
rect 2160 -1146 2166 -1140
rect 2160 -1152 2166 -1146
rect 2160 -1158 2166 -1152
rect 2160 -1164 2166 -1158
rect 2160 -1170 2166 -1164
rect 2160 -1176 2166 -1170
rect 2160 -1182 2166 -1176
rect 2160 -1188 2166 -1182
rect 2160 -1194 2166 -1188
rect 2160 -1200 2166 -1194
rect 2160 -1206 2166 -1200
rect 2160 -1212 2166 -1206
rect 2160 -1218 2166 -1212
rect 2160 -1224 2166 -1218
rect 2160 -1230 2166 -1224
rect 2160 -1236 2166 -1230
rect 2160 -1242 2166 -1236
rect 2160 -1248 2166 -1242
rect 2160 -1254 2166 -1248
rect 2160 -1260 2166 -1254
rect 2160 -1266 2166 -1260
rect 2160 -1272 2166 -1266
rect 2160 -1278 2166 -1272
rect 2160 -1284 2166 -1278
rect 2160 -1290 2166 -1284
rect 2160 -1296 2166 -1290
rect 2160 -1302 2166 -1296
rect 2160 -1308 2166 -1302
rect 2160 -1314 2166 -1308
rect 2160 -1320 2166 -1314
rect 2160 -1326 2166 -1320
rect 2160 -1332 2166 -1326
rect 2160 -1338 2166 -1332
rect 2160 -1590 2166 -1584
rect 2160 -1596 2166 -1590
rect 2160 -1602 2166 -1596
rect 2160 -1608 2166 -1602
rect 2160 -1614 2166 -1608
rect 2160 -1620 2166 -1614
rect 2160 -1626 2166 -1620
rect 2160 -1632 2166 -1626
rect 2160 -1638 2166 -1632
rect 2160 -1644 2166 -1638
rect 2160 -1650 2166 -1644
rect 2160 -1656 2166 -1650
rect 2160 -1662 2166 -1656
rect 2160 -1668 2166 -1662
rect 2160 -1674 2166 -1668
rect 2160 -1680 2166 -1674
rect 2160 -1686 2166 -1680
rect 2160 -1692 2166 -1686
rect 2160 -1698 2166 -1692
rect 2160 -1704 2166 -1698
rect 2160 -1710 2166 -1704
rect 2160 -1716 2166 -1710
rect 2160 -1722 2166 -1716
rect 2160 -1728 2166 -1722
rect 2160 -1734 2166 -1728
rect 2160 -1740 2166 -1734
rect 2160 -1746 2166 -1740
rect 2160 -1752 2166 -1746
rect 2160 -1758 2166 -1752
rect 2160 -1764 2166 -1758
rect 2160 -1770 2166 -1764
rect 2160 -1776 2166 -1770
rect 2160 -1782 2166 -1776
rect 2160 -1788 2166 -1782
rect 2160 -1794 2166 -1788
rect 2160 -1800 2166 -1794
rect 2160 -1806 2166 -1800
rect 2160 -1812 2166 -1806
rect 2160 -1818 2166 -1812
rect 2160 -1824 2166 -1818
rect 2160 -1830 2166 -1824
rect 2160 -1836 2166 -1830
rect 2160 -1842 2166 -1836
rect 2160 -1848 2166 -1842
rect 2160 -1854 2166 -1848
rect 2160 -1860 2166 -1854
rect 2160 -1866 2166 -1860
rect 2160 -1872 2166 -1866
rect 2160 -1878 2166 -1872
rect 2160 -1884 2166 -1878
rect 2160 -1890 2166 -1884
rect 2160 -1896 2166 -1890
rect 2160 -1902 2166 -1896
rect 2160 -1908 2166 -1902
rect 2160 -1914 2166 -1908
rect 2160 -1920 2166 -1914
rect 2160 -1926 2166 -1920
rect 2160 -1932 2166 -1926
rect 2160 -1938 2166 -1932
rect 2160 -1944 2166 -1938
rect 2160 -1950 2166 -1944
rect 2160 -1956 2166 -1950
rect 2160 -1962 2166 -1956
rect 2160 -1968 2166 -1962
rect 2160 -1974 2166 -1968
rect 2160 -1980 2166 -1974
rect 2160 -1986 2166 -1980
rect 2160 -1992 2166 -1986
rect 2160 -1998 2166 -1992
rect 2160 -2004 2166 -1998
rect 2160 -2010 2166 -2004
rect 2160 -2016 2166 -2010
rect 2160 -2022 2166 -2016
rect 2160 -2028 2166 -2022
rect 2160 -2034 2166 -2028
rect 2160 -2040 2166 -2034
rect 2160 -2046 2166 -2040
rect 2160 -2052 2166 -2046
rect 2160 -2058 2166 -2052
rect 2160 -2064 2166 -2058
rect 2160 -2070 2166 -2064
rect 2160 -2076 2166 -2070
rect 2160 -2082 2166 -2076
rect 2160 -2088 2166 -2082
rect 2160 -2094 2166 -2088
rect 2160 -2100 2166 -2094
rect 2160 -2106 2166 -2100
rect 2160 -2112 2166 -2106
rect 2160 -2118 2166 -2112
rect 2160 -2124 2166 -2118
rect 2160 -2130 2166 -2124
rect 2160 -2136 2166 -2130
rect 2160 -2142 2166 -2136
rect 2160 -2148 2166 -2142
rect 2160 -2154 2166 -2148
rect 2160 -2160 2166 -2154
rect 2160 -2166 2166 -2160
rect 2160 -2172 2166 -2166
rect 2160 -2178 2166 -2172
rect 2160 -2184 2166 -2178
rect 2160 -2190 2166 -2184
rect 2160 -2196 2166 -2190
rect 2160 -2202 2166 -2196
rect 2160 -2208 2166 -2202
rect 2160 -2214 2166 -2208
rect 2160 -2220 2166 -2214
rect 2160 -2226 2166 -2220
rect 2160 -2232 2166 -2226
rect 2160 -2238 2166 -2232
rect 2160 -2244 2166 -2238
rect 2160 -2250 2166 -2244
rect 2160 -2256 2166 -2250
rect 2160 -2262 2166 -2256
rect 2160 -2268 2166 -2262
rect 2160 -2274 2166 -2268
rect 2160 -2280 2166 -2274
rect 2160 -2286 2166 -2280
rect 2160 -2292 2166 -2286
rect 2160 -2298 2166 -2292
rect 2160 -2304 2166 -2298
rect 2160 -2310 2166 -2304
rect 2160 -2316 2166 -2310
rect 2160 -2322 2166 -2316
rect 2160 -2328 2166 -2322
rect 2160 -2334 2166 -2328
rect 2160 -2340 2166 -2334
rect 2160 -2346 2166 -2340
rect 2160 -2352 2166 -2346
rect 2160 -2358 2166 -2352
rect 2160 -2364 2166 -2358
rect 2160 -2370 2166 -2364
rect 2160 -2376 2166 -2370
rect 2160 -2382 2166 -2376
rect 2160 -2388 2166 -2382
rect 2160 -2394 2166 -2388
rect 2160 -2550 2166 -2544
rect 2160 -2556 2166 -2550
rect 2160 -2562 2166 -2556
rect 2160 -2568 2166 -2562
rect 2160 -2574 2166 -2568
rect 2160 -2580 2166 -2574
rect 2160 -2586 2166 -2580
rect 2160 -2592 2166 -2586
rect 2160 -2598 2166 -2592
rect 2160 -2604 2166 -2598
rect 2160 -2610 2166 -2604
rect 2160 -2616 2166 -2610
rect 2160 -2622 2166 -2616
rect 2160 -2628 2166 -2622
rect 2160 -2634 2166 -2628
rect 2160 -2640 2166 -2634
rect 2160 -2646 2166 -2640
rect 2160 -2652 2166 -2646
rect 2160 -2658 2166 -2652
rect 2160 -2664 2166 -2658
rect 2160 -2670 2166 -2664
rect 2160 -2676 2166 -2670
rect 2160 -2682 2166 -2676
rect 2160 -2688 2166 -2682
rect 2160 -2694 2166 -2688
rect 2160 -2700 2166 -2694
rect 2160 -2706 2166 -2700
rect 2160 -2712 2166 -2706
rect 2160 -2718 2166 -2712
rect 2160 -2724 2166 -2718
rect 2160 -2730 2166 -2724
rect 2160 -2736 2166 -2730
rect 2160 -2742 2166 -2736
rect 2160 -2748 2166 -2742
rect 2160 -2754 2166 -2748
rect 2160 -2760 2166 -2754
rect 2160 -2766 2166 -2760
rect 2160 -2772 2166 -2766
rect 2160 -2778 2166 -2772
rect 2160 -2784 2166 -2778
rect 2160 -2790 2166 -2784
rect 2160 -2796 2166 -2790
rect 2160 -2802 2166 -2796
rect 2160 -2808 2166 -2802
rect 2160 -2814 2166 -2808
rect 2160 -2820 2166 -2814
rect 2160 -2826 2166 -2820
rect 2160 -2832 2166 -2826
rect 2160 -2838 2166 -2832
rect 2160 -2844 2166 -2838
rect 2160 -2850 2166 -2844
rect 2160 -2856 2166 -2850
rect 2160 -2862 2166 -2856
rect 2160 -2868 2166 -2862
rect 2160 -2874 2166 -2868
rect 2160 -2880 2166 -2874
rect 2160 -2886 2166 -2880
rect 2160 -2892 2166 -2886
rect 2160 -2898 2166 -2892
rect 2160 -2904 2166 -2898
rect 2160 -2910 2166 -2904
rect 2160 -2916 2166 -2910
rect 2160 -2922 2166 -2916
rect 2160 -2928 2166 -2922
rect 2160 -2934 2166 -2928
rect 2160 -2940 2166 -2934
rect 2160 -2946 2166 -2940
rect 2160 -2952 2166 -2946
rect 2160 -2958 2166 -2952
rect 2160 -2964 2166 -2958
rect 2160 -2970 2166 -2964
rect 2160 -2976 2166 -2970
rect 2160 -2982 2166 -2976
rect 2160 -2988 2166 -2982
rect 2160 -2994 2166 -2988
rect 2160 -3000 2166 -2994
rect 2160 -3006 2166 -3000
rect 2160 -3012 2166 -3006
rect 2160 -3018 2166 -3012
rect 2160 -3024 2166 -3018
rect 2160 -3030 2166 -3024
rect 2166 -240 2172 -234
rect 2166 -246 2172 -240
rect 2166 -252 2172 -246
rect 2166 -258 2172 -252
rect 2166 -264 2172 -258
rect 2166 -270 2172 -264
rect 2166 -276 2172 -270
rect 2166 -282 2172 -276
rect 2166 -288 2172 -282
rect 2166 -294 2172 -288
rect 2166 -300 2172 -294
rect 2166 -306 2172 -300
rect 2166 -312 2172 -306
rect 2166 -318 2172 -312
rect 2166 -324 2172 -318
rect 2166 -330 2172 -324
rect 2166 -336 2172 -330
rect 2166 -342 2172 -336
rect 2166 -348 2172 -342
rect 2166 -354 2172 -348
rect 2166 -360 2172 -354
rect 2166 -366 2172 -360
rect 2166 -372 2172 -366
rect 2166 -378 2172 -372
rect 2166 -384 2172 -378
rect 2166 -390 2172 -384
rect 2166 -396 2172 -390
rect 2166 -402 2172 -396
rect 2166 -408 2172 -402
rect 2166 -414 2172 -408
rect 2166 -420 2172 -414
rect 2166 -426 2172 -420
rect 2166 -432 2172 -426
rect 2166 -438 2172 -432
rect 2166 -444 2172 -438
rect 2166 -450 2172 -444
rect 2166 -456 2172 -450
rect 2166 -462 2172 -456
rect 2166 -468 2172 -462
rect 2166 -474 2172 -468
rect 2166 -480 2172 -474
rect 2166 -486 2172 -480
rect 2166 -492 2172 -486
rect 2166 -498 2172 -492
rect 2166 -504 2172 -498
rect 2166 -510 2172 -504
rect 2166 -516 2172 -510
rect 2166 -522 2172 -516
rect 2166 -528 2172 -522
rect 2166 -534 2172 -528
rect 2166 -540 2172 -534
rect 2166 -546 2172 -540
rect 2166 -552 2172 -546
rect 2166 -558 2172 -552
rect 2166 -564 2172 -558
rect 2166 -570 2172 -564
rect 2166 -576 2172 -570
rect 2166 -582 2172 -576
rect 2166 -588 2172 -582
rect 2166 -594 2172 -588
rect 2166 -600 2172 -594
rect 2166 -606 2172 -600
rect 2166 -612 2172 -606
rect 2166 -618 2172 -612
rect 2166 -624 2172 -618
rect 2166 -630 2172 -624
rect 2166 -636 2172 -630
rect 2166 -642 2172 -636
rect 2166 -648 2172 -642
rect 2166 -654 2172 -648
rect 2166 -660 2172 -654
rect 2166 -666 2172 -660
rect 2166 -672 2172 -666
rect 2166 -678 2172 -672
rect 2166 -684 2172 -678
rect 2166 -690 2172 -684
rect 2166 -696 2172 -690
rect 2166 -702 2172 -696
rect 2166 -708 2172 -702
rect 2166 -714 2172 -708
rect 2166 -720 2172 -714
rect 2166 -726 2172 -720
rect 2166 -732 2172 -726
rect 2166 -738 2172 -732
rect 2166 -744 2172 -738
rect 2166 -750 2172 -744
rect 2166 -756 2172 -750
rect 2166 -762 2172 -756
rect 2166 -768 2172 -762
rect 2166 -774 2172 -768
rect 2166 -780 2172 -774
rect 2166 -786 2172 -780
rect 2166 -792 2172 -786
rect 2166 -798 2172 -792
rect 2166 -804 2172 -798
rect 2166 -810 2172 -804
rect 2166 -816 2172 -810
rect 2166 -822 2172 -816
rect 2166 -828 2172 -822
rect 2166 -834 2172 -828
rect 2166 -840 2172 -834
rect 2166 -846 2172 -840
rect 2166 -852 2172 -846
rect 2166 -858 2172 -852
rect 2166 -864 2172 -858
rect 2166 -870 2172 -864
rect 2166 -876 2172 -870
rect 2166 -882 2172 -876
rect 2166 -888 2172 -882
rect 2166 -894 2172 -888
rect 2166 -900 2172 -894
rect 2166 -906 2172 -900
rect 2166 -912 2172 -906
rect 2166 -918 2172 -912
rect 2166 -924 2172 -918
rect 2166 -930 2172 -924
rect 2166 -936 2172 -930
rect 2166 -942 2172 -936
rect 2166 -948 2172 -942
rect 2166 -954 2172 -948
rect 2166 -960 2172 -954
rect 2166 -966 2172 -960
rect 2166 -972 2172 -966
rect 2166 -978 2172 -972
rect 2166 -984 2172 -978
rect 2166 -990 2172 -984
rect 2166 -996 2172 -990
rect 2166 -1002 2172 -996
rect 2166 -1008 2172 -1002
rect 2166 -1014 2172 -1008
rect 2166 -1020 2172 -1014
rect 2166 -1026 2172 -1020
rect 2166 -1032 2172 -1026
rect 2166 -1038 2172 -1032
rect 2166 -1044 2172 -1038
rect 2166 -1050 2172 -1044
rect 2166 -1056 2172 -1050
rect 2166 -1062 2172 -1056
rect 2166 -1068 2172 -1062
rect 2166 -1074 2172 -1068
rect 2166 -1080 2172 -1074
rect 2166 -1086 2172 -1080
rect 2166 -1092 2172 -1086
rect 2166 -1098 2172 -1092
rect 2166 -1104 2172 -1098
rect 2166 -1110 2172 -1104
rect 2166 -1116 2172 -1110
rect 2166 -1122 2172 -1116
rect 2166 -1128 2172 -1122
rect 2166 -1134 2172 -1128
rect 2166 -1140 2172 -1134
rect 2166 -1146 2172 -1140
rect 2166 -1152 2172 -1146
rect 2166 -1158 2172 -1152
rect 2166 -1164 2172 -1158
rect 2166 -1170 2172 -1164
rect 2166 -1176 2172 -1170
rect 2166 -1182 2172 -1176
rect 2166 -1188 2172 -1182
rect 2166 -1194 2172 -1188
rect 2166 -1200 2172 -1194
rect 2166 -1206 2172 -1200
rect 2166 -1212 2172 -1206
rect 2166 -1218 2172 -1212
rect 2166 -1224 2172 -1218
rect 2166 -1230 2172 -1224
rect 2166 -1236 2172 -1230
rect 2166 -1242 2172 -1236
rect 2166 -1248 2172 -1242
rect 2166 -1254 2172 -1248
rect 2166 -1260 2172 -1254
rect 2166 -1266 2172 -1260
rect 2166 -1272 2172 -1266
rect 2166 -1278 2172 -1272
rect 2166 -1284 2172 -1278
rect 2166 -1290 2172 -1284
rect 2166 -1296 2172 -1290
rect 2166 -1302 2172 -1296
rect 2166 -1308 2172 -1302
rect 2166 -1314 2172 -1308
rect 2166 -1320 2172 -1314
rect 2166 -1326 2172 -1320
rect 2166 -1584 2172 -1578
rect 2166 -1590 2172 -1584
rect 2166 -1596 2172 -1590
rect 2166 -1602 2172 -1596
rect 2166 -1608 2172 -1602
rect 2166 -1614 2172 -1608
rect 2166 -1620 2172 -1614
rect 2166 -1626 2172 -1620
rect 2166 -1632 2172 -1626
rect 2166 -1638 2172 -1632
rect 2166 -1644 2172 -1638
rect 2166 -1650 2172 -1644
rect 2166 -1656 2172 -1650
rect 2166 -1662 2172 -1656
rect 2166 -1668 2172 -1662
rect 2166 -1674 2172 -1668
rect 2166 -1680 2172 -1674
rect 2166 -1686 2172 -1680
rect 2166 -1692 2172 -1686
rect 2166 -1698 2172 -1692
rect 2166 -1704 2172 -1698
rect 2166 -1710 2172 -1704
rect 2166 -1716 2172 -1710
rect 2166 -1722 2172 -1716
rect 2166 -1728 2172 -1722
rect 2166 -1734 2172 -1728
rect 2166 -1740 2172 -1734
rect 2166 -1746 2172 -1740
rect 2166 -1752 2172 -1746
rect 2166 -1758 2172 -1752
rect 2166 -1764 2172 -1758
rect 2166 -1770 2172 -1764
rect 2166 -1776 2172 -1770
rect 2166 -1782 2172 -1776
rect 2166 -1788 2172 -1782
rect 2166 -1794 2172 -1788
rect 2166 -1800 2172 -1794
rect 2166 -1806 2172 -1800
rect 2166 -1812 2172 -1806
rect 2166 -1818 2172 -1812
rect 2166 -1824 2172 -1818
rect 2166 -1830 2172 -1824
rect 2166 -1836 2172 -1830
rect 2166 -1842 2172 -1836
rect 2166 -1848 2172 -1842
rect 2166 -1854 2172 -1848
rect 2166 -1860 2172 -1854
rect 2166 -1866 2172 -1860
rect 2166 -1872 2172 -1866
rect 2166 -1878 2172 -1872
rect 2166 -1884 2172 -1878
rect 2166 -1890 2172 -1884
rect 2166 -1896 2172 -1890
rect 2166 -1902 2172 -1896
rect 2166 -1908 2172 -1902
rect 2166 -1914 2172 -1908
rect 2166 -1920 2172 -1914
rect 2166 -1926 2172 -1920
rect 2166 -1932 2172 -1926
rect 2166 -1938 2172 -1932
rect 2166 -1944 2172 -1938
rect 2166 -1950 2172 -1944
rect 2166 -1956 2172 -1950
rect 2166 -1962 2172 -1956
rect 2166 -1968 2172 -1962
rect 2166 -1974 2172 -1968
rect 2166 -1980 2172 -1974
rect 2166 -1986 2172 -1980
rect 2166 -1992 2172 -1986
rect 2166 -1998 2172 -1992
rect 2166 -2004 2172 -1998
rect 2166 -2010 2172 -2004
rect 2166 -2016 2172 -2010
rect 2166 -2022 2172 -2016
rect 2166 -2028 2172 -2022
rect 2166 -2034 2172 -2028
rect 2166 -2040 2172 -2034
rect 2166 -2046 2172 -2040
rect 2166 -2052 2172 -2046
rect 2166 -2058 2172 -2052
rect 2166 -2064 2172 -2058
rect 2166 -2070 2172 -2064
rect 2166 -2076 2172 -2070
rect 2166 -2082 2172 -2076
rect 2166 -2088 2172 -2082
rect 2166 -2094 2172 -2088
rect 2166 -2100 2172 -2094
rect 2166 -2106 2172 -2100
rect 2166 -2112 2172 -2106
rect 2166 -2118 2172 -2112
rect 2166 -2124 2172 -2118
rect 2166 -2130 2172 -2124
rect 2166 -2136 2172 -2130
rect 2166 -2142 2172 -2136
rect 2166 -2148 2172 -2142
rect 2166 -2154 2172 -2148
rect 2166 -2160 2172 -2154
rect 2166 -2166 2172 -2160
rect 2166 -2172 2172 -2166
rect 2166 -2178 2172 -2172
rect 2166 -2184 2172 -2178
rect 2166 -2190 2172 -2184
rect 2166 -2196 2172 -2190
rect 2166 -2202 2172 -2196
rect 2166 -2208 2172 -2202
rect 2166 -2214 2172 -2208
rect 2166 -2220 2172 -2214
rect 2166 -2226 2172 -2220
rect 2166 -2232 2172 -2226
rect 2166 -2238 2172 -2232
rect 2166 -2244 2172 -2238
rect 2166 -2250 2172 -2244
rect 2166 -2256 2172 -2250
rect 2166 -2262 2172 -2256
rect 2166 -2268 2172 -2262
rect 2166 -2274 2172 -2268
rect 2166 -2280 2172 -2274
rect 2166 -2286 2172 -2280
rect 2166 -2292 2172 -2286
rect 2166 -2298 2172 -2292
rect 2166 -2304 2172 -2298
rect 2166 -2310 2172 -2304
rect 2166 -2316 2172 -2310
rect 2166 -2322 2172 -2316
rect 2166 -2328 2172 -2322
rect 2166 -2334 2172 -2328
rect 2166 -2340 2172 -2334
rect 2166 -2346 2172 -2340
rect 2166 -2352 2172 -2346
rect 2166 -2358 2172 -2352
rect 2166 -2364 2172 -2358
rect 2166 -2370 2172 -2364
rect 2166 -2376 2172 -2370
rect 2166 -2382 2172 -2376
rect 2166 -2550 2172 -2544
rect 2166 -2556 2172 -2550
rect 2166 -2562 2172 -2556
rect 2166 -2568 2172 -2562
rect 2166 -2574 2172 -2568
rect 2166 -2580 2172 -2574
rect 2166 -2586 2172 -2580
rect 2166 -2592 2172 -2586
rect 2166 -2598 2172 -2592
rect 2166 -2604 2172 -2598
rect 2166 -2610 2172 -2604
rect 2166 -2616 2172 -2610
rect 2166 -2622 2172 -2616
rect 2166 -2628 2172 -2622
rect 2166 -2634 2172 -2628
rect 2166 -2640 2172 -2634
rect 2166 -2646 2172 -2640
rect 2166 -2652 2172 -2646
rect 2166 -2658 2172 -2652
rect 2166 -2664 2172 -2658
rect 2166 -2670 2172 -2664
rect 2166 -2676 2172 -2670
rect 2166 -2682 2172 -2676
rect 2166 -2688 2172 -2682
rect 2166 -2694 2172 -2688
rect 2166 -2700 2172 -2694
rect 2166 -2706 2172 -2700
rect 2166 -2712 2172 -2706
rect 2166 -2718 2172 -2712
rect 2166 -2724 2172 -2718
rect 2166 -2730 2172 -2724
rect 2166 -2736 2172 -2730
rect 2166 -2742 2172 -2736
rect 2166 -2748 2172 -2742
rect 2166 -2754 2172 -2748
rect 2166 -2760 2172 -2754
rect 2166 -2766 2172 -2760
rect 2166 -2772 2172 -2766
rect 2166 -2778 2172 -2772
rect 2166 -2784 2172 -2778
rect 2166 -2790 2172 -2784
rect 2166 -2796 2172 -2790
rect 2166 -2802 2172 -2796
rect 2166 -2808 2172 -2802
rect 2166 -2814 2172 -2808
rect 2166 -2820 2172 -2814
rect 2166 -2826 2172 -2820
rect 2166 -2832 2172 -2826
rect 2166 -2838 2172 -2832
rect 2166 -2844 2172 -2838
rect 2166 -2850 2172 -2844
rect 2166 -2856 2172 -2850
rect 2166 -2862 2172 -2856
rect 2166 -2868 2172 -2862
rect 2166 -2874 2172 -2868
rect 2166 -2880 2172 -2874
rect 2166 -2886 2172 -2880
rect 2166 -2892 2172 -2886
rect 2166 -2898 2172 -2892
rect 2166 -2904 2172 -2898
rect 2166 -2910 2172 -2904
rect 2166 -2916 2172 -2910
rect 2166 -2922 2172 -2916
rect 2166 -2928 2172 -2922
rect 2166 -2934 2172 -2928
rect 2166 -2940 2172 -2934
rect 2166 -2946 2172 -2940
rect 2166 -2952 2172 -2946
rect 2166 -2958 2172 -2952
rect 2166 -2964 2172 -2958
rect 2166 -2970 2172 -2964
rect 2166 -2976 2172 -2970
rect 2166 -2982 2172 -2976
rect 2166 -2988 2172 -2982
rect 2166 -2994 2172 -2988
rect 2166 -3000 2172 -2994
rect 2166 -3006 2172 -3000
rect 2166 -3012 2172 -3006
rect 2166 -3018 2172 -3012
rect 2166 -3024 2172 -3018
rect 2172 -234 2178 -228
rect 2172 -240 2178 -234
rect 2172 -246 2178 -240
rect 2172 -252 2178 -246
rect 2172 -258 2178 -252
rect 2172 -264 2178 -258
rect 2172 -270 2178 -264
rect 2172 -276 2178 -270
rect 2172 -282 2178 -276
rect 2172 -288 2178 -282
rect 2172 -294 2178 -288
rect 2172 -300 2178 -294
rect 2172 -306 2178 -300
rect 2172 -312 2178 -306
rect 2172 -318 2178 -312
rect 2172 -324 2178 -318
rect 2172 -330 2178 -324
rect 2172 -336 2178 -330
rect 2172 -342 2178 -336
rect 2172 -348 2178 -342
rect 2172 -354 2178 -348
rect 2172 -360 2178 -354
rect 2172 -366 2178 -360
rect 2172 -372 2178 -366
rect 2172 -378 2178 -372
rect 2172 -384 2178 -378
rect 2172 -390 2178 -384
rect 2172 -396 2178 -390
rect 2172 -402 2178 -396
rect 2172 -408 2178 -402
rect 2172 -414 2178 -408
rect 2172 -420 2178 -414
rect 2172 -426 2178 -420
rect 2172 -432 2178 -426
rect 2172 -438 2178 -432
rect 2172 -444 2178 -438
rect 2172 -450 2178 -444
rect 2172 -456 2178 -450
rect 2172 -462 2178 -456
rect 2172 -468 2178 -462
rect 2172 -474 2178 -468
rect 2172 -480 2178 -474
rect 2172 -486 2178 -480
rect 2172 -492 2178 -486
rect 2172 -498 2178 -492
rect 2172 -504 2178 -498
rect 2172 -510 2178 -504
rect 2172 -516 2178 -510
rect 2172 -522 2178 -516
rect 2172 -528 2178 -522
rect 2172 -534 2178 -528
rect 2172 -540 2178 -534
rect 2172 -546 2178 -540
rect 2172 -552 2178 -546
rect 2172 -558 2178 -552
rect 2172 -564 2178 -558
rect 2172 -570 2178 -564
rect 2172 -576 2178 -570
rect 2172 -582 2178 -576
rect 2172 -588 2178 -582
rect 2172 -594 2178 -588
rect 2172 -600 2178 -594
rect 2172 -606 2178 -600
rect 2172 -612 2178 -606
rect 2172 -618 2178 -612
rect 2172 -624 2178 -618
rect 2172 -630 2178 -624
rect 2172 -636 2178 -630
rect 2172 -642 2178 -636
rect 2172 -648 2178 -642
rect 2172 -654 2178 -648
rect 2172 -660 2178 -654
rect 2172 -666 2178 -660
rect 2172 -672 2178 -666
rect 2172 -678 2178 -672
rect 2172 -684 2178 -678
rect 2172 -690 2178 -684
rect 2172 -696 2178 -690
rect 2172 -702 2178 -696
rect 2172 -708 2178 -702
rect 2172 -714 2178 -708
rect 2172 -720 2178 -714
rect 2172 -726 2178 -720
rect 2172 -732 2178 -726
rect 2172 -738 2178 -732
rect 2172 -744 2178 -738
rect 2172 -750 2178 -744
rect 2172 -756 2178 -750
rect 2172 -762 2178 -756
rect 2172 -768 2178 -762
rect 2172 -774 2178 -768
rect 2172 -780 2178 -774
rect 2172 -786 2178 -780
rect 2172 -792 2178 -786
rect 2172 -798 2178 -792
rect 2172 -804 2178 -798
rect 2172 -810 2178 -804
rect 2172 -816 2178 -810
rect 2172 -822 2178 -816
rect 2172 -828 2178 -822
rect 2172 -834 2178 -828
rect 2172 -840 2178 -834
rect 2172 -846 2178 -840
rect 2172 -852 2178 -846
rect 2172 -858 2178 -852
rect 2172 -864 2178 -858
rect 2172 -870 2178 -864
rect 2172 -876 2178 -870
rect 2172 -882 2178 -876
rect 2172 -888 2178 -882
rect 2172 -894 2178 -888
rect 2172 -900 2178 -894
rect 2172 -906 2178 -900
rect 2172 -912 2178 -906
rect 2172 -918 2178 -912
rect 2172 -924 2178 -918
rect 2172 -930 2178 -924
rect 2172 -936 2178 -930
rect 2172 -942 2178 -936
rect 2172 -948 2178 -942
rect 2172 -954 2178 -948
rect 2172 -960 2178 -954
rect 2172 -966 2178 -960
rect 2172 -972 2178 -966
rect 2172 -978 2178 -972
rect 2172 -984 2178 -978
rect 2172 -990 2178 -984
rect 2172 -996 2178 -990
rect 2172 -1002 2178 -996
rect 2172 -1008 2178 -1002
rect 2172 -1014 2178 -1008
rect 2172 -1020 2178 -1014
rect 2172 -1026 2178 -1020
rect 2172 -1032 2178 -1026
rect 2172 -1038 2178 -1032
rect 2172 -1044 2178 -1038
rect 2172 -1050 2178 -1044
rect 2172 -1056 2178 -1050
rect 2172 -1062 2178 -1056
rect 2172 -1068 2178 -1062
rect 2172 -1074 2178 -1068
rect 2172 -1080 2178 -1074
rect 2172 -1086 2178 -1080
rect 2172 -1092 2178 -1086
rect 2172 -1098 2178 -1092
rect 2172 -1104 2178 -1098
rect 2172 -1110 2178 -1104
rect 2172 -1116 2178 -1110
rect 2172 -1122 2178 -1116
rect 2172 -1128 2178 -1122
rect 2172 -1134 2178 -1128
rect 2172 -1140 2178 -1134
rect 2172 -1146 2178 -1140
rect 2172 -1152 2178 -1146
rect 2172 -1158 2178 -1152
rect 2172 -1164 2178 -1158
rect 2172 -1170 2178 -1164
rect 2172 -1176 2178 -1170
rect 2172 -1182 2178 -1176
rect 2172 -1188 2178 -1182
rect 2172 -1194 2178 -1188
rect 2172 -1200 2178 -1194
rect 2172 -1206 2178 -1200
rect 2172 -1212 2178 -1206
rect 2172 -1218 2178 -1212
rect 2172 -1224 2178 -1218
rect 2172 -1230 2178 -1224
rect 2172 -1236 2178 -1230
rect 2172 -1242 2178 -1236
rect 2172 -1248 2178 -1242
rect 2172 -1254 2178 -1248
rect 2172 -1260 2178 -1254
rect 2172 -1266 2178 -1260
rect 2172 -1272 2178 -1266
rect 2172 -1278 2178 -1272
rect 2172 -1284 2178 -1278
rect 2172 -1290 2178 -1284
rect 2172 -1296 2178 -1290
rect 2172 -1302 2178 -1296
rect 2172 -1308 2178 -1302
rect 2172 -1314 2178 -1308
rect 2172 -1578 2178 -1572
rect 2172 -1584 2178 -1578
rect 2172 -1590 2178 -1584
rect 2172 -1596 2178 -1590
rect 2172 -1602 2178 -1596
rect 2172 -1608 2178 -1602
rect 2172 -1614 2178 -1608
rect 2172 -1620 2178 -1614
rect 2172 -1626 2178 -1620
rect 2172 -1632 2178 -1626
rect 2172 -1638 2178 -1632
rect 2172 -1644 2178 -1638
rect 2172 -1650 2178 -1644
rect 2172 -1656 2178 -1650
rect 2172 -1662 2178 -1656
rect 2172 -1668 2178 -1662
rect 2172 -1674 2178 -1668
rect 2172 -1680 2178 -1674
rect 2172 -1686 2178 -1680
rect 2172 -1692 2178 -1686
rect 2172 -1698 2178 -1692
rect 2172 -1704 2178 -1698
rect 2172 -1710 2178 -1704
rect 2172 -1716 2178 -1710
rect 2172 -1722 2178 -1716
rect 2172 -1728 2178 -1722
rect 2172 -1734 2178 -1728
rect 2172 -1740 2178 -1734
rect 2172 -1746 2178 -1740
rect 2172 -1752 2178 -1746
rect 2172 -1758 2178 -1752
rect 2172 -1764 2178 -1758
rect 2172 -1770 2178 -1764
rect 2172 -1776 2178 -1770
rect 2172 -1782 2178 -1776
rect 2172 -1788 2178 -1782
rect 2172 -1794 2178 -1788
rect 2172 -1800 2178 -1794
rect 2172 -1806 2178 -1800
rect 2172 -1812 2178 -1806
rect 2172 -1818 2178 -1812
rect 2172 -1824 2178 -1818
rect 2172 -1830 2178 -1824
rect 2172 -1836 2178 -1830
rect 2172 -1842 2178 -1836
rect 2172 -1848 2178 -1842
rect 2172 -1854 2178 -1848
rect 2172 -1860 2178 -1854
rect 2172 -1866 2178 -1860
rect 2172 -1872 2178 -1866
rect 2172 -1878 2178 -1872
rect 2172 -1884 2178 -1878
rect 2172 -1890 2178 -1884
rect 2172 -1896 2178 -1890
rect 2172 -1902 2178 -1896
rect 2172 -1908 2178 -1902
rect 2172 -1914 2178 -1908
rect 2172 -1920 2178 -1914
rect 2172 -1926 2178 -1920
rect 2172 -1932 2178 -1926
rect 2172 -1938 2178 -1932
rect 2172 -1944 2178 -1938
rect 2172 -1950 2178 -1944
rect 2172 -1956 2178 -1950
rect 2172 -1962 2178 -1956
rect 2172 -1968 2178 -1962
rect 2172 -1974 2178 -1968
rect 2172 -1980 2178 -1974
rect 2172 -1986 2178 -1980
rect 2172 -1992 2178 -1986
rect 2172 -1998 2178 -1992
rect 2172 -2004 2178 -1998
rect 2172 -2010 2178 -2004
rect 2172 -2016 2178 -2010
rect 2172 -2022 2178 -2016
rect 2172 -2028 2178 -2022
rect 2172 -2034 2178 -2028
rect 2172 -2040 2178 -2034
rect 2172 -2046 2178 -2040
rect 2172 -2052 2178 -2046
rect 2172 -2058 2178 -2052
rect 2172 -2064 2178 -2058
rect 2172 -2070 2178 -2064
rect 2172 -2076 2178 -2070
rect 2172 -2082 2178 -2076
rect 2172 -2088 2178 -2082
rect 2172 -2094 2178 -2088
rect 2172 -2100 2178 -2094
rect 2172 -2106 2178 -2100
rect 2172 -2112 2178 -2106
rect 2172 -2118 2178 -2112
rect 2172 -2124 2178 -2118
rect 2172 -2130 2178 -2124
rect 2172 -2136 2178 -2130
rect 2172 -2142 2178 -2136
rect 2172 -2148 2178 -2142
rect 2172 -2154 2178 -2148
rect 2172 -2160 2178 -2154
rect 2172 -2166 2178 -2160
rect 2172 -2172 2178 -2166
rect 2172 -2178 2178 -2172
rect 2172 -2184 2178 -2178
rect 2172 -2190 2178 -2184
rect 2172 -2196 2178 -2190
rect 2172 -2202 2178 -2196
rect 2172 -2208 2178 -2202
rect 2172 -2214 2178 -2208
rect 2172 -2220 2178 -2214
rect 2172 -2226 2178 -2220
rect 2172 -2232 2178 -2226
rect 2172 -2238 2178 -2232
rect 2172 -2244 2178 -2238
rect 2172 -2250 2178 -2244
rect 2172 -2256 2178 -2250
rect 2172 -2262 2178 -2256
rect 2172 -2268 2178 -2262
rect 2172 -2274 2178 -2268
rect 2172 -2280 2178 -2274
rect 2172 -2286 2178 -2280
rect 2172 -2292 2178 -2286
rect 2172 -2298 2178 -2292
rect 2172 -2304 2178 -2298
rect 2172 -2310 2178 -2304
rect 2172 -2316 2178 -2310
rect 2172 -2322 2178 -2316
rect 2172 -2328 2178 -2322
rect 2172 -2334 2178 -2328
rect 2172 -2340 2178 -2334
rect 2172 -2346 2178 -2340
rect 2172 -2352 2178 -2346
rect 2172 -2358 2178 -2352
rect 2172 -2364 2178 -2358
rect 2172 -2370 2178 -2364
rect 2172 -2376 2178 -2370
rect 2172 -2550 2178 -2544
rect 2172 -2556 2178 -2550
rect 2172 -2562 2178 -2556
rect 2172 -2568 2178 -2562
rect 2172 -2574 2178 -2568
rect 2172 -2580 2178 -2574
rect 2172 -2586 2178 -2580
rect 2172 -2592 2178 -2586
rect 2172 -2598 2178 -2592
rect 2172 -2604 2178 -2598
rect 2172 -2610 2178 -2604
rect 2172 -2616 2178 -2610
rect 2172 -2622 2178 -2616
rect 2172 -2628 2178 -2622
rect 2172 -2634 2178 -2628
rect 2172 -2640 2178 -2634
rect 2172 -2646 2178 -2640
rect 2172 -2652 2178 -2646
rect 2172 -2658 2178 -2652
rect 2172 -2664 2178 -2658
rect 2172 -2670 2178 -2664
rect 2172 -2676 2178 -2670
rect 2172 -2682 2178 -2676
rect 2172 -2688 2178 -2682
rect 2172 -2694 2178 -2688
rect 2172 -2700 2178 -2694
rect 2172 -2706 2178 -2700
rect 2172 -2712 2178 -2706
rect 2172 -2718 2178 -2712
rect 2172 -2724 2178 -2718
rect 2172 -2730 2178 -2724
rect 2172 -2736 2178 -2730
rect 2172 -2742 2178 -2736
rect 2172 -2748 2178 -2742
rect 2172 -2754 2178 -2748
rect 2172 -2760 2178 -2754
rect 2172 -2766 2178 -2760
rect 2172 -2772 2178 -2766
rect 2172 -2778 2178 -2772
rect 2172 -2784 2178 -2778
rect 2172 -2790 2178 -2784
rect 2172 -2796 2178 -2790
rect 2172 -2802 2178 -2796
rect 2172 -2808 2178 -2802
rect 2172 -2814 2178 -2808
rect 2172 -2820 2178 -2814
rect 2172 -2826 2178 -2820
rect 2172 -2832 2178 -2826
rect 2172 -2838 2178 -2832
rect 2172 -2844 2178 -2838
rect 2172 -2850 2178 -2844
rect 2172 -2856 2178 -2850
rect 2172 -2862 2178 -2856
rect 2172 -2868 2178 -2862
rect 2172 -2874 2178 -2868
rect 2172 -2880 2178 -2874
rect 2172 -2886 2178 -2880
rect 2172 -2892 2178 -2886
rect 2172 -2898 2178 -2892
rect 2172 -2904 2178 -2898
rect 2172 -2910 2178 -2904
rect 2172 -2916 2178 -2910
rect 2172 -2922 2178 -2916
rect 2172 -2928 2178 -2922
rect 2172 -2934 2178 -2928
rect 2172 -2940 2178 -2934
rect 2172 -2946 2178 -2940
rect 2172 -2952 2178 -2946
rect 2172 -2958 2178 -2952
rect 2172 -2964 2178 -2958
rect 2172 -2970 2178 -2964
rect 2172 -2976 2178 -2970
rect 2172 -2982 2178 -2976
rect 2172 -2988 2178 -2982
rect 2172 -2994 2178 -2988
rect 2172 -3000 2178 -2994
rect 2172 -3006 2178 -3000
rect 2172 -3012 2178 -3006
rect 2172 -3018 2178 -3012
rect 2172 -3024 2178 -3018
rect 2178 -228 2184 -222
rect 2178 -234 2184 -228
rect 2178 -240 2184 -234
rect 2178 -246 2184 -240
rect 2178 -252 2184 -246
rect 2178 -258 2184 -252
rect 2178 -264 2184 -258
rect 2178 -270 2184 -264
rect 2178 -276 2184 -270
rect 2178 -282 2184 -276
rect 2178 -288 2184 -282
rect 2178 -294 2184 -288
rect 2178 -300 2184 -294
rect 2178 -306 2184 -300
rect 2178 -312 2184 -306
rect 2178 -318 2184 -312
rect 2178 -324 2184 -318
rect 2178 -330 2184 -324
rect 2178 -336 2184 -330
rect 2178 -342 2184 -336
rect 2178 -348 2184 -342
rect 2178 -354 2184 -348
rect 2178 -360 2184 -354
rect 2178 -366 2184 -360
rect 2178 -372 2184 -366
rect 2178 -378 2184 -372
rect 2178 -384 2184 -378
rect 2178 -390 2184 -384
rect 2178 -396 2184 -390
rect 2178 -402 2184 -396
rect 2178 -408 2184 -402
rect 2178 -414 2184 -408
rect 2178 -420 2184 -414
rect 2178 -426 2184 -420
rect 2178 -432 2184 -426
rect 2178 -438 2184 -432
rect 2178 -444 2184 -438
rect 2178 -450 2184 -444
rect 2178 -456 2184 -450
rect 2178 -462 2184 -456
rect 2178 -468 2184 -462
rect 2178 -474 2184 -468
rect 2178 -480 2184 -474
rect 2178 -486 2184 -480
rect 2178 -492 2184 -486
rect 2178 -498 2184 -492
rect 2178 -504 2184 -498
rect 2178 -510 2184 -504
rect 2178 -516 2184 -510
rect 2178 -522 2184 -516
rect 2178 -528 2184 -522
rect 2178 -534 2184 -528
rect 2178 -540 2184 -534
rect 2178 -546 2184 -540
rect 2178 -552 2184 -546
rect 2178 -558 2184 -552
rect 2178 -564 2184 -558
rect 2178 -570 2184 -564
rect 2178 -576 2184 -570
rect 2178 -582 2184 -576
rect 2178 -588 2184 -582
rect 2178 -594 2184 -588
rect 2178 -600 2184 -594
rect 2178 -606 2184 -600
rect 2178 -612 2184 -606
rect 2178 -618 2184 -612
rect 2178 -624 2184 -618
rect 2178 -630 2184 -624
rect 2178 -636 2184 -630
rect 2178 -642 2184 -636
rect 2178 -648 2184 -642
rect 2178 -654 2184 -648
rect 2178 -660 2184 -654
rect 2178 -666 2184 -660
rect 2178 -672 2184 -666
rect 2178 -678 2184 -672
rect 2178 -684 2184 -678
rect 2178 -690 2184 -684
rect 2178 -696 2184 -690
rect 2178 -702 2184 -696
rect 2178 -708 2184 -702
rect 2178 -714 2184 -708
rect 2178 -720 2184 -714
rect 2178 -726 2184 -720
rect 2178 -732 2184 -726
rect 2178 -738 2184 -732
rect 2178 -744 2184 -738
rect 2178 -750 2184 -744
rect 2178 -756 2184 -750
rect 2178 -762 2184 -756
rect 2178 -768 2184 -762
rect 2178 -774 2184 -768
rect 2178 -780 2184 -774
rect 2178 -786 2184 -780
rect 2178 -792 2184 -786
rect 2178 -798 2184 -792
rect 2178 -804 2184 -798
rect 2178 -810 2184 -804
rect 2178 -816 2184 -810
rect 2178 -822 2184 -816
rect 2178 -828 2184 -822
rect 2178 -834 2184 -828
rect 2178 -840 2184 -834
rect 2178 -846 2184 -840
rect 2178 -852 2184 -846
rect 2178 -858 2184 -852
rect 2178 -864 2184 -858
rect 2178 -870 2184 -864
rect 2178 -876 2184 -870
rect 2178 -882 2184 -876
rect 2178 -888 2184 -882
rect 2178 -894 2184 -888
rect 2178 -900 2184 -894
rect 2178 -906 2184 -900
rect 2178 -912 2184 -906
rect 2178 -918 2184 -912
rect 2178 -924 2184 -918
rect 2178 -930 2184 -924
rect 2178 -936 2184 -930
rect 2178 -942 2184 -936
rect 2178 -948 2184 -942
rect 2178 -954 2184 -948
rect 2178 -960 2184 -954
rect 2178 -966 2184 -960
rect 2178 -972 2184 -966
rect 2178 -978 2184 -972
rect 2178 -984 2184 -978
rect 2178 -990 2184 -984
rect 2178 -996 2184 -990
rect 2178 -1002 2184 -996
rect 2178 -1008 2184 -1002
rect 2178 -1014 2184 -1008
rect 2178 -1020 2184 -1014
rect 2178 -1026 2184 -1020
rect 2178 -1032 2184 -1026
rect 2178 -1038 2184 -1032
rect 2178 -1044 2184 -1038
rect 2178 -1050 2184 -1044
rect 2178 -1056 2184 -1050
rect 2178 -1062 2184 -1056
rect 2178 -1068 2184 -1062
rect 2178 -1074 2184 -1068
rect 2178 -1080 2184 -1074
rect 2178 -1086 2184 -1080
rect 2178 -1092 2184 -1086
rect 2178 -1098 2184 -1092
rect 2178 -1104 2184 -1098
rect 2178 -1110 2184 -1104
rect 2178 -1116 2184 -1110
rect 2178 -1122 2184 -1116
rect 2178 -1128 2184 -1122
rect 2178 -1134 2184 -1128
rect 2178 -1140 2184 -1134
rect 2178 -1146 2184 -1140
rect 2178 -1152 2184 -1146
rect 2178 -1158 2184 -1152
rect 2178 -1164 2184 -1158
rect 2178 -1170 2184 -1164
rect 2178 -1176 2184 -1170
rect 2178 -1182 2184 -1176
rect 2178 -1188 2184 -1182
rect 2178 -1194 2184 -1188
rect 2178 -1200 2184 -1194
rect 2178 -1206 2184 -1200
rect 2178 -1212 2184 -1206
rect 2178 -1218 2184 -1212
rect 2178 -1224 2184 -1218
rect 2178 -1230 2184 -1224
rect 2178 -1236 2184 -1230
rect 2178 -1242 2184 -1236
rect 2178 -1248 2184 -1242
rect 2178 -1254 2184 -1248
rect 2178 -1260 2184 -1254
rect 2178 -1266 2184 -1260
rect 2178 -1272 2184 -1266
rect 2178 -1278 2184 -1272
rect 2178 -1284 2184 -1278
rect 2178 -1290 2184 -1284
rect 2178 -1296 2184 -1290
rect 2178 -1572 2184 -1566
rect 2178 -1578 2184 -1572
rect 2178 -1584 2184 -1578
rect 2178 -1590 2184 -1584
rect 2178 -1596 2184 -1590
rect 2178 -1602 2184 -1596
rect 2178 -1608 2184 -1602
rect 2178 -1614 2184 -1608
rect 2178 -1620 2184 -1614
rect 2178 -1626 2184 -1620
rect 2178 -1632 2184 -1626
rect 2178 -1638 2184 -1632
rect 2178 -1644 2184 -1638
rect 2178 -1650 2184 -1644
rect 2178 -1656 2184 -1650
rect 2178 -1662 2184 -1656
rect 2178 -1668 2184 -1662
rect 2178 -1674 2184 -1668
rect 2178 -1680 2184 -1674
rect 2178 -1686 2184 -1680
rect 2178 -1692 2184 -1686
rect 2178 -1698 2184 -1692
rect 2178 -1704 2184 -1698
rect 2178 -1710 2184 -1704
rect 2178 -1716 2184 -1710
rect 2178 -1722 2184 -1716
rect 2178 -1728 2184 -1722
rect 2178 -1734 2184 -1728
rect 2178 -1740 2184 -1734
rect 2178 -1746 2184 -1740
rect 2178 -1752 2184 -1746
rect 2178 -1758 2184 -1752
rect 2178 -1764 2184 -1758
rect 2178 -1770 2184 -1764
rect 2178 -1776 2184 -1770
rect 2178 -1782 2184 -1776
rect 2178 -1788 2184 -1782
rect 2178 -1794 2184 -1788
rect 2178 -1800 2184 -1794
rect 2178 -1806 2184 -1800
rect 2178 -1812 2184 -1806
rect 2178 -1818 2184 -1812
rect 2178 -1824 2184 -1818
rect 2178 -1830 2184 -1824
rect 2178 -1836 2184 -1830
rect 2178 -1842 2184 -1836
rect 2178 -1848 2184 -1842
rect 2178 -1854 2184 -1848
rect 2178 -1860 2184 -1854
rect 2178 -1866 2184 -1860
rect 2178 -1872 2184 -1866
rect 2178 -1878 2184 -1872
rect 2178 -1884 2184 -1878
rect 2178 -1890 2184 -1884
rect 2178 -1896 2184 -1890
rect 2178 -1902 2184 -1896
rect 2178 -1908 2184 -1902
rect 2178 -1914 2184 -1908
rect 2178 -1920 2184 -1914
rect 2178 -1926 2184 -1920
rect 2178 -1932 2184 -1926
rect 2178 -1938 2184 -1932
rect 2178 -1944 2184 -1938
rect 2178 -1950 2184 -1944
rect 2178 -1956 2184 -1950
rect 2178 -1962 2184 -1956
rect 2178 -1968 2184 -1962
rect 2178 -1974 2184 -1968
rect 2178 -1980 2184 -1974
rect 2178 -1986 2184 -1980
rect 2178 -1992 2184 -1986
rect 2178 -1998 2184 -1992
rect 2178 -2004 2184 -1998
rect 2178 -2010 2184 -2004
rect 2178 -2016 2184 -2010
rect 2178 -2022 2184 -2016
rect 2178 -2028 2184 -2022
rect 2178 -2034 2184 -2028
rect 2178 -2040 2184 -2034
rect 2178 -2046 2184 -2040
rect 2178 -2052 2184 -2046
rect 2178 -2058 2184 -2052
rect 2178 -2064 2184 -2058
rect 2178 -2070 2184 -2064
rect 2178 -2076 2184 -2070
rect 2178 -2082 2184 -2076
rect 2178 -2088 2184 -2082
rect 2178 -2094 2184 -2088
rect 2178 -2100 2184 -2094
rect 2178 -2106 2184 -2100
rect 2178 -2112 2184 -2106
rect 2178 -2118 2184 -2112
rect 2178 -2124 2184 -2118
rect 2178 -2130 2184 -2124
rect 2178 -2136 2184 -2130
rect 2178 -2142 2184 -2136
rect 2178 -2148 2184 -2142
rect 2178 -2154 2184 -2148
rect 2178 -2160 2184 -2154
rect 2178 -2166 2184 -2160
rect 2178 -2172 2184 -2166
rect 2178 -2178 2184 -2172
rect 2178 -2184 2184 -2178
rect 2178 -2190 2184 -2184
rect 2178 -2196 2184 -2190
rect 2178 -2202 2184 -2196
rect 2178 -2208 2184 -2202
rect 2178 -2214 2184 -2208
rect 2178 -2220 2184 -2214
rect 2178 -2226 2184 -2220
rect 2178 -2232 2184 -2226
rect 2178 -2238 2184 -2232
rect 2178 -2244 2184 -2238
rect 2178 -2250 2184 -2244
rect 2178 -2256 2184 -2250
rect 2178 -2262 2184 -2256
rect 2178 -2268 2184 -2262
rect 2178 -2274 2184 -2268
rect 2178 -2280 2184 -2274
rect 2178 -2286 2184 -2280
rect 2178 -2292 2184 -2286
rect 2178 -2298 2184 -2292
rect 2178 -2304 2184 -2298
rect 2178 -2310 2184 -2304
rect 2178 -2316 2184 -2310
rect 2178 -2322 2184 -2316
rect 2178 -2328 2184 -2322
rect 2178 -2334 2184 -2328
rect 2178 -2340 2184 -2334
rect 2178 -2346 2184 -2340
rect 2178 -2352 2184 -2346
rect 2178 -2358 2184 -2352
rect 2178 -2364 2184 -2358
rect 2178 -2370 2184 -2364
rect 2178 -2544 2184 -2538
rect 2178 -2550 2184 -2544
rect 2178 -2556 2184 -2550
rect 2178 -2562 2184 -2556
rect 2178 -2568 2184 -2562
rect 2178 -2574 2184 -2568
rect 2178 -2580 2184 -2574
rect 2178 -2586 2184 -2580
rect 2178 -2592 2184 -2586
rect 2178 -2598 2184 -2592
rect 2178 -2604 2184 -2598
rect 2178 -2610 2184 -2604
rect 2178 -2616 2184 -2610
rect 2178 -2622 2184 -2616
rect 2178 -2628 2184 -2622
rect 2178 -2634 2184 -2628
rect 2178 -2640 2184 -2634
rect 2178 -2646 2184 -2640
rect 2178 -2652 2184 -2646
rect 2178 -2658 2184 -2652
rect 2178 -2664 2184 -2658
rect 2178 -2670 2184 -2664
rect 2178 -2676 2184 -2670
rect 2178 -2682 2184 -2676
rect 2178 -2688 2184 -2682
rect 2178 -2694 2184 -2688
rect 2178 -2700 2184 -2694
rect 2178 -2706 2184 -2700
rect 2178 -2712 2184 -2706
rect 2178 -2718 2184 -2712
rect 2178 -2724 2184 -2718
rect 2178 -2730 2184 -2724
rect 2178 -2736 2184 -2730
rect 2178 -2742 2184 -2736
rect 2178 -2748 2184 -2742
rect 2178 -2754 2184 -2748
rect 2178 -2760 2184 -2754
rect 2178 -2766 2184 -2760
rect 2178 -2772 2184 -2766
rect 2178 -2778 2184 -2772
rect 2178 -2784 2184 -2778
rect 2178 -2790 2184 -2784
rect 2178 -2796 2184 -2790
rect 2178 -2802 2184 -2796
rect 2178 -2808 2184 -2802
rect 2178 -2814 2184 -2808
rect 2178 -2820 2184 -2814
rect 2178 -2826 2184 -2820
rect 2178 -2832 2184 -2826
rect 2178 -2838 2184 -2832
rect 2178 -2844 2184 -2838
rect 2178 -2850 2184 -2844
rect 2178 -2856 2184 -2850
rect 2178 -2862 2184 -2856
rect 2178 -2868 2184 -2862
rect 2178 -2874 2184 -2868
rect 2178 -2880 2184 -2874
rect 2178 -2886 2184 -2880
rect 2178 -2892 2184 -2886
rect 2178 -2898 2184 -2892
rect 2178 -2904 2184 -2898
rect 2178 -2910 2184 -2904
rect 2178 -2916 2184 -2910
rect 2178 -2922 2184 -2916
rect 2178 -2928 2184 -2922
rect 2178 -2934 2184 -2928
rect 2178 -2940 2184 -2934
rect 2178 -2946 2184 -2940
rect 2178 -2952 2184 -2946
rect 2178 -2958 2184 -2952
rect 2178 -2964 2184 -2958
rect 2178 -2970 2184 -2964
rect 2178 -2976 2184 -2970
rect 2178 -2982 2184 -2976
rect 2178 -2988 2184 -2982
rect 2178 -2994 2184 -2988
rect 2178 -3000 2184 -2994
rect 2178 -3006 2184 -3000
rect 2178 -3012 2184 -3006
rect 2178 -3018 2184 -3012
rect 2184 -216 2190 -210
rect 2184 -222 2190 -216
rect 2184 -228 2190 -222
rect 2184 -234 2190 -228
rect 2184 -240 2190 -234
rect 2184 -246 2190 -240
rect 2184 -252 2190 -246
rect 2184 -258 2190 -252
rect 2184 -264 2190 -258
rect 2184 -270 2190 -264
rect 2184 -276 2190 -270
rect 2184 -282 2190 -276
rect 2184 -288 2190 -282
rect 2184 -294 2190 -288
rect 2184 -300 2190 -294
rect 2184 -306 2190 -300
rect 2184 -312 2190 -306
rect 2184 -318 2190 -312
rect 2184 -324 2190 -318
rect 2184 -330 2190 -324
rect 2184 -336 2190 -330
rect 2184 -342 2190 -336
rect 2184 -348 2190 -342
rect 2184 -354 2190 -348
rect 2184 -360 2190 -354
rect 2184 -366 2190 -360
rect 2184 -372 2190 -366
rect 2184 -378 2190 -372
rect 2184 -384 2190 -378
rect 2184 -390 2190 -384
rect 2184 -396 2190 -390
rect 2184 -402 2190 -396
rect 2184 -408 2190 -402
rect 2184 -414 2190 -408
rect 2184 -420 2190 -414
rect 2184 -426 2190 -420
rect 2184 -432 2190 -426
rect 2184 -438 2190 -432
rect 2184 -444 2190 -438
rect 2184 -450 2190 -444
rect 2184 -456 2190 -450
rect 2184 -462 2190 -456
rect 2184 -468 2190 -462
rect 2184 -474 2190 -468
rect 2184 -480 2190 -474
rect 2184 -486 2190 -480
rect 2184 -492 2190 -486
rect 2184 -498 2190 -492
rect 2184 -504 2190 -498
rect 2184 -510 2190 -504
rect 2184 -516 2190 -510
rect 2184 -522 2190 -516
rect 2184 -528 2190 -522
rect 2184 -534 2190 -528
rect 2184 -540 2190 -534
rect 2184 -546 2190 -540
rect 2184 -552 2190 -546
rect 2184 -558 2190 -552
rect 2184 -564 2190 -558
rect 2184 -570 2190 -564
rect 2184 -576 2190 -570
rect 2184 -582 2190 -576
rect 2184 -588 2190 -582
rect 2184 -594 2190 -588
rect 2184 -600 2190 -594
rect 2184 -606 2190 -600
rect 2184 -612 2190 -606
rect 2184 -618 2190 -612
rect 2184 -624 2190 -618
rect 2184 -630 2190 -624
rect 2184 -636 2190 -630
rect 2184 -642 2190 -636
rect 2184 -648 2190 -642
rect 2184 -654 2190 -648
rect 2184 -660 2190 -654
rect 2184 -666 2190 -660
rect 2184 -672 2190 -666
rect 2184 -678 2190 -672
rect 2184 -684 2190 -678
rect 2184 -690 2190 -684
rect 2184 -696 2190 -690
rect 2184 -702 2190 -696
rect 2184 -708 2190 -702
rect 2184 -714 2190 -708
rect 2184 -720 2190 -714
rect 2184 -726 2190 -720
rect 2184 -732 2190 -726
rect 2184 -738 2190 -732
rect 2184 -744 2190 -738
rect 2184 -750 2190 -744
rect 2184 -756 2190 -750
rect 2184 -762 2190 -756
rect 2184 -768 2190 -762
rect 2184 -774 2190 -768
rect 2184 -780 2190 -774
rect 2184 -786 2190 -780
rect 2184 -792 2190 -786
rect 2184 -798 2190 -792
rect 2184 -804 2190 -798
rect 2184 -810 2190 -804
rect 2184 -816 2190 -810
rect 2184 -822 2190 -816
rect 2184 -828 2190 -822
rect 2184 -834 2190 -828
rect 2184 -840 2190 -834
rect 2184 -846 2190 -840
rect 2184 -852 2190 -846
rect 2184 -858 2190 -852
rect 2184 -864 2190 -858
rect 2184 -870 2190 -864
rect 2184 -876 2190 -870
rect 2184 -882 2190 -876
rect 2184 -888 2190 -882
rect 2184 -894 2190 -888
rect 2184 -900 2190 -894
rect 2184 -906 2190 -900
rect 2184 -912 2190 -906
rect 2184 -918 2190 -912
rect 2184 -924 2190 -918
rect 2184 -930 2190 -924
rect 2184 -936 2190 -930
rect 2184 -942 2190 -936
rect 2184 -948 2190 -942
rect 2184 -954 2190 -948
rect 2184 -960 2190 -954
rect 2184 -966 2190 -960
rect 2184 -972 2190 -966
rect 2184 -978 2190 -972
rect 2184 -984 2190 -978
rect 2184 -990 2190 -984
rect 2184 -996 2190 -990
rect 2184 -1002 2190 -996
rect 2184 -1008 2190 -1002
rect 2184 -1014 2190 -1008
rect 2184 -1020 2190 -1014
rect 2184 -1026 2190 -1020
rect 2184 -1032 2190 -1026
rect 2184 -1038 2190 -1032
rect 2184 -1044 2190 -1038
rect 2184 -1050 2190 -1044
rect 2184 -1056 2190 -1050
rect 2184 -1062 2190 -1056
rect 2184 -1068 2190 -1062
rect 2184 -1074 2190 -1068
rect 2184 -1080 2190 -1074
rect 2184 -1086 2190 -1080
rect 2184 -1092 2190 -1086
rect 2184 -1098 2190 -1092
rect 2184 -1104 2190 -1098
rect 2184 -1110 2190 -1104
rect 2184 -1116 2190 -1110
rect 2184 -1122 2190 -1116
rect 2184 -1128 2190 -1122
rect 2184 -1134 2190 -1128
rect 2184 -1140 2190 -1134
rect 2184 -1146 2190 -1140
rect 2184 -1152 2190 -1146
rect 2184 -1158 2190 -1152
rect 2184 -1164 2190 -1158
rect 2184 -1170 2190 -1164
rect 2184 -1176 2190 -1170
rect 2184 -1182 2190 -1176
rect 2184 -1188 2190 -1182
rect 2184 -1194 2190 -1188
rect 2184 -1200 2190 -1194
rect 2184 -1206 2190 -1200
rect 2184 -1212 2190 -1206
rect 2184 -1218 2190 -1212
rect 2184 -1224 2190 -1218
rect 2184 -1230 2190 -1224
rect 2184 -1236 2190 -1230
rect 2184 -1242 2190 -1236
rect 2184 -1248 2190 -1242
rect 2184 -1254 2190 -1248
rect 2184 -1260 2190 -1254
rect 2184 -1266 2190 -1260
rect 2184 -1272 2190 -1266
rect 2184 -1278 2190 -1272
rect 2184 -1284 2190 -1278
rect 2184 -1566 2190 -1560
rect 2184 -1572 2190 -1566
rect 2184 -1578 2190 -1572
rect 2184 -1584 2190 -1578
rect 2184 -1590 2190 -1584
rect 2184 -1596 2190 -1590
rect 2184 -1602 2190 -1596
rect 2184 -1608 2190 -1602
rect 2184 -1614 2190 -1608
rect 2184 -1620 2190 -1614
rect 2184 -1626 2190 -1620
rect 2184 -1632 2190 -1626
rect 2184 -1638 2190 -1632
rect 2184 -1644 2190 -1638
rect 2184 -1650 2190 -1644
rect 2184 -1656 2190 -1650
rect 2184 -1662 2190 -1656
rect 2184 -1668 2190 -1662
rect 2184 -1674 2190 -1668
rect 2184 -1680 2190 -1674
rect 2184 -1686 2190 -1680
rect 2184 -1692 2190 -1686
rect 2184 -1698 2190 -1692
rect 2184 -1704 2190 -1698
rect 2184 -1710 2190 -1704
rect 2184 -1716 2190 -1710
rect 2184 -1722 2190 -1716
rect 2184 -1728 2190 -1722
rect 2184 -1734 2190 -1728
rect 2184 -1740 2190 -1734
rect 2184 -1746 2190 -1740
rect 2184 -1752 2190 -1746
rect 2184 -1758 2190 -1752
rect 2184 -1764 2190 -1758
rect 2184 -1770 2190 -1764
rect 2184 -1776 2190 -1770
rect 2184 -1782 2190 -1776
rect 2184 -1788 2190 -1782
rect 2184 -1794 2190 -1788
rect 2184 -1800 2190 -1794
rect 2184 -1806 2190 -1800
rect 2184 -1812 2190 -1806
rect 2184 -1818 2190 -1812
rect 2184 -1824 2190 -1818
rect 2184 -1830 2190 -1824
rect 2184 -1836 2190 -1830
rect 2184 -1842 2190 -1836
rect 2184 -1848 2190 -1842
rect 2184 -1854 2190 -1848
rect 2184 -1860 2190 -1854
rect 2184 -1866 2190 -1860
rect 2184 -1872 2190 -1866
rect 2184 -1878 2190 -1872
rect 2184 -1884 2190 -1878
rect 2184 -1890 2190 -1884
rect 2184 -1896 2190 -1890
rect 2184 -1902 2190 -1896
rect 2184 -1908 2190 -1902
rect 2184 -1914 2190 -1908
rect 2184 -1920 2190 -1914
rect 2184 -1926 2190 -1920
rect 2184 -1932 2190 -1926
rect 2184 -1938 2190 -1932
rect 2184 -1944 2190 -1938
rect 2184 -1950 2190 -1944
rect 2184 -1956 2190 -1950
rect 2184 -1962 2190 -1956
rect 2184 -1968 2190 -1962
rect 2184 -1974 2190 -1968
rect 2184 -1980 2190 -1974
rect 2184 -1986 2190 -1980
rect 2184 -1992 2190 -1986
rect 2184 -1998 2190 -1992
rect 2184 -2004 2190 -1998
rect 2184 -2010 2190 -2004
rect 2184 -2016 2190 -2010
rect 2184 -2022 2190 -2016
rect 2184 -2028 2190 -2022
rect 2184 -2034 2190 -2028
rect 2184 -2040 2190 -2034
rect 2184 -2046 2190 -2040
rect 2184 -2052 2190 -2046
rect 2184 -2058 2190 -2052
rect 2184 -2064 2190 -2058
rect 2184 -2070 2190 -2064
rect 2184 -2076 2190 -2070
rect 2184 -2082 2190 -2076
rect 2184 -2088 2190 -2082
rect 2184 -2094 2190 -2088
rect 2184 -2100 2190 -2094
rect 2184 -2106 2190 -2100
rect 2184 -2112 2190 -2106
rect 2184 -2118 2190 -2112
rect 2184 -2124 2190 -2118
rect 2184 -2130 2190 -2124
rect 2184 -2136 2190 -2130
rect 2184 -2142 2190 -2136
rect 2184 -2148 2190 -2142
rect 2184 -2154 2190 -2148
rect 2184 -2160 2190 -2154
rect 2184 -2166 2190 -2160
rect 2184 -2172 2190 -2166
rect 2184 -2178 2190 -2172
rect 2184 -2184 2190 -2178
rect 2184 -2190 2190 -2184
rect 2184 -2196 2190 -2190
rect 2184 -2202 2190 -2196
rect 2184 -2208 2190 -2202
rect 2184 -2214 2190 -2208
rect 2184 -2220 2190 -2214
rect 2184 -2226 2190 -2220
rect 2184 -2232 2190 -2226
rect 2184 -2238 2190 -2232
rect 2184 -2244 2190 -2238
rect 2184 -2250 2190 -2244
rect 2184 -2256 2190 -2250
rect 2184 -2262 2190 -2256
rect 2184 -2268 2190 -2262
rect 2184 -2274 2190 -2268
rect 2184 -2280 2190 -2274
rect 2184 -2286 2190 -2280
rect 2184 -2292 2190 -2286
rect 2184 -2298 2190 -2292
rect 2184 -2304 2190 -2298
rect 2184 -2310 2190 -2304
rect 2184 -2316 2190 -2310
rect 2184 -2322 2190 -2316
rect 2184 -2328 2190 -2322
rect 2184 -2334 2190 -2328
rect 2184 -2340 2190 -2334
rect 2184 -2346 2190 -2340
rect 2184 -2352 2190 -2346
rect 2184 -2358 2190 -2352
rect 2184 -2364 2190 -2358
rect 2184 -2544 2190 -2538
rect 2184 -2550 2190 -2544
rect 2184 -2556 2190 -2550
rect 2184 -2562 2190 -2556
rect 2184 -2568 2190 -2562
rect 2184 -2574 2190 -2568
rect 2184 -2580 2190 -2574
rect 2184 -2586 2190 -2580
rect 2184 -2592 2190 -2586
rect 2184 -2598 2190 -2592
rect 2184 -2604 2190 -2598
rect 2184 -2610 2190 -2604
rect 2184 -2616 2190 -2610
rect 2184 -2622 2190 -2616
rect 2184 -2628 2190 -2622
rect 2184 -2634 2190 -2628
rect 2184 -2640 2190 -2634
rect 2184 -2646 2190 -2640
rect 2184 -2652 2190 -2646
rect 2184 -2658 2190 -2652
rect 2184 -2664 2190 -2658
rect 2184 -2670 2190 -2664
rect 2184 -2676 2190 -2670
rect 2184 -2682 2190 -2676
rect 2184 -2688 2190 -2682
rect 2184 -2694 2190 -2688
rect 2184 -2700 2190 -2694
rect 2184 -2706 2190 -2700
rect 2184 -2712 2190 -2706
rect 2184 -2718 2190 -2712
rect 2184 -2724 2190 -2718
rect 2184 -2730 2190 -2724
rect 2184 -2736 2190 -2730
rect 2184 -2742 2190 -2736
rect 2184 -2748 2190 -2742
rect 2184 -2754 2190 -2748
rect 2184 -2760 2190 -2754
rect 2184 -2766 2190 -2760
rect 2184 -2772 2190 -2766
rect 2184 -2778 2190 -2772
rect 2184 -2784 2190 -2778
rect 2184 -2790 2190 -2784
rect 2184 -2796 2190 -2790
rect 2184 -2802 2190 -2796
rect 2184 -2808 2190 -2802
rect 2184 -2814 2190 -2808
rect 2184 -2820 2190 -2814
rect 2184 -2826 2190 -2820
rect 2184 -2832 2190 -2826
rect 2184 -2838 2190 -2832
rect 2184 -2844 2190 -2838
rect 2184 -2850 2190 -2844
rect 2184 -2856 2190 -2850
rect 2184 -2862 2190 -2856
rect 2184 -2868 2190 -2862
rect 2184 -2874 2190 -2868
rect 2184 -2880 2190 -2874
rect 2184 -2886 2190 -2880
rect 2184 -2892 2190 -2886
rect 2184 -2898 2190 -2892
rect 2184 -2904 2190 -2898
rect 2184 -2910 2190 -2904
rect 2184 -2916 2190 -2910
rect 2184 -2922 2190 -2916
rect 2184 -2928 2190 -2922
rect 2184 -2934 2190 -2928
rect 2184 -2940 2190 -2934
rect 2184 -2946 2190 -2940
rect 2184 -2952 2190 -2946
rect 2184 -2958 2190 -2952
rect 2184 -2964 2190 -2958
rect 2184 -2970 2190 -2964
rect 2184 -2976 2190 -2970
rect 2184 -2982 2190 -2976
rect 2184 -2988 2190 -2982
rect 2184 -2994 2190 -2988
rect 2184 -3000 2190 -2994
rect 2184 -3006 2190 -3000
rect 2184 -3012 2190 -3006
rect 2184 -3018 2190 -3012
rect 2190 -210 2196 -204
rect 2190 -216 2196 -210
rect 2190 -222 2196 -216
rect 2190 -228 2196 -222
rect 2190 -234 2196 -228
rect 2190 -240 2196 -234
rect 2190 -246 2196 -240
rect 2190 -252 2196 -246
rect 2190 -258 2196 -252
rect 2190 -264 2196 -258
rect 2190 -270 2196 -264
rect 2190 -276 2196 -270
rect 2190 -282 2196 -276
rect 2190 -288 2196 -282
rect 2190 -294 2196 -288
rect 2190 -300 2196 -294
rect 2190 -306 2196 -300
rect 2190 -312 2196 -306
rect 2190 -318 2196 -312
rect 2190 -324 2196 -318
rect 2190 -330 2196 -324
rect 2190 -336 2196 -330
rect 2190 -342 2196 -336
rect 2190 -348 2196 -342
rect 2190 -354 2196 -348
rect 2190 -360 2196 -354
rect 2190 -366 2196 -360
rect 2190 -372 2196 -366
rect 2190 -378 2196 -372
rect 2190 -384 2196 -378
rect 2190 -390 2196 -384
rect 2190 -396 2196 -390
rect 2190 -402 2196 -396
rect 2190 -408 2196 -402
rect 2190 -414 2196 -408
rect 2190 -420 2196 -414
rect 2190 -426 2196 -420
rect 2190 -432 2196 -426
rect 2190 -438 2196 -432
rect 2190 -444 2196 -438
rect 2190 -450 2196 -444
rect 2190 -456 2196 -450
rect 2190 -462 2196 -456
rect 2190 -468 2196 -462
rect 2190 -474 2196 -468
rect 2190 -480 2196 -474
rect 2190 -486 2196 -480
rect 2190 -492 2196 -486
rect 2190 -498 2196 -492
rect 2190 -504 2196 -498
rect 2190 -510 2196 -504
rect 2190 -516 2196 -510
rect 2190 -522 2196 -516
rect 2190 -528 2196 -522
rect 2190 -534 2196 -528
rect 2190 -540 2196 -534
rect 2190 -546 2196 -540
rect 2190 -552 2196 -546
rect 2190 -558 2196 -552
rect 2190 -564 2196 -558
rect 2190 -570 2196 -564
rect 2190 -576 2196 -570
rect 2190 -582 2196 -576
rect 2190 -588 2196 -582
rect 2190 -594 2196 -588
rect 2190 -600 2196 -594
rect 2190 -606 2196 -600
rect 2190 -612 2196 -606
rect 2190 -618 2196 -612
rect 2190 -624 2196 -618
rect 2190 -630 2196 -624
rect 2190 -636 2196 -630
rect 2190 -642 2196 -636
rect 2190 -648 2196 -642
rect 2190 -654 2196 -648
rect 2190 -660 2196 -654
rect 2190 -666 2196 -660
rect 2190 -672 2196 -666
rect 2190 -678 2196 -672
rect 2190 -684 2196 -678
rect 2190 -690 2196 -684
rect 2190 -696 2196 -690
rect 2190 -702 2196 -696
rect 2190 -708 2196 -702
rect 2190 -714 2196 -708
rect 2190 -720 2196 -714
rect 2190 -726 2196 -720
rect 2190 -732 2196 -726
rect 2190 -738 2196 -732
rect 2190 -744 2196 -738
rect 2190 -750 2196 -744
rect 2190 -756 2196 -750
rect 2190 -762 2196 -756
rect 2190 -768 2196 -762
rect 2190 -774 2196 -768
rect 2190 -780 2196 -774
rect 2190 -786 2196 -780
rect 2190 -792 2196 -786
rect 2190 -798 2196 -792
rect 2190 -804 2196 -798
rect 2190 -810 2196 -804
rect 2190 -816 2196 -810
rect 2190 -822 2196 -816
rect 2190 -828 2196 -822
rect 2190 -834 2196 -828
rect 2190 -840 2196 -834
rect 2190 -846 2196 -840
rect 2190 -852 2196 -846
rect 2190 -858 2196 -852
rect 2190 -864 2196 -858
rect 2190 -870 2196 -864
rect 2190 -876 2196 -870
rect 2190 -882 2196 -876
rect 2190 -888 2196 -882
rect 2190 -894 2196 -888
rect 2190 -900 2196 -894
rect 2190 -906 2196 -900
rect 2190 -912 2196 -906
rect 2190 -918 2196 -912
rect 2190 -924 2196 -918
rect 2190 -930 2196 -924
rect 2190 -936 2196 -930
rect 2190 -942 2196 -936
rect 2190 -948 2196 -942
rect 2190 -954 2196 -948
rect 2190 -960 2196 -954
rect 2190 -966 2196 -960
rect 2190 -972 2196 -966
rect 2190 -978 2196 -972
rect 2190 -984 2196 -978
rect 2190 -990 2196 -984
rect 2190 -996 2196 -990
rect 2190 -1002 2196 -996
rect 2190 -1008 2196 -1002
rect 2190 -1014 2196 -1008
rect 2190 -1020 2196 -1014
rect 2190 -1026 2196 -1020
rect 2190 -1032 2196 -1026
rect 2190 -1038 2196 -1032
rect 2190 -1044 2196 -1038
rect 2190 -1050 2196 -1044
rect 2190 -1056 2196 -1050
rect 2190 -1062 2196 -1056
rect 2190 -1068 2196 -1062
rect 2190 -1074 2196 -1068
rect 2190 -1080 2196 -1074
rect 2190 -1086 2196 -1080
rect 2190 -1092 2196 -1086
rect 2190 -1098 2196 -1092
rect 2190 -1104 2196 -1098
rect 2190 -1110 2196 -1104
rect 2190 -1116 2196 -1110
rect 2190 -1122 2196 -1116
rect 2190 -1128 2196 -1122
rect 2190 -1134 2196 -1128
rect 2190 -1140 2196 -1134
rect 2190 -1146 2196 -1140
rect 2190 -1152 2196 -1146
rect 2190 -1158 2196 -1152
rect 2190 -1164 2196 -1158
rect 2190 -1170 2196 -1164
rect 2190 -1176 2196 -1170
rect 2190 -1182 2196 -1176
rect 2190 -1188 2196 -1182
rect 2190 -1194 2196 -1188
rect 2190 -1200 2196 -1194
rect 2190 -1206 2196 -1200
rect 2190 -1212 2196 -1206
rect 2190 -1218 2196 -1212
rect 2190 -1224 2196 -1218
rect 2190 -1230 2196 -1224
rect 2190 -1236 2196 -1230
rect 2190 -1242 2196 -1236
rect 2190 -1248 2196 -1242
rect 2190 -1254 2196 -1248
rect 2190 -1260 2196 -1254
rect 2190 -1266 2196 -1260
rect 2190 -1560 2196 -1554
rect 2190 -1566 2196 -1560
rect 2190 -1572 2196 -1566
rect 2190 -1578 2196 -1572
rect 2190 -1584 2196 -1578
rect 2190 -1590 2196 -1584
rect 2190 -1596 2196 -1590
rect 2190 -1602 2196 -1596
rect 2190 -1608 2196 -1602
rect 2190 -1614 2196 -1608
rect 2190 -1620 2196 -1614
rect 2190 -1626 2196 -1620
rect 2190 -1632 2196 -1626
rect 2190 -1638 2196 -1632
rect 2190 -1644 2196 -1638
rect 2190 -1650 2196 -1644
rect 2190 -1656 2196 -1650
rect 2190 -1662 2196 -1656
rect 2190 -1668 2196 -1662
rect 2190 -1674 2196 -1668
rect 2190 -1680 2196 -1674
rect 2190 -1686 2196 -1680
rect 2190 -1692 2196 -1686
rect 2190 -1698 2196 -1692
rect 2190 -1704 2196 -1698
rect 2190 -1710 2196 -1704
rect 2190 -1716 2196 -1710
rect 2190 -1722 2196 -1716
rect 2190 -1728 2196 -1722
rect 2190 -1734 2196 -1728
rect 2190 -1740 2196 -1734
rect 2190 -1746 2196 -1740
rect 2190 -1752 2196 -1746
rect 2190 -1758 2196 -1752
rect 2190 -1764 2196 -1758
rect 2190 -1770 2196 -1764
rect 2190 -1776 2196 -1770
rect 2190 -1782 2196 -1776
rect 2190 -1788 2196 -1782
rect 2190 -1794 2196 -1788
rect 2190 -1800 2196 -1794
rect 2190 -1806 2196 -1800
rect 2190 -1812 2196 -1806
rect 2190 -1818 2196 -1812
rect 2190 -1824 2196 -1818
rect 2190 -1830 2196 -1824
rect 2190 -1836 2196 -1830
rect 2190 -1842 2196 -1836
rect 2190 -1848 2196 -1842
rect 2190 -1854 2196 -1848
rect 2190 -1860 2196 -1854
rect 2190 -1866 2196 -1860
rect 2190 -1872 2196 -1866
rect 2190 -1878 2196 -1872
rect 2190 -1884 2196 -1878
rect 2190 -1890 2196 -1884
rect 2190 -1896 2196 -1890
rect 2190 -1902 2196 -1896
rect 2190 -1908 2196 -1902
rect 2190 -1914 2196 -1908
rect 2190 -1920 2196 -1914
rect 2190 -1926 2196 -1920
rect 2190 -1932 2196 -1926
rect 2190 -1938 2196 -1932
rect 2190 -1944 2196 -1938
rect 2190 -1950 2196 -1944
rect 2190 -1956 2196 -1950
rect 2190 -1962 2196 -1956
rect 2190 -1968 2196 -1962
rect 2190 -1974 2196 -1968
rect 2190 -1980 2196 -1974
rect 2190 -1986 2196 -1980
rect 2190 -1992 2196 -1986
rect 2190 -1998 2196 -1992
rect 2190 -2004 2196 -1998
rect 2190 -2010 2196 -2004
rect 2190 -2016 2196 -2010
rect 2190 -2022 2196 -2016
rect 2190 -2028 2196 -2022
rect 2190 -2034 2196 -2028
rect 2190 -2040 2196 -2034
rect 2190 -2046 2196 -2040
rect 2190 -2052 2196 -2046
rect 2190 -2058 2196 -2052
rect 2190 -2064 2196 -2058
rect 2190 -2070 2196 -2064
rect 2190 -2076 2196 -2070
rect 2190 -2082 2196 -2076
rect 2190 -2088 2196 -2082
rect 2190 -2094 2196 -2088
rect 2190 -2100 2196 -2094
rect 2190 -2106 2196 -2100
rect 2190 -2112 2196 -2106
rect 2190 -2118 2196 -2112
rect 2190 -2124 2196 -2118
rect 2190 -2130 2196 -2124
rect 2190 -2136 2196 -2130
rect 2190 -2142 2196 -2136
rect 2190 -2148 2196 -2142
rect 2190 -2154 2196 -2148
rect 2190 -2160 2196 -2154
rect 2190 -2166 2196 -2160
rect 2190 -2172 2196 -2166
rect 2190 -2178 2196 -2172
rect 2190 -2184 2196 -2178
rect 2190 -2190 2196 -2184
rect 2190 -2196 2196 -2190
rect 2190 -2202 2196 -2196
rect 2190 -2208 2196 -2202
rect 2190 -2214 2196 -2208
rect 2190 -2220 2196 -2214
rect 2190 -2226 2196 -2220
rect 2190 -2232 2196 -2226
rect 2190 -2238 2196 -2232
rect 2190 -2244 2196 -2238
rect 2190 -2250 2196 -2244
rect 2190 -2256 2196 -2250
rect 2190 -2262 2196 -2256
rect 2190 -2268 2196 -2262
rect 2190 -2274 2196 -2268
rect 2190 -2280 2196 -2274
rect 2190 -2286 2196 -2280
rect 2190 -2292 2196 -2286
rect 2190 -2298 2196 -2292
rect 2190 -2304 2196 -2298
rect 2190 -2310 2196 -2304
rect 2190 -2316 2196 -2310
rect 2190 -2322 2196 -2316
rect 2190 -2328 2196 -2322
rect 2190 -2334 2196 -2328
rect 2190 -2340 2196 -2334
rect 2190 -2346 2196 -2340
rect 2190 -2352 2196 -2346
rect 2190 -2358 2196 -2352
rect 2190 -2544 2196 -2538
rect 2190 -2550 2196 -2544
rect 2190 -2556 2196 -2550
rect 2190 -2562 2196 -2556
rect 2190 -2568 2196 -2562
rect 2190 -2574 2196 -2568
rect 2190 -2580 2196 -2574
rect 2190 -2586 2196 -2580
rect 2190 -2592 2196 -2586
rect 2190 -2598 2196 -2592
rect 2190 -2604 2196 -2598
rect 2190 -2610 2196 -2604
rect 2190 -2616 2196 -2610
rect 2190 -2622 2196 -2616
rect 2190 -2628 2196 -2622
rect 2190 -2634 2196 -2628
rect 2190 -2640 2196 -2634
rect 2190 -2646 2196 -2640
rect 2190 -2652 2196 -2646
rect 2190 -2658 2196 -2652
rect 2190 -2664 2196 -2658
rect 2190 -2670 2196 -2664
rect 2190 -2676 2196 -2670
rect 2190 -2682 2196 -2676
rect 2190 -2688 2196 -2682
rect 2190 -2694 2196 -2688
rect 2190 -2700 2196 -2694
rect 2190 -2706 2196 -2700
rect 2190 -2712 2196 -2706
rect 2190 -2718 2196 -2712
rect 2190 -2724 2196 -2718
rect 2190 -2730 2196 -2724
rect 2190 -2736 2196 -2730
rect 2190 -2742 2196 -2736
rect 2190 -2748 2196 -2742
rect 2190 -2754 2196 -2748
rect 2190 -2760 2196 -2754
rect 2190 -2766 2196 -2760
rect 2190 -2772 2196 -2766
rect 2190 -2778 2196 -2772
rect 2190 -2784 2196 -2778
rect 2190 -2790 2196 -2784
rect 2190 -2796 2196 -2790
rect 2190 -2802 2196 -2796
rect 2190 -2808 2196 -2802
rect 2190 -2814 2196 -2808
rect 2190 -2820 2196 -2814
rect 2190 -2826 2196 -2820
rect 2190 -2832 2196 -2826
rect 2190 -2838 2196 -2832
rect 2190 -2844 2196 -2838
rect 2190 -2850 2196 -2844
rect 2190 -2856 2196 -2850
rect 2190 -2862 2196 -2856
rect 2190 -2868 2196 -2862
rect 2190 -2874 2196 -2868
rect 2190 -2880 2196 -2874
rect 2190 -2886 2196 -2880
rect 2190 -2892 2196 -2886
rect 2190 -2898 2196 -2892
rect 2190 -2904 2196 -2898
rect 2190 -2910 2196 -2904
rect 2190 -2916 2196 -2910
rect 2190 -2922 2196 -2916
rect 2190 -2928 2196 -2922
rect 2190 -2934 2196 -2928
rect 2190 -2940 2196 -2934
rect 2190 -2946 2196 -2940
rect 2190 -2952 2196 -2946
rect 2190 -2958 2196 -2952
rect 2190 -2964 2196 -2958
rect 2190 -2970 2196 -2964
rect 2190 -2976 2196 -2970
rect 2190 -2982 2196 -2976
rect 2190 -2988 2196 -2982
rect 2190 -2994 2196 -2988
rect 2190 -3000 2196 -2994
rect 2190 -3006 2196 -3000
rect 2190 -3012 2196 -3006
rect 2196 -204 2202 -198
rect 2196 -210 2202 -204
rect 2196 -216 2202 -210
rect 2196 -222 2202 -216
rect 2196 -228 2202 -222
rect 2196 -234 2202 -228
rect 2196 -240 2202 -234
rect 2196 -246 2202 -240
rect 2196 -252 2202 -246
rect 2196 -258 2202 -252
rect 2196 -264 2202 -258
rect 2196 -270 2202 -264
rect 2196 -276 2202 -270
rect 2196 -282 2202 -276
rect 2196 -288 2202 -282
rect 2196 -294 2202 -288
rect 2196 -300 2202 -294
rect 2196 -306 2202 -300
rect 2196 -312 2202 -306
rect 2196 -318 2202 -312
rect 2196 -324 2202 -318
rect 2196 -330 2202 -324
rect 2196 -336 2202 -330
rect 2196 -342 2202 -336
rect 2196 -348 2202 -342
rect 2196 -354 2202 -348
rect 2196 -360 2202 -354
rect 2196 -366 2202 -360
rect 2196 -372 2202 -366
rect 2196 -378 2202 -372
rect 2196 -384 2202 -378
rect 2196 -390 2202 -384
rect 2196 -396 2202 -390
rect 2196 -402 2202 -396
rect 2196 -408 2202 -402
rect 2196 -414 2202 -408
rect 2196 -420 2202 -414
rect 2196 -426 2202 -420
rect 2196 -432 2202 -426
rect 2196 -438 2202 -432
rect 2196 -444 2202 -438
rect 2196 -450 2202 -444
rect 2196 -456 2202 -450
rect 2196 -462 2202 -456
rect 2196 -468 2202 -462
rect 2196 -474 2202 -468
rect 2196 -480 2202 -474
rect 2196 -486 2202 -480
rect 2196 -492 2202 -486
rect 2196 -498 2202 -492
rect 2196 -504 2202 -498
rect 2196 -510 2202 -504
rect 2196 -516 2202 -510
rect 2196 -522 2202 -516
rect 2196 -528 2202 -522
rect 2196 -534 2202 -528
rect 2196 -540 2202 -534
rect 2196 -546 2202 -540
rect 2196 -552 2202 -546
rect 2196 -558 2202 -552
rect 2196 -564 2202 -558
rect 2196 -570 2202 -564
rect 2196 -576 2202 -570
rect 2196 -582 2202 -576
rect 2196 -588 2202 -582
rect 2196 -594 2202 -588
rect 2196 -600 2202 -594
rect 2196 -606 2202 -600
rect 2196 -612 2202 -606
rect 2196 -618 2202 -612
rect 2196 -624 2202 -618
rect 2196 -630 2202 -624
rect 2196 -636 2202 -630
rect 2196 -642 2202 -636
rect 2196 -648 2202 -642
rect 2196 -654 2202 -648
rect 2196 -660 2202 -654
rect 2196 -666 2202 -660
rect 2196 -672 2202 -666
rect 2196 -678 2202 -672
rect 2196 -684 2202 -678
rect 2196 -690 2202 -684
rect 2196 -696 2202 -690
rect 2196 -702 2202 -696
rect 2196 -708 2202 -702
rect 2196 -714 2202 -708
rect 2196 -720 2202 -714
rect 2196 -726 2202 -720
rect 2196 -732 2202 -726
rect 2196 -738 2202 -732
rect 2196 -744 2202 -738
rect 2196 -750 2202 -744
rect 2196 -756 2202 -750
rect 2196 -762 2202 -756
rect 2196 -768 2202 -762
rect 2196 -774 2202 -768
rect 2196 -780 2202 -774
rect 2196 -786 2202 -780
rect 2196 -792 2202 -786
rect 2196 -798 2202 -792
rect 2196 -804 2202 -798
rect 2196 -810 2202 -804
rect 2196 -816 2202 -810
rect 2196 -822 2202 -816
rect 2196 -828 2202 -822
rect 2196 -834 2202 -828
rect 2196 -840 2202 -834
rect 2196 -846 2202 -840
rect 2196 -852 2202 -846
rect 2196 -858 2202 -852
rect 2196 -864 2202 -858
rect 2196 -870 2202 -864
rect 2196 -876 2202 -870
rect 2196 -882 2202 -876
rect 2196 -888 2202 -882
rect 2196 -894 2202 -888
rect 2196 -900 2202 -894
rect 2196 -906 2202 -900
rect 2196 -912 2202 -906
rect 2196 -918 2202 -912
rect 2196 -924 2202 -918
rect 2196 -930 2202 -924
rect 2196 -936 2202 -930
rect 2196 -942 2202 -936
rect 2196 -948 2202 -942
rect 2196 -954 2202 -948
rect 2196 -960 2202 -954
rect 2196 -966 2202 -960
rect 2196 -972 2202 -966
rect 2196 -978 2202 -972
rect 2196 -984 2202 -978
rect 2196 -990 2202 -984
rect 2196 -996 2202 -990
rect 2196 -1002 2202 -996
rect 2196 -1008 2202 -1002
rect 2196 -1014 2202 -1008
rect 2196 -1020 2202 -1014
rect 2196 -1026 2202 -1020
rect 2196 -1032 2202 -1026
rect 2196 -1038 2202 -1032
rect 2196 -1044 2202 -1038
rect 2196 -1050 2202 -1044
rect 2196 -1056 2202 -1050
rect 2196 -1062 2202 -1056
rect 2196 -1068 2202 -1062
rect 2196 -1074 2202 -1068
rect 2196 -1080 2202 -1074
rect 2196 -1086 2202 -1080
rect 2196 -1092 2202 -1086
rect 2196 -1098 2202 -1092
rect 2196 -1104 2202 -1098
rect 2196 -1110 2202 -1104
rect 2196 -1116 2202 -1110
rect 2196 -1122 2202 -1116
rect 2196 -1128 2202 -1122
rect 2196 -1134 2202 -1128
rect 2196 -1140 2202 -1134
rect 2196 -1146 2202 -1140
rect 2196 -1152 2202 -1146
rect 2196 -1158 2202 -1152
rect 2196 -1164 2202 -1158
rect 2196 -1170 2202 -1164
rect 2196 -1176 2202 -1170
rect 2196 -1182 2202 -1176
rect 2196 -1188 2202 -1182
rect 2196 -1194 2202 -1188
rect 2196 -1200 2202 -1194
rect 2196 -1206 2202 -1200
rect 2196 -1212 2202 -1206
rect 2196 -1218 2202 -1212
rect 2196 -1224 2202 -1218
rect 2196 -1230 2202 -1224
rect 2196 -1236 2202 -1230
rect 2196 -1242 2202 -1236
rect 2196 -1248 2202 -1242
rect 2196 -1254 2202 -1248
rect 2196 -1554 2202 -1548
rect 2196 -1560 2202 -1554
rect 2196 -1566 2202 -1560
rect 2196 -1572 2202 -1566
rect 2196 -1578 2202 -1572
rect 2196 -1584 2202 -1578
rect 2196 -1590 2202 -1584
rect 2196 -1596 2202 -1590
rect 2196 -1602 2202 -1596
rect 2196 -1608 2202 -1602
rect 2196 -1614 2202 -1608
rect 2196 -1620 2202 -1614
rect 2196 -1626 2202 -1620
rect 2196 -1632 2202 -1626
rect 2196 -1638 2202 -1632
rect 2196 -1644 2202 -1638
rect 2196 -1650 2202 -1644
rect 2196 -1656 2202 -1650
rect 2196 -1662 2202 -1656
rect 2196 -1668 2202 -1662
rect 2196 -1674 2202 -1668
rect 2196 -1680 2202 -1674
rect 2196 -1686 2202 -1680
rect 2196 -1692 2202 -1686
rect 2196 -1698 2202 -1692
rect 2196 -1704 2202 -1698
rect 2196 -1710 2202 -1704
rect 2196 -1716 2202 -1710
rect 2196 -1722 2202 -1716
rect 2196 -1728 2202 -1722
rect 2196 -1734 2202 -1728
rect 2196 -1740 2202 -1734
rect 2196 -1746 2202 -1740
rect 2196 -1752 2202 -1746
rect 2196 -1758 2202 -1752
rect 2196 -1764 2202 -1758
rect 2196 -1770 2202 -1764
rect 2196 -1776 2202 -1770
rect 2196 -1782 2202 -1776
rect 2196 -1788 2202 -1782
rect 2196 -1794 2202 -1788
rect 2196 -1800 2202 -1794
rect 2196 -1806 2202 -1800
rect 2196 -1812 2202 -1806
rect 2196 -1818 2202 -1812
rect 2196 -1824 2202 -1818
rect 2196 -1830 2202 -1824
rect 2196 -1836 2202 -1830
rect 2196 -1842 2202 -1836
rect 2196 -1848 2202 -1842
rect 2196 -1854 2202 -1848
rect 2196 -1860 2202 -1854
rect 2196 -1866 2202 -1860
rect 2196 -1872 2202 -1866
rect 2196 -1878 2202 -1872
rect 2196 -1884 2202 -1878
rect 2196 -1890 2202 -1884
rect 2196 -1896 2202 -1890
rect 2196 -1902 2202 -1896
rect 2196 -1908 2202 -1902
rect 2196 -1914 2202 -1908
rect 2196 -1920 2202 -1914
rect 2196 -1926 2202 -1920
rect 2196 -1932 2202 -1926
rect 2196 -1938 2202 -1932
rect 2196 -1944 2202 -1938
rect 2196 -1950 2202 -1944
rect 2196 -1956 2202 -1950
rect 2196 -1962 2202 -1956
rect 2196 -1968 2202 -1962
rect 2196 -1974 2202 -1968
rect 2196 -1980 2202 -1974
rect 2196 -1986 2202 -1980
rect 2196 -1992 2202 -1986
rect 2196 -1998 2202 -1992
rect 2196 -2004 2202 -1998
rect 2196 -2010 2202 -2004
rect 2196 -2016 2202 -2010
rect 2196 -2022 2202 -2016
rect 2196 -2028 2202 -2022
rect 2196 -2034 2202 -2028
rect 2196 -2040 2202 -2034
rect 2196 -2046 2202 -2040
rect 2196 -2052 2202 -2046
rect 2196 -2058 2202 -2052
rect 2196 -2064 2202 -2058
rect 2196 -2070 2202 -2064
rect 2196 -2076 2202 -2070
rect 2196 -2082 2202 -2076
rect 2196 -2088 2202 -2082
rect 2196 -2094 2202 -2088
rect 2196 -2100 2202 -2094
rect 2196 -2106 2202 -2100
rect 2196 -2112 2202 -2106
rect 2196 -2118 2202 -2112
rect 2196 -2124 2202 -2118
rect 2196 -2130 2202 -2124
rect 2196 -2136 2202 -2130
rect 2196 -2142 2202 -2136
rect 2196 -2148 2202 -2142
rect 2196 -2154 2202 -2148
rect 2196 -2160 2202 -2154
rect 2196 -2166 2202 -2160
rect 2196 -2172 2202 -2166
rect 2196 -2178 2202 -2172
rect 2196 -2184 2202 -2178
rect 2196 -2190 2202 -2184
rect 2196 -2196 2202 -2190
rect 2196 -2202 2202 -2196
rect 2196 -2208 2202 -2202
rect 2196 -2214 2202 -2208
rect 2196 -2220 2202 -2214
rect 2196 -2226 2202 -2220
rect 2196 -2232 2202 -2226
rect 2196 -2238 2202 -2232
rect 2196 -2244 2202 -2238
rect 2196 -2250 2202 -2244
rect 2196 -2256 2202 -2250
rect 2196 -2262 2202 -2256
rect 2196 -2268 2202 -2262
rect 2196 -2274 2202 -2268
rect 2196 -2280 2202 -2274
rect 2196 -2286 2202 -2280
rect 2196 -2292 2202 -2286
rect 2196 -2298 2202 -2292
rect 2196 -2304 2202 -2298
rect 2196 -2310 2202 -2304
rect 2196 -2316 2202 -2310
rect 2196 -2322 2202 -2316
rect 2196 -2328 2202 -2322
rect 2196 -2334 2202 -2328
rect 2196 -2340 2202 -2334
rect 2196 -2346 2202 -2340
rect 2196 -2538 2202 -2532
rect 2196 -2544 2202 -2538
rect 2196 -2550 2202 -2544
rect 2196 -2556 2202 -2550
rect 2196 -2562 2202 -2556
rect 2196 -2568 2202 -2562
rect 2196 -2574 2202 -2568
rect 2196 -2580 2202 -2574
rect 2196 -2586 2202 -2580
rect 2196 -2592 2202 -2586
rect 2196 -2598 2202 -2592
rect 2196 -2604 2202 -2598
rect 2196 -2610 2202 -2604
rect 2196 -2616 2202 -2610
rect 2196 -2622 2202 -2616
rect 2196 -2628 2202 -2622
rect 2196 -2634 2202 -2628
rect 2196 -2640 2202 -2634
rect 2196 -2646 2202 -2640
rect 2196 -2652 2202 -2646
rect 2196 -2658 2202 -2652
rect 2196 -2664 2202 -2658
rect 2196 -2670 2202 -2664
rect 2196 -2676 2202 -2670
rect 2196 -2682 2202 -2676
rect 2196 -2688 2202 -2682
rect 2196 -2694 2202 -2688
rect 2196 -2700 2202 -2694
rect 2196 -2706 2202 -2700
rect 2196 -2712 2202 -2706
rect 2196 -2718 2202 -2712
rect 2196 -2724 2202 -2718
rect 2196 -2730 2202 -2724
rect 2196 -2736 2202 -2730
rect 2196 -2742 2202 -2736
rect 2196 -2748 2202 -2742
rect 2196 -2754 2202 -2748
rect 2196 -2760 2202 -2754
rect 2196 -2766 2202 -2760
rect 2196 -2772 2202 -2766
rect 2196 -2778 2202 -2772
rect 2196 -2784 2202 -2778
rect 2196 -2790 2202 -2784
rect 2196 -2796 2202 -2790
rect 2196 -2802 2202 -2796
rect 2196 -2808 2202 -2802
rect 2196 -2814 2202 -2808
rect 2196 -2820 2202 -2814
rect 2196 -2826 2202 -2820
rect 2196 -2832 2202 -2826
rect 2196 -2838 2202 -2832
rect 2196 -2844 2202 -2838
rect 2196 -2850 2202 -2844
rect 2196 -2856 2202 -2850
rect 2196 -2862 2202 -2856
rect 2196 -2868 2202 -2862
rect 2196 -2874 2202 -2868
rect 2196 -2880 2202 -2874
rect 2196 -2886 2202 -2880
rect 2196 -2892 2202 -2886
rect 2196 -2898 2202 -2892
rect 2196 -2904 2202 -2898
rect 2196 -2910 2202 -2904
rect 2196 -2916 2202 -2910
rect 2196 -2922 2202 -2916
rect 2196 -2928 2202 -2922
rect 2196 -2934 2202 -2928
rect 2196 -2940 2202 -2934
rect 2196 -2946 2202 -2940
rect 2196 -2952 2202 -2946
rect 2196 -2958 2202 -2952
rect 2196 -2964 2202 -2958
rect 2196 -2970 2202 -2964
rect 2196 -2976 2202 -2970
rect 2196 -2982 2202 -2976
rect 2196 -2988 2202 -2982
rect 2196 -2994 2202 -2988
rect 2196 -3000 2202 -2994
rect 2196 -3006 2202 -3000
rect 2202 -198 2208 -192
rect 2202 -204 2208 -198
rect 2202 -210 2208 -204
rect 2202 -216 2208 -210
rect 2202 -222 2208 -216
rect 2202 -228 2208 -222
rect 2202 -234 2208 -228
rect 2202 -240 2208 -234
rect 2202 -246 2208 -240
rect 2202 -252 2208 -246
rect 2202 -258 2208 -252
rect 2202 -264 2208 -258
rect 2202 -270 2208 -264
rect 2202 -276 2208 -270
rect 2202 -282 2208 -276
rect 2202 -288 2208 -282
rect 2202 -294 2208 -288
rect 2202 -300 2208 -294
rect 2202 -306 2208 -300
rect 2202 -312 2208 -306
rect 2202 -318 2208 -312
rect 2202 -324 2208 -318
rect 2202 -330 2208 -324
rect 2202 -336 2208 -330
rect 2202 -342 2208 -336
rect 2202 -348 2208 -342
rect 2202 -354 2208 -348
rect 2202 -360 2208 -354
rect 2202 -366 2208 -360
rect 2202 -372 2208 -366
rect 2202 -378 2208 -372
rect 2202 -384 2208 -378
rect 2202 -390 2208 -384
rect 2202 -396 2208 -390
rect 2202 -402 2208 -396
rect 2202 -408 2208 -402
rect 2202 -414 2208 -408
rect 2202 -420 2208 -414
rect 2202 -426 2208 -420
rect 2202 -432 2208 -426
rect 2202 -438 2208 -432
rect 2202 -444 2208 -438
rect 2202 -450 2208 -444
rect 2202 -456 2208 -450
rect 2202 -462 2208 -456
rect 2202 -468 2208 -462
rect 2202 -474 2208 -468
rect 2202 -480 2208 -474
rect 2202 -486 2208 -480
rect 2202 -492 2208 -486
rect 2202 -498 2208 -492
rect 2202 -504 2208 -498
rect 2202 -510 2208 -504
rect 2202 -516 2208 -510
rect 2202 -522 2208 -516
rect 2202 -528 2208 -522
rect 2202 -534 2208 -528
rect 2202 -540 2208 -534
rect 2202 -546 2208 -540
rect 2202 -552 2208 -546
rect 2202 -558 2208 -552
rect 2202 -564 2208 -558
rect 2202 -570 2208 -564
rect 2202 -576 2208 -570
rect 2202 -582 2208 -576
rect 2202 -588 2208 -582
rect 2202 -594 2208 -588
rect 2202 -600 2208 -594
rect 2202 -606 2208 -600
rect 2202 -612 2208 -606
rect 2202 -618 2208 -612
rect 2202 -624 2208 -618
rect 2202 -630 2208 -624
rect 2202 -636 2208 -630
rect 2202 -642 2208 -636
rect 2202 -648 2208 -642
rect 2202 -654 2208 -648
rect 2202 -660 2208 -654
rect 2202 -666 2208 -660
rect 2202 -672 2208 -666
rect 2202 -678 2208 -672
rect 2202 -684 2208 -678
rect 2202 -690 2208 -684
rect 2202 -696 2208 -690
rect 2202 -702 2208 -696
rect 2202 -708 2208 -702
rect 2202 -714 2208 -708
rect 2202 -720 2208 -714
rect 2202 -726 2208 -720
rect 2202 -732 2208 -726
rect 2202 -738 2208 -732
rect 2202 -744 2208 -738
rect 2202 -750 2208 -744
rect 2202 -756 2208 -750
rect 2202 -762 2208 -756
rect 2202 -768 2208 -762
rect 2202 -774 2208 -768
rect 2202 -780 2208 -774
rect 2202 -786 2208 -780
rect 2202 -792 2208 -786
rect 2202 -798 2208 -792
rect 2202 -804 2208 -798
rect 2202 -810 2208 -804
rect 2202 -816 2208 -810
rect 2202 -822 2208 -816
rect 2202 -828 2208 -822
rect 2202 -834 2208 -828
rect 2202 -840 2208 -834
rect 2202 -846 2208 -840
rect 2202 -852 2208 -846
rect 2202 -858 2208 -852
rect 2202 -864 2208 -858
rect 2202 -870 2208 -864
rect 2202 -876 2208 -870
rect 2202 -882 2208 -876
rect 2202 -888 2208 -882
rect 2202 -894 2208 -888
rect 2202 -900 2208 -894
rect 2202 -906 2208 -900
rect 2202 -912 2208 -906
rect 2202 -918 2208 -912
rect 2202 -924 2208 -918
rect 2202 -930 2208 -924
rect 2202 -936 2208 -930
rect 2202 -942 2208 -936
rect 2202 -948 2208 -942
rect 2202 -954 2208 -948
rect 2202 -960 2208 -954
rect 2202 -966 2208 -960
rect 2202 -972 2208 -966
rect 2202 -978 2208 -972
rect 2202 -984 2208 -978
rect 2202 -990 2208 -984
rect 2202 -996 2208 -990
rect 2202 -1002 2208 -996
rect 2202 -1008 2208 -1002
rect 2202 -1014 2208 -1008
rect 2202 -1020 2208 -1014
rect 2202 -1026 2208 -1020
rect 2202 -1032 2208 -1026
rect 2202 -1038 2208 -1032
rect 2202 -1044 2208 -1038
rect 2202 -1050 2208 -1044
rect 2202 -1056 2208 -1050
rect 2202 -1062 2208 -1056
rect 2202 -1068 2208 -1062
rect 2202 -1074 2208 -1068
rect 2202 -1080 2208 -1074
rect 2202 -1086 2208 -1080
rect 2202 -1092 2208 -1086
rect 2202 -1098 2208 -1092
rect 2202 -1104 2208 -1098
rect 2202 -1110 2208 -1104
rect 2202 -1116 2208 -1110
rect 2202 -1122 2208 -1116
rect 2202 -1128 2208 -1122
rect 2202 -1134 2208 -1128
rect 2202 -1140 2208 -1134
rect 2202 -1146 2208 -1140
rect 2202 -1152 2208 -1146
rect 2202 -1158 2208 -1152
rect 2202 -1164 2208 -1158
rect 2202 -1170 2208 -1164
rect 2202 -1176 2208 -1170
rect 2202 -1182 2208 -1176
rect 2202 -1188 2208 -1182
rect 2202 -1194 2208 -1188
rect 2202 -1200 2208 -1194
rect 2202 -1206 2208 -1200
rect 2202 -1212 2208 -1206
rect 2202 -1218 2208 -1212
rect 2202 -1224 2208 -1218
rect 2202 -1230 2208 -1224
rect 2202 -1236 2208 -1230
rect 2202 -1242 2208 -1236
rect 2202 -1548 2208 -1542
rect 2202 -1554 2208 -1548
rect 2202 -1560 2208 -1554
rect 2202 -1566 2208 -1560
rect 2202 -1572 2208 -1566
rect 2202 -1578 2208 -1572
rect 2202 -1584 2208 -1578
rect 2202 -1590 2208 -1584
rect 2202 -1596 2208 -1590
rect 2202 -1602 2208 -1596
rect 2202 -1608 2208 -1602
rect 2202 -1614 2208 -1608
rect 2202 -1620 2208 -1614
rect 2202 -1626 2208 -1620
rect 2202 -1632 2208 -1626
rect 2202 -1638 2208 -1632
rect 2202 -1644 2208 -1638
rect 2202 -1650 2208 -1644
rect 2202 -1656 2208 -1650
rect 2202 -1662 2208 -1656
rect 2202 -1668 2208 -1662
rect 2202 -1674 2208 -1668
rect 2202 -1680 2208 -1674
rect 2202 -1686 2208 -1680
rect 2202 -1692 2208 -1686
rect 2202 -1698 2208 -1692
rect 2202 -1704 2208 -1698
rect 2202 -1710 2208 -1704
rect 2202 -1716 2208 -1710
rect 2202 -1722 2208 -1716
rect 2202 -1728 2208 -1722
rect 2202 -1734 2208 -1728
rect 2202 -1740 2208 -1734
rect 2202 -1746 2208 -1740
rect 2202 -1752 2208 -1746
rect 2202 -1758 2208 -1752
rect 2202 -1764 2208 -1758
rect 2202 -1770 2208 -1764
rect 2202 -1776 2208 -1770
rect 2202 -1782 2208 -1776
rect 2202 -1788 2208 -1782
rect 2202 -1794 2208 -1788
rect 2202 -1800 2208 -1794
rect 2202 -1806 2208 -1800
rect 2202 -1812 2208 -1806
rect 2202 -1818 2208 -1812
rect 2202 -1824 2208 -1818
rect 2202 -1830 2208 -1824
rect 2202 -1836 2208 -1830
rect 2202 -1842 2208 -1836
rect 2202 -1848 2208 -1842
rect 2202 -1854 2208 -1848
rect 2202 -1860 2208 -1854
rect 2202 -1866 2208 -1860
rect 2202 -1872 2208 -1866
rect 2202 -1878 2208 -1872
rect 2202 -1884 2208 -1878
rect 2202 -1890 2208 -1884
rect 2202 -1896 2208 -1890
rect 2202 -1902 2208 -1896
rect 2202 -1908 2208 -1902
rect 2202 -1914 2208 -1908
rect 2202 -1920 2208 -1914
rect 2202 -1926 2208 -1920
rect 2202 -1932 2208 -1926
rect 2202 -1938 2208 -1932
rect 2202 -1944 2208 -1938
rect 2202 -1950 2208 -1944
rect 2202 -1956 2208 -1950
rect 2202 -1962 2208 -1956
rect 2202 -1968 2208 -1962
rect 2202 -1974 2208 -1968
rect 2202 -1980 2208 -1974
rect 2202 -1986 2208 -1980
rect 2202 -1992 2208 -1986
rect 2202 -1998 2208 -1992
rect 2202 -2004 2208 -1998
rect 2202 -2010 2208 -2004
rect 2202 -2016 2208 -2010
rect 2202 -2022 2208 -2016
rect 2202 -2028 2208 -2022
rect 2202 -2034 2208 -2028
rect 2202 -2040 2208 -2034
rect 2202 -2046 2208 -2040
rect 2202 -2052 2208 -2046
rect 2202 -2058 2208 -2052
rect 2202 -2064 2208 -2058
rect 2202 -2070 2208 -2064
rect 2202 -2076 2208 -2070
rect 2202 -2082 2208 -2076
rect 2202 -2088 2208 -2082
rect 2202 -2094 2208 -2088
rect 2202 -2100 2208 -2094
rect 2202 -2106 2208 -2100
rect 2202 -2112 2208 -2106
rect 2202 -2118 2208 -2112
rect 2202 -2124 2208 -2118
rect 2202 -2130 2208 -2124
rect 2202 -2136 2208 -2130
rect 2202 -2142 2208 -2136
rect 2202 -2148 2208 -2142
rect 2202 -2154 2208 -2148
rect 2202 -2160 2208 -2154
rect 2202 -2166 2208 -2160
rect 2202 -2172 2208 -2166
rect 2202 -2178 2208 -2172
rect 2202 -2184 2208 -2178
rect 2202 -2190 2208 -2184
rect 2202 -2196 2208 -2190
rect 2202 -2202 2208 -2196
rect 2202 -2208 2208 -2202
rect 2202 -2214 2208 -2208
rect 2202 -2220 2208 -2214
rect 2202 -2226 2208 -2220
rect 2202 -2232 2208 -2226
rect 2202 -2238 2208 -2232
rect 2202 -2244 2208 -2238
rect 2202 -2250 2208 -2244
rect 2202 -2256 2208 -2250
rect 2202 -2262 2208 -2256
rect 2202 -2268 2208 -2262
rect 2202 -2274 2208 -2268
rect 2202 -2280 2208 -2274
rect 2202 -2286 2208 -2280
rect 2202 -2292 2208 -2286
rect 2202 -2298 2208 -2292
rect 2202 -2304 2208 -2298
rect 2202 -2310 2208 -2304
rect 2202 -2316 2208 -2310
rect 2202 -2322 2208 -2316
rect 2202 -2328 2208 -2322
rect 2202 -2334 2208 -2328
rect 2202 -2340 2208 -2334
rect 2202 -2478 2208 -2472
rect 2202 -2538 2208 -2532
rect 2202 -2544 2208 -2538
rect 2202 -2550 2208 -2544
rect 2202 -2556 2208 -2550
rect 2202 -2562 2208 -2556
rect 2202 -2568 2208 -2562
rect 2202 -2574 2208 -2568
rect 2202 -2580 2208 -2574
rect 2202 -2586 2208 -2580
rect 2202 -2592 2208 -2586
rect 2202 -2598 2208 -2592
rect 2202 -2604 2208 -2598
rect 2202 -2610 2208 -2604
rect 2202 -2616 2208 -2610
rect 2202 -2622 2208 -2616
rect 2202 -2628 2208 -2622
rect 2202 -2634 2208 -2628
rect 2202 -2640 2208 -2634
rect 2202 -2646 2208 -2640
rect 2202 -2652 2208 -2646
rect 2202 -2658 2208 -2652
rect 2202 -2664 2208 -2658
rect 2202 -2670 2208 -2664
rect 2202 -2676 2208 -2670
rect 2202 -2682 2208 -2676
rect 2202 -2688 2208 -2682
rect 2202 -2694 2208 -2688
rect 2202 -2700 2208 -2694
rect 2202 -2706 2208 -2700
rect 2202 -2712 2208 -2706
rect 2202 -2718 2208 -2712
rect 2202 -2724 2208 -2718
rect 2202 -2730 2208 -2724
rect 2202 -2736 2208 -2730
rect 2202 -2742 2208 -2736
rect 2202 -2748 2208 -2742
rect 2202 -2754 2208 -2748
rect 2202 -2760 2208 -2754
rect 2202 -2766 2208 -2760
rect 2202 -2772 2208 -2766
rect 2202 -2778 2208 -2772
rect 2202 -2784 2208 -2778
rect 2202 -2790 2208 -2784
rect 2202 -2796 2208 -2790
rect 2202 -2802 2208 -2796
rect 2202 -2808 2208 -2802
rect 2202 -2814 2208 -2808
rect 2202 -2820 2208 -2814
rect 2202 -2826 2208 -2820
rect 2202 -2832 2208 -2826
rect 2202 -2838 2208 -2832
rect 2202 -2844 2208 -2838
rect 2202 -2850 2208 -2844
rect 2202 -2856 2208 -2850
rect 2202 -2862 2208 -2856
rect 2202 -2868 2208 -2862
rect 2202 -2874 2208 -2868
rect 2202 -2880 2208 -2874
rect 2202 -2886 2208 -2880
rect 2202 -2892 2208 -2886
rect 2202 -2898 2208 -2892
rect 2202 -2904 2208 -2898
rect 2202 -2910 2208 -2904
rect 2202 -2916 2208 -2910
rect 2202 -2922 2208 -2916
rect 2202 -2928 2208 -2922
rect 2202 -2934 2208 -2928
rect 2202 -2940 2208 -2934
rect 2202 -2946 2208 -2940
rect 2202 -2952 2208 -2946
rect 2202 -2958 2208 -2952
rect 2202 -2964 2208 -2958
rect 2202 -2970 2208 -2964
rect 2202 -2976 2208 -2970
rect 2202 -2982 2208 -2976
rect 2202 -2988 2208 -2982
rect 2202 -2994 2208 -2988
rect 2202 -3000 2208 -2994
rect 2202 -3006 2208 -3000
rect 2208 -186 2214 -180
rect 2208 -192 2214 -186
rect 2208 -198 2214 -192
rect 2208 -204 2214 -198
rect 2208 -210 2214 -204
rect 2208 -216 2214 -210
rect 2208 -222 2214 -216
rect 2208 -228 2214 -222
rect 2208 -234 2214 -228
rect 2208 -240 2214 -234
rect 2208 -246 2214 -240
rect 2208 -252 2214 -246
rect 2208 -258 2214 -252
rect 2208 -264 2214 -258
rect 2208 -270 2214 -264
rect 2208 -276 2214 -270
rect 2208 -282 2214 -276
rect 2208 -288 2214 -282
rect 2208 -294 2214 -288
rect 2208 -300 2214 -294
rect 2208 -306 2214 -300
rect 2208 -312 2214 -306
rect 2208 -318 2214 -312
rect 2208 -324 2214 -318
rect 2208 -330 2214 -324
rect 2208 -336 2214 -330
rect 2208 -342 2214 -336
rect 2208 -348 2214 -342
rect 2208 -354 2214 -348
rect 2208 -360 2214 -354
rect 2208 -366 2214 -360
rect 2208 -372 2214 -366
rect 2208 -378 2214 -372
rect 2208 -384 2214 -378
rect 2208 -390 2214 -384
rect 2208 -396 2214 -390
rect 2208 -402 2214 -396
rect 2208 -408 2214 -402
rect 2208 -414 2214 -408
rect 2208 -420 2214 -414
rect 2208 -426 2214 -420
rect 2208 -432 2214 -426
rect 2208 -438 2214 -432
rect 2208 -444 2214 -438
rect 2208 -450 2214 -444
rect 2208 -456 2214 -450
rect 2208 -462 2214 -456
rect 2208 -468 2214 -462
rect 2208 -474 2214 -468
rect 2208 -480 2214 -474
rect 2208 -486 2214 -480
rect 2208 -492 2214 -486
rect 2208 -498 2214 -492
rect 2208 -504 2214 -498
rect 2208 -510 2214 -504
rect 2208 -516 2214 -510
rect 2208 -522 2214 -516
rect 2208 -528 2214 -522
rect 2208 -534 2214 -528
rect 2208 -540 2214 -534
rect 2208 -546 2214 -540
rect 2208 -552 2214 -546
rect 2208 -558 2214 -552
rect 2208 -564 2214 -558
rect 2208 -570 2214 -564
rect 2208 -576 2214 -570
rect 2208 -582 2214 -576
rect 2208 -588 2214 -582
rect 2208 -594 2214 -588
rect 2208 -600 2214 -594
rect 2208 -606 2214 -600
rect 2208 -612 2214 -606
rect 2208 -618 2214 -612
rect 2208 -624 2214 -618
rect 2208 -630 2214 -624
rect 2208 -636 2214 -630
rect 2208 -642 2214 -636
rect 2208 -648 2214 -642
rect 2208 -654 2214 -648
rect 2208 -660 2214 -654
rect 2208 -666 2214 -660
rect 2208 -672 2214 -666
rect 2208 -678 2214 -672
rect 2208 -684 2214 -678
rect 2208 -690 2214 -684
rect 2208 -696 2214 -690
rect 2208 -702 2214 -696
rect 2208 -708 2214 -702
rect 2208 -714 2214 -708
rect 2208 -720 2214 -714
rect 2208 -726 2214 -720
rect 2208 -732 2214 -726
rect 2208 -738 2214 -732
rect 2208 -744 2214 -738
rect 2208 -750 2214 -744
rect 2208 -756 2214 -750
rect 2208 -762 2214 -756
rect 2208 -768 2214 -762
rect 2208 -774 2214 -768
rect 2208 -780 2214 -774
rect 2208 -786 2214 -780
rect 2208 -792 2214 -786
rect 2208 -798 2214 -792
rect 2208 -804 2214 -798
rect 2208 -810 2214 -804
rect 2208 -816 2214 -810
rect 2208 -822 2214 -816
rect 2208 -828 2214 -822
rect 2208 -834 2214 -828
rect 2208 -840 2214 -834
rect 2208 -846 2214 -840
rect 2208 -852 2214 -846
rect 2208 -858 2214 -852
rect 2208 -864 2214 -858
rect 2208 -870 2214 -864
rect 2208 -876 2214 -870
rect 2208 -882 2214 -876
rect 2208 -888 2214 -882
rect 2208 -894 2214 -888
rect 2208 -900 2214 -894
rect 2208 -906 2214 -900
rect 2208 -912 2214 -906
rect 2208 -918 2214 -912
rect 2208 -924 2214 -918
rect 2208 -930 2214 -924
rect 2208 -936 2214 -930
rect 2208 -942 2214 -936
rect 2208 -948 2214 -942
rect 2208 -954 2214 -948
rect 2208 -960 2214 -954
rect 2208 -966 2214 -960
rect 2208 -972 2214 -966
rect 2208 -978 2214 -972
rect 2208 -984 2214 -978
rect 2208 -990 2214 -984
rect 2208 -996 2214 -990
rect 2208 -1002 2214 -996
rect 2208 -1008 2214 -1002
rect 2208 -1014 2214 -1008
rect 2208 -1020 2214 -1014
rect 2208 -1026 2214 -1020
rect 2208 -1032 2214 -1026
rect 2208 -1038 2214 -1032
rect 2208 -1044 2214 -1038
rect 2208 -1050 2214 -1044
rect 2208 -1056 2214 -1050
rect 2208 -1062 2214 -1056
rect 2208 -1068 2214 -1062
rect 2208 -1074 2214 -1068
rect 2208 -1080 2214 -1074
rect 2208 -1086 2214 -1080
rect 2208 -1092 2214 -1086
rect 2208 -1098 2214 -1092
rect 2208 -1104 2214 -1098
rect 2208 -1110 2214 -1104
rect 2208 -1116 2214 -1110
rect 2208 -1122 2214 -1116
rect 2208 -1128 2214 -1122
rect 2208 -1134 2214 -1128
rect 2208 -1140 2214 -1134
rect 2208 -1146 2214 -1140
rect 2208 -1152 2214 -1146
rect 2208 -1158 2214 -1152
rect 2208 -1164 2214 -1158
rect 2208 -1170 2214 -1164
rect 2208 -1176 2214 -1170
rect 2208 -1182 2214 -1176
rect 2208 -1188 2214 -1182
rect 2208 -1194 2214 -1188
rect 2208 -1200 2214 -1194
rect 2208 -1206 2214 -1200
rect 2208 -1212 2214 -1206
rect 2208 -1218 2214 -1212
rect 2208 -1224 2214 -1218
rect 2208 -1548 2214 -1542
rect 2208 -1554 2214 -1548
rect 2208 -1560 2214 -1554
rect 2208 -1566 2214 -1560
rect 2208 -1572 2214 -1566
rect 2208 -1578 2214 -1572
rect 2208 -1584 2214 -1578
rect 2208 -1590 2214 -1584
rect 2208 -1596 2214 -1590
rect 2208 -1602 2214 -1596
rect 2208 -1608 2214 -1602
rect 2208 -1614 2214 -1608
rect 2208 -1620 2214 -1614
rect 2208 -1626 2214 -1620
rect 2208 -1632 2214 -1626
rect 2208 -1638 2214 -1632
rect 2208 -1644 2214 -1638
rect 2208 -1650 2214 -1644
rect 2208 -1656 2214 -1650
rect 2208 -1662 2214 -1656
rect 2208 -1668 2214 -1662
rect 2208 -1674 2214 -1668
rect 2208 -1680 2214 -1674
rect 2208 -1686 2214 -1680
rect 2208 -1692 2214 -1686
rect 2208 -1698 2214 -1692
rect 2208 -1704 2214 -1698
rect 2208 -1710 2214 -1704
rect 2208 -1716 2214 -1710
rect 2208 -1722 2214 -1716
rect 2208 -1728 2214 -1722
rect 2208 -1734 2214 -1728
rect 2208 -1740 2214 -1734
rect 2208 -1746 2214 -1740
rect 2208 -1752 2214 -1746
rect 2208 -1758 2214 -1752
rect 2208 -1764 2214 -1758
rect 2208 -1770 2214 -1764
rect 2208 -1776 2214 -1770
rect 2208 -1782 2214 -1776
rect 2208 -1788 2214 -1782
rect 2208 -1794 2214 -1788
rect 2208 -1800 2214 -1794
rect 2208 -1806 2214 -1800
rect 2208 -1812 2214 -1806
rect 2208 -1818 2214 -1812
rect 2208 -1824 2214 -1818
rect 2208 -1830 2214 -1824
rect 2208 -1836 2214 -1830
rect 2208 -1842 2214 -1836
rect 2208 -1848 2214 -1842
rect 2208 -1854 2214 -1848
rect 2208 -1860 2214 -1854
rect 2208 -1866 2214 -1860
rect 2208 -1872 2214 -1866
rect 2208 -1878 2214 -1872
rect 2208 -1884 2214 -1878
rect 2208 -1890 2214 -1884
rect 2208 -1896 2214 -1890
rect 2208 -1902 2214 -1896
rect 2208 -1908 2214 -1902
rect 2208 -1914 2214 -1908
rect 2208 -1920 2214 -1914
rect 2208 -1926 2214 -1920
rect 2208 -1932 2214 -1926
rect 2208 -1938 2214 -1932
rect 2208 -1944 2214 -1938
rect 2208 -1950 2214 -1944
rect 2208 -1956 2214 -1950
rect 2208 -1962 2214 -1956
rect 2208 -1968 2214 -1962
rect 2208 -1974 2214 -1968
rect 2208 -1980 2214 -1974
rect 2208 -1986 2214 -1980
rect 2208 -1992 2214 -1986
rect 2208 -1998 2214 -1992
rect 2208 -2004 2214 -1998
rect 2208 -2010 2214 -2004
rect 2208 -2016 2214 -2010
rect 2208 -2022 2214 -2016
rect 2208 -2028 2214 -2022
rect 2208 -2034 2214 -2028
rect 2208 -2040 2214 -2034
rect 2208 -2046 2214 -2040
rect 2208 -2052 2214 -2046
rect 2208 -2058 2214 -2052
rect 2208 -2064 2214 -2058
rect 2208 -2070 2214 -2064
rect 2208 -2076 2214 -2070
rect 2208 -2082 2214 -2076
rect 2208 -2088 2214 -2082
rect 2208 -2094 2214 -2088
rect 2208 -2100 2214 -2094
rect 2208 -2106 2214 -2100
rect 2208 -2112 2214 -2106
rect 2208 -2118 2214 -2112
rect 2208 -2124 2214 -2118
rect 2208 -2130 2214 -2124
rect 2208 -2136 2214 -2130
rect 2208 -2142 2214 -2136
rect 2208 -2148 2214 -2142
rect 2208 -2154 2214 -2148
rect 2208 -2160 2214 -2154
rect 2208 -2166 2214 -2160
rect 2208 -2172 2214 -2166
rect 2208 -2178 2214 -2172
rect 2208 -2184 2214 -2178
rect 2208 -2190 2214 -2184
rect 2208 -2196 2214 -2190
rect 2208 -2202 2214 -2196
rect 2208 -2208 2214 -2202
rect 2208 -2214 2214 -2208
rect 2208 -2220 2214 -2214
rect 2208 -2226 2214 -2220
rect 2208 -2232 2214 -2226
rect 2208 -2238 2214 -2232
rect 2208 -2244 2214 -2238
rect 2208 -2250 2214 -2244
rect 2208 -2256 2214 -2250
rect 2208 -2262 2214 -2256
rect 2208 -2268 2214 -2262
rect 2208 -2274 2214 -2268
rect 2208 -2280 2214 -2274
rect 2208 -2286 2214 -2280
rect 2208 -2292 2214 -2286
rect 2208 -2298 2214 -2292
rect 2208 -2304 2214 -2298
rect 2208 -2310 2214 -2304
rect 2208 -2316 2214 -2310
rect 2208 -2322 2214 -2316
rect 2208 -2328 2214 -2322
rect 2208 -2334 2214 -2328
rect 2208 -2400 2214 -2394
rect 2208 -2406 2214 -2400
rect 2208 -2412 2214 -2406
rect 2208 -2418 2214 -2412
rect 2208 -2424 2214 -2418
rect 2208 -2430 2214 -2424
rect 2208 -2436 2214 -2430
rect 2208 -2442 2214 -2436
rect 2208 -2448 2214 -2442
rect 2208 -2454 2214 -2448
rect 2208 -2460 2214 -2454
rect 2208 -2466 2214 -2460
rect 2208 -2472 2214 -2466
rect 2208 -2478 2214 -2472
rect 2208 -2538 2214 -2532
rect 2208 -2544 2214 -2538
rect 2208 -2550 2214 -2544
rect 2208 -2556 2214 -2550
rect 2208 -2562 2214 -2556
rect 2208 -2568 2214 -2562
rect 2208 -2574 2214 -2568
rect 2208 -2580 2214 -2574
rect 2208 -2586 2214 -2580
rect 2208 -2592 2214 -2586
rect 2208 -2598 2214 -2592
rect 2208 -2604 2214 -2598
rect 2208 -2610 2214 -2604
rect 2208 -2616 2214 -2610
rect 2208 -2622 2214 -2616
rect 2208 -2628 2214 -2622
rect 2208 -2634 2214 -2628
rect 2208 -2640 2214 -2634
rect 2208 -2646 2214 -2640
rect 2208 -2652 2214 -2646
rect 2208 -2658 2214 -2652
rect 2208 -2664 2214 -2658
rect 2208 -2670 2214 -2664
rect 2208 -2676 2214 -2670
rect 2208 -2682 2214 -2676
rect 2208 -2688 2214 -2682
rect 2208 -2694 2214 -2688
rect 2208 -2700 2214 -2694
rect 2208 -2706 2214 -2700
rect 2208 -2712 2214 -2706
rect 2208 -2718 2214 -2712
rect 2208 -2724 2214 -2718
rect 2208 -2730 2214 -2724
rect 2208 -2736 2214 -2730
rect 2208 -2742 2214 -2736
rect 2208 -2748 2214 -2742
rect 2208 -2754 2214 -2748
rect 2208 -2760 2214 -2754
rect 2208 -2766 2214 -2760
rect 2208 -2772 2214 -2766
rect 2208 -2778 2214 -2772
rect 2208 -2784 2214 -2778
rect 2208 -2790 2214 -2784
rect 2208 -2796 2214 -2790
rect 2208 -2802 2214 -2796
rect 2208 -2808 2214 -2802
rect 2208 -2814 2214 -2808
rect 2208 -2820 2214 -2814
rect 2208 -2826 2214 -2820
rect 2208 -2832 2214 -2826
rect 2208 -2838 2214 -2832
rect 2208 -2844 2214 -2838
rect 2208 -2850 2214 -2844
rect 2208 -2856 2214 -2850
rect 2208 -2862 2214 -2856
rect 2208 -2868 2214 -2862
rect 2208 -2874 2214 -2868
rect 2208 -2880 2214 -2874
rect 2208 -2886 2214 -2880
rect 2208 -2892 2214 -2886
rect 2208 -2898 2214 -2892
rect 2208 -2904 2214 -2898
rect 2208 -2910 2214 -2904
rect 2208 -2916 2214 -2910
rect 2208 -2922 2214 -2916
rect 2208 -2928 2214 -2922
rect 2208 -2934 2214 -2928
rect 2208 -2940 2214 -2934
rect 2208 -2946 2214 -2940
rect 2208 -2952 2214 -2946
rect 2208 -2958 2214 -2952
rect 2208 -2964 2214 -2958
rect 2208 -2970 2214 -2964
rect 2208 -2976 2214 -2970
rect 2208 -2982 2214 -2976
rect 2208 -2988 2214 -2982
rect 2208 -2994 2214 -2988
rect 2208 -3000 2214 -2994
rect 2214 -180 2220 -174
rect 2214 -186 2220 -180
rect 2214 -192 2220 -186
rect 2214 -198 2220 -192
rect 2214 -204 2220 -198
rect 2214 -210 2220 -204
rect 2214 -216 2220 -210
rect 2214 -222 2220 -216
rect 2214 -228 2220 -222
rect 2214 -234 2220 -228
rect 2214 -240 2220 -234
rect 2214 -246 2220 -240
rect 2214 -252 2220 -246
rect 2214 -258 2220 -252
rect 2214 -264 2220 -258
rect 2214 -270 2220 -264
rect 2214 -276 2220 -270
rect 2214 -282 2220 -276
rect 2214 -288 2220 -282
rect 2214 -294 2220 -288
rect 2214 -300 2220 -294
rect 2214 -306 2220 -300
rect 2214 -312 2220 -306
rect 2214 -318 2220 -312
rect 2214 -324 2220 -318
rect 2214 -330 2220 -324
rect 2214 -336 2220 -330
rect 2214 -342 2220 -336
rect 2214 -348 2220 -342
rect 2214 -354 2220 -348
rect 2214 -360 2220 -354
rect 2214 -366 2220 -360
rect 2214 -372 2220 -366
rect 2214 -378 2220 -372
rect 2214 -384 2220 -378
rect 2214 -390 2220 -384
rect 2214 -396 2220 -390
rect 2214 -402 2220 -396
rect 2214 -408 2220 -402
rect 2214 -414 2220 -408
rect 2214 -420 2220 -414
rect 2214 -426 2220 -420
rect 2214 -432 2220 -426
rect 2214 -438 2220 -432
rect 2214 -444 2220 -438
rect 2214 -450 2220 -444
rect 2214 -456 2220 -450
rect 2214 -462 2220 -456
rect 2214 -468 2220 -462
rect 2214 -474 2220 -468
rect 2214 -480 2220 -474
rect 2214 -486 2220 -480
rect 2214 -492 2220 -486
rect 2214 -498 2220 -492
rect 2214 -504 2220 -498
rect 2214 -510 2220 -504
rect 2214 -516 2220 -510
rect 2214 -522 2220 -516
rect 2214 -528 2220 -522
rect 2214 -534 2220 -528
rect 2214 -540 2220 -534
rect 2214 -546 2220 -540
rect 2214 -552 2220 -546
rect 2214 -558 2220 -552
rect 2214 -564 2220 -558
rect 2214 -570 2220 -564
rect 2214 -576 2220 -570
rect 2214 -582 2220 -576
rect 2214 -588 2220 -582
rect 2214 -594 2220 -588
rect 2214 -600 2220 -594
rect 2214 -606 2220 -600
rect 2214 -612 2220 -606
rect 2214 -618 2220 -612
rect 2214 -624 2220 -618
rect 2214 -630 2220 -624
rect 2214 -636 2220 -630
rect 2214 -642 2220 -636
rect 2214 -648 2220 -642
rect 2214 -654 2220 -648
rect 2214 -660 2220 -654
rect 2214 -666 2220 -660
rect 2214 -672 2220 -666
rect 2214 -678 2220 -672
rect 2214 -684 2220 -678
rect 2214 -690 2220 -684
rect 2214 -696 2220 -690
rect 2214 -702 2220 -696
rect 2214 -708 2220 -702
rect 2214 -714 2220 -708
rect 2214 -720 2220 -714
rect 2214 -726 2220 -720
rect 2214 -732 2220 -726
rect 2214 -738 2220 -732
rect 2214 -744 2220 -738
rect 2214 -750 2220 -744
rect 2214 -756 2220 -750
rect 2214 -762 2220 -756
rect 2214 -768 2220 -762
rect 2214 -774 2220 -768
rect 2214 -780 2220 -774
rect 2214 -786 2220 -780
rect 2214 -792 2220 -786
rect 2214 -798 2220 -792
rect 2214 -804 2220 -798
rect 2214 -810 2220 -804
rect 2214 -816 2220 -810
rect 2214 -822 2220 -816
rect 2214 -828 2220 -822
rect 2214 -834 2220 -828
rect 2214 -840 2220 -834
rect 2214 -846 2220 -840
rect 2214 -852 2220 -846
rect 2214 -858 2220 -852
rect 2214 -864 2220 -858
rect 2214 -870 2220 -864
rect 2214 -876 2220 -870
rect 2214 -882 2220 -876
rect 2214 -888 2220 -882
rect 2214 -894 2220 -888
rect 2214 -900 2220 -894
rect 2214 -906 2220 -900
rect 2214 -912 2220 -906
rect 2214 -918 2220 -912
rect 2214 -924 2220 -918
rect 2214 -930 2220 -924
rect 2214 -936 2220 -930
rect 2214 -942 2220 -936
rect 2214 -948 2220 -942
rect 2214 -954 2220 -948
rect 2214 -960 2220 -954
rect 2214 -966 2220 -960
rect 2214 -972 2220 -966
rect 2214 -978 2220 -972
rect 2214 -984 2220 -978
rect 2214 -990 2220 -984
rect 2214 -996 2220 -990
rect 2214 -1002 2220 -996
rect 2214 -1008 2220 -1002
rect 2214 -1014 2220 -1008
rect 2214 -1020 2220 -1014
rect 2214 -1026 2220 -1020
rect 2214 -1032 2220 -1026
rect 2214 -1038 2220 -1032
rect 2214 -1044 2220 -1038
rect 2214 -1050 2220 -1044
rect 2214 -1056 2220 -1050
rect 2214 -1062 2220 -1056
rect 2214 -1068 2220 -1062
rect 2214 -1074 2220 -1068
rect 2214 -1080 2220 -1074
rect 2214 -1086 2220 -1080
rect 2214 -1092 2220 -1086
rect 2214 -1098 2220 -1092
rect 2214 -1104 2220 -1098
rect 2214 -1110 2220 -1104
rect 2214 -1116 2220 -1110
rect 2214 -1122 2220 -1116
rect 2214 -1128 2220 -1122
rect 2214 -1134 2220 -1128
rect 2214 -1140 2220 -1134
rect 2214 -1146 2220 -1140
rect 2214 -1152 2220 -1146
rect 2214 -1158 2220 -1152
rect 2214 -1164 2220 -1158
rect 2214 -1170 2220 -1164
rect 2214 -1176 2220 -1170
rect 2214 -1182 2220 -1176
rect 2214 -1188 2220 -1182
rect 2214 -1194 2220 -1188
rect 2214 -1200 2220 -1194
rect 2214 -1206 2220 -1200
rect 2214 -1212 2220 -1206
rect 2214 -1542 2220 -1536
rect 2214 -1548 2220 -1542
rect 2214 -1554 2220 -1548
rect 2214 -1560 2220 -1554
rect 2214 -1566 2220 -1560
rect 2214 -1572 2220 -1566
rect 2214 -1578 2220 -1572
rect 2214 -1584 2220 -1578
rect 2214 -1590 2220 -1584
rect 2214 -1596 2220 -1590
rect 2214 -1602 2220 -1596
rect 2214 -1608 2220 -1602
rect 2214 -1614 2220 -1608
rect 2214 -1620 2220 -1614
rect 2214 -1626 2220 -1620
rect 2214 -1632 2220 -1626
rect 2214 -1638 2220 -1632
rect 2214 -1644 2220 -1638
rect 2214 -1650 2220 -1644
rect 2214 -1656 2220 -1650
rect 2214 -1662 2220 -1656
rect 2214 -1668 2220 -1662
rect 2214 -1674 2220 -1668
rect 2214 -1680 2220 -1674
rect 2214 -1686 2220 -1680
rect 2214 -1692 2220 -1686
rect 2214 -1698 2220 -1692
rect 2214 -1704 2220 -1698
rect 2214 -1710 2220 -1704
rect 2214 -1716 2220 -1710
rect 2214 -1722 2220 -1716
rect 2214 -1728 2220 -1722
rect 2214 -1734 2220 -1728
rect 2214 -1740 2220 -1734
rect 2214 -1746 2220 -1740
rect 2214 -1752 2220 -1746
rect 2214 -1758 2220 -1752
rect 2214 -1764 2220 -1758
rect 2214 -1770 2220 -1764
rect 2214 -1776 2220 -1770
rect 2214 -1782 2220 -1776
rect 2214 -1788 2220 -1782
rect 2214 -1794 2220 -1788
rect 2214 -1800 2220 -1794
rect 2214 -1806 2220 -1800
rect 2214 -1812 2220 -1806
rect 2214 -1818 2220 -1812
rect 2214 -1824 2220 -1818
rect 2214 -1830 2220 -1824
rect 2214 -1836 2220 -1830
rect 2214 -1842 2220 -1836
rect 2214 -1848 2220 -1842
rect 2214 -1854 2220 -1848
rect 2214 -1860 2220 -1854
rect 2214 -1866 2220 -1860
rect 2214 -1872 2220 -1866
rect 2214 -1878 2220 -1872
rect 2214 -1884 2220 -1878
rect 2214 -1890 2220 -1884
rect 2214 -1896 2220 -1890
rect 2214 -1902 2220 -1896
rect 2214 -1908 2220 -1902
rect 2214 -1914 2220 -1908
rect 2214 -1920 2220 -1914
rect 2214 -1926 2220 -1920
rect 2214 -1932 2220 -1926
rect 2214 -1938 2220 -1932
rect 2214 -1944 2220 -1938
rect 2214 -1950 2220 -1944
rect 2214 -1956 2220 -1950
rect 2214 -1962 2220 -1956
rect 2214 -1968 2220 -1962
rect 2214 -1974 2220 -1968
rect 2214 -1980 2220 -1974
rect 2214 -1986 2220 -1980
rect 2214 -1992 2220 -1986
rect 2214 -1998 2220 -1992
rect 2214 -2004 2220 -1998
rect 2214 -2010 2220 -2004
rect 2214 -2016 2220 -2010
rect 2214 -2022 2220 -2016
rect 2214 -2028 2220 -2022
rect 2214 -2034 2220 -2028
rect 2214 -2040 2220 -2034
rect 2214 -2046 2220 -2040
rect 2214 -2052 2220 -2046
rect 2214 -2058 2220 -2052
rect 2214 -2064 2220 -2058
rect 2214 -2070 2220 -2064
rect 2214 -2076 2220 -2070
rect 2214 -2082 2220 -2076
rect 2214 -2088 2220 -2082
rect 2214 -2094 2220 -2088
rect 2214 -2100 2220 -2094
rect 2214 -2106 2220 -2100
rect 2214 -2112 2220 -2106
rect 2214 -2118 2220 -2112
rect 2214 -2124 2220 -2118
rect 2214 -2130 2220 -2124
rect 2214 -2136 2220 -2130
rect 2214 -2142 2220 -2136
rect 2214 -2148 2220 -2142
rect 2214 -2154 2220 -2148
rect 2214 -2160 2220 -2154
rect 2214 -2166 2220 -2160
rect 2214 -2172 2220 -2166
rect 2214 -2178 2220 -2172
rect 2214 -2184 2220 -2178
rect 2214 -2190 2220 -2184
rect 2214 -2196 2220 -2190
rect 2214 -2202 2220 -2196
rect 2214 -2208 2220 -2202
rect 2214 -2214 2220 -2208
rect 2214 -2220 2220 -2214
rect 2214 -2226 2220 -2220
rect 2214 -2232 2220 -2226
rect 2214 -2238 2220 -2232
rect 2214 -2244 2220 -2238
rect 2214 -2250 2220 -2244
rect 2214 -2256 2220 -2250
rect 2214 -2262 2220 -2256
rect 2214 -2268 2220 -2262
rect 2214 -2274 2220 -2268
rect 2214 -2280 2220 -2274
rect 2214 -2286 2220 -2280
rect 2214 -2292 2220 -2286
rect 2214 -2298 2220 -2292
rect 2214 -2304 2220 -2298
rect 2214 -2310 2220 -2304
rect 2214 -2316 2220 -2310
rect 2214 -2322 2220 -2316
rect 2214 -2328 2220 -2322
rect 2214 -2394 2220 -2388
rect 2214 -2400 2220 -2394
rect 2214 -2406 2220 -2400
rect 2214 -2412 2220 -2406
rect 2214 -2418 2220 -2412
rect 2214 -2424 2220 -2418
rect 2214 -2430 2220 -2424
rect 2214 -2436 2220 -2430
rect 2214 -2442 2220 -2436
rect 2214 -2448 2220 -2442
rect 2214 -2454 2220 -2448
rect 2214 -2460 2220 -2454
rect 2214 -2466 2220 -2460
rect 2214 -2472 2220 -2466
rect 2214 -2532 2220 -2526
rect 2214 -2538 2220 -2532
rect 2214 -2544 2220 -2538
rect 2214 -2550 2220 -2544
rect 2214 -2556 2220 -2550
rect 2214 -2562 2220 -2556
rect 2214 -2568 2220 -2562
rect 2214 -2574 2220 -2568
rect 2214 -2580 2220 -2574
rect 2214 -2586 2220 -2580
rect 2214 -2592 2220 -2586
rect 2214 -2598 2220 -2592
rect 2214 -2604 2220 -2598
rect 2214 -2610 2220 -2604
rect 2214 -2616 2220 -2610
rect 2214 -2622 2220 -2616
rect 2214 -2628 2220 -2622
rect 2214 -2634 2220 -2628
rect 2214 -2640 2220 -2634
rect 2214 -2646 2220 -2640
rect 2214 -2652 2220 -2646
rect 2214 -2658 2220 -2652
rect 2214 -2664 2220 -2658
rect 2214 -2670 2220 -2664
rect 2214 -2676 2220 -2670
rect 2214 -2682 2220 -2676
rect 2214 -2688 2220 -2682
rect 2214 -2694 2220 -2688
rect 2214 -2700 2220 -2694
rect 2214 -2706 2220 -2700
rect 2214 -2712 2220 -2706
rect 2214 -2718 2220 -2712
rect 2214 -2724 2220 -2718
rect 2214 -2730 2220 -2724
rect 2214 -2736 2220 -2730
rect 2214 -2742 2220 -2736
rect 2214 -2748 2220 -2742
rect 2214 -2754 2220 -2748
rect 2214 -2760 2220 -2754
rect 2214 -2766 2220 -2760
rect 2214 -2772 2220 -2766
rect 2214 -2778 2220 -2772
rect 2214 -2784 2220 -2778
rect 2214 -2790 2220 -2784
rect 2214 -2796 2220 -2790
rect 2214 -2802 2220 -2796
rect 2214 -2808 2220 -2802
rect 2214 -2814 2220 -2808
rect 2214 -2820 2220 -2814
rect 2214 -2826 2220 -2820
rect 2214 -2832 2220 -2826
rect 2214 -2838 2220 -2832
rect 2214 -2844 2220 -2838
rect 2214 -2850 2220 -2844
rect 2214 -2856 2220 -2850
rect 2214 -2862 2220 -2856
rect 2214 -2868 2220 -2862
rect 2214 -2874 2220 -2868
rect 2214 -2880 2220 -2874
rect 2214 -2886 2220 -2880
rect 2214 -2892 2220 -2886
rect 2214 -2898 2220 -2892
rect 2214 -2904 2220 -2898
rect 2214 -2910 2220 -2904
rect 2214 -2916 2220 -2910
rect 2214 -2922 2220 -2916
rect 2214 -2928 2220 -2922
rect 2214 -2934 2220 -2928
rect 2214 -2940 2220 -2934
rect 2214 -2946 2220 -2940
rect 2214 -2952 2220 -2946
rect 2214 -2958 2220 -2952
rect 2214 -2964 2220 -2958
rect 2214 -2970 2220 -2964
rect 2214 -2976 2220 -2970
rect 2214 -2982 2220 -2976
rect 2214 -2988 2220 -2982
rect 2214 -2994 2220 -2988
rect 2214 -3000 2220 -2994
rect 2220 -174 2226 -168
rect 2220 -180 2226 -174
rect 2220 -186 2226 -180
rect 2220 -192 2226 -186
rect 2220 -198 2226 -192
rect 2220 -204 2226 -198
rect 2220 -210 2226 -204
rect 2220 -216 2226 -210
rect 2220 -222 2226 -216
rect 2220 -228 2226 -222
rect 2220 -234 2226 -228
rect 2220 -240 2226 -234
rect 2220 -246 2226 -240
rect 2220 -252 2226 -246
rect 2220 -258 2226 -252
rect 2220 -264 2226 -258
rect 2220 -270 2226 -264
rect 2220 -276 2226 -270
rect 2220 -282 2226 -276
rect 2220 -288 2226 -282
rect 2220 -294 2226 -288
rect 2220 -300 2226 -294
rect 2220 -306 2226 -300
rect 2220 -312 2226 -306
rect 2220 -318 2226 -312
rect 2220 -324 2226 -318
rect 2220 -330 2226 -324
rect 2220 -336 2226 -330
rect 2220 -342 2226 -336
rect 2220 -348 2226 -342
rect 2220 -354 2226 -348
rect 2220 -360 2226 -354
rect 2220 -366 2226 -360
rect 2220 -372 2226 -366
rect 2220 -378 2226 -372
rect 2220 -384 2226 -378
rect 2220 -390 2226 -384
rect 2220 -396 2226 -390
rect 2220 -402 2226 -396
rect 2220 -408 2226 -402
rect 2220 -414 2226 -408
rect 2220 -420 2226 -414
rect 2220 -426 2226 -420
rect 2220 -432 2226 -426
rect 2220 -438 2226 -432
rect 2220 -444 2226 -438
rect 2220 -450 2226 -444
rect 2220 -456 2226 -450
rect 2220 -462 2226 -456
rect 2220 -468 2226 -462
rect 2220 -474 2226 -468
rect 2220 -480 2226 -474
rect 2220 -486 2226 -480
rect 2220 -492 2226 -486
rect 2220 -498 2226 -492
rect 2220 -504 2226 -498
rect 2220 -510 2226 -504
rect 2220 -516 2226 -510
rect 2220 -522 2226 -516
rect 2220 -528 2226 -522
rect 2220 -534 2226 -528
rect 2220 -540 2226 -534
rect 2220 -546 2226 -540
rect 2220 -552 2226 -546
rect 2220 -558 2226 -552
rect 2220 -564 2226 -558
rect 2220 -570 2226 -564
rect 2220 -576 2226 -570
rect 2220 -582 2226 -576
rect 2220 -588 2226 -582
rect 2220 -594 2226 -588
rect 2220 -600 2226 -594
rect 2220 -606 2226 -600
rect 2220 -612 2226 -606
rect 2220 -618 2226 -612
rect 2220 -624 2226 -618
rect 2220 -630 2226 -624
rect 2220 -636 2226 -630
rect 2220 -642 2226 -636
rect 2220 -648 2226 -642
rect 2220 -654 2226 -648
rect 2220 -660 2226 -654
rect 2220 -666 2226 -660
rect 2220 -672 2226 -666
rect 2220 -678 2226 -672
rect 2220 -684 2226 -678
rect 2220 -690 2226 -684
rect 2220 -696 2226 -690
rect 2220 -702 2226 -696
rect 2220 -708 2226 -702
rect 2220 -714 2226 -708
rect 2220 -720 2226 -714
rect 2220 -726 2226 -720
rect 2220 -732 2226 -726
rect 2220 -738 2226 -732
rect 2220 -744 2226 -738
rect 2220 -750 2226 -744
rect 2220 -756 2226 -750
rect 2220 -762 2226 -756
rect 2220 -768 2226 -762
rect 2220 -774 2226 -768
rect 2220 -780 2226 -774
rect 2220 -786 2226 -780
rect 2220 -792 2226 -786
rect 2220 -798 2226 -792
rect 2220 -804 2226 -798
rect 2220 -810 2226 -804
rect 2220 -816 2226 -810
rect 2220 -822 2226 -816
rect 2220 -828 2226 -822
rect 2220 -834 2226 -828
rect 2220 -840 2226 -834
rect 2220 -846 2226 -840
rect 2220 -852 2226 -846
rect 2220 -858 2226 -852
rect 2220 -864 2226 -858
rect 2220 -870 2226 -864
rect 2220 -876 2226 -870
rect 2220 -882 2226 -876
rect 2220 -888 2226 -882
rect 2220 -894 2226 -888
rect 2220 -900 2226 -894
rect 2220 -906 2226 -900
rect 2220 -912 2226 -906
rect 2220 -918 2226 -912
rect 2220 -924 2226 -918
rect 2220 -930 2226 -924
rect 2220 -936 2226 -930
rect 2220 -942 2226 -936
rect 2220 -948 2226 -942
rect 2220 -954 2226 -948
rect 2220 -960 2226 -954
rect 2220 -966 2226 -960
rect 2220 -972 2226 -966
rect 2220 -978 2226 -972
rect 2220 -984 2226 -978
rect 2220 -990 2226 -984
rect 2220 -996 2226 -990
rect 2220 -1002 2226 -996
rect 2220 -1008 2226 -1002
rect 2220 -1014 2226 -1008
rect 2220 -1020 2226 -1014
rect 2220 -1026 2226 -1020
rect 2220 -1032 2226 -1026
rect 2220 -1038 2226 -1032
rect 2220 -1044 2226 -1038
rect 2220 -1050 2226 -1044
rect 2220 -1056 2226 -1050
rect 2220 -1062 2226 -1056
rect 2220 -1068 2226 -1062
rect 2220 -1074 2226 -1068
rect 2220 -1080 2226 -1074
rect 2220 -1086 2226 -1080
rect 2220 -1092 2226 -1086
rect 2220 -1098 2226 -1092
rect 2220 -1104 2226 -1098
rect 2220 -1110 2226 -1104
rect 2220 -1116 2226 -1110
rect 2220 -1122 2226 -1116
rect 2220 -1128 2226 -1122
rect 2220 -1134 2226 -1128
rect 2220 -1140 2226 -1134
rect 2220 -1146 2226 -1140
rect 2220 -1152 2226 -1146
rect 2220 -1158 2226 -1152
rect 2220 -1164 2226 -1158
rect 2220 -1170 2226 -1164
rect 2220 -1176 2226 -1170
rect 2220 -1182 2226 -1176
rect 2220 -1188 2226 -1182
rect 2220 -1194 2226 -1188
rect 2220 -1536 2226 -1530
rect 2220 -1542 2226 -1536
rect 2220 -1548 2226 -1542
rect 2220 -1554 2226 -1548
rect 2220 -1560 2226 -1554
rect 2220 -1566 2226 -1560
rect 2220 -1572 2226 -1566
rect 2220 -1578 2226 -1572
rect 2220 -1584 2226 -1578
rect 2220 -1590 2226 -1584
rect 2220 -1596 2226 -1590
rect 2220 -1602 2226 -1596
rect 2220 -1608 2226 -1602
rect 2220 -1614 2226 -1608
rect 2220 -1620 2226 -1614
rect 2220 -1626 2226 -1620
rect 2220 -1632 2226 -1626
rect 2220 -1638 2226 -1632
rect 2220 -1644 2226 -1638
rect 2220 -1650 2226 -1644
rect 2220 -1656 2226 -1650
rect 2220 -1662 2226 -1656
rect 2220 -1668 2226 -1662
rect 2220 -1674 2226 -1668
rect 2220 -1680 2226 -1674
rect 2220 -1686 2226 -1680
rect 2220 -1692 2226 -1686
rect 2220 -1698 2226 -1692
rect 2220 -1704 2226 -1698
rect 2220 -1710 2226 -1704
rect 2220 -1716 2226 -1710
rect 2220 -1722 2226 -1716
rect 2220 -1728 2226 -1722
rect 2220 -1734 2226 -1728
rect 2220 -1740 2226 -1734
rect 2220 -1746 2226 -1740
rect 2220 -1752 2226 -1746
rect 2220 -1758 2226 -1752
rect 2220 -1764 2226 -1758
rect 2220 -1770 2226 -1764
rect 2220 -1776 2226 -1770
rect 2220 -1782 2226 -1776
rect 2220 -1788 2226 -1782
rect 2220 -1794 2226 -1788
rect 2220 -1800 2226 -1794
rect 2220 -1806 2226 -1800
rect 2220 -1812 2226 -1806
rect 2220 -1818 2226 -1812
rect 2220 -1824 2226 -1818
rect 2220 -1830 2226 -1824
rect 2220 -1836 2226 -1830
rect 2220 -1842 2226 -1836
rect 2220 -1848 2226 -1842
rect 2220 -1854 2226 -1848
rect 2220 -1860 2226 -1854
rect 2220 -1866 2226 -1860
rect 2220 -1872 2226 -1866
rect 2220 -1878 2226 -1872
rect 2220 -1884 2226 -1878
rect 2220 -1890 2226 -1884
rect 2220 -1896 2226 -1890
rect 2220 -1902 2226 -1896
rect 2220 -1908 2226 -1902
rect 2220 -1914 2226 -1908
rect 2220 -1920 2226 -1914
rect 2220 -1926 2226 -1920
rect 2220 -1932 2226 -1926
rect 2220 -1938 2226 -1932
rect 2220 -1944 2226 -1938
rect 2220 -1950 2226 -1944
rect 2220 -1956 2226 -1950
rect 2220 -1962 2226 -1956
rect 2220 -1968 2226 -1962
rect 2220 -1974 2226 -1968
rect 2220 -1980 2226 -1974
rect 2220 -1986 2226 -1980
rect 2220 -1992 2226 -1986
rect 2220 -1998 2226 -1992
rect 2220 -2004 2226 -1998
rect 2220 -2010 2226 -2004
rect 2220 -2016 2226 -2010
rect 2220 -2022 2226 -2016
rect 2220 -2028 2226 -2022
rect 2220 -2034 2226 -2028
rect 2220 -2040 2226 -2034
rect 2220 -2046 2226 -2040
rect 2220 -2052 2226 -2046
rect 2220 -2058 2226 -2052
rect 2220 -2064 2226 -2058
rect 2220 -2070 2226 -2064
rect 2220 -2076 2226 -2070
rect 2220 -2082 2226 -2076
rect 2220 -2088 2226 -2082
rect 2220 -2094 2226 -2088
rect 2220 -2100 2226 -2094
rect 2220 -2106 2226 -2100
rect 2220 -2112 2226 -2106
rect 2220 -2118 2226 -2112
rect 2220 -2124 2226 -2118
rect 2220 -2130 2226 -2124
rect 2220 -2136 2226 -2130
rect 2220 -2142 2226 -2136
rect 2220 -2148 2226 -2142
rect 2220 -2154 2226 -2148
rect 2220 -2160 2226 -2154
rect 2220 -2166 2226 -2160
rect 2220 -2172 2226 -2166
rect 2220 -2178 2226 -2172
rect 2220 -2184 2226 -2178
rect 2220 -2190 2226 -2184
rect 2220 -2196 2226 -2190
rect 2220 -2202 2226 -2196
rect 2220 -2208 2226 -2202
rect 2220 -2214 2226 -2208
rect 2220 -2220 2226 -2214
rect 2220 -2226 2226 -2220
rect 2220 -2232 2226 -2226
rect 2220 -2238 2226 -2232
rect 2220 -2244 2226 -2238
rect 2220 -2250 2226 -2244
rect 2220 -2256 2226 -2250
rect 2220 -2262 2226 -2256
rect 2220 -2268 2226 -2262
rect 2220 -2274 2226 -2268
rect 2220 -2280 2226 -2274
rect 2220 -2286 2226 -2280
rect 2220 -2292 2226 -2286
rect 2220 -2298 2226 -2292
rect 2220 -2304 2226 -2298
rect 2220 -2310 2226 -2304
rect 2220 -2316 2226 -2310
rect 2220 -2388 2226 -2382
rect 2220 -2394 2226 -2388
rect 2220 -2400 2226 -2394
rect 2220 -2406 2226 -2400
rect 2220 -2412 2226 -2406
rect 2220 -2418 2226 -2412
rect 2220 -2424 2226 -2418
rect 2220 -2430 2226 -2424
rect 2220 -2436 2226 -2430
rect 2220 -2442 2226 -2436
rect 2220 -2448 2226 -2442
rect 2220 -2454 2226 -2448
rect 2220 -2460 2226 -2454
rect 2220 -2466 2226 -2460
rect 2220 -2472 2226 -2466
rect 2220 -2532 2226 -2526
rect 2220 -2538 2226 -2532
rect 2220 -2544 2226 -2538
rect 2220 -2550 2226 -2544
rect 2220 -2556 2226 -2550
rect 2220 -2562 2226 -2556
rect 2220 -2568 2226 -2562
rect 2220 -2574 2226 -2568
rect 2220 -2580 2226 -2574
rect 2220 -2586 2226 -2580
rect 2220 -2592 2226 -2586
rect 2220 -2598 2226 -2592
rect 2220 -2604 2226 -2598
rect 2220 -2610 2226 -2604
rect 2220 -2616 2226 -2610
rect 2220 -2622 2226 -2616
rect 2220 -2628 2226 -2622
rect 2220 -2634 2226 -2628
rect 2220 -2640 2226 -2634
rect 2220 -2646 2226 -2640
rect 2220 -2652 2226 -2646
rect 2220 -2658 2226 -2652
rect 2220 -2664 2226 -2658
rect 2220 -2670 2226 -2664
rect 2220 -2676 2226 -2670
rect 2220 -2682 2226 -2676
rect 2220 -2688 2226 -2682
rect 2220 -2694 2226 -2688
rect 2220 -2700 2226 -2694
rect 2220 -2706 2226 -2700
rect 2220 -2712 2226 -2706
rect 2220 -2718 2226 -2712
rect 2220 -2724 2226 -2718
rect 2220 -2730 2226 -2724
rect 2220 -2736 2226 -2730
rect 2220 -2742 2226 -2736
rect 2220 -2748 2226 -2742
rect 2220 -2754 2226 -2748
rect 2220 -2760 2226 -2754
rect 2220 -2766 2226 -2760
rect 2220 -2772 2226 -2766
rect 2220 -2778 2226 -2772
rect 2220 -2784 2226 -2778
rect 2220 -2790 2226 -2784
rect 2220 -2796 2226 -2790
rect 2220 -2802 2226 -2796
rect 2220 -2808 2226 -2802
rect 2220 -2814 2226 -2808
rect 2220 -2820 2226 -2814
rect 2220 -2826 2226 -2820
rect 2220 -2832 2226 -2826
rect 2220 -2838 2226 -2832
rect 2220 -2844 2226 -2838
rect 2220 -2850 2226 -2844
rect 2220 -2856 2226 -2850
rect 2220 -2862 2226 -2856
rect 2220 -2868 2226 -2862
rect 2220 -2874 2226 -2868
rect 2220 -2880 2226 -2874
rect 2220 -2886 2226 -2880
rect 2220 -2892 2226 -2886
rect 2220 -2898 2226 -2892
rect 2220 -2904 2226 -2898
rect 2220 -2910 2226 -2904
rect 2220 -2916 2226 -2910
rect 2220 -2922 2226 -2916
rect 2220 -2928 2226 -2922
rect 2220 -2934 2226 -2928
rect 2220 -2940 2226 -2934
rect 2220 -2946 2226 -2940
rect 2220 -2952 2226 -2946
rect 2220 -2958 2226 -2952
rect 2220 -2964 2226 -2958
rect 2220 -2970 2226 -2964
rect 2220 -2976 2226 -2970
rect 2220 -2982 2226 -2976
rect 2220 -2988 2226 -2982
rect 2220 -2994 2226 -2988
rect 2226 -168 2232 -162
rect 2226 -174 2232 -168
rect 2226 -180 2232 -174
rect 2226 -186 2232 -180
rect 2226 -192 2232 -186
rect 2226 -198 2232 -192
rect 2226 -204 2232 -198
rect 2226 -210 2232 -204
rect 2226 -216 2232 -210
rect 2226 -222 2232 -216
rect 2226 -228 2232 -222
rect 2226 -234 2232 -228
rect 2226 -240 2232 -234
rect 2226 -246 2232 -240
rect 2226 -252 2232 -246
rect 2226 -258 2232 -252
rect 2226 -264 2232 -258
rect 2226 -270 2232 -264
rect 2226 -276 2232 -270
rect 2226 -282 2232 -276
rect 2226 -288 2232 -282
rect 2226 -294 2232 -288
rect 2226 -300 2232 -294
rect 2226 -306 2232 -300
rect 2226 -312 2232 -306
rect 2226 -318 2232 -312
rect 2226 -324 2232 -318
rect 2226 -330 2232 -324
rect 2226 -336 2232 -330
rect 2226 -342 2232 -336
rect 2226 -348 2232 -342
rect 2226 -354 2232 -348
rect 2226 -360 2232 -354
rect 2226 -366 2232 -360
rect 2226 -372 2232 -366
rect 2226 -378 2232 -372
rect 2226 -384 2232 -378
rect 2226 -390 2232 -384
rect 2226 -396 2232 -390
rect 2226 -402 2232 -396
rect 2226 -408 2232 -402
rect 2226 -414 2232 -408
rect 2226 -420 2232 -414
rect 2226 -426 2232 -420
rect 2226 -432 2232 -426
rect 2226 -438 2232 -432
rect 2226 -444 2232 -438
rect 2226 -450 2232 -444
rect 2226 -456 2232 -450
rect 2226 -462 2232 -456
rect 2226 -468 2232 -462
rect 2226 -474 2232 -468
rect 2226 -480 2232 -474
rect 2226 -486 2232 -480
rect 2226 -492 2232 -486
rect 2226 -498 2232 -492
rect 2226 -504 2232 -498
rect 2226 -510 2232 -504
rect 2226 -516 2232 -510
rect 2226 -522 2232 -516
rect 2226 -528 2232 -522
rect 2226 -534 2232 -528
rect 2226 -540 2232 -534
rect 2226 -546 2232 -540
rect 2226 -552 2232 -546
rect 2226 -558 2232 -552
rect 2226 -564 2232 -558
rect 2226 -570 2232 -564
rect 2226 -576 2232 -570
rect 2226 -582 2232 -576
rect 2226 -588 2232 -582
rect 2226 -594 2232 -588
rect 2226 -600 2232 -594
rect 2226 -606 2232 -600
rect 2226 -612 2232 -606
rect 2226 -618 2232 -612
rect 2226 -624 2232 -618
rect 2226 -630 2232 -624
rect 2226 -636 2232 -630
rect 2226 -642 2232 -636
rect 2226 -648 2232 -642
rect 2226 -654 2232 -648
rect 2226 -660 2232 -654
rect 2226 -666 2232 -660
rect 2226 -672 2232 -666
rect 2226 -678 2232 -672
rect 2226 -684 2232 -678
rect 2226 -690 2232 -684
rect 2226 -696 2232 -690
rect 2226 -702 2232 -696
rect 2226 -708 2232 -702
rect 2226 -714 2232 -708
rect 2226 -720 2232 -714
rect 2226 -726 2232 -720
rect 2226 -732 2232 -726
rect 2226 -738 2232 -732
rect 2226 -744 2232 -738
rect 2226 -750 2232 -744
rect 2226 -756 2232 -750
rect 2226 -762 2232 -756
rect 2226 -768 2232 -762
rect 2226 -774 2232 -768
rect 2226 -780 2232 -774
rect 2226 -786 2232 -780
rect 2226 -792 2232 -786
rect 2226 -798 2232 -792
rect 2226 -804 2232 -798
rect 2226 -810 2232 -804
rect 2226 -816 2232 -810
rect 2226 -822 2232 -816
rect 2226 -828 2232 -822
rect 2226 -834 2232 -828
rect 2226 -840 2232 -834
rect 2226 -846 2232 -840
rect 2226 -852 2232 -846
rect 2226 -858 2232 -852
rect 2226 -864 2232 -858
rect 2226 -870 2232 -864
rect 2226 -876 2232 -870
rect 2226 -882 2232 -876
rect 2226 -888 2232 -882
rect 2226 -894 2232 -888
rect 2226 -900 2232 -894
rect 2226 -906 2232 -900
rect 2226 -912 2232 -906
rect 2226 -918 2232 -912
rect 2226 -924 2232 -918
rect 2226 -930 2232 -924
rect 2226 -936 2232 -930
rect 2226 -942 2232 -936
rect 2226 -948 2232 -942
rect 2226 -954 2232 -948
rect 2226 -960 2232 -954
rect 2226 -966 2232 -960
rect 2226 -972 2232 -966
rect 2226 -978 2232 -972
rect 2226 -984 2232 -978
rect 2226 -990 2232 -984
rect 2226 -996 2232 -990
rect 2226 -1002 2232 -996
rect 2226 -1008 2232 -1002
rect 2226 -1014 2232 -1008
rect 2226 -1020 2232 -1014
rect 2226 -1026 2232 -1020
rect 2226 -1032 2232 -1026
rect 2226 -1038 2232 -1032
rect 2226 -1044 2232 -1038
rect 2226 -1050 2232 -1044
rect 2226 -1056 2232 -1050
rect 2226 -1062 2232 -1056
rect 2226 -1068 2232 -1062
rect 2226 -1074 2232 -1068
rect 2226 -1080 2232 -1074
rect 2226 -1086 2232 -1080
rect 2226 -1092 2232 -1086
rect 2226 -1098 2232 -1092
rect 2226 -1104 2232 -1098
rect 2226 -1110 2232 -1104
rect 2226 -1116 2232 -1110
rect 2226 -1122 2232 -1116
rect 2226 -1128 2232 -1122
rect 2226 -1134 2232 -1128
rect 2226 -1140 2232 -1134
rect 2226 -1146 2232 -1140
rect 2226 -1152 2232 -1146
rect 2226 -1158 2232 -1152
rect 2226 -1164 2232 -1158
rect 2226 -1170 2232 -1164
rect 2226 -1176 2232 -1170
rect 2226 -1182 2232 -1176
rect 2226 -1530 2232 -1524
rect 2226 -1536 2232 -1530
rect 2226 -1542 2232 -1536
rect 2226 -1548 2232 -1542
rect 2226 -1554 2232 -1548
rect 2226 -1560 2232 -1554
rect 2226 -1566 2232 -1560
rect 2226 -1572 2232 -1566
rect 2226 -1578 2232 -1572
rect 2226 -1584 2232 -1578
rect 2226 -1590 2232 -1584
rect 2226 -1596 2232 -1590
rect 2226 -1602 2232 -1596
rect 2226 -1608 2232 -1602
rect 2226 -1614 2232 -1608
rect 2226 -1620 2232 -1614
rect 2226 -1626 2232 -1620
rect 2226 -1632 2232 -1626
rect 2226 -1638 2232 -1632
rect 2226 -1644 2232 -1638
rect 2226 -1650 2232 -1644
rect 2226 -1656 2232 -1650
rect 2226 -1662 2232 -1656
rect 2226 -1668 2232 -1662
rect 2226 -1674 2232 -1668
rect 2226 -1680 2232 -1674
rect 2226 -1686 2232 -1680
rect 2226 -1692 2232 -1686
rect 2226 -1698 2232 -1692
rect 2226 -1704 2232 -1698
rect 2226 -1710 2232 -1704
rect 2226 -1716 2232 -1710
rect 2226 -1722 2232 -1716
rect 2226 -1728 2232 -1722
rect 2226 -1734 2232 -1728
rect 2226 -1740 2232 -1734
rect 2226 -1746 2232 -1740
rect 2226 -1752 2232 -1746
rect 2226 -1758 2232 -1752
rect 2226 -1764 2232 -1758
rect 2226 -1770 2232 -1764
rect 2226 -1776 2232 -1770
rect 2226 -1782 2232 -1776
rect 2226 -1788 2232 -1782
rect 2226 -1794 2232 -1788
rect 2226 -1800 2232 -1794
rect 2226 -1806 2232 -1800
rect 2226 -1812 2232 -1806
rect 2226 -1818 2232 -1812
rect 2226 -1824 2232 -1818
rect 2226 -1830 2232 -1824
rect 2226 -1836 2232 -1830
rect 2226 -1842 2232 -1836
rect 2226 -1848 2232 -1842
rect 2226 -1854 2232 -1848
rect 2226 -1860 2232 -1854
rect 2226 -1866 2232 -1860
rect 2226 -1872 2232 -1866
rect 2226 -1878 2232 -1872
rect 2226 -1884 2232 -1878
rect 2226 -1890 2232 -1884
rect 2226 -1896 2232 -1890
rect 2226 -1902 2232 -1896
rect 2226 -1908 2232 -1902
rect 2226 -1914 2232 -1908
rect 2226 -1920 2232 -1914
rect 2226 -1926 2232 -1920
rect 2226 -1932 2232 -1926
rect 2226 -1938 2232 -1932
rect 2226 -1944 2232 -1938
rect 2226 -1950 2232 -1944
rect 2226 -1956 2232 -1950
rect 2226 -1962 2232 -1956
rect 2226 -1968 2232 -1962
rect 2226 -1974 2232 -1968
rect 2226 -1980 2232 -1974
rect 2226 -1986 2232 -1980
rect 2226 -1992 2232 -1986
rect 2226 -1998 2232 -1992
rect 2226 -2004 2232 -1998
rect 2226 -2010 2232 -2004
rect 2226 -2016 2232 -2010
rect 2226 -2022 2232 -2016
rect 2226 -2028 2232 -2022
rect 2226 -2034 2232 -2028
rect 2226 -2040 2232 -2034
rect 2226 -2046 2232 -2040
rect 2226 -2052 2232 -2046
rect 2226 -2058 2232 -2052
rect 2226 -2064 2232 -2058
rect 2226 -2070 2232 -2064
rect 2226 -2076 2232 -2070
rect 2226 -2082 2232 -2076
rect 2226 -2088 2232 -2082
rect 2226 -2094 2232 -2088
rect 2226 -2100 2232 -2094
rect 2226 -2106 2232 -2100
rect 2226 -2112 2232 -2106
rect 2226 -2118 2232 -2112
rect 2226 -2124 2232 -2118
rect 2226 -2130 2232 -2124
rect 2226 -2136 2232 -2130
rect 2226 -2142 2232 -2136
rect 2226 -2148 2232 -2142
rect 2226 -2154 2232 -2148
rect 2226 -2160 2232 -2154
rect 2226 -2166 2232 -2160
rect 2226 -2172 2232 -2166
rect 2226 -2178 2232 -2172
rect 2226 -2184 2232 -2178
rect 2226 -2190 2232 -2184
rect 2226 -2196 2232 -2190
rect 2226 -2202 2232 -2196
rect 2226 -2208 2232 -2202
rect 2226 -2214 2232 -2208
rect 2226 -2220 2232 -2214
rect 2226 -2226 2232 -2220
rect 2226 -2232 2232 -2226
rect 2226 -2238 2232 -2232
rect 2226 -2244 2232 -2238
rect 2226 -2250 2232 -2244
rect 2226 -2256 2232 -2250
rect 2226 -2262 2232 -2256
rect 2226 -2268 2232 -2262
rect 2226 -2274 2232 -2268
rect 2226 -2280 2232 -2274
rect 2226 -2286 2232 -2280
rect 2226 -2292 2232 -2286
rect 2226 -2298 2232 -2292
rect 2226 -2304 2232 -2298
rect 2226 -2310 2232 -2304
rect 2226 -2376 2232 -2370
rect 2226 -2382 2232 -2376
rect 2226 -2388 2232 -2382
rect 2226 -2394 2232 -2388
rect 2226 -2400 2232 -2394
rect 2226 -2406 2232 -2400
rect 2226 -2412 2232 -2406
rect 2226 -2418 2232 -2412
rect 2226 -2424 2232 -2418
rect 2226 -2430 2232 -2424
rect 2226 -2436 2232 -2430
rect 2226 -2442 2232 -2436
rect 2226 -2448 2232 -2442
rect 2226 -2454 2232 -2448
rect 2226 -2460 2232 -2454
rect 2226 -2466 2232 -2460
rect 2226 -2472 2232 -2466
rect 2226 -2532 2232 -2526
rect 2226 -2538 2232 -2532
rect 2226 -2544 2232 -2538
rect 2226 -2550 2232 -2544
rect 2226 -2556 2232 -2550
rect 2226 -2562 2232 -2556
rect 2226 -2568 2232 -2562
rect 2226 -2574 2232 -2568
rect 2226 -2580 2232 -2574
rect 2226 -2586 2232 -2580
rect 2226 -2592 2232 -2586
rect 2226 -2598 2232 -2592
rect 2226 -2604 2232 -2598
rect 2226 -2610 2232 -2604
rect 2226 -2616 2232 -2610
rect 2226 -2622 2232 -2616
rect 2226 -2628 2232 -2622
rect 2226 -2634 2232 -2628
rect 2226 -2640 2232 -2634
rect 2226 -2646 2232 -2640
rect 2226 -2652 2232 -2646
rect 2226 -2658 2232 -2652
rect 2226 -2664 2232 -2658
rect 2226 -2670 2232 -2664
rect 2226 -2676 2232 -2670
rect 2226 -2682 2232 -2676
rect 2226 -2688 2232 -2682
rect 2226 -2694 2232 -2688
rect 2226 -2700 2232 -2694
rect 2226 -2706 2232 -2700
rect 2226 -2712 2232 -2706
rect 2226 -2718 2232 -2712
rect 2226 -2724 2232 -2718
rect 2226 -2730 2232 -2724
rect 2226 -2736 2232 -2730
rect 2226 -2742 2232 -2736
rect 2226 -2748 2232 -2742
rect 2226 -2754 2232 -2748
rect 2226 -2760 2232 -2754
rect 2226 -2766 2232 -2760
rect 2226 -2772 2232 -2766
rect 2226 -2778 2232 -2772
rect 2226 -2784 2232 -2778
rect 2226 -2790 2232 -2784
rect 2226 -2796 2232 -2790
rect 2226 -2802 2232 -2796
rect 2226 -2808 2232 -2802
rect 2226 -2814 2232 -2808
rect 2226 -2820 2232 -2814
rect 2226 -2826 2232 -2820
rect 2226 -2832 2232 -2826
rect 2226 -2838 2232 -2832
rect 2226 -2844 2232 -2838
rect 2226 -2850 2232 -2844
rect 2226 -2856 2232 -2850
rect 2226 -2862 2232 -2856
rect 2226 -2868 2232 -2862
rect 2226 -2874 2232 -2868
rect 2226 -2880 2232 -2874
rect 2226 -2886 2232 -2880
rect 2226 -2892 2232 -2886
rect 2226 -2898 2232 -2892
rect 2226 -2904 2232 -2898
rect 2226 -2910 2232 -2904
rect 2226 -2916 2232 -2910
rect 2226 -2922 2232 -2916
rect 2226 -2928 2232 -2922
rect 2226 -2934 2232 -2928
rect 2226 -2940 2232 -2934
rect 2226 -2946 2232 -2940
rect 2226 -2952 2232 -2946
rect 2226 -2958 2232 -2952
rect 2226 -2964 2232 -2958
rect 2226 -2970 2232 -2964
rect 2226 -2976 2232 -2970
rect 2226 -2982 2232 -2976
rect 2226 -2988 2232 -2982
rect 2232 -156 2238 -150
rect 2232 -162 2238 -156
rect 2232 -168 2238 -162
rect 2232 -174 2238 -168
rect 2232 -180 2238 -174
rect 2232 -186 2238 -180
rect 2232 -192 2238 -186
rect 2232 -198 2238 -192
rect 2232 -204 2238 -198
rect 2232 -210 2238 -204
rect 2232 -216 2238 -210
rect 2232 -222 2238 -216
rect 2232 -228 2238 -222
rect 2232 -234 2238 -228
rect 2232 -240 2238 -234
rect 2232 -246 2238 -240
rect 2232 -252 2238 -246
rect 2232 -258 2238 -252
rect 2232 -264 2238 -258
rect 2232 -270 2238 -264
rect 2232 -276 2238 -270
rect 2232 -282 2238 -276
rect 2232 -288 2238 -282
rect 2232 -294 2238 -288
rect 2232 -300 2238 -294
rect 2232 -306 2238 -300
rect 2232 -312 2238 -306
rect 2232 -318 2238 -312
rect 2232 -324 2238 -318
rect 2232 -330 2238 -324
rect 2232 -336 2238 -330
rect 2232 -342 2238 -336
rect 2232 -348 2238 -342
rect 2232 -354 2238 -348
rect 2232 -360 2238 -354
rect 2232 -366 2238 -360
rect 2232 -372 2238 -366
rect 2232 -378 2238 -372
rect 2232 -384 2238 -378
rect 2232 -390 2238 -384
rect 2232 -396 2238 -390
rect 2232 -402 2238 -396
rect 2232 -408 2238 -402
rect 2232 -414 2238 -408
rect 2232 -420 2238 -414
rect 2232 -426 2238 -420
rect 2232 -432 2238 -426
rect 2232 -438 2238 -432
rect 2232 -444 2238 -438
rect 2232 -450 2238 -444
rect 2232 -456 2238 -450
rect 2232 -462 2238 -456
rect 2232 -468 2238 -462
rect 2232 -474 2238 -468
rect 2232 -480 2238 -474
rect 2232 -486 2238 -480
rect 2232 -492 2238 -486
rect 2232 -498 2238 -492
rect 2232 -504 2238 -498
rect 2232 -510 2238 -504
rect 2232 -516 2238 -510
rect 2232 -522 2238 -516
rect 2232 -528 2238 -522
rect 2232 -534 2238 -528
rect 2232 -540 2238 -534
rect 2232 -546 2238 -540
rect 2232 -552 2238 -546
rect 2232 -558 2238 -552
rect 2232 -564 2238 -558
rect 2232 -570 2238 -564
rect 2232 -576 2238 -570
rect 2232 -582 2238 -576
rect 2232 -588 2238 -582
rect 2232 -594 2238 -588
rect 2232 -600 2238 -594
rect 2232 -606 2238 -600
rect 2232 -612 2238 -606
rect 2232 -618 2238 -612
rect 2232 -624 2238 -618
rect 2232 -630 2238 -624
rect 2232 -636 2238 -630
rect 2232 -642 2238 -636
rect 2232 -648 2238 -642
rect 2232 -654 2238 -648
rect 2232 -660 2238 -654
rect 2232 -666 2238 -660
rect 2232 -672 2238 -666
rect 2232 -678 2238 -672
rect 2232 -684 2238 -678
rect 2232 -690 2238 -684
rect 2232 -696 2238 -690
rect 2232 -702 2238 -696
rect 2232 -708 2238 -702
rect 2232 -714 2238 -708
rect 2232 -720 2238 -714
rect 2232 -726 2238 -720
rect 2232 -732 2238 -726
rect 2232 -738 2238 -732
rect 2232 -744 2238 -738
rect 2232 -750 2238 -744
rect 2232 -756 2238 -750
rect 2232 -762 2238 -756
rect 2232 -768 2238 -762
rect 2232 -774 2238 -768
rect 2232 -780 2238 -774
rect 2232 -786 2238 -780
rect 2232 -792 2238 -786
rect 2232 -798 2238 -792
rect 2232 -804 2238 -798
rect 2232 -810 2238 -804
rect 2232 -816 2238 -810
rect 2232 -822 2238 -816
rect 2232 -828 2238 -822
rect 2232 -834 2238 -828
rect 2232 -840 2238 -834
rect 2232 -846 2238 -840
rect 2232 -852 2238 -846
rect 2232 -858 2238 -852
rect 2232 -864 2238 -858
rect 2232 -870 2238 -864
rect 2232 -876 2238 -870
rect 2232 -882 2238 -876
rect 2232 -888 2238 -882
rect 2232 -894 2238 -888
rect 2232 -900 2238 -894
rect 2232 -906 2238 -900
rect 2232 -912 2238 -906
rect 2232 -918 2238 -912
rect 2232 -924 2238 -918
rect 2232 -930 2238 -924
rect 2232 -936 2238 -930
rect 2232 -942 2238 -936
rect 2232 -948 2238 -942
rect 2232 -954 2238 -948
rect 2232 -960 2238 -954
rect 2232 -966 2238 -960
rect 2232 -972 2238 -966
rect 2232 -978 2238 -972
rect 2232 -984 2238 -978
rect 2232 -990 2238 -984
rect 2232 -996 2238 -990
rect 2232 -1002 2238 -996
rect 2232 -1008 2238 -1002
rect 2232 -1014 2238 -1008
rect 2232 -1020 2238 -1014
rect 2232 -1026 2238 -1020
rect 2232 -1032 2238 -1026
rect 2232 -1038 2238 -1032
rect 2232 -1044 2238 -1038
rect 2232 -1050 2238 -1044
rect 2232 -1056 2238 -1050
rect 2232 -1062 2238 -1056
rect 2232 -1068 2238 -1062
rect 2232 -1074 2238 -1068
rect 2232 -1080 2238 -1074
rect 2232 -1086 2238 -1080
rect 2232 -1092 2238 -1086
rect 2232 -1098 2238 -1092
rect 2232 -1104 2238 -1098
rect 2232 -1110 2238 -1104
rect 2232 -1116 2238 -1110
rect 2232 -1122 2238 -1116
rect 2232 -1128 2238 -1122
rect 2232 -1134 2238 -1128
rect 2232 -1140 2238 -1134
rect 2232 -1146 2238 -1140
rect 2232 -1152 2238 -1146
rect 2232 -1158 2238 -1152
rect 2232 -1164 2238 -1158
rect 2232 -1524 2238 -1518
rect 2232 -1530 2238 -1524
rect 2232 -1536 2238 -1530
rect 2232 -1542 2238 -1536
rect 2232 -1548 2238 -1542
rect 2232 -1554 2238 -1548
rect 2232 -1560 2238 -1554
rect 2232 -1566 2238 -1560
rect 2232 -1572 2238 -1566
rect 2232 -1578 2238 -1572
rect 2232 -1584 2238 -1578
rect 2232 -1590 2238 -1584
rect 2232 -1596 2238 -1590
rect 2232 -1602 2238 -1596
rect 2232 -1608 2238 -1602
rect 2232 -1614 2238 -1608
rect 2232 -1620 2238 -1614
rect 2232 -1626 2238 -1620
rect 2232 -1632 2238 -1626
rect 2232 -1638 2238 -1632
rect 2232 -1644 2238 -1638
rect 2232 -1650 2238 -1644
rect 2232 -1656 2238 -1650
rect 2232 -1662 2238 -1656
rect 2232 -1668 2238 -1662
rect 2232 -1674 2238 -1668
rect 2232 -1680 2238 -1674
rect 2232 -1686 2238 -1680
rect 2232 -1692 2238 -1686
rect 2232 -1698 2238 -1692
rect 2232 -1704 2238 -1698
rect 2232 -1710 2238 -1704
rect 2232 -1716 2238 -1710
rect 2232 -1722 2238 -1716
rect 2232 -1728 2238 -1722
rect 2232 -1734 2238 -1728
rect 2232 -1740 2238 -1734
rect 2232 -1746 2238 -1740
rect 2232 -1752 2238 -1746
rect 2232 -1758 2238 -1752
rect 2232 -1764 2238 -1758
rect 2232 -1770 2238 -1764
rect 2232 -1776 2238 -1770
rect 2232 -1782 2238 -1776
rect 2232 -1788 2238 -1782
rect 2232 -1794 2238 -1788
rect 2232 -1800 2238 -1794
rect 2232 -1806 2238 -1800
rect 2232 -1812 2238 -1806
rect 2232 -1818 2238 -1812
rect 2232 -1824 2238 -1818
rect 2232 -1830 2238 -1824
rect 2232 -1836 2238 -1830
rect 2232 -1842 2238 -1836
rect 2232 -1848 2238 -1842
rect 2232 -1854 2238 -1848
rect 2232 -1860 2238 -1854
rect 2232 -1866 2238 -1860
rect 2232 -1872 2238 -1866
rect 2232 -1878 2238 -1872
rect 2232 -1884 2238 -1878
rect 2232 -1890 2238 -1884
rect 2232 -1896 2238 -1890
rect 2232 -1902 2238 -1896
rect 2232 -1908 2238 -1902
rect 2232 -1914 2238 -1908
rect 2232 -1920 2238 -1914
rect 2232 -1926 2238 -1920
rect 2232 -1932 2238 -1926
rect 2232 -1938 2238 -1932
rect 2232 -1944 2238 -1938
rect 2232 -1950 2238 -1944
rect 2232 -1956 2238 -1950
rect 2232 -1962 2238 -1956
rect 2232 -1968 2238 -1962
rect 2232 -1974 2238 -1968
rect 2232 -1980 2238 -1974
rect 2232 -1986 2238 -1980
rect 2232 -1992 2238 -1986
rect 2232 -1998 2238 -1992
rect 2232 -2004 2238 -1998
rect 2232 -2010 2238 -2004
rect 2232 -2016 2238 -2010
rect 2232 -2022 2238 -2016
rect 2232 -2028 2238 -2022
rect 2232 -2034 2238 -2028
rect 2232 -2040 2238 -2034
rect 2232 -2046 2238 -2040
rect 2232 -2052 2238 -2046
rect 2232 -2058 2238 -2052
rect 2232 -2064 2238 -2058
rect 2232 -2070 2238 -2064
rect 2232 -2076 2238 -2070
rect 2232 -2082 2238 -2076
rect 2232 -2088 2238 -2082
rect 2232 -2094 2238 -2088
rect 2232 -2100 2238 -2094
rect 2232 -2106 2238 -2100
rect 2232 -2112 2238 -2106
rect 2232 -2118 2238 -2112
rect 2232 -2124 2238 -2118
rect 2232 -2130 2238 -2124
rect 2232 -2136 2238 -2130
rect 2232 -2142 2238 -2136
rect 2232 -2148 2238 -2142
rect 2232 -2154 2238 -2148
rect 2232 -2160 2238 -2154
rect 2232 -2166 2238 -2160
rect 2232 -2172 2238 -2166
rect 2232 -2178 2238 -2172
rect 2232 -2184 2238 -2178
rect 2232 -2190 2238 -2184
rect 2232 -2196 2238 -2190
rect 2232 -2202 2238 -2196
rect 2232 -2208 2238 -2202
rect 2232 -2214 2238 -2208
rect 2232 -2220 2238 -2214
rect 2232 -2226 2238 -2220
rect 2232 -2232 2238 -2226
rect 2232 -2238 2238 -2232
rect 2232 -2244 2238 -2238
rect 2232 -2250 2238 -2244
rect 2232 -2256 2238 -2250
rect 2232 -2262 2238 -2256
rect 2232 -2268 2238 -2262
rect 2232 -2274 2238 -2268
rect 2232 -2280 2238 -2274
rect 2232 -2286 2238 -2280
rect 2232 -2292 2238 -2286
rect 2232 -2298 2238 -2292
rect 2232 -2304 2238 -2298
rect 2232 -2370 2238 -2364
rect 2232 -2376 2238 -2370
rect 2232 -2382 2238 -2376
rect 2232 -2388 2238 -2382
rect 2232 -2394 2238 -2388
rect 2232 -2400 2238 -2394
rect 2232 -2406 2238 -2400
rect 2232 -2412 2238 -2406
rect 2232 -2418 2238 -2412
rect 2232 -2424 2238 -2418
rect 2232 -2430 2238 -2424
rect 2232 -2436 2238 -2430
rect 2232 -2442 2238 -2436
rect 2232 -2448 2238 -2442
rect 2232 -2454 2238 -2448
rect 2232 -2460 2238 -2454
rect 2232 -2466 2238 -2460
rect 2232 -2526 2238 -2520
rect 2232 -2532 2238 -2526
rect 2232 -2538 2238 -2532
rect 2232 -2544 2238 -2538
rect 2232 -2550 2238 -2544
rect 2232 -2556 2238 -2550
rect 2232 -2562 2238 -2556
rect 2232 -2568 2238 -2562
rect 2232 -2574 2238 -2568
rect 2232 -2580 2238 -2574
rect 2232 -2586 2238 -2580
rect 2232 -2592 2238 -2586
rect 2232 -2598 2238 -2592
rect 2232 -2604 2238 -2598
rect 2232 -2610 2238 -2604
rect 2232 -2616 2238 -2610
rect 2232 -2622 2238 -2616
rect 2232 -2628 2238 -2622
rect 2232 -2634 2238 -2628
rect 2232 -2640 2238 -2634
rect 2232 -2646 2238 -2640
rect 2232 -2652 2238 -2646
rect 2232 -2658 2238 -2652
rect 2232 -2664 2238 -2658
rect 2232 -2670 2238 -2664
rect 2232 -2676 2238 -2670
rect 2232 -2682 2238 -2676
rect 2232 -2688 2238 -2682
rect 2232 -2694 2238 -2688
rect 2232 -2700 2238 -2694
rect 2232 -2706 2238 -2700
rect 2232 -2712 2238 -2706
rect 2232 -2718 2238 -2712
rect 2232 -2724 2238 -2718
rect 2232 -2730 2238 -2724
rect 2232 -2736 2238 -2730
rect 2232 -2742 2238 -2736
rect 2232 -2748 2238 -2742
rect 2232 -2754 2238 -2748
rect 2232 -2760 2238 -2754
rect 2232 -2766 2238 -2760
rect 2232 -2772 2238 -2766
rect 2232 -2778 2238 -2772
rect 2232 -2784 2238 -2778
rect 2232 -2790 2238 -2784
rect 2232 -2796 2238 -2790
rect 2232 -2802 2238 -2796
rect 2232 -2808 2238 -2802
rect 2232 -2814 2238 -2808
rect 2232 -2820 2238 -2814
rect 2232 -2826 2238 -2820
rect 2232 -2832 2238 -2826
rect 2232 -2838 2238 -2832
rect 2232 -2844 2238 -2838
rect 2232 -2850 2238 -2844
rect 2232 -2856 2238 -2850
rect 2232 -2862 2238 -2856
rect 2232 -2868 2238 -2862
rect 2232 -2874 2238 -2868
rect 2232 -2880 2238 -2874
rect 2232 -2886 2238 -2880
rect 2232 -2892 2238 -2886
rect 2232 -2898 2238 -2892
rect 2232 -2904 2238 -2898
rect 2232 -2910 2238 -2904
rect 2232 -2916 2238 -2910
rect 2232 -2922 2238 -2916
rect 2232 -2928 2238 -2922
rect 2232 -2934 2238 -2928
rect 2232 -2940 2238 -2934
rect 2232 -2946 2238 -2940
rect 2232 -2952 2238 -2946
rect 2232 -2958 2238 -2952
rect 2232 -2964 2238 -2958
rect 2232 -2970 2238 -2964
rect 2232 -2976 2238 -2970
rect 2232 -2982 2238 -2976
rect 2232 -2988 2238 -2982
rect 2238 -150 2244 -144
rect 2238 -156 2244 -150
rect 2238 -162 2244 -156
rect 2238 -168 2244 -162
rect 2238 -174 2244 -168
rect 2238 -180 2244 -174
rect 2238 -186 2244 -180
rect 2238 -192 2244 -186
rect 2238 -198 2244 -192
rect 2238 -204 2244 -198
rect 2238 -210 2244 -204
rect 2238 -216 2244 -210
rect 2238 -222 2244 -216
rect 2238 -228 2244 -222
rect 2238 -234 2244 -228
rect 2238 -240 2244 -234
rect 2238 -246 2244 -240
rect 2238 -252 2244 -246
rect 2238 -258 2244 -252
rect 2238 -264 2244 -258
rect 2238 -270 2244 -264
rect 2238 -276 2244 -270
rect 2238 -282 2244 -276
rect 2238 -288 2244 -282
rect 2238 -294 2244 -288
rect 2238 -300 2244 -294
rect 2238 -306 2244 -300
rect 2238 -312 2244 -306
rect 2238 -318 2244 -312
rect 2238 -324 2244 -318
rect 2238 -330 2244 -324
rect 2238 -336 2244 -330
rect 2238 -342 2244 -336
rect 2238 -348 2244 -342
rect 2238 -354 2244 -348
rect 2238 -360 2244 -354
rect 2238 -366 2244 -360
rect 2238 -372 2244 -366
rect 2238 -378 2244 -372
rect 2238 -384 2244 -378
rect 2238 -390 2244 -384
rect 2238 -396 2244 -390
rect 2238 -402 2244 -396
rect 2238 -408 2244 -402
rect 2238 -414 2244 -408
rect 2238 -420 2244 -414
rect 2238 -426 2244 -420
rect 2238 -432 2244 -426
rect 2238 -438 2244 -432
rect 2238 -444 2244 -438
rect 2238 -450 2244 -444
rect 2238 -456 2244 -450
rect 2238 -462 2244 -456
rect 2238 -468 2244 -462
rect 2238 -474 2244 -468
rect 2238 -480 2244 -474
rect 2238 -486 2244 -480
rect 2238 -492 2244 -486
rect 2238 -498 2244 -492
rect 2238 -504 2244 -498
rect 2238 -510 2244 -504
rect 2238 -516 2244 -510
rect 2238 -522 2244 -516
rect 2238 -528 2244 -522
rect 2238 -534 2244 -528
rect 2238 -540 2244 -534
rect 2238 -546 2244 -540
rect 2238 -552 2244 -546
rect 2238 -558 2244 -552
rect 2238 -564 2244 -558
rect 2238 -570 2244 -564
rect 2238 -576 2244 -570
rect 2238 -582 2244 -576
rect 2238 -588 2244 -582
rect 2238 -594 2244 -588
rect 2238 -600 2244 -594
rect 2238 -606 2244 -600
rect 2238 -612 2244 -606
rect 2238 -618 2244 -612
rect 2238 -624 2244 -618
rect 2238 -630 2244 -624
rect 2238 -636 2244 -630
rect 2238 -642 2244 -636
rect 2238 -648 2244 -642
rect 2238 -654 2244 -648
rect 2238 -660 2244 -654
rect 2238 -666 2244 -660
rect 2238 -672 2244 -666
rect 2238 -678 2244 -672
rect 2238 -684 2244 -678
rect 2238 -690 2244 -684
rect 2238 -696 2244 -690
rect 2238 -702 2244 -696
rect 2238 -708 2244 -702
rect 2238 -714 2244 -708
rect 2238 -720 2244 -714
rect 2238 -726 2244 -720
rect 2238 -732 2244 -726
rect 2238 -738 2244 -732
rect 2238 -744 2244 -738
rect 2238 -750 2244 -744
rect 2238 -756 2244 -750
rect 2238 -762 2244 -756
rect 2238 -768 2244 -762
rect 2238 -774 2244 -768
rect 2238 -780 2244 -774
rect 2238 -786 2244 -780
rect 2238 -792 2244 -786
rect 2238 -798 2244 -792
rect 2238 -804 2244 -798
rect 2238 -810 2244 -804
rect 2238 -816 2244 -810
rect 2238 -822 2244 -816
rect 2238 -828 2244 -822
rect 2238 -834 2244 -828
rect 2238 -840 2244 -834
rect 2238 -846 2244 -840
rect 2238 -852 2244 -846
rect 2238 -858 2244 -852
rect 2238 -864 2244 -858
rect 2238 -870 2244 -864
rect 2238 -876 2244 -870
rect 2238 -882 2244 -876
rect 2238 -888 2244 -882
rect 2238 -894 2244 -888
rect 2238 -900 2244 -894
rect 2238 -906 2244 -900
rect 2238 -912 2244 -906
rect 2238 -918 2244 -912
rect 2238 -924 2244 -918
rect 2238 -930 2244 -924
rect 2238 -936 2244 -930
rect 2238 -942 2244 -936
rect 2238 -948 2244 -942
rect 2238 -954 2244 -948
rect 2238 -960 2244 -954
rect 2238 -966 2244 -960
rect 2238 -972 2244 -966
rect 2238 -978 2244 -972
rect 2238 -984 2244 -978
rect 2238 -990 2244 -984
rect 2238 -996 2244 -990
rect 2238 -1002 2244 -996
rect 2238 -1008 2244 -1002
rect 2238 -1014 2244 -1008
rect 2238 -1020 2244 -1014
rect 2238 -1026 2244 -1020
rect 2238 -1032 2244 -1026
rect 2238 -1038 2244 -1032
rect 2238 -1044 2244 -1038
rect 2238 -1050 2244 -1044
rect 2238 -1056 2244 -1050
rect 2238 -1062 2244 -1056
rect 2238 -1068 2244 -1062
rect 2238 -1074 2244 -1068
rect 2238 -1080 2244 -1074
rect 2238 -1086 2244 -1080
rect 2238 -1092 2244 -1086
rect 2238 -1098 2244 -1092
rect 2238 -1104 2244 -1098
rect 2238 -1110 2244 -1104
rect 2238 -1116 2244 -1110
rect 2238 -1122 2244 -1116
rect 2238 -1128 2244 -1122
rect 2238 -1134 2244 -1128
rect 2238 -1140 2244 -1134
rect 2238 -1146 2244 -1140
rect 2238 -1152 2244 -1146
rect 2238 -1518 2244 -1512
rect 2238 -1524 2244 -1518
rect 2238 -1530 2244 -1524
rect 2238 -1536 2244 -1530
rect 2238 -1542 2244 -1536
rect 2238 -1548 2244 -1542
rect 2238 -1554 2244 -1548
rect 2238 -1560 2244 -1554
rect 2238 -1566 2244 -1560
rect 2238 -1572 2244 -1566
rect 2238 -1578 2244 -1572
rect 2238 -1584 2244 -1578
rect 2238 -1590 2244 -1584
rect 2238 -1596 2244 -1590
rect 2238 -1602 2244 -1596
rect 2238 -1608 2244 -1602
rect 2238 -1614 2244 -1608
rect 2238 -1620 2244 -1614
rect 2238 -1626 2244 -1620
rect 2238 -1632 2244 -1626
rect 2238 -1638 2244 -1632
rect 2238 -1644 2244 -1638
rect 2238 -1650 2244 -1644
rect 2238 -1656 2244 -1650
rect 2238 -1662 2244 -1656
rect 2238 -1668 2244 -1662
rect 2238 -1674 2244 -1668
rect 2238 -1680 2244 -1674
rect 2238 -1686 2244 -1680
rect 2238 -1692 2244 -1686
rect 2238 -1698 2244 -1692
rect 2238 -1704 2244 -1698
rect 2238 -1710 2244 -1704
rect 2238 -1716 2244 -1710
rect 2238 -1722 2244 -1716
rect 2238 -1728 2244 -1722
rect 2238 -1734 2244 -1728
rect 2238 -1740 2244 -1734
rect 2238 -1746 2244 -1740
rect 2238 -1752 2244 -1746
rect 2238 -1758 2244 -1752
rect 2238 -1764 2244 -1758
rect 2238 -1770 2244 -1764
rect 2238 -1776 2244 -1770
rect 2238 -1782 2244 -1776
rect 2238 -1788 2244 -1782
rect 2238 -1794 2244 -1788
rect 2238 -1800 2244 -1794
rect 2238 -1806 2244 -1800
rect 2238 -1812 2244 -1806
rect 2238 -1818 2244 -1812
rect 2238 -1824 2244 -1818
rect 2238 -1830 2244 -1824
rect 2238 -1836 2244 -1830
rect 2238 -1842 2244 -1836
rect 2238 -1848 2244 -1842
rect 2238 -1854 2244 -1848
rect 2238 -1860 2244 -1854
rect 2238 -1866 2244 -1860
rect 2238 -1872 2244 -1866
rect 2238 -1878 2244 -1872
rect 2238 -1884 2244 -1878
rect 2238 -1890 2244 -1884
rect 2238 -1896 2244 -1890
rect 2238 -1902 2244 -1896
rect 2238 -1908 2244 -1902
rect 2238 -1914 2244 -1908
rect 2238 -1920 2244 -1914
rect 2238 -1926 2244 -1920
rect 2238 -1932 2244 -1926
rect 2238 -1938 2244 -1932
rect 2238 -1944 2244 -1938
rect 2238 -1950 2244 -1944
rect 2238 -1956 2244 -1950
rect 2238 -1962 2244 -1956
rect 2238 -1968 2244 -1962
rect 2238 -1974 2244 -1968
rect 2238 -1980 2244 -1974
rect 2238 -1986 2244 -1980
rect 2238 -1992 2244 -1986
rect 2238 -1998 2244 -1992
rect 2238 -2004 2244 -1998
rect 2238 -2010 2244 -2004
rect 2238 -2016 2244 -2010
rect 2238 -2022 2244 -2016
rect 2238 -2028 2244 -2022
rect 2238 -2034 2244 -2028
rect 2238 -2040 2244 -2034
rect 2238 -2046 2244 -2040
rect 2238 -2052 2244 -2046
rect 2238 -2058 2244 -2052
rect 2238 -2064 2244 -2058
rect 2238 -2070 2244 -2064
rect 2238 -2076 2244 -2070
rect 2238 -2082 2244 -2076
rect 2238 -2088 2244 -2082
rect 2238 -2094 2244 -2088
rect 2238 -2100 2244 -2094
rect 2238 -2106 2244 -2100
rect 2238 -2112 2244 -2106
rect 2238 -2118 2244 -2112
rect 2238 -2124 2244 -2118
rect 2238 -2130 2244 -2124
rect 2238 -2136 2244 -2130
rect 2238 -2142 2244 -2136
rect 2238 -2148 2244 -2142
rect 2238 -2154 2244 -2148
rect 2238 -2160 2244 -2154
rect 2238 -2166 2244 -2160
rect 2238 -2172 2244 -2166
rect 2238 -2178 2244 -2172
rect 2238 -2184 2244 -2178
rect 2238 -2190 2244 -2184
rect 2238 -2196 2244 -2190
rect 2238 -2202 2244 -2196
rect 2238 -2208 2244 -2202
rect 2238 -2214 2244 -2208
rect 2238 -2220 2244 -2214
rect 2238 -2226 2244 -2220
rect 2238 -2232 2244 -2226
rect 2238 -2238 2244 -2232
rect 2238 -2244 2244 -2238
rect 2238 -2250 2244 -2244
rect 2238 -2256 2244 -2250
rect 2238 -2262 2244 -2256
rect 2238 -2268 2244 -2262
rect 2238 -2274 2244 -2268
rect 2238 -2280 2244 -2274
rect 2238 -2286 2244 -2280
rect 2238 -2292 2244 -2286
rect 2238 -2298 2244 -2292
rect 2238 -2364 2244 -2358
rect 2238 -2370 2244 -2364
rect 2238 -2376 2244 -2370
rect 2238 -2382 2244 -2376
rect 2238 -2388 2244 -2382
rect 2238 -2394 2244 -2388
rect 2238 -2400 2244 -2394
rect 2238 -2406 2244 -2400
rect 2238 -2412 2244 -2406
rect 2238 -2418 2244 -2412
rect 2238 -2424 2244 -2418
rect 2238 -2430 2244 -2424
rect 2238 -2436 2244 -2430
rect 2238 -2442 2244 -2436
rect 2238 -2448 2244 -2442
rect 2238 -2454 2244 -2448
rect 2238 -2460 2244 -2454
rect 2238 -2466 2244 -2460
rect 2238 -2526 2244 -2520
rect 2238 -2532 2244 -2526
rect 2238 -2538 2244 -2532
rect 2238 -2544 2244 -2538
rect 2238 -2550 2244 -2544
rect 2238 -2556 2244 -2550
rect 2238 -2562 2244 -2556
rect 2238 -2568 2244 -2562
rect 2238 -2574 2244 -2568
rect 2238 -2580 2244 -2574
rect 2238 -2586 2244 -2580
rect 2238 -2592 2244 -2586
rect 2238 -2598 2244 -2592
rect 2238 -2604 2244 -2598
rect 2238 -2610 2244 -2604
rect 2238 -2616 2244 -2610
rect 2238 -2622 2244 -2616
rect 2238 -2628 2244 -2622
rect 2238 -2634 2244 -2628
rect 2238 -2640 2244 -2634
rect 2238 -2646 2244 -2640
rect 2238 -2652 2244 -2646
rect 2238 -2658 2244 -2652
rect 2238 -2664 2244 -2658
rect 2238 -2670 2244 -2664
rect 2238 -2676 2244 -2670
rect 2238 -2682 2244 -2676
rect 2238 -2688 2244 -2682
rect 2238 -2694 2244 -2688
rect 2238 -2700 2244 -2694
rect 2238 -2706 2244 -2700
rect 2238 -2712 2244 -2706
rect 2238 -2718 2244 -2712
rect 2238 -2724 2244 -2718
rect 2238 -2730 2244 -2724
rect 2238 -2736 2244 -2730
rect 2238 -2742 2244 -2736
rect 2238 -2748 2244 -2742
rect 2238 -2754 2244 -2748
rect 2238 -2760 2244 -2754
rect 2238 -2766 2244 -2760
rect 2238 -2772 2244 -2766
rect 2238 -2778 2244 -2772
rect 2238 -2784 2244 -2778
rect 2238 -2790 2244 -2784
rect 2238 -2796 2244 -2790
rect 2238 -2802 2244 -2796
rect 2238 -2808 2244 -2802
rect 2238 -2814 2244 -2808
rect 2238 -2820 2244 -2814
rect 2238 -2826 2244 -2820
rect 2238 -2832 2244 -2826
rect 2238 -2838 2244 -2832
rect 2238 -2844 2244 -2838
rect 2238 -2850 2244 -2844
rect 2238 -2856 2244 -2850
rect 2238 -2862 2244 -2856
rect 2238 -2868 2244 -2862
rect 2238 -2874 2244 -2868
rect 2238 -2880 2244 -2874
rect 2238 -2886 2244 -2880
rect 2238 -2892 2244 -2886
rect 2238 -2898 2244 -2892
rect 2238 -2904 2244 -2898
rect 2238 -2910 2244 -2904
rect 2238 -2916 2244 -2910
rect 2238 -2922 2244 -2916
rect 2238 -2928 2244 -2922
rect 2238 -2934 2244 -2928
rect 2238 -2940 2244 -2934
rect 2238 -2946 2244 -2940
rect 2238 -2952 2244 -2946
rect 2238 -2958 2244 -2952
rect 2238 -2964 2244 -2958
rect 2238 -2970 2244 -2964
rect 2238 -2976 2244 -2970
rect 2238 -2982 2244 -2976
rect 2244 -144 2250 -138
rect 2244 -150 2250 -144
rect 2244 -156 2250 -150
rect 2244 -162 2250 -156
rect 2244 -168 2250 -162
rect 2244 -174 2250 -168
rect 2244 -180 2250 -174
rect 2244 -186 2250 -180
rect 2244 -192 2250 -186
rect 2244 -198 2250 -192
rect 2244 -204 2250 -198
rect 2244 -210 2250 -204
rect 2244 -216 2250 -210
rect 2244 -222 2250 -216
rect 2244 -228 2250 -222
rect 2244 -234 2250 -228
rect 2244 -240 2250 -234
rect 2244 -246 2250 -240
rect 2244 -252 2250 -246
rect 2244 -258 2250 -252
rect 2244 -264 2250 -258
rect 2244 -270 2250 -264
rect 2244 -276 2250 -270
rect 2244 -282 2250 -276
rect 2244 -288 2250 -282
rect 2244 -294 2250 -288
rect 2244 -300 2250 -294
rect 2244 -306 2250 -300
rect 2244 -312 2250 -306
rect 2244 -318 2250 -312
rect 2244 -324 2250 -318
rect 2244 -330 2250 -324
rect 2244 -336 2250 -330
rect 2244 -342 2250 -336
rect 2244 -348 2250 -342
rect 2244 -354 2250 -348
rect 2244 -360 2250 -354
rect 2244 -366 2250 -360
rect 2244 -372 2250 -366
rect 2244 -378 2250 -372
rect 2244 -384 2250 -378
rect 2244 -390 2250 -384
rect 2244 -396 2250 -390
rect 2244 -402 2250 -396
rect 2244 -408 2250 -402
rect 2244 -414 2250 -408
rect 2244 -420 2250 -414
rect 2244 -426 2250 -420
rect 2244 -432 2250 -426
rect 2244 -438 2250 -432
rect 2244 -444 2250 -438
rect 2244 -450 2250 -444
rect 2244 -456 2250 -450
rect 2244 -462 2250 -456
rect 2244 -468 2250 -462
rect 2244 -474 2250 -468
rect 2244 -480 2250 -474
rect 2244 -486 2250 -480
rect 2244 -492 2250 -486
rect 2244 -498 2250 -492
rect 2244 -504 2250 -498
rect 2244 -510 2250 -504
rect 2244 -516 2250 -510
rect 2244 -522 2250 -516
rect 2244 -528 2250 -522
rect 2244 -534 2250 -528
rect 2244 -540 2250 -534
rect 2244 -546 2250 -540
rect 2244 -552 2250 -546
rect 2244 -558 2250 -552
rect 2244 -564 2250 -558
rect 2244 -570 2250 -564
rect 2244 -576 2250 -570
rect 2244 -582 2250 -576
rect 2244 -588 2250 -582
rect 2244 -594 2250 -588
rect 2244 -600 2250 -594
rect 2244 -606 2250 -600
rect 2244 -612 2250 -606
rect 2244 -618 2250 -612
rect 2244 -624 2250 -618
rect 2244 -630 2250 -624
rect 2244 -636 2250 -630
rect 2244 -642 2250 -636
rect 2244 -648 2250 -642
rect 2244 -654 2250 -648
rect 2244 -660 2250 -654
rect 2244 -666 2250 -660
rect 2244 -672 2250 -666
rect 2244 -678 2250 -672
rect 2244 -684 2250 -678
rect 2244 -690 2250 -684
rect 2244 -696 2250 -690
rect 2244 -702 2250 -696
rect 2244 -708 2250 -702
rect 2244 -714 2250 -708
rect 2244 -720 2250 -714
rect 2244 -726 2250 -720
rect 2244 -732 2250 -726
rect 2244 -738 2250 -732
rect 2244 -744 2250 -738
rect 2244 -750 2250 -744
rect 2244 -756 2250 -750
rect 2244 -762 2250 -756
rect 2244 -768 2250 -762
rect 2244 -774 2250 -768
rect 2244 -780 2250 -774
rect 2244 -786 2250 -780
rect 2244 -792 2250 -786
rect 2244 -798 2250 -792
rect 2244 -804 2250 -798
rect 2244 -810 2250 -804
rect 2244 -816 2250 -810
rect 2244 -822 2250 -816
rect 2244 -828 2250 -822
rect 2244 -834 2250 -828
rect 2244 -840 2250 -834
rect 2244 -846 2250 -840
rect 2244 -852 2250 -846
rect 2244 -858 2250 -852
rect 2244 -864 2250 -858
rect 2244 -870 2250 -864
rect 2244 -876 2250 -870
rect 2244 -882 2250 -876
rect 2244 -888 2250 -882
rect 2244 -894 2250 -888
rect 2244 -900 2250 -894
rect 2244 -906 2250 -900
rect 2244 -912 2250 -906
rect 2244 -918 2250 -912
rect 2244 -924 2250 -918
rect 2244 -930 2250 -924
rect 2244 -936 2250 -930
rect 2244 -942 2250 -936
rect 2244 -948 2250 -942
rect 2244 -954 2250 -948
rect 2244 -960 2250 -954
rect 2244 -966 2250 -960
rect 2244 -972 2250 -966
rect 2244 -978 2250 -972
rect 2244 -984 2250 -978
rect 2244 -990 2250 -984
rect 2244 -996 2250 -990
rect 2244 -1002 2250 -996
rect 2244 -1008 2250 -1002
rect 2244 -1014 2250 -1008
rect 2244 -1020 2250 -1014
rect 2244 -1026 2250 -1020
rect 2244 -1032 2250 -1026
rect 2244 -1038 2250 -1032
rect 2244 -1044 2250 -1038
rect 2244 -1050 2250 -1044
rect 2244 -1056 2250 -1050
rect 2244 -1062 2250 -1056
rect 2244 -1068 2250 -1062
rect 2244 -1074 2250 -1068
rect 2244 -1080 2250 -1074
rect 2244 -1086 2250 -1080
rect 2244 -1092 2250 -1086
rect 2244 -1098 2250 -1092
rect 2244 -1104 2250 -1098
rect 2244 -1110 2250 -1104
rect 2244 -1116 2250 -1110
rect 2244 -1122 2250 -1116
rect 2244 -1128 2250 -1122
rect 2244 -1134 2250 -1128
rect 2244 -1518 2250 -1512
rect 2244 -1524 2250 -1518
rect 2244 -1530 2250 -1524
rect 2244 -1536 2250 -1530
rect 2244 -1542 2250 -1536
rect 2244 -1548 2250 -1542
rect 2244 -1554 2250 -1548
rect 2244 -1560 2250 -1554
rect 2244 -1566 2250 -1560
rect 2244 -1572 2250 -1566
rect 2244 -1578 2250 -1572
rect 2244 -1584 2250 -1578
rect 2244 -1590 2250 -1584
rect 2244 -1596 2250 -1590
rect 2244 -1602 2250 -1596
rect 2244 -1608 2250 -1602
rect 2244 -1614 2250 -1608
rect 2244 -1620 2250 -1614
rect 2244 -1626 2250 -1620
rect 2244 -1632 2250 -1626
rect 2244 -1638 2250 -1632
rect 2244 -1644 2250 -1638
rect 2244 -1650 2250 -1644
rect 2244 -1656 2250 -1650
rect 2244 -1662 2250 -1656
rect 2244 -1668 2250 -1662
rect 2244 -1674 2250 -1668
rect 2244 -1680 2250 -1674
rect 2244 -1686 2250 -1680
rect 2244 -1692 2250 -1686
rect 2244 -1698 2250 -1692
rect 2244 -1704 2250 -1698
rect 2244 -1710 2250 -1704
rect 2244 -1716 2250 -1710
rect 2244 -1722 2250 -1716
rect 2244 -1728 2250 -1722
rect 2244 -1734 2250 -1728
rect 2244 -1740 2250 -1734
rect 2244 -1746 2250 -1740
rect 2244 -1752 2250 -1746
rect 2244 -1758 2250 -1752
rect 2244 -1764 2250 -1758
rect 2244 -1770 2250 -1764
rect 2244 -1776 2250 -1770
rect 2244 -1782 2250 -1776
rect 2244 -1788 2250 -1782
rect 2244 -1794 2250 -1788
rect 2244 -1800 2250 -1794
rect 2244 -1806 2250 -1800
rect 2244 -1812 2250 -1806
rect 2244 -1818 2250 -1812
rect 2244 -1824 2250 -1818
rect 2244 -1830 2250 -1824
rect 2244 -1836 2250 -1830
rect 2244 -1842 2250 -1836
rect 2244 -1848 2250 -1842
rect 2244 -1854 2250 -1848
rect 2244 -1860 2250 -1854
rect 2244 -1866 2250 -1860
rect 2244 -1872 2250 -1866
rect 2244 -1878 2250 -1872
rect 2244 -1884 2250 -1878
rect 2244 -1890 2250 -1884
rect 2244 -1896 2250 -1890
rect 2244 -1902 2250 -1896
rect 2244 -1908 2250 -1902
rect 2244 -1914 2250 -1908
rect 2244 -1920 2250 -1914
rect 2244 -1926 2250 -1920
rect 2244 -1932 2250 -1926
rect 2244 -1938 2250 -1932
rect 2244 -1944 2250 -1938
rect 2244 -1950 2250 -1944
rect 2244 -1956 2250 -1950
rect 2244 -1962 2250 -1956
rect 2244 -1968 2250 -1962
rect 2244 -1974 2250 -1968
rect 2244 -1980 2250 -1974
rect 2244 -1986 2250 -1980
rect 2244 -1992 2250 -1986
rect 2244 -1998 2250 -1992
rect 2244 -2004 2250 -1998
rect 2244 -2010 2250 -2004
rect 2244 -2016 2250 -2010
rect 2244 -2022 2250 -2016
rect 2244 -2028 2250 -2022
rect 2244 -2034 2250 -2028
rect 2244 -2040 2250 -2034
rect 2244 -2046 2250 -2040
rect 2244 -2052 2250 -2046
rect 2244 -2058 2250 -2052
rect 2244 -2064 2250 -2058
rect 2244 -2070 2250 -2064
rect 2244 -2076 2250 -2070
rect 2244 -2082 2250 -2076
rect 2244 -2088 2250 -2082
rect 2244 -2094 2250 -2088
rect 2244 -2100 2250 -2094
rect 2244 -2106 2250 -2100
rect 2244 -2112 2250 -2106
rect 2244 -2118 2250 -2112
rect 2244 -2124 2250 -2118
rect 2244 -2130 2250 -2124
rect 2244 -2136 2250 -2130
rect 2244 -2142 2250 -2136
rect 2244 -2148 2250 -2142
rect 2244 -2154 2250 -2148
rect 2244 -2160 2250 -2154
rect 2244 -2166 2250 -2160
rect 2244 -2172 2250 -2166
rect 2244 -2178 2250 -2172
rect 2244 -2184 2250 -2178
rect 2244 -2190 2250 -2184
rect 2244 -2196 2250 -2190
rect 2244 -2202 2250 -2196
rect 2244 -2208 2250 -2202
rect 2244 -2214 2250 -2208
rect 2244 -2220 2250 -2214
rect 2244 -2226 2250 -2220
rect 2244 -2232 2250 -2226
rect 2244 -2238 2250 -2232
rect 2244 -2244 2250 -2238
rect 2244 -2250 2250 -2244
rect 2244 -2256 2250 -2250
rect 2244 -2262 2250 -2256
rect 2244 -2268 2250 -2262
rect 2244 -2274 2250 -2268
rect 2244 -2280 2250 -2274
rect 2244 -2286 2250 -2280
rect 2244 -2292 2250 -2286
rect 2244 -2358 2250 -2352
rect 2244 -2364 2250 -2358
rect 2244 -2370 2250 -2364
rect 2244 -2376 2250 -2370
rect 2244 -2382 2250 -2376
rect 2244 -2388 2250 -2382
rect 2244 -2394 2250 -2388
rect 2244 -2400 2250 -2394
rect 2244 -2406 2250 -2400
rect 2244 -2412 2250 -2406
rect 2244 -2418 2250 -2412
rect 2244 -2424 2250 -2418
rect 2244 -2430 2250 -2424
rect 2244 -2436 2250 -2430
rect 2244 -2442 2250 -2436
rect 2244 -2448 2250 -2442
rect 2244 -2454 2250 -2448
rect 2244 -2460 2250 -2454
rect 2244 -2466 2250 -2460
rect 2244 -2526 2250 -2520
rect 2244 -2532 2250 -2526
rect 2244 -2538 2250 -2532
rect 2244 -2544 2250 -2538
rect 2244 -2550 2250 -2544
rect 2244 -2556 2250 -2550
rect 2244 -2562 2250 -2556
rect 2244 -2568 2250 -2562
rect 2244 -2574 2250 -2568
rect 2244 -2580 2250 -2574
rect 2244 -2586 2250 -2580
rect 2244 -2592 2250 -2586
rect 2244 -2598 2250 -2592
rect 2244 -2604 2250 -2598
rect 2244 -2610 2250 -2604
rect 2244 -2616 2250 -2610
rect 2244 -2622 2250 -2616
rect 2244 -2628 2250 -2622
rect 2244 -2634 2250 -2628
rect 2244 -2640 2250 -2634
rect 2244 -2646 2250 -2640
rect 2244 -2652 2250 -2646
rect 2244 -2658 2250 -2652
rect 2244 -2664 2250 -2658
rect 2244 -2670 2250 -2664
rect 2244 -2676 2250 -2670
rect 2244 -2682 2250 -2676
rect 2244 -2688 2250 -2682
rect 2244 -2694 2250 -2688
rect 2244 -2700 2250 -2694
rect 2244 -2706 2250 -2700
rect 2244 -2712 2250 -2706
rect 2244 -2718 2250 -2712
rect 2244 -2724 2250 -2718
rect 2244 -2730 2250 -2724
rect 2244 -2736 2250 -2730
rect 2244 -2742 2250 -2736
rect 2244 -2748 2250 -2742
rect 2244 -2754 2250 -2748
rect 2244 -2760 2250 -2754
rect 2244 -2766 2250 -2760
rect 2244 -2772 2250 -2766
rect 2244 -2778 2250 -2772
rect 2244 -2784 2250 -2778
rect 2244 -2790 2250 -2784
rect 2244 -2796 2250 -2790
rect 2244 -2802 2250 -2796
rect 2244 -2808 2250 -2802
rect 2244 -2814 2250 -2808
rect 2244 -2820 2250 -2814
rect 2244 -2826 2250 -2820
rect 2244 -2832 2250 -2826
rect 2244 -2838 2250 -2832
rect 2244 -2844 2250 -2838
rect 2244 -2850 2250 -2844
rect 2244 -2856 2250 -2850
rect 2244 -2862 2250 -2856
rect 2244 -2868 2250 -2862
rect 2244 -2874 2250 -2868
rect 2244 -2880 2250 -2874
rect 2244 -2886 2250 -2880
rect 2244 -2892 2250 -2886
rect 2244 -2898 2250 -2892
rect 2244 -2904 2250 -2898
rect 2244 -2910 2250 -2904
rect 2244 -2916 2250 -2910
rect 2244 -2922 2250 -2916
rect 2244 -2928 2250 -2922
rect 2244 -2934 2250 -2928
rect 2244 -2940 2250 -2934
rect 2244 -2946 2250 -2940
rect 2244 -2952 2250 -2946
rect 2244 -2958 2250 -2952
rect 2244 -2964 2250 -2958
rect 2244 -2970 2250 -2964
rect 2244 -2976 2250 -2970
rect 2244 -2982 2250 -2976
rect 2250 -138 2256 -132
rect 2250 -144 2256 -138
rect 2250 -150 2256 -144
rect 2250 -156 2256 -150
rect 2250 -162 2256 -156
rect 2250 -168 2256 -162
rect 2250 -174 2256 -168
rect 2250 -180 2256 -174
rect 2250 -186 2256 -180
rect 2250 -192 2256 -186
rect 2250 -198 2256 -192
rect 2250 -204 2256 -198
rect 2250 -210 2256 -204
rect 2250 -216 2256 -210
rect 2250 -222 2256 -216
rect 2250 -228 2256 -222
rect 2250 -234 2256 -228
rect 2250 -240 2256 -234
rect 2250 -246 2256 -240
rect 2250 -252 2256 -246
rect 2250 -258 2256 -252
rect 2250 -264 2256 -258
rect 2250 -270 2256 -264
rect 2250 -276 2256 -270
rect 2250 -282 2256 -276
rect 2250 -288 2256 -282
rect 2250 -294 2256 -288
rect 2250 -300 2256 -294
rect 2250 -306 2256 -300
rect 2250 -312 2256 -306
rect 2250 -318 2256 -312
rect 2250 -324 2256 -318
rect 2250 -330 2256 -324
rect 2250 -336 2256 -330
rect 2250 -342 2256 -336
rect 2250 -348 2256 -342
rect 2250 -354 2256 -348
rect 2250 -360 2256 -354
rect 2250 -366 2256 -360
rect 2250 -372 2256 -366
rect 2250 -378 2256 -372
rect 2250 -384 2256 -378
rect 2250 -390 2256 -384
rect 2250 -396 2256 -390
rect 2250 -402 2256 -396
rect 2250 -408 2256 -402
rect 2250 -414 2256 -408
rect 2250 -420 2256 -414
rect 2250 -426 2256 -420
rect 2250 -432 2256 -426
rect 2250 -438 2256 -432
rect 2250 -444 2256 -438
rect 2250 -450 2256 -444
rect 2250 -456 2256 -450
rect 2250 -462 2256 -456
rect 2250 -468 2256 -462
rect 2250 -474 2256 -468
rect 2250 -480 2256 -474
rect 2250 -486 2256 -480
rect 2250 -492 2256 -486
rect 2250 -498 2256 -492
rect 2250 -504 2256 -498
rect 2250 -510 2256 -504
rect 2250 -516 2256 -510
rect 2250 -522 2256 -516
rect 2250 -528 2256 -522
rect 2250 -534 2256 -528
rect 2250 -540 2256 -534
rect 2250 -546 2256 -540
rect 2250 -552 2256 -546
rect 2250 -558 2256 -552
rect 2250 -564 2256 -558
rect 2250 -570 2256 -564
rect 2250 -576 2256 -570
rect 2250 -582 2256 -576
rect 2250 -588 2256 -582
rect 2250 -594 2256 -588
rect 2250 -600 2256 -594
rect 2250 -606 2256 -600
rect 2250 -612 2256 -606
rect 2250 -618 2256 -612
rect 2250 -624 2256 -618
rect 2250 -630 2256 -624
rect 2250 -636 2256 -630
rect 2250 -642 2256 -636
rect 2250 -648 2256 -642
rect 2250 -654 2256 -648
rect 2250 -660 2256 -654
rect 2250 -666 2256 -660
rect 2250 -672 2256 -666
rect 2250 -678 2256 -672
rect 2250 -684 2256 -678
rect 2250 -690 2256 -684
rect 2250 -696 2256 -690
rect 2250 -702 2256 -696
rect 2250 -708 2256 -702
rect 2250 -714 2256 -708
rect 2250 -720 2256 -714
rect 2250 -726 2256 -720
rect 2250 -732 2256 -726
rect 2250 -738 2256 -732
rect 2250 -744 2256 -738
rect 2250 -750 2256 -744
rect 2250 -756 2256 -750
rect 2250 -762 2256 -756
rect 2250 -768 2256 -762
rect 2250 -774 2256 -768
rect 2250 -780 2256 -774
rect 2250 -786 2256 -780
rect 2250 -792 2256 -786
rect 2250 -798 2256 -792
rect 2250 -804 2256 -798
rect 2250 -810 2256 -804
rect 2250 -816 2256 -810
rect 2250 -822 2256 -816
rect 2250 -828 2256 -822
rect 2250 -834 2256 -828
rect 2250 -840 2256 -834
rect 2250 -846 2256 -840
rect 2250 -852 2256 -846
rect 2250 -858 2256 -852
rect 2250 -864 2256 -858
rect 2250 -870 2256 -864
rect 2250 -876 2256 -870
rect 2250 -882 2256 -876
rect 2250 -888 2256 -882
rect 2250 -894 2256 -888
rect 2250 -900 2256 -894
rect 2250 -906 2256 -900
rect 2250 -912 2256 -906
rect 2250 -918 2256 -912
rect 2250 -924 2256 -918
rect 2250 -930 2256 -924
rect 2250 -936 2256 -930
rect 2250 -942 2256 -936
rect 2250 -948 2256 -942
rect 2250 -954 2256 -948
rect 2250 -960 2256 -954
rect 2250 -966 2256 -960
rect 2250 -972 2256 -966
rect 2250 -978 2256 -972
rect 2250 -984 2256 -978
rect 2250 -990 2256 -984
rect 2250 -996 2256 -990
rect 2250 -1002 2256 -996
rect 2250 -1008 2256 -1002
rect 2250 -1014 2256 -1008
rect 2250 -1020 2256 -1014
rect 2250 -1026 2256 -1020
rect 2250 -1032 2256 -1026
rect 2250 -1038 2256 -1032
rect 2250 -1044 2256 -1038
rect 2250 -1050 2256 -1044
rect 2250 -1056 2256 -1050
rect 2250 -1062 2256 -1056
rect 2250 -1068 2256 -1062
rect 2250 -1074 2256 -1068
rect 2250 -1080 2256 -1074
rect 2250 -1086 2256 -1080
rect 2250 -1092 2256 -1086
rect 2250 -1098 2256 -1092
rect 2250 -1104 2256 -1098
rect 2250 -1110 2256 -1104
rect 2250 -1116 2256 -1110
rect 2250 -1122 2256 -1116
rect 2250 -1512 2256 -1506
rect 2250 -1518 2256 -1512
rect 2250 -1524 2256 -1518
rect 2250 -1530 2256 -1524
rect 2250 -1536 2256 -1530
rect 2250 -1542 2256 -1536
rect 2250 -1548 2256 -1542
rect 2250 -1554 2256 -1548
rect 2250 -1560 2256 -1554
rect 2250 -1566 2256 -1560
rect 2250 -1572 2256 -1566
rect 2250 -1578 2256 -1572
rect 2250 -1584 2256 -1578
rect 2250 -1590 2256 -1584
rect 2250 -1596 2256 -1590
rect 2250 -1602 2256 -1596
rect 2250 -1608 2256 -1602
rect 2250 -1614 2256 -1608
rect 2250 -1620 2256 -1614
rect 2250 -1626 2256 -1620
rect 2250 -1632 2256 -1626
rect 2250 -1638 2256 -1632
rect 2250 -1644 2256 -1638
rect 2250 -1650 2256 -1644
rect 2250 -1656 2256 -1650
rect 2250 -1662 2256 -1656
rect 2250 -1668 2256 -1662
rect 2250 -1674 2256 -1668
rect 2250 -1680 2256 -1674
rect 2250 -1686 2256 -1680
rect 2250 -1692 2256 -1686
rect 2250 -1698 2256 -1692
rect 2250 -1704 2256 -1698
rect 2250 -1710 2256 -1704
rect 2250 -1716 2256 -1710
rect 2250 -1722 2256 -1716
rect 2250 -1728 2256 -1722
rect 2250 -1734 2256 -1728
rect 2250 -1740 2256 -1734
rect 2250 -1746 2256 -1740
rect 2250 -1752 2256 -1746
rect 2250 -1758 2256 -1752
rect 2250 -1764 2256 -1758
rect 2250 -1770 2256 -1764
rect 2250 -1776 2256 -1770
rect 2250 -1782 2256 -1776
rect 2250 -1788 2256 -1782
rect 2250 -1794 2256 -1788
rect 2250 -1800 2256 -1794
rect 2250 -1806 2256 -1800
rect 2250 -1812 2256 -1806
rect 2250 -1818 2256 -1812
rect 2250 -1824 2256 -1818
rect 2250 -1830 2256 -1824
rect 2250 -1836 2256 -1830
rect 2250 -1842 2256 -1836
rect 2250 -1848 2256 -1842
rect 2250 -1854 2256 -1848
rect 2250 -1860 2256 -1854
rect 2250 -1866 2256 -1860
rect 2250 -1872 2256 -1866
rect 2250 -1878 2256 -1872
rect 2250 -1884 2256 -1878
rect 2250 -1890 2256 -1884
rect 2250 -1896 2256 -1890
rect 2250 -1902 2256 -1896
rect 2250 -1908 2256 -1902
rect 2250 -1914 2256 -1908
rect 2250 -1920 2256 -1914
rect 2250 -1926 2256 -1920
rect 2250 -1932 2256 -1926
rect 2250 -1938 2256 -1932
rect 2250 -1944 2256 -1938
rect 2250 -1950 2256 -1944
rect 2250 -1956 2256 -1950
rect 2250 -1962 2256 -1956
rect 2250 -1968 2256 -1962
rect 2250 -1974 2256 -1968
rect 2250 -1980 2256 -1974
rect 2250 -1986 2256 -1980
rect 2250 -1992 2256 -1986
rect 2250 -1998 2256 -1992
rect 2250 -2004 2256 -1998
rect 2250 -2010 2256 -2004
rect 2250 -2016 2256 -2010
rect 2250 -2022 2256 -2016
rect 2250 -2028 2256 -2022
rect 2250 -2034 2256 -2028
rect 2250 -2040 2256 -2034
rect 2250 -2046 2256 -2040
rect 2250 -2052 2256 -2046
rect 2250 -2058 2256 -2052
rect 2250 -2064 2256 -2058
rect 2250 -2070 2256 -2064
rect 2250 -2076 2256 -2070
rect 2250 -2082 2256 -2076
rect 2250 -2088 2256 -2082
rect 2250 -2094 2256 -2088
rect 2250 -2100 2256 -2094
rect 2250 -2106 2256 -2100
rect 2250 -2112 2256 -2106
rect 2250 -2118 2256 -2112
rect 2250 -2124 2256 -2118
rect 2250 -2130 2256 -2124
rect 2250 -2136 2256 -2130
rect 2250 -2142 2256 -2136
rect 2250 -2148 2256 -2142
rect 2250 -2154 2256 -2148
rect 2250 -2160 2256 -2154
rect 2250 -2166 2256 -2160
rect 2250 -2172 2256 -2166
rect 2250 -2178 2256 -2172
rect 2250 -2184 2256 -2178
rect 2250 -2190 2256 -2184
rect 2250 -2196 2256 -2190
rect 2250 -2202 2256 -2196
rect 2250 -2208 2256 -2202
rect 2250 -2214 2256 -2208
rect 2250 -2220 2256 -2214
rect 2250 -2226 2256 -2220
rect 2250 -2232 2256 -2226
rect 2250 -2238 2256 -2232
rect 2250 -2244 2256 -2238
rect 2250 -2250 2256 -2244
rect 2250 -2256 2256 -2250
rect 2250 -2262 2256 -2256
rect 2250 -2268 2256 -2262
rect 2250 -2274 2256 -2268
rect 2250 -2280 2256 -2274
rect 2250 -2352 2256 -2346
rect 2250 -2358 2256 -2352
rect 2250 -2364 2256 -2358
rect 2250 -2370 2256 -2364
rect 2250 -2376 2256 -2370
rect 2250 -2382 2256 -2376
rect 2250 -2388 2256 -2382
rect 2250 -2394 2256 -2388
rect 2250 -2400 2256 -2394
rect 2250 -2406 2256 -2400
rect 2250 -2412 2256 -2406
rect 2250 -2418 2256 -2412
rect 2250 -2424 2256 -2418
rect 2250 -2430 2256 -2424
rect 2250 -2436 2256 -2430
rect 2250 -2442 2256 -2436
rect 2250 -2448 2256 -2442
rect 2250 -2454 2256 -2448
rect 2250 -2460 2256 -2454
rect 2250 -2520 2256 -2514
rect 2250 -2526 2256 -2520
rect 2250 -2532 2256 -2526
rect 2250 -2538 2256 -2532
rect 2250 -2544 2256 -2538
rect 2250 -2550 2256 -2544
rect 2250 -2556 2256 -2550
rect 2250 -2562 2256 -2556
rect 2250 -2568 2256 -2562
rect 2250 -2574 2256 -2568
rect 2250 -2580 2256 -2574
rect 2250 -2586 2256 -2580
rect 2250 -2592 2256 -2586
rect 2250 -2598 2256 -2592
rect 2250 -2604 2256 -2598
rect 2250 -2610 2256 -2604
rect 2250 -2616 2256 -2610
rect 2250 -2622 2256 -2616
rect 2250 -2628 2256 -2622
rect 2250 -2634 2256 -2628
rect 2250 -2640 2256 -2634
rect 2250 -2646 2256 -2640
rect 2250 -2652 2256 -2646
rect 2250 -2658 2256 -2652
rect 2250 -2664 2256 -2658
rect 2250 -2670 2256 -2664
rect 2250 -2676 2256 -2670
rect 2250 -2682 2256 -2676
rect 2250 -2688 2256 -2682
rect 2250 -2694 2256 -2688
rect 2250 -2700 2256 -2694
rect 2250 -2706 2256 -2700
rect 2250 -2712 2256 -2706
rect 2250 -2718 2256 -2712
rect 2250 -2724 2256 -2718
rect 2250 -2730 2256 -2724
rect 2250 -2736 2256 -2730
rect 2250 -2742 2256 -2736
rect 2250 -2748 2256 -2742
rect 2250 -2754 2256 -2748
rect 2250 -2760 2256 -2754
rect 2250 -2766 2256 -2760
rect 2250 -2772 2256 -2766
rect 2250 -2778 2256 -2772
rect 2250 -2784 2256 -2778
rect 2250 -2790 2256 -2784
rect 2250 -2796 2256 -2790
rect 2250 -2802 2256 -2796
rect 2250 -2808 2256 -2802
rect 2250 -2814 2256 -2808
rect 2250 -2820 2256 -2814
rect 2250 -2826 2256 -2820
rect 2250 -2832 2256 -2826
rect 2250 -2838 2256 -2832
rect 2250 -2844 2256 -2838
rect 2250 -2850 2256 -2844
rect 2250 -2856 2256 -2850
rect 2250 -2862 2256 -2856
rect 2250 -2868 2256 -2862
rect 2250 -2874 2256 -2868
rect 2250 -2880 2256 -2874
rect 2250 -2886 2256 -2880
rect 2250 -2892 2256 -2886
rect 2250 -2898 2256 -2892
rect 2250 -2904 2256 -2898
rect 2250 -2910 2256 -2904
rect 2250 -2916 2256 -2910
rect 2250 -2922 2256 -2916
rect 2250 -2928 2256 -2922
rect 2250 -2934 2256 -2928
rect 2250 -2940 2256 -2934
rect 2250 -2946 2256 -2940
rect 2250 -2952 2256 -2946
rect 2250 -2958 2256 -2952
rect 2250 -2964 2256 -2958
rect 2250 -2970 2256 -2964
rect 2250 -2976 2256 -2970
rect 2256 -126 2262 -120
rect 2256 -132 2262 -126
rect 2256 -138 2262 -132
rect 2256 -144 2262 -138
rect 2256 -150 2262 -144
rect 2256 -156 2262 -150
rect 2256 -162 2262 -156
rect 2256 -168 2262 -162
rect 2256 -174 2262 -168
rect 2256 -180 2262 -174
rect 2256 -186 2262 -180
rect 2256 -192 2262 -186
rect 2256 -198 2262 -192
rect 2256 -204 2262 -198
rect 2256 -210 2262 -204
rect 2256 -216 2262 -210
rect 2256 -222 2262 -216
rect 2256 -228 2262 -222
rect 2256 -234 2262 -228
rect 2256 -240 2262 -234
rect 2256 -246 2262 -240
rect 2256 -252 2262 -246
rect 2256 -258 2262 -252
rect 2256 -264 2262 -258
rect 2256 -270 2262 -264
rect 2256 -276 2262 -270
rect 2256 -282 2262 -276
rect 2256 -288 2262 -282
rect 2256 -294 2262 -288
rect 2256 -300 2262 -294
rect 2256 -306 2262 -300
rect 2256 -312 2262 -306
rect 2256 -318 2262 -312
rect 2256 -324 2262 -318
rect 2256 -330 2262 -324
rect 2256 -336 2262 -330
rect 2256 -342 2262 -336
rect 2256 -348 2262 -342
rect 2256 -354 2262 -348
rect 2256 -360 2262 -354
rect 2256 -366 2262 -360
rect 2256 -372 2262 -366
rect 2256 -378 2262 -372
rect 2256 -384 2262 -378
rect 2256 -390 2262 -384
rect 2256 -396 2262 -390
rect 2256 -402 2262 -396
rect 2256 -408 2262 -402
rect 2256 -414 2262 -408
rect 2256 -420 2262 -414
rect 2256 -426 2262 -420
rect 2256 -432 2262 -426
rect 2256 -438 2262 -432
rect 2256 -444 2262 -438
rect 2256 -450 2262 -444
rect 2256 -456 2262 -450
rect 2256 -462 2262 -456
rect 2256 -468 2262 -462
rect 2256 -474 2262 -468
rect 2256 -480 2262 -474
rect 2256 -486 2262 -480
rect 2256 -492 2262 -486
rect 2256 -498 2262 -492
rect 2256 -504 2262 -498
rect 2256 -510 2262 -504
rect 2256 -516 2262 -510
rect 2256 -522 2262 -516
rect 2256 -528 2262 -522
rect 2256 -534 2262 -528
rect 2256 -540 2262 -534
rect 2256 -546 2262 -540
rect 2256 -552 2262 -546
rect 2256 -558 2262 -552
rect 2256 -564 2262 -558
rect 2256 -570 2262 -564
rect 2256 -576 2262 -570
rect 2256 -582 2262 -576
rect 2256 -588 2262 -582
rect 2256 -594 2262 -588
rect 2256 -600 2262 -594
rect 2256 -606 2262 -600
rect 2256 -612 2262 -606
rect 2256 -618 2262 -612
rect 2256 -624 2262 -618
rect 2256 -630 2262 -624
rect 2256 -636 2262 -630
rect 2256 -642 2262 -636
rect 2256 -648 2262 -642
rect 2256 -654 2262 -648
rect 2256 -660 2262 -654
rect 2256 -666 2262 -660
rect 2256 -672 2262 -666
rect 2256 -678 2262 -672
rect 2256 -684 2262 -678
rect 2256 -690 2262 -684
rect 2256 -696 2262 -690
rect 2256 -702 2262 -696
rect 2256 -708 2262 -702
rect 2256 -714 2262 -708
rect 2256 -720 2262 -714
rect 2256 -726 2262 -720
rect 2256 -732 2262 -726
rect 2256 -738 2262 -732
rect 2256 -744 2262 -738
rect 2256 -750 2262 -744
rect 2256 -756 2262 -750
rect 2256 -762 2262 -756
rect 2256 -768 2262 -762
rect 2256 -774 2262 -768
rect 2256 -780 2262 -774
rect 2256 -786 2262 -780
rect 2256 -792 2262 -786
rect 2256 -798 2262 -792
rect 2256 -804 2262 -798
rect 2256 -810 2262 -804
rect 2256 -816 2262 -810
rect 2256 -822 2262 -816
rect 2256 -828 2262 -822
rect 2256 -834 2262 -828
rect 2256 -840 2262 -834
rect 2256 -846 2262 -840
rect 2256 -852 2262 -846
rect 2256 -858 2262 -852
rect 2256 -864 2262 -858
rect 2256 -870 2262 -864
rect 2256 -876 2262 -870
rect 2256 -882 2262 -876
rect 2256 -888 2262 -882
rect 2256 -894 2262 -888
rect 2256 -900 2262 -894
rect 2256 -906 2262 -900
rect 2256 -912 2262 -906
rect 2256 -918 2262 -912
rect 2256 -924 2262 -918
rect 2256 -930 2262 -924
rect 2256 -936 2262 -930
rect 2256 -942 2262 -936
rect 2256 -948 2262 -942
rect 2256 -954 2262 -948
rect 2256 -960 2262 -954
rect 2256 -966 2262 -960
rect 2256 -972 2262 -966
rect 2256 -978 2262 -972
rect 2256 -984 2262 -978
rect 2256 -990 2262 -984
rect 2256 -996 2262 -990
rect 2256 -1002 2262 -996
rect 2256 -1008 2262 -1002
rect 2256 -1014 2262 -1008
rect 2256 -1020 2262 -1014
rect 2256 -1026 2262 -1020
rect 2256 -1032 2262 -1026
rect 2256 -1038 2262 -1032
rect 2256 -1044 2262 -1038
rect 2256 -1050 2262 -1044
rect 2256 -1056 2262 -1050
rect 2256 -1062 2262 -1056
rect 2256 -1068 2262 -1062
rect 2256 -1074 2262 -1068
rect 2256 -1080 2262 -1074
rect 2256 -1086 2262 -1080
rect 2256 -1092 2262 -1086
rect 2256 -1098 2262 -1092
rect 2256 -1104 2262 -1098
rect 2256 -1506 2262 -1500
rect 2256 -1512 2262 -1506
rect 2256 -1518 2262 -1512
rect 2256 -1524 2262 -1518
rect 2256 -1530 2262 -1524
rect 2256 -1536 2262 -1530
rect 2256 -1542 2262 -1536
rect 2256 -1548 2262 -1542
rect 2256 -1554 2262 -1548
rect 2256 -1560 2262 -1554
rect 2256 -1566 2262 -1560
rect 2256 -1572 2262 -1566
rect 2256 -1578 2262 -1572
rect 2256 -1584 2262 -1578
rect 2256 -1590 2262 -1584
rect 2256 -1596 2262 -1590
rect 2256 -1602 2262 -1596
rect 2256 -1608 2262 -1602
rect 2256 -1614 2262 -1608
rect 2256 -1620 2262 -1614
rect 2256 -1626 2262 -1620
rect 2256 -1632 2262 -1626
rect 2256 -1638 2262 -1632
rect 2256 -1644 2262 -1638
rect 2256 -1650 2262 -1644
rect 2256 -1656 2262 -1650
rect 2256 -1662 2262 -1656
rect 2256 -1668 2262 -1662
rect 2256 -1674 2262 -1668
rect 2256 -1680 2262 -1674
rect 2256 -1686 2262 -1680
rect 2256 -1692 2262 -1686
rect 2256 -1698 2262 -1692
rect 2256 -1704 2262 -1698
rect 2256 -1710 2262 -1704
rect 2256 -1716 2262 -1710
rect 2256 -1722 2262 -1716
rect 2256 -1728 2262 -1722
rect 2256 -1734 2262 -1728
rect 2256 -1740 2262 -1734
rect 2256 -1746 2262 -1740
rect 2256 -1752 2262 -1746
rect 2256 -1758 2262 -1752
rect 2256 -1764 2262 -1758
rect 2256 -1770 2262 -1764
rect 2256 -1776 2262 -1770
rect 2256 -1782 2262 -1776
rect 2256 -1788 2262 -1782
rect 2256 -1794 2262 -1788
rect 2256 -1800 2262 -1794
rect 2256 -1806 2262 -1800
rect 2256 -1812 2262 -1806
rect 2256 -1818 2262 -1812
rect 2256 -1824 2262 -1818
rect 2256 -1830 2262 -1824
rect 2256 -1836 2262 -1830
rect 2256 -1842 2262 -1836
rect 2256 -1848 2262 -1842
rect 2256 -1854 2262 -1848
rect 2256 -1860 2262 -1854
rect 2256 -1866 2262 -1860
rect 2256 -1872 2262 -1866
rect 2256 -1878 2262 -1872
rect 2256 -1884 2262 -1878
rect 2256 -1890 2262 -1884
rect 2256 -1896 2262 -1890
rect 2256 -1902 2262 -1896
rect 2256 -1908 2262 -1902
rect 2256 -1914 2262 -1908
rect 2256 -1920 2262 -1914
rect 2256 -1926 2262 -1920
rect 2256 -1932 2262 -1926
rect 2256 -1938 2262 -1932
rect 2256 -1944 2262 -1938
rect 2256 -1950 2262 -1944
rect 2256 -1956 2262 -1950
rect 2256 -1962 2262 -1956
rect 2256 -1968 2262 -1962
rect 2256 -1974 2262 -1968
rect 2256 -1980 2262 -1974
rect 2256 -1986 2262 -1980
rect 2256 -1992 2262 -1986
rect 2256 -1998 2262 -1992
rect 2256 -2004 2262 -1998
rect 2256 -2010 2262 -2004
rect 2256 -2016 2262 -2010
rect 2256 -2022 2262 -2016
rect 2256 -2028 2262 -2022
rect 2256 -2034 2262 -2028
rect 2256 -2040 2262 -2034
rect 2256 -2046 2262 -2040
rect 2256 -2052 2262 -2046
rect 2256 -2058 2262 -2052
rect 2256 -2064 2262 -2058
rect 2256 -2070 2262 -2064
rect 2256 -2076 2262 -2070
rect 2256 -2082 2262 -2076
rect 2256 -2088 2262 -2082
rect 2256 -2094 2262 -2088
rect 2256 -2100 2262 -2094
rect 2256 -2106 2262 -2100
rect 2256 -2112 2262 -2106
rect 2256 -2118 2262 -2112
rect 2256 -2124 2262 -2118
rect 2256 -2130 2262 -2124
rect 2256 -2136 2262 -2130
rect 2256 -2142 2262 -2136
rect 2256 -2148 2262 -2142
rect 2256 -2154 2262 -2148
rect 2256 -2160 2262 -2154
rect 2256 -2166 2262 -2160
rect 2256 -2172 2262 -2166
rect 2256 -2178 2262 -2172
rect 2256 -2184 2262 -2178
rect 2256 -2190 2262 -2184
rect 2256 -2196 2262 -2190
rect 2256 -2202 2262 -2196
rect 2256 -2208 2262 -2202
rect 2256 -2214 2262 -2208
rect 2256 -2220 2262 -2214
rect 2256 -2226 2262 -2220
rect 2256 -2232 2262 -2226
rect 2256 -2238 2262 -2232
rect 2256 -2244 2262 -2238
rect 2256 -2250 2262 -2244
rect 2256 -2256 2262 -2250
rect 2256 -2262 2262 -2256
rect 2256 -2268 2262 -2262
rect 2256 -2274 2262 -2268
rect 2256 -2346 2262 -2340
rect 2256 -2352 2262 -2346
rect 2256 -2358 2262 -2352
rect 2256 -2364 2262 -2358
rect 2256 -2370 2262 -2364
rect 2256 -2376 2262 -2370
rect 2256 -2382 2262 -2376
rect 2256 -2388 2262 -2382
rect 2256 -2394 2262 -2388
rect 2256 -2400 2262 -2394
rect 2256 -2406 2262 -2400
rect 2256 -2412 2262 -2406
rect 2256 -2418 2262 -2412
rect 2256 -2424 2262 -2418
rect 2256 -2430 2262 -2424
rect 2256 -2436 2262 -2430
rect 2256 -2442 2262 -2436
rect 2256 -2448 2262 -2442
rect 2256 -2454 2262 -2448
rect 2256 -2460 2262 -2454
rect 2256 -2520 2262 -2514
rect 2256 -2526 2262 -2520
rect 2256 -2532 2262 -2526
rect 2256 -2538 2262 -2532
rect 2256 -2544 2262 -2538
rect 2256 -2550 2262 -2544
rect 2256 -2556 2262 -2550
rect 2256 -2562 2262 -2556
rect 2256 -2568 2262 -2562
rect 2256 -2574 2262 -2568
rect 2256 -2580 2262 -2574
rect 2256 -2586 2262 -2580
rect 2256 -2592 2262 -2586
rect 2256 -2598 2262 -2592
rect 2256 -2604 2262 -2598
rect 2256 -2610 2262 -2604
rect 2256 -2616 2262 -2610
rect 2256 -2622 2262 -2616
rect 2256 -2628 2262 -2622
rect 2256 -2634 2262 -2628
rect 2256 -2640 2262 -2634
rect 2256 -2646 2262 -2640
rect 2256 -2652 2262 -2646
rect 2256 -2658 2262 -2652
rect 2256 -2664 2262 -2658
rect 2256 -2670 2262 -2664
rect 2256 -2676 2262 -2670
rect 2256 -2682 2262 -2676
rect 2256 -2688 2262 -2682
rect 2256 -2694 2262 -2688
rect 2256 -2700 2262 -2694
rect 2256 -2706 2262 -2700
rect 2256 -2712 2262 -2706
rect 2256 -2718 2262 -2712
rect 2256 -2724 2262 -2718
rect 2256 -2730 2262 -2724
rect 2256 -2736 2262 -2730
rect 2256 -2742 2262 -2736
rect 2256 -2748 2262 -2742
rect 2256 -2754 2262 -2748
rect 2256 -2760 2262 -2754
rect 2256 -2766 2262 -2760
rect 2256 -2772 2262 -2766
rect 2256 -2778 2262 -2772
rect 2256 -2784 2262 -2778
rect 2256 -2790 2262 -2784
rect 2256 -2796 2262 -2790
rect 2256 -2802 2262 -2796
rect 2256 -2808 2262 -2802
rect 2256 -2814 2262 -2808
rect 2256 -2820 2262 -2814
rect 2256 -2826 2262 -2820
rect 2256 -2832 2262 -2826
rect 2256 -2838 2262 -2832
rect 2256 -2844 2262 -2838
rect 2256 -2850 2262 -2844
rect 2256 -2856 2262 -2850
rect 2256 -2862 2262 -2856
rect 2256 -2868 2262 -2862
rect 2256 -2874 2262 -2868
rect 2256 -2880 2262 -2874
rect 2256 -2886 2262 -2880
rect 2256 -2892 2262 -2886
rect 2256 -2898 2262 -2892
rect 2256 -2904 2262 -2898
rect 2256 -2910 2262 -2904
rect 2256 -2916 2262 -2910
rect 2256 -2922 2262 -2916
rect 2256 -2928 2262 -2922
rect 2256 -2934 2262 -2928
rect 2256 -2940 2262 -2934
rect 2256 -2946 2262 -2940
rect 2256 -2952 2262 -2946
rect 2256 -2958 2262 -2952
rect 2256 -2964 2262 -2958
rect 2256 -2970 2262 -2964
rect 2262 -120 2268 -114
rect 2262 -126 2268 -120
rect 2262 -132 2268 -126
rect 2262 -138 2268 -132
rect 2262 -144 2268 -138
rect 2262 -150 2268 -144
rect 2262 -156 2268 -150
rect 2262 -162 2268 -156
rect 2262 -168 2268 -162
rect 2262 -174 2268 -168
rect 2262 -180 2268 -174
rect 2262 -186 2268 -180
rect 2262 -192 2268 -186
rect 2262 -198 2268 -192
rect 2262 -204 2268 -198
rect 2262 -210 2268 -204
rect 2262 -216 2268 -210
rect 2262 -222 2268 -216
rect 2262 -228 2268 -222
rect 2262 -234 2268 -228
rect 2262 -240 2268 -234
rect 2262 -246 2268 -240
rect 2262 -252 2268 -246
rect 2262 -258 2268 -252
rect 2262 -264 2268 -258
rect 2262 -270 2268 -264
rect 2262 -276 2268 -270
rect 2262 -282 2268 -276
rect 2262 -288 2268 -282
rect 2262 -294 2268 -288
rect 2262 -300 2268 -294
rect 2262 -306 2268 -300
rect 2262 -312 2268 -306
rect 2262 -318 2268 -312
rect 2262 -324 2268 -318
rect 2262 -330 2268 -324
rect 2262 -336 2268 -330
rect 2262 -342 2268 -336
rect 2262 -348 2268 -342
rect 2262 -354 2268 -348
rect 2262 -360 2268 -354
rect 2262 -366 2268 -360
rect 2262 -372 2268 -366
rect 2262 -378 2268 -372
rect 2262 -384 2268 -378
rect 2262 -390 2268 -384
rect 2262 -396 2268 -390
rect 2262 -402 2268 -396
rect 2262 -408 2268 -402
rect 2262 -414 2268 -408
rect 2262 -420 2268 -414
rect 2262 -426 2268 -420
rect 2262 -432 2268 -426
rect 2262 -438 2268 -432
rect 2262 -444 2268 -438
rect 2262 -450 2268 -444
rect 2262 -456 2268 -450
rect 2262 -462 2268 -456
rect 2262 -468 2268 -462
rect 2262 -474 2268 -468
rect 2262 -480 2268 -474
rect 2262 -486 2268 -480
rect 2262 -492 2268 -486
rect 2262 -498 2268 -492
rect 2262 -504 2268 -498
rect 2262 -510 2268 -504
rect 2262 -516 2268 -510
rect 2262 -522 2268 -516
rect 2262 -528 2268 -522
rect 2262 -534 2268 -528
rect 2262 -540 2268 -534
rect 2262 -546 2268 -540
rect 2262 -552 2268 -546
rect 2262 -558 2268 -552
rect 2262 -564 2268 -558
rect 2262 -570 2268 -564
rect 2262 -576 2268 -570
rect 2262 -582 2268 -576
rect 2262 -588 2268 -582
rect 2262 -594 2268 -588
rect 2262 -600 2268 -594
rect 2262 -606 2268 -600
rect 2262 -612 2268 -606
rect 2262 -618 2268 -612
rect 2262 -624 2268 -618
rect 2262 -630 2268 -624
rect 2262 -636 2268 -630
rect 2262 -642 2268 -636
rect 2262 -648 2268 -642
rect 2262 -654 2268 -648
rect 2262 -660 2268 -654
rect 2262 -666 2268 -660
rect 2262 -672 2268 -666
rect 2262 -678 2268 -672
rect 2262 -684 2268 -678
rect 2262 -690 2268 -684
rect 2262 -696 2268 -690
rect 2262 -702 2268 -696
rect 2262 -708 2268 -702
rect 2262 -714 2268 -708
rect 2262 -720 2268 -714
rect 2262 -726 2268 -720
rect 2262 -732 2268 -726
rect 2262 -738 2268 -732
rect 2262 -744 2268 -738
rect 2262 -750 2268 -744
rect 2262 -756 2268 -750
rect 2262 -762 2268 -756
rect 2262 -768 2268 -762
rect 2262 -774 2268 -768
rect 2262 -780 2268 -774
rect 2262 -786 2268 -780
rect 2262 -792 2268 -786
rect 2262 -798 2268 -792
rect 2262 -804 2268 -798
rect 2262 -810 2268 -804
rect 2262 -816 2268 -810
rect 2262 -822 2268 -816
rect 2262 -828 2268 -822
rect 2262 -834 2268 -828
rect 2262 -840 2268 -834
rect 2262 -846 2268 -840
rect 2262 -852 2268 -846
rect 2262 -858 2268 -852
rect 2262 -864 2268 -858
rect 2262 -870 2268 -864
rect 2262 -876 2268 -870
rect 2262 -882 2268 -876
rect 2262 -888 2268 -882
rect 2262 -894 2268 -888
rect 2262 -900 2268 -894
rect 2262 -906 2268 -900
rect 2262 -912 2268 -906
rect 2262 -918 2268 -912
rect 2262 -924 2268 -918
rect 2262 -930 2268 -924
rect 2262 -936 2268 -930
rect 2262 -942 2268 -936
rect 2262 -948 2268 -942
rect 2262 -954 2268 -948
rect 2262 -960 2268 -954
rect 2262 -966 2268 -960
rect 2262 -972 2268 -966
rect 2262 -978 2268 -972
rect 2262 -984 2268 -978
rect 2262 -990 2268 -984
rect 2262 -996 2268 -990
rect 2262 -1002 2268 -996
rect 2262 -1008 2268 -1002
rect 2262 -1014 2268 -1008
rect 2262 -1020 2268 -1014
rect 2262 -1026 2268 -1020
rect 2262 -1032 2268 -1026
rect 2262 -1038 2268 -1032
rect 2262 -1044 2268 -1038
rect 2262 -1050 2268 -1044
rect 2262 -1056 2268 -1050
rect 2262 -1062 2268 -1056
rect 2262 -1068 2268 -1062
rect 2262 -1074 2268 -1068
rect 2262 -1080 2268 -1074
rect 2262 -1086 2268 -1080
rect 2262 -1092 2268 -1086
rect 2262 -1500 2268 -1494
rect 2262 -1506 2268 -1500
rect 2262 -1512 2268 -1506
rect 2262 -1518 2268 -1512
rect 2262 -1524 2268 -1518
rect 2262 -1530 2268 -1524
rect 2262 -1536 2268 -1530
rect 2262 -1542 2268 -1536
rect 2262 -1548 2268 -1542
rect 2262 -1554 2268 -1548
rect 2262 -1560 2268 -1554
rect 2262 -1566 2268 -1560
rect 2262 -1572 2268 -1566
rect 2262 -1578 2268 -1572
rect 2262 -1584 2268 -1578
rect 2262 -1590 2268 -1584
rect 2262 -1596 2268 -1590
rect 2262 -1602 2268 -1596
rect 2262 -1608 2268 -1602
rect 2262 -1614 2268 -1608
rect 2262 -1620 2268 -1614
rect 2262 -1626 2268 -1620
rect 2262 -1632 2268 -1626
rect 2262 -1638 2268 -1632
rect 2262 -1644 2268 -1638
rect 2262 -1650 2268 -1644
rect 2262 -1656 2268 -1650
rect 2262 -1662 2268 -1656
rect 2262 -1668 2268 -1662
rect 2262 -1674 2268 -1668
rect 2262 -1680 2268 -1674
rect 2262 -1686 2268 -1680
rect 2262 -1692 2268 -1686
rect 2262 -1698 2268 -1692
rect 2262 -1704 2268 -1698
rect 2262 -1710 2268 -1704
rect 2262 -1716 2268 -1710
rect 2262 -1722 2268 -1716
rect 2262 -1728 2268 -1722
rect 2262 -1734 2268 -1728
rect 2262 -1740 2268 -1734
rect 2262 -1746 2268 -1740
rect 2262 -1752 2268 -1746
rect 2262 -1758 2268 -1752
rect 2262 -1764 2268 -1758
rect 2262 -1770 2268 -1764
rect 2262 -1776 2268 -1770
rect 2262 -1782 2268 -1776
rect 2262 -1788 2268 -1782
rect 2262 -1794 2268 -1788
rect 2262 -1800 2268 -1794
rect 2262 -1806 2268 -1800
rect 2262 -1812 2268 -1806
rect 2262 -1818 2268 -1812
rect 2262 -1824 2268 -1818
rect 2262 -1830 2268 -1824
rect 2262 -1836 2268 -1830
rect 2262 -1842 2268 -1836
rect 2262 -1848 2268 -1842
rect 2262 -1854 2268 -1848
rect 2262 -1860 2268 -1854
rect 2262 -1866 2268 -1860
rect 2262 -1872 2268 -1866
rect 2262 -1878 2268 -1872
rect 2262 -1884 2268 -1878
rect 2262 -1890 2268 -1884
rect 2262 -1896 2268 -1890
rect 2262 -1902 2268 -1896
rect 2262 -1908 2268 -1902
rect 2262 -1914 2268 -1908
rect 2262 -1920 2268 -1914
rect 2262 -1926 2268 -1920
rect 2262 -1932 2268 -1926
rect 2262 -1938 2268 -1932
rect 2262 -1944 2268 -1938
rect 2262 -1950 2268 -1944
rect 2262 -1956 2268 -1950
rect 2262 -1962 2268 -1956
rect 2262 -1968 2268 -1962
rect 2262 -1974 2268 -1968
rect 2262 -1980 2268 -1974
rect 2262 -1986 2268 -1980
rect 2262 -1992 2268 -1986
rect 2262 -1998 2268 -1992
rect 2262 -2004 2268 -1998
rect 2262 -2010 2268 -2004
rect 2262 -2016 2268 -2010
rect 2262 -2022 2268 -2016
rect 2262 -2028 2268 -2022
rect 2262 -2034 2268 -2028
rect 2262 -2040 2268 -2034
rect 2262 -2046 2268 -2040
rect 2262 -2052 2268 -2046
rect 2262 -2058 2268 -2052
rect 2262 -2064 2268 -2058
rect 2262 -2070 2268 -2064
rect 2262 -2076 2268 -2070
rect 2262 -2082 2268 -2076
rect 2262 -2088 2268 -2082
rect 2262 -2094 2268 -2088
rect 2262 -2100 2268 -2094
rect 2262 -2106 2268 -2100
rect 2262 -2112 2268 -2106
rect 2262 -2118 2268 -2112
rect 2262 -2124 2268 -2118
rect 2262 -2130 2268 -2124
rect 2262 -2136 2268 -2130
rect 2262 -2142 2268 -2136
rect 2262 -2148 2268 -2142
rect 2262 -2154 2268 -2148
rect 2262 -2160 2268 -2154
rect 2262 -2166 2268 -2160
rect 2262 -2172 2268 -2166
rect 2262 -2178 2268 -2172
rect 2262 -2184 2268 -2178
rect 2262 -2190 2268 -2184
rect 2262 -2196 2268 -2190
rect 2262 -2202 2268 -2196
rect 2262 -2208 2268 -2202
rect 2262 -2214 2268 -2208
rect 2262 -2220 2268 -2214
rect 2262 -2226 2268 -2220
rect 2262 -2232 2268 -2226
rect 2262 -2238 2268 -2232
rect 2262 -2244 2268 -2238
rect 2262 -2250 2268 -2244
rect 2262 -2256 2268 -2250
rect 2262 -2262 2268 -2256
rect 2262 -2268 2268 -2262
rect 2262 -2334 2268 -2328
rect 2262 -2340 2268 -2334
rect 2262 -2346 2268 -2340
rect 2262 -2352 2268 -2346
rect 2262 -2358 2268 -2352
rect 2262 -2364 2268 -2358
rect 2262 -2370 2268 -2364
rect 2262 -2376 2268 -2370
rect 2262 -2382 2268 -2376
rect 2262 -2388 2268 -2382
rect 2262 -2394 2268 -2388
rect 2262 -2400 2268 -2394
rect 2262 -2406 2268 -2400
rect 2262 -2412 2268 -2406
rect 2262 -2418 2268 -2412
rect 2262 -2424 2268 -2418
rect 2262 -2430 2268 -2424
rect 2262 -2436 2268 -2430
rect 2262 -2442 2268 -2436
rect 2262 -2448 2268 -2442
rect 2262 -2454 2268 -2448
rect 2262 -2460 2268 -2454
rect 2262 -2520 2268 -2514
rect 2262 -2526 2268 -2520
rect 2262 -2532 2268 -2526
rect 2262 -2538 2268 -2532
rect 2262 -2544 2268 -2538
rect 2262 -2550 2268 -2544
rect 2262 -2556 2268 -2550
rect 2262 -2562 2268 -2556
rect 2262 -2568 2268 -2562
rect 2262 -2574 2268 -2568
rect 2262 -2580 2268 -2574
rect 2262 -2586 2268 -2580
rect 2262 -2592 2268 -2586
rect 2262 -2598 2268 -2592
rect 2262 -2604 2268 -2598
rect 2262 -2610 2268 -2604
rect 2262 -2616 2268 -2610
rect 2262 -2622 2268 -2616
rect 2262 -2628 2268 -2622
rect 2262 -2634 2268 -2628
rect 2262 -2640 2268 -2634
rect 2262 -2646 2268 -2640
rect 2262 -2652 2268 -2646
rect 2262 -2658 2268 -2652
rect 2262 -2664 2268 -2658
rect 2262 -2670 2268 -2664
rect 2262 -2676 2268 -2670
rect 2262 -2682 2268 -2676
rect 2262 -2688 2268 -2682
rect 2262 -2694 2268 -2688
rect 2262 -2700 2268 -2694
rect 2262 -2706 2268 -2700
rect 2262 -2712 2268 -2706
rect 2262 -2718 2268 -2712
rect 2262 -2724 2268 -2718
rect 2262 -2730 2268 -2724
rect 2262 -2736 2268 -2730
rect 2262 -2742 2268 -2736
rect 2262 -2748 2268 -2742
rect 2262 -2754 2268 -2748
rect 2262 -2760 2268 -2754
rect 2262 -2766 2268 -2760
rect 2262 -2772 2268 -2766
rect 2262 -2778 2268 -2772
rect 2262 -2784 2268 -2778
rect 2262 -2790 2268 -2784
rect 2262 -2796 2268 -2790
rect 2262 -2802 2268 -2796
rect 2262 -2808 2268 -2802
rect 2262 -2814 2268 -2808
rect 2262 -2820 2268 -2814
rect 2262 -2826 2268 -2820
rect 2262 -2832 2268 -2826
rect 2262 -2838 2268 -2832
rect 2262 -2844 2268 -2838
rect 2262 -2850 2268 -2844
rect 2262 -2856 2268 -2850
rect 2262 -2862 2268 -2856
rect 2262 -2868 2268 -2862
rect 2262 -2874 2268 -2868
rect 2262 -2880 2268 -2874
rect 2262 -2886 2268 -2880
rect 2262 -2892 2268 -2886
rect 2262 -2898 2268 -2892
rect 2262 -2904 2268 -2898
rect 2262 -2910 2268 -2904
rect 2262 -2916 2268 -2910
rect 2262 -2922 2268 -2916
rect 2262 -2928 2268 -2922
rect 2262 -2934 2268 -2928
rect 2262 -2940 2268 -2934
rect 2262 -2946 2268 -2940
rect 2262 -2952 2268 -2946
rect 2262 -2958 2268 -2952
rect 2262 -2964 2268 -2958
rect 2262 -2970 2268 -2964
rect 2268 -114 2274 -108
rect 2268 -120 2274 -114
rect 2268 -126 2274 -120
rect 2268 -132 2274 -126
rect 2268 -138 2274 -132
rect 2268 -144 2274 -138
rect 2268 -150 2274 -144
rect 2268 -156 2274 -150
rect 2268 -162 2274 -156
rect 2268 -168 2274 -162
rect 2268 -174 2274 -168
rect 2268 -180 2274 -174
rect 2268 -186 2274 -180
rect 2268 -192 2274 -186
rect 2268 -198 2274 -192
rect 2268 -204 2274 -198
rect 2268 -210 2274 -204
rect 2268 -216 2274 -210
rect 2268 -222 2274 -216
rect 2268 -228 2274 -222
rect 2268 -234 2274 -228
rect 2268 -240 2274 -234
rect 2268 -246 2274 -240
rect 2268 -252 2274 -246
rect 2268 -258 2274 -252
rect 2268 -264 2274 -258
rect 2268 -270 2274 -264
rect 2268 -276 2274 -270
rect 2268 -282 2274 -276
rect 2268 -288 2274 -282
rect 2268 -294 2274 -288
rect 2268 -300 2274 -294
rect 2268 -306 2274 -300
rect 2268 -312 2274 -306
rect 2268 -318 2274 -312
rect 2268 -324 2274 -318
rect 2268 -330 2274 -324
rect 2268 -336 2274 -330
rect 2268 -342 2274 -336
rect 2268 -348 2274 -342
rect 2268 -354 2274 -348
rect 2268 -360 2274 -354
rect 2268 -366 2274 -360
rect 2268 -372 2274 -366
rect 2268 -378 2274 -372
rect 2268 -384 2274 -378
rect 2268 -390 2274 -384
rect 2268 -396 2274 -390
rect 2268 -402 2274 -396
rect 2268 -408 2274 -402
rect 2268 -414 2274 -408
rect 2268 -420 2274 -414
rect 2268 -426 2274 -420
rect 2268 -432 2274 -426
rect 2268 -438 2274 -432
rect 2268 -444 2274 -438
rect 2268 -450 2274 -444
rect 2268 -456 2274 -450
rect 2268 -462 2274 -456
rect 2268 -468 2274 -462
rect 2268 -474 2274 -468
rect 2268 -480 2274 -474
rect 2268 -486 2274 -480
rect 2268 -492 2274 -486
rect 2268 -498 2274 -492
rect 2268 -504 2274 -498
rect 2268 -510 2274 -504
rect 2268 -516 2274 -510
rect 2268 -522 2274 -516
rect 2268 -528 2274 -522
rect 2268 -534 2274 -528
rect 2268 -540 2274 -534
rect 2268 -546 2274 -540
rect 2268 -552 2274 -546
rect 2268 -558 2274 -552
rect 2268 -564 2274 -558
rect 2268 -570 2274 -564
rect 2268 -576 2274 -570
rect 2268 -582 2274 -576
rect 2268 -588 2274 -582
rect 2268 -594 2274 -588
rect 2268 -600 2274 -594
rect 2268 -606 2274 -600
rect 2268 -612 2274 -606
rect 2268 -618 2274 -612
rect 2268 -624 2274 -618
rect 2268 -630 2274 -624
rect 2268 -636 2274 -630
rect 2268 -642 2274 -636
rect 2268 -648 2274 -642
rect 2268 -654 2274 -648
rect 2268 -660 2274 -654
rect 2268 -666 2274 -660
rect 2268 -672 2274 -666
rect 2268 -678 2274 -672
rect 2268 -684 2274 -678
rect 2268 -690 2274 -684
rect 2268 -696 2274 -690
rect 2268 -702 2274 -696
rect 2268 -708 2274 -702
rect 2268 -714 2274 -708
rect 2268 -720 2274 -714
rect 2268 -726 2274 -720
rect 2268 -732 2274 -726
rect 2268 -738 2274 -732
rect 2268 -744 2274 -738
rect 2268 -750 2274 -744
rect 2268 -756 2274 -750
rect 2268 -762 2274 -756
rect 2268 -768 2274 -762
rect 2268 -774 2274 -768
rect 2268 -780 2274 -774
rect 2268 -786 2274 -780
rect 2268 -792 2274 -786
rect 2268 -798 2274 -792
rect 2268 -804 2274 -798
rect 2268 -810 2274 -804
rect 2268 -816 2274 -810
rect 2268 -822 2274 -816
rect 2268 -828 2274 -822
rect 2268 -834 2274 -828
rect 2268 -840 2274 -834
rect 2268 -846 2274 -840
rect 2268 -852 2274 -846
rect 2268 -858 2274 -852
rect 2268 -864 2274 -858
rect 2268 -870 2274 -864
rect 2268 -876 2274 -870
rect 2268 -882 2274 -876
rect 2268 -888 2274 -882
rect 2268 -894 2274 -888
rect 2268 -900 2274 -894
rect 2268 -906 2274 -900
rect 2268 -912 2274 -906
rect 2268 -918 2274 -912
rect 2268 -924 2274 -918
rect 2268 -930 2274 -924
rect 2268 -936 2274 -930
rect 2268 -942 2274 -936
rect 2268 -948 2274 -942
rect 2268 -954 2274 -948
rect 2268 -960 2274 -954
rect 2268 -966 2274 -960
rect 2268 -972 2274 -966
rect 2268 -978 2274 -972
rect 2268 -984 2274 -978
rect 2268 -990 2274 -984
rect 2268 -996 2274 -990
rect 2268 -1002 2274 -996
rect 2268 -1008 2274 -1002
rect 2268 -1014 2274 -1008
rect 2268 -1020 2274 -1014
rect 2268 -1026 2274 -1020
rect 2268 -1032 2274 -1026
rect 2268 -1038 2274 -1032
rect 2268 -1044 2274 -1038
rect 2268 -1050 2274 -1044
rect 2268 -1056 2274 -1050
rect 2268 -1062 2274 -1056
rect 2268 -1068 2274 -1062
rect 2268 -1074 2274 -1068
rect 2268 -1494 2274 -1488
rect 2268 -1500 2274 -1494
rect 2268 -1506 2274 -1500
rect 2268 -1512 2274 -1506
rect 2268 -1518 2274 -1512
rect 2268 -1524 2274 -1518
rect 2268 -1530 2274 -1524
rect 2268 -1536 2274 -1530
rect 2268 -1542 2274 -1536
rect 2268 -1548 2274 -1542
rect 2268 -1554 2274 -1548
rect 2268 -1560 2274 -1554
rect 2268 -1566 2274 -1560
rect 2268 -1572 2274 -1566
rect 2268 -1578 2274 -1572
rect 2268 -1584 2274 -1578
rect 2268 -1590 2274 -1584
rect 2268 -1596 2274 -1590
rect 2268 -1602 2274 -1596
rect 2268 -1608 2274 -1602
rect 2268 -1614 2274 -1608
rect 2268 -1620 2274 -1614
rect 2268 -1626 2274 -1620
rect 2268 -1632 2274 -1626
rect 2268 -1638 2274 -1632
rect 2268 -1644 2274 -1638
rect 2268 -1650 2274 -1644
rect 2268 -1656 2274 -1650
rect 2268 -1662 2274 -1656
rect 2268 -1668 2274 -1662
rect 2268 -1674 2274 -1668
rect 2268 -1680 2274 -1674
rect 2268 -1686 2274 -1680
rect 2268 -1692 2274 -1686
rect 2268 -1698 2274 -1692
rect 2268 -1704 2274 -1698
rect 2268 -1710 2274 -1704
rect 2268 -1716 2274 -1710
rect 2268 -1722 2274 -1716
rect 2268 -1728 2274 -1722
rect 2268 -1734 2274 -1728
rect 2268 -1740 2274 -1734
rect 2268 -1746 2274 -1740
rect 2268 -1752 2274 -1746
rect 2268 -1758 2274 -1752
rect 2268 -1764 2274 -1758
rect 2268 -1770 2274 -1764
rect 2268 -1776 2274 -1770
rect 2268 -1782 2274 -1776
rect 2268 -1788 2274 -1782
rect 2268 -1794 2274 -1788
rect 2268 -1800 2274 -1794
rect 2268 -1806 2274 -1800
rect 2268 -1812 2274 -1806
rect 2268 -1818 2274 -1812
rect 2268 -1824 2274 -1818
rect 2268 -1830 2274 -1824
rect 2268 -1836 2274 -1830
rect 2268 -1842 2274 -1836
rect 2268 -1848 2274 -1842
rect 2268 -1854 2274 -1848
rect 2268 -1860 2274 -1854
rect 2268 -1866 2274 -1860
rect 2268 -1872 2274 -1866
rect 2268 -1878 2274 -1872
rect 2268 -1884 2274 -1878
rect 2268 -1890 2274 -1884
rect 2268 -1896 2274 -1890
rect 2268 -1902 2274 -1896
rect 2268 -1908 2274 -1902
rect 2268 -1914 2274 -1908
rect 2268 -1920 2274 -1914
rect 2268 -1926 2274 -1920
rect 2268 -1932 2274 -1926
rect 2268 -1938 2274 -1932
rect 2268 -1944 2274 -1938
rect 2268 -1950 2274 -1944
rect 2268 -1956 2274 -1950
rect 2268 -1962 2274 -1956
rect 2268 -1968 2274 -1962
rect 2268 -1974 2274 -1968
rect 2268 -1980 2274 -1974
rect 2268 -1986 2274 -1980
rect 2268 -1992 2274 -1986
rect 2268 -1998 2274 -1992
rect 2268 -2004 2274 -1998
rect 2268 -2010 2274 -2004
rect 2268 -2016 2274 -2010
rect 2268 -2022 2274 -2016
rect 2268 -2028 2274 -2022
rect 2268 -2034 2274 -2028
rect 2268 -2040 2274 -2034
rect 2268 -2046 2274 -2040
rect 2268 -2052 2274 -2046
rect 2268 -2058 2274 -2052
rect 2268 -2064 2274 -2058
rect 2268 -2070 2274 -2064
rect 2268 -2076 2274 -2070
rect 2268 -2082 2274 -2076
rect 2268 -2088 2274 -2082
rect 2268 -2094 2274 -2088
rect 2268 -2100 2274 -2094
rect 2268 -2106 2274 -2100
rect 2268 -2112 2274 -2106
rect 2268 -2118 2274 -2112
rect 2268 -2124 2274 -2118
rect 2268 -2130 2274 -2124
rect 2268 -2136 2274 -2130
rect 2268 -2142 2274 -2136
rect 2268 -2148 2274 -2142
rect 2268 -2154 2274 -2148
rect 2268 -2160 2274 -2154
rect 2268 -2166 2274 -2160
rect 2268 -2172 2274 -2166
rect 2268 -2178 2274 -2172
rect 2268 -2184 2274 -2178
rect 2268 -2190 2274 -2184
rect 2268 -2196 2274 -2190
rect 2268 -2202 2274 -2196
rect 2268 -2208 2274 -2202
rect 2268 -2214 2274 -2208
rect 2268 -2220 2274 -2214
rect 2268 -2226 2274 -2220
rect 2268 -2232 2274 -2226
rect 2268 -2238 2274 -2232
rect 2268 -2244 2274 -2238
rect 2268 -2250 2274 -2244
rect 2268 -2256 2274 -2250
rect 2268 -2262 2274 -2256
rect 2268 -2328 2274 -2322
rect 2268 -2334 2274 -2328
rect 2268 -2340 2274 -2334
rect 2268 -2346 2274 -2340
rect 2268 -2352 2274 -2346
rect 2268 -2358 2274 -2352
rect 2268 -2364 2274 -2358
rect 2268 -2370 2274 -2364
rect 2268 -2376 2274 -2370
rect 2268 -2382 2274 -2376
rect 2268 -2388 2274 -2382
rect 2268 -2394 2274 -2388
rect 2268 -2400 2274 -2394
rect 2268 -2406 2274 -2400
rect 2268 -2412 2274 -2406
rect 2268 -2418 2274 -2412
rect 2268 -2424 2274 -2418
rect 2268 -2430 2274 -2424
rect 2268 -2436 2274 -2430
rect 2268 -2442 2274 -2436
rect 2268 -2448 2274 -2442
rect 2268 -2454 2274 -2448
rect 2268 -2514 2274 -2508
rect 2268 -2520 2274 -2514
rect 2268 -2526 2274 -2520
rect 2268 -2532 2274 -2526
rect 2268 -2538 2274 -2532
rect 2268 -2544 2274 -2538
rect 2268 -2550 2274 -2544
rect 2268 -2556 2274 -2550
rect 2268 -2562 2274 -2556
rect 2268 -2568 2274 -2562
rect 2268 -2574 2274 -2568
rect 2268 -2580 2274 -2574
rect 2268 -2586 2274 -2580
rect 2268 -2592 2274 -2586
rect 2268 -2598 2274 -2592
rect 2268 -2604 2274 -2598
rect 2268 -2610 2274 -2604
rect 2268 -2616 2274 -2610
rect 2268 -2622 2274 -2616
rect 2268 -2628 2274 -2622
rect 2268 -2634 2274 -2628
rect 2268 -2640 2274 -2634
rect 2268 -2646 2274 -2640
rect 2268 -2652 2274 -2646
rect 2268 -2658 2274 -2652
rect 2268 -2664 2274 -2658
rect 2268 -2670 2274 -2664
rect 2268 -2676 2274 -2670
rect 2268 -2682 2274 -2676
rect 2268 -2688 2274 -2682
rect 2268 -2694 2274 -2688
rect 2268 -2700 2274 -2694
rect 2268 -2706 2274 -2700
rect 2268 -2712 2274 -2706
rect 2268 -2718 2274 -2712
rect 2268 -2724 2274 -2718
rect 2268 -2730 2274 -2724
rect 2268 -2736 2274 -2730
rect 2268 -2742 2274 -2736
rect 2268 -2748 2274 -2742
rect 2268 -2754 2274 -2748
rect 2268 -2760 2274 -2754
rect 2268 -2766 2274 -2760
rect 2268 -2772 2274 -2766
rect 2268 -2778 2274 -2772
rect 2268 -2784 2274 -2778
rect 2268 -2790 2274 -2784
rect 2268 -2796 2274 -2790
rect 2268 -2802 2274 -2796
rect 2268 -2808 2274 -2802
rect 2268 -2814 2274 -2808
rect 2268 -2820 2274 -2814
rect 2268 -2826 2274 -2820
rect 2268 -2832 2274 -2826
rect 2268 -2838 2274 -2832
rect 2268 -2844 2274 -2838
rect 2268 -2850 2274 -2844
rect 2268 -2856 2274 -2850
rect 2268 -2862 2274 -2856
rect 2268 -2868 2274 -2862
rect 2268 -2874 2274 -2868
rect 2268 -2880 2274 -2874
rect 2268 -2886 2274 -2880
rect 2268 -2892 2274 -2886
rect 2268 -2898 2274 -2892
rect 2268 -2904 2274 -2898
rect 2268 -2910 2274 -2904
rect 2268 -2916 2274 -2910
rect 2268 -2922 2274 -2916
rect 2268 -2928 2274 -2922
rect 2268 -2934 2274 -2928
rect 2268 -2940 2274 -2934
rect 2268 -2946 2274 -2940
rect 2268 -2952 2274 -2946
rect 2268 -2958 2274 -2952
rect 2268 -2964 2274 -2958
rect 2274 -108 2280 -102
rect 2274 -114 2280 -108
rect 2274 -120 2280 -114
rect 2274 -126 2280 -120
rect 2274 -132 2280 -126
rect 2274 -138 2280 -132
rect 2274 -144 2280 -138
rect 2274 -150 2280 -144
rect 2274 -156 2280 -150
rect 2274 -162 2280 -156
rect 2274 -168 2280 -162
rect 2274 -174 2280 -168
rect 2274 -180 2280 -174
rect 2274 -186 2280 -180
rect 2274 -192 2280 -186
rect 2274 -198 2280 -192
rect 2274 -204 2280 -198
rect 2274 -210 2280 -204
rect 2274 -216 2280 -210
rect 2274 -222 2280 -216
rect 2274 -228 2280 -222
rect 2274 -234 2280 -228
rect 2274 -240 2280 -234
rect 2274 -246 2280 -240
rect 2274 -252 2280 -246
rect 2274 -258 2280 -252
rect 2274 -264 2280 -258
rect 2274 -270 2280 -264
rect 2274 -276 2280 -270
rect 2274 -282 2280 -276
rect 2274 -288 2280 -282
rect 2274 -294 2280 -288
rect 2274 -300 2280 -294
rect 2274 -306 2280 -300
rect 2274 -312 2280 -306
rect 2274 -318 2280 -312
rect 2274 -324 2280 -318
rect 2274 -330 2280 -324
rect 2274 -336 2280 -330
rect 2274 -342 2280 -336
rect 2274 -348 2280 -342
rect 2274 -354 2280 -348
rect 2274 -360 2280 -354
rect 2274 -366 2280 -360
rect 2274 -372 2280 -366
rect 2274 -378 2280 -372
rect 2274 -384 2280 -378
rect 2274 -390 2280 -384
rect 2274 -396 2280 -390
rect 2274 -402 2280 -396
rect 2274 -408 2280 -402
rect 2274 -414 2280 -408
rect 2274 -420 2280 -414
rect 2274 -426 2280 -420
rect 2274 -432 2280 -426
rect 2274 -438 2280 -432
rect 2274 -444 2280 -438
rect 2274 -450 2280 -444
rect 2274 -456 2280 -450
rect 2274 -462 2280 -456
rect 2274 -468 2280 -462
rect 2274 -474 2280 -468
rect 2274 -480 2280 -474
rect 2274 -486 2280 -480
rect 2274 -492 2280 -486
rect 2274 -498 2280 -492
rect 2274 -504 2280 -498
rect 2274 -510 2280 -504
rect 2274 -516 2280 -510
rect 2274 -522 2280 -516
rect 2274 -528 2280 -522
rect 2274 -534 2280 -528
rect 2274 -540 2280 -534
rect 2274 -546 2280 -540
rect 2274 -552 2280 -546
rect 2274 -558 2280 -552
rect 2274 -564 2280 -558
rect 2274 -570 2280 -564
rect 2274 -576 2280 -570
rect 2274 -582 2280 -576
rect 2274 -588 2280 -582
rect 2274 -594 2280 -588
rect 2274 -600 2280 -594
rect 2274 -606 2280 -600
rect 2274 -612 2280 -606
rect 2274 -618 2280 -612
rect 2274 -624 2280 -618
rect 2274 -630 2280 -624
rect 2274 -636 2280 -630
rect 2274 -642 2280 -636
rect 2274 -648 2280 -642
rect 2274 -654 2280 -648
rect 2274 -660 2280 -654
rect 2274 -666 2280 -660
rect 2274 -672 2280 -666
rect 2274 -678 2280 -672
rect 2274 -684 2280 -678
rect 2274 -690 2280 -684
rect 2274 -696 2280 -690
rect 2274 -702 2280 -696
rect 2274 -708 2280 -702
rect 2274 -714 2280 -708
rect 2274 -720 2280 -714
rect 2274 -726 2280 -720
rect 2274 -732 2280 -726
rect 2274 -738 2280 -732
rect 2274 -744 2280 -738
rect 2274 -750 2280 -744
rect 2274 -756 2280 -750
rect 2274 -762 2280 -756
rect 2274 -768 2280 -762
rect 2274 -774 2280 -768
rect 2274 -780 2280 -774
rect 2274 -786 2280 -780
rect 2274 -792 2280 -786
rect 2274 -798 2280 -792
rect 2274 -804 2280 -798
rect 2274 -810 2280 -804
rect 2274 -816 2280 -810
rect 2274 -822 2280 -816
rect 2274 -828 2280 -822
rect 2274 -834 2280 -828
rect 2274 -840 2280 -834
rect 2274 -846 2280 -840
rect 2274 -852 2280 -846
rect 2274 -858 2280 -852
rect 2274 -864 2280 -858
rect 2274 -870 2280 -864
rect 2274 -876 2280 -870
rect 2274 -882 2280 -876
rect 2274 -888 2280 -882
rect 2274 -894 2280 -888
rect 2274 -900 2280 -894
rect 2274 -906 2280 -900
rect 2274 -912 2280 -906
rect 2274 -918 2280 -912
rect 2274 -924 2280 -918
rect 2274 -930 2280 -924
rect 2274 -936 2280 -930
rect 2274 -942 2280 -936
rect 2274 -948 2280 -942
rect 2274 -954 2280 -948
rect 2274 -960 2280 -954
rect 2274 -966 2280 -960
rect 2274 -972 2280 -966
rect 2274 -978 2280 -972
rect 2274 -984 2280 -978
rect 2274 -990 2280 -984
rect 2274 -996 2280 -990
rect 2274 -1002 2280 -996
rect 2274 -1008 2280 -1002
rect 2274 -1014 2280 -1008
rect 2274 -1020 2280 -1014
rect 2274 -1026 2280 -1020
rect 2274 -1032 2280 -1026
rect 2274 -1038 2280 -1032
rect 2274 -1044 2280 -1038
rect 2274 -1050 2280 -1044
rect 2274 -1056 2280 -1050
rect 2274 -1062 2280 -1056
rect 2274 -1488 2280 -1482
rect 2274 -1494 2280 -1488
rect 2274 -1500 2280 -1494
rect 2274 -1506 2280 -1500
rect 2274 -1512 2280 -1506
rect 2274 -1518 2280 -1512
rect 2274 -1524 2280 -1518
rect 2274 -1530 2280 -1524
rect 2274 -1536 2280 -1530
rect 2274 -1542 2280 -1536
rect 2274 -1548 2280 -1542
rect 2274 -1554 2280 -1548
rect 2274 -1560 2280 -1554
rect 2274 -1566 2280 -1560
rect 2274 -1572 2280 -1566
rect 2274 -1578 2280 -1572
rect 2274 -1584 2280 -1578
rect 2274 -1590 2280 -1584
rect 2274 -1596 2280 -1590
rect 2274 -1602 2280 -1596
rect 2274 -1608 2280 -1602
rect 2274 -1614 2280 -1608
rect 2274 -1620 2280 -1614
rect 2274 -1626 2280 -1620
rect 2274 -1632 2280 -1626
rect 2274 -1638 2280 -1632
rect 2274 -1644 2280 -1638
rect 2274 -1650 2280 -1644
rect 2274 -1656 2280 -1650
rect 2274 -1662 2280 -1656
rect 2274 -1668 2280 -1662
rect 2274 -1674 2280 -1668
rect 2274 -1680 2280 -1674
rect 2274 -1686 2280 -1680
rect 2274 -1692 2280 -1686
rect 2274 -1698 2280 -1692
rect 2274 -1704 2280 -1698
rect 2274 -1710 2280 -1704
rect 2274 -1716 2280 -1710
rect 2274 -1722 2280 -1716
rect 2274 -1728 2280 -1722
rect 2274 -1734 2280 -1728
rect 2274 -1740 2280 -1734
rect 2274 -1746 2280 -1740
rect 2274 -1752 2280 -1746
rect 2274 -1758 2280 -1752
rect 2274 -1764 2280 -1758
rect 2274 -1770 2280 -1764
rect 2274 -1776 2280 -1770
rect 2274 -1782 2280 -1776
rect 2274 -1788 2280 -1782
rect 2274 -1794 2280 -1788
rect 2274 -1800 2280 -1794
rect 2274 -1806 2280 -1800
rect 2274 -1812 2280 -1806
rect 2274 -1818 2280 -1812
rect 2274 -1824 2280 -1818
rect 2274 -1830 2280 -1824
rect 2274 -1836 2280 -1830
rect 2274 -1842 2280 -1836
rect 2274 -1848 2280 -1842
rect 2274 -1854 2280 -1848
rect 2274 -1860 2280 -1854
rect 2274 -1866 2280 -1860
rect 2274 -1872 2280 -1866
rect 2274 -1878 2280 -1872
rect 2274 -1884 2280 -1878
rect 2274 -1890 2280 -1884
rect 2274 -1896 2280 -1890
rect 2274 -1902 2280 -1896
rect 2274 -1908 2280 -1902
rect 2274 -1914 2280 -1908
rect 2274 -1920 2280 -1914
rect 2274 -1926 2280 -1920
rect 2274 -1932 2280 -1926
rect 2274 -1938 2280 -1932
rect 2274 -1944 2280 -1938
rect 2274 -1950 2280 -1944
rect 2274 -1956 2280 -1950
rect 2274 -1962 2280 -1956
rect 2274 -1968 2280 -1962
rect 2274 -1974 2280 -1968
rect 2274 -1980 2280 -1974
rect 2274 -1986 2280 -1980
rect 2274 -1992 2280 -1986
rect 2274 -1998 2280 -1992
rect 2274 -2004 2280 -1998
rect 2274 -2010 2280 -2004
rect 2274 -2016 2280 -2010
rect 2274 -2022 2280 -2016
rect 2274 -2028 2280 -2022
rect 2274 -2034 2280 -2028
rect 2274 -2040 2280 -2034
rect 2274 -2046 2280 -2040
rect 2274 -2052 2280 -2046
rect 2274 -2058 2280 -2052
rect 2274 -2064 2280 -2058
rect 2274 -2070 2280 -2064
rect 2274 -2076 2280 -2070
rect 2274 -2082 2280 -2076
rect 2274 -2088 2280 -2082
rect 2274 -2094 2280 -2088
rect 2274 -2100 2280 -2094
rect 2274 -2106 2280 -2100
rect 2274 -2112 2280 -2106
rect 2274 -2118 2280 -2112
rect 2274 -2124 2280 -2118
rect 2274 -2130 2280 -2124
rect 2274 -2136 2280 -2130
rect 2274 -2142 2280 -2136
rect 2274 -2148 2280 -2142
rect 2274 -2154 2280 -2148
rect 2274 -2160 2280 -2154
rect 2274 -2166 2280 -2160
rect 2274 -2172 2280 -2166
rect 2274 -2178 2280 -2172
rect 2274 -2184 2280 -2178
rect 2274 -2190 2280 -2184
rect 2274 -2196 2280 -2190
rect 2274 -2202 2280 -2196
rect 2274 -2208 2280 -2202
rect 2274 -2214 2280 -2208
rect 2274 -2220 2280 -2214
rect 2274 -2226 2280 -2220
rect 2274 -2232 2280 -2226
rect 2274 -2238 2280 -2232
rect 2274 -2244 2280 -2238
rect 2274 -2250 2280 -2244
rect 2274 -2322 2280 -2316
rect 2274 -2328 2280 -2322
rect 2274 -2334 2280 -2328
rect 2274 -2340 2280 -2334
rect 2274 -2346 2280 -2340
rect 2274 -2352 2280 -2346
rect 2274 -2358 2280 -2352
rect 2274 -2364 2280 -2358
rect 2274 -2370 2280 -2364
rect 2274 -2376 2280 -2370
rect 2274 -2382 2280 -2376
rect 2274 -2388 2280 -2382
rect 2274 -2394 2280 -2388
rect 2274 -2400 2280 -2394
rect 2274 -2406 2280 -2400
rect 2274 -2412 2280 -2406
rect 2274 -2418 2280 -2412
rect 2274 -2424 2280 -2418
rect 2274 -2430 2280 -2424
rect 2274 -2436 2280 -2430
rect 2274 -2442 2280 -2436
rect 2274 -2448 2280 -2442
rect 2274 -2454 2280 -2448
rect 2274 -2514 2280 -2508
rect 2274 -2520 2280 -2514
rect 2274 -2526 2280 -2520
rect 2274 -2532 2280 -2526
rect 2274 -2538 2280 -2532
rect 2274 -2544 2280 -2538
rect 2274 -2550 2280 -2544
rect 2274 -2556 2280 -2550
rect 2274 -2562 2280 -2556
rect 2274 -2568 2280 -2562
rect 2274 -2574 2280 -2568
rect 2274 -2580 2280 -2574
rect 2274 -2586 2280 -2580
rect 2274 -2592 2280 -2586
rect 2274 -2598 2280 -2592
rect 2274 -2604 2280 -2598
rect 2274 -2610 2280 -2604
rect 2274 -2616 2280 -2610
rect 2274 -2622 2280 -2616
rect 2274 -2628 2280 -2622
rect 2274 -2634 2280 -2628
rect 2274 -2640 2280 -2634
rect 2274 -2646 2280 -2640
rect 2274 -2652 2280 -2646
rect 2274 -2658 2280 -2652
rect 2274 -2664 2280 -2658
rect 2274 -2670 2280 -2664
rect 2274 -2676 2280 -2670
rect 2274 -2682 2280 -2676
rect 2274 -2688 2280 -2682
rect 2274 -2694 2280 -2688
rect 2274 -2700 2280 -2694
rect 2274 -2706 2280 -2700
rect 2274 -2712 2280 -2706
rect 2274 -2718 2280 -2712
rect 2274 -2724 2280 -2718
rect 2274 -2730 2280 -2724
rect 2274 -2736 2280 -2730
rect 2274 -2742 2280 -2736
rect 2274 -2748 2280 -2742
rect 2274 -2754 2280 -2748
rect 2274 -2760 2280 -2754
rect 2274 -2766 2280 -2760
rect 2274 -2772 2280 -2766
rect 2274 -2778 2280 -2772
rect 2274 -2784 2280 -2778
rect 2274 -2790 2280 -2784
rect 2274 -2796 2280 -2790
rect 2274 -2802 2280 -2796
rect 2274 -2808 2280 -2802
rect 2274 -2814 2280 -2808
rect 2274 -2820 2280 -2814
rect 2274 -2826 2280 -2820
rect 2274 -2832 2280 -2826
rect 2274 -2838 2280 -2832
rect 2274 -2844 2280 -2838
rect 2274 -2850 2280 -2844
rect 2274 -2856 2280 -2850
rect 2274 -2862 2280 -2856
rect 2274 -2868 2280 -2862
rect 2274 -2874 2280 -2868
rect 2274 -2880 2280 -2874
rect 2274 -2886 2280 -2880
rect 2274 -2892 2280 -2886
rect 2274 -2898 2280 -2892
rect 2274 -2904 2280 -2898
rect 2274 -2910 2280 -2904
rect 2274 -2916 2280 -2910
rect 2274 -2922 2280 -2916
rect 2274 -2928 2280 -2922
rect 2274 -2934 2280 -2928
rect 2274 -2940 2280 -2934
rect 2274 -2946 2280 -2940
rect 2274 -2952 2280 -2946
rect 2274 -2958 2280 -2952
rect 2274 -2964 2280 -2958
rect 2280 -102 2286 -96
rect 2280 -108 2286 -102
rect 2280 -114 2286 -108
rect 2280 -120 2286 -114
rect 2280 -126 2286 -120
rect 2280 -132 2286 -126
rect 2280 -138 2286 -132
rect 2280 -144 2286 -138
rect 2280 -150 2286 -144
rect 2280 -156 2286 -150
rect 2280 -162 2286 -156
rect 2280 -168 2286 -162
rect 2280 -174 2286 -168
rect 2280 -180 2286 -174
rect 2280 -186 2286 -180
rect 2280 -192 2286 -186
rect 2280 -198 2286 -192
rect 2280 -204 2286 -198
rect 2280 -210 2286 -204
rect 2280 -216 2286 -210
rect 2280 -222 2286 -216
rect 2280 -228 2286 -222
rect 2280 -234 2286 -228
rect 2280 -240 2286 -234
rect 2280 -246 2286 -240
rect 2280 -252 2286 -246
rect 2280 -258 2286 -252
rect 2280 -264 2286 -258
rect 2280 -270 2286 -264
rect 2280 -276 2286 -270
rect 2280 -282 2286 -276
rect 2280 -288 2286 -282
rect 2280 -294 2286 -288
rect 2280 -300 2286 -294
rect 2280 -306 2286 -300
rect 2280 -312 2286 -306
rect 2280 -318 2286 -312
rect 2280 -324 2286 -318
rect 2280 -330 2286 -324
rect 2280 -336 2286 -330
rect 2280 -342 2286 -336
rect 2280 -348 2286 -342
rect 2280 -354 2286 -348
rect 2280 -360 2286 -354
rect 2280 -366 2286 -360
rect 2280 -372 2286 -366
rect 2280 -378 2286 -372
rect 2280 -384 2286 -378
rect 2280 -390 2286 -384
rect 2280 -396 2286 -390
rect 2280 -402 2286 -396
rect 2280 -408 2286 -402
rect 2280 -414 2286 -408
rect 2280 -420 2286 -414
rect 2280 -426 2286 -420
rect 2280 -432 2286 -426
rect 2280 -438 2286 -432
rect 2280 -444 2286 -438
rect 2280 -450 2286 -444
rect 2280 -456 2286 -450
rect 2280 -462 2286 -456
rect 2280 -468 2286 -462
rect 2280 -474 2286 -468
rect 2280 -480 2286 -474
rect 2280 -486 2286 -480
rect 2280 -492 2286 -486
rect 2280 -498 2286 -492
rect 2280 -504 2286 -498
rect 2280 -510 2286 -504
rect 2280 -516 2286 -510
rect 2280 -522 2286 -516
rect 2280 -528 2286 -522
rect 2280 -534 2286 -528
rect 2280 -540 2286 -534
rect 2280 -546 2286 -540
rect 2280 -552 2286 -546
rect 2280 -558 2286 -552
rect 2280 -564 2286 -558
rect 2280 -570 2286 -564
rect 2280 -576 2286 -570
rect 2280 -582 2286 -576
rect 2280 -588 2286 -582
rect 2280 -594 2286 -588
rect 2280 -600 2286 -594
rect 2280 -606 2286 -600
rect 2280 -612 2286 -606
rect 2280 -618 2286 -612
rect 2280 -624 2286 -618
rect 2280 -630 2286 -624
rect 2280 -636 2286 -630
rect 2280 -642 2286 -636
rect 2280 -648 2286 -642
rect 2280 -654 2286 -648
rect 2280 -660 2286 -654
rect 2280 -666 2286 -660
rect 2280 -672 2286 -666
rect 2280 -678 2286 -672
rect 2280 -684 2286 -678
rect 2280 -690 2286 -684
rect 2280 -696 2286 -690
rect 2280 -702 2286 -696
rect 2280 -708 2286 -702
rect 2280 -714 2286 -708
rect 2280 -720 2286 -714
rect 2280 -726 2286 -720
rect 2280 -732 2286 -726
rect 2280 -738 2286 -732
rect 2280 -744 2286 -738
rect 2280 -750 2286 -744
rect 2280 -756 2286 -750
rect 2280 -762 2286 -756
rect 2280 -768 2286 -762
rect 2280 -774 2286 -768
rect 2280 -780 2286 -774
rect 2280 -786 2286 -780
rect 2280 -792 2286 -786
rect 2280 -798 2286 -792
rect 2280 -804 2286 -798
rect 2280 -810 2286 -804
rect 2280 -816 2286 -810
rect 2280 -822 2286 -816
rect 2280 -828 2286 -822
rect 2280 -834 2286 -828
rect 2280 -840 2286 -834
rect 2280 -846 2286 -840
rect 2280 -852 2286 -846
rect 2280 -858 2286 -852
rect 2280 -864 2286 -858
rect 2280 -870 2286 -864
rect 2280 -876 2286 -870
rect 2280 -882 2286 -876
rect 2280 -888 2286 -882
rect 2280 -894 2286 -888
rect 2280 -900 2286 -894
rect 2280 -906 2286 -900
rect 2280 -912 2286 -906
rect 2280 -918 2286 -912
rect 2280 -924 2286 -918
rect 2280 -930 2286 -924
rect 2280 -936 2286 -930
rect 2280 -942 2286 -936
rect 2280 -948 2286 -942
rect 2280 -954 2286 -948
rect 2280 -960 2286 -954
rect 2280 -966 2286 -960
rect 2280 -972 2286 -966
rect 2280 -978 2286 -972
rect 2280 -984 2286 -978
rect 2280 -990 2286 -984
rect 2280 -996 2286 -990
rect 2280 -1002 2286 -996
rect 2280 -1008 2286 -1002
rect 2280 -1014 2286 -1008
rect 2280 -1020 2286 -1014
rect 2280 -1026 2286 -1020
rect 2280 -1032 2286 -1026
rect 2280 -1038 2286 -1032
rect 2280 -1044 2286 -1038
rect 2280 -1482 2286 -1476
rect 2280 -1488 2286 -1482
rect 2280 -1494 2286 -1488
rect 2280 -1500 2286 -1494
rect 2280 -1506 2286 -1500
rect 2280 -1512 2286 -1506
rect 2280 -1518 2286 -1512
rect 2280 -1524 2286 -1518
rect 2280 -1530 2286 -1524
rect 2280 -1536 2286 -1530
rect 2280 -1542 2286 -1536
rect 2280 -1548 2286 -1542
rect 2280 -1554 2286 -1548
rect 2280 -1560 2286 -1554
rect 2280 -1566 2286 -1560
rect 2280 -1572 2286 -1566
rect 2280 -1578 2286 -1572
rect 2280 -1584 2286 -1578
rect 2280 -1590 2286 -1584
rect 2280 -1596 2286 -1590
rect 2280 -1602 2286 -1596
rect 2280 -1608 2286 -1602
rect 2280 -1614 2286 -1608
rect 2280 -1620 2286 -1614
rect 2280 -1626 2286 -1620
rect 2280 -1632 2286 -1626
rect 2280 -1638 2286 -1632
rect 2280 -1644 2286 -1638
rect 2280 -1650 2286 -1644
rect 2280 -1656 2286 -1650
rect 2280 -1662 2286 -1656
rect 2280 -1668 2286 -1662
rect 2280 -1674 2286 -1668
rect 2280 -1680 2286 -1674
rect 2280 -1686 2286 -1680
rect 2280 -1692 2286 -1686
rect 2280 -1698 2286 -1692
rect 2280 -1704 2286 -1698
rect 2280 -1710 2286 -1704
rect 2280 -1716 2286 -1710
rect 2280 -1722 2286 -1716
rect 2280 -1728 2286 -1722
rect 2280 -1734 2286 -1728
rect 2280 -1740 2286 -1734
rect 2280 -1746 2286 -1740
rect 2280 -1752 2286 -1746
rect 2280 -1758 2286 -1752
rect 2280 -1764 2286 -1758
rect 2280 -1770 2286 -1764
rect 2280 -1776 2286 -1770
rect 2280 -1782 2286 -1776
rect 2280 -1788 2286 -1782
rect 2280 -1794 2286 -1788
rect 2280 -1800 2286 -1794
rect 2280 -1806 2286 -1800
rect 2280 -1812 2286 -1806
rect 2280 -1818 2286 -1812
rect 2280 -1824 2286 -1818
rect 2280 -1830 2286 -1824
rect 2280 -1836 2286 -1830
rect 2280 -1842 2286 -1836
rect 2280 -1848 2286 -1842
rect 2280 -1854 2286 -1848
rect 2280 -1860 2286 -1854
rect 2280 -1866 2286 -1860
rect 2280 -1872 2286 -1866
rect 2280 -1878 2286 -1872
rect 2280 -1884 2286 -1878
rect 2280 -1890 2286 -1884
rect 2280 -1896 2286 -1890
rect 2280 -1902 2286 -1896
rect 2280 -1908 2286 -1902
rect 2280 -1914 2286 -1908
rect 2280 -1920 2286 -1914
rect 2280 -1926 2286 -1920
rect 2280 -1932 2286 -1926
rect 2280 -1938 2286 -1932
rect 2280 -1944 2286 -1938
rect 2280 -1950 2286 -1944
rect 2280 -1956 2286 -1950
rect 2280 -1962 2286 -1956
rect 2280 -1968 2286 -1962
rect 2280 -1974 2286 -1968
rect 2280 -1980 2286 -1974
rect 2280 -1986 2286 -1980
rect 2280 -1992 2286 -1986
rect 2280 -1998 2286 -1992
rect 2280 -2004 2286 -1998
rect 2280 -2010 2286 -2004
rect 2280 -2016 2286 -2010
rect 2280 -2022 2286 -2016
rect 2280 -2028 2286 -2022
rect 2280 -2034 2286 -2028
rect 2280 -2040 2286 -2034
rect 2280 -2046 2286 -2040
rect 2280 -2052 2286 -2046
rect 2280 -2058 2286 -2052
rect 2280 -2064 2286 -2058
rect 2280 -2070 2286 -2064
rect 2280 -2076 2286 -2070
rect 2280 -2082 2286 -2076
rect 2280 -2088 2286 -2082
rect 2280 -2094 2286 -2088
rect 2280 -2100 2286 -2094
rect 2280 -2106 2286 -2100
rect 2280 -2112 2286 -2106
rect 2280 -2118 2286 -2112
rect 2280 -2124 2286 -2118
rect 2280 -2130 2286 -2124
rect 2280 -2136 2286 -2130
rect 2280 -2142 2286 -2136
rect 2280 -2148 2286 -2142
rect 2280 -2154 2286 -2148
rect 2280 -2160 2286 -2154
rect 2280 -2166 2286 -2160
rect 2280 -2172 2286 -2166
rect 2280 -2178 2286 -2172
rect 2280 -2184 2286 -2178
rect 2280 -2190 2286 -2184
rect 2280 -2196 2286 -2190
rect 2280 -2202 2286 -2196
rect 2280 -2208 2286 -2202
rect 2280 -2214 2286 -2208
rect 2280 -2220 2286 -2214
rect 2280 -2226 2286 -2220
rect 2280 -2232 2286 -2226
rect 2280 -2238 2286 -2232
rect 2280 -2244 2286 -2238
rect 2280 -2316 2286 -2310
rect 2280 -2322 2286 -2316
rect 2280 -2328 2286 -2322
rect 2280 -2334 2286 -2328
rect 2280 -2340 2286 -2334
rect 2280 -2346 2286 -2340
rect 2280 -2352 2286 -2346
rect 2280 -2358 2286 -2352
rect 2280 -2364 2286 -2358
rect 2280 -2370 2286 -2364
rect 2280 -2376 2286 -2370
rect 2280 -2382 2286 -2376
rect 2280 -2388 2286 -2382
rect 2280 -2394 2286 -2388
rect 2280 -2400 2286 -2394
rect 2280 -2406 2286 -2400
rect 2280 -2412 2286 -2406
rect 2280 -2418 2286 -2412
rect 2280 -2424 2286 -2418
rect 2280 -2430 2286 -2424
rect 2280 -2436 2286 -2430
rect 2280 -2442 2286 -2436
rect 2280 -2448 2286 -2442
rect 2280 -2514 2286 -2508
rect 2280 -2520 2286 -2514
rect 2280 -2526 2286 -2520
rect 2280 -2532 2286 -2526
rect 2280 -2538 2286 -2532
rect 2280 -2544 2286 -2538
rect 2280 -2550 2286 -2544
rect 2280 -2556 2286 -2550
rect 2280 -2562 2286 -2556
rect 2280 -2568 2286 -2562
rect 2280 -2574 2286 -2568
rect 2280 -2580 2286 -2574
rect 2280 -2586 2286 -2580
rect 2280 -2592 2286 -2586
rect 2280 -2598 2286 -2592
rect 2280 -2604 2286 -2598
rect 2280 -2610 2286 -2604
rect 2280 -2616 2286 -2610
rect 2280 -2622 2286 -2616
rect 2280 -2628 2286 -2622
rect 2280 -2634 2286 -2628
rect 2280 -2640 2286 -2634
rect 2280 -2646 2286 -2640
rect 2280 -2652 2286 -2646
rect 2280 -2658 2286 -2652
rect 2280 -2664 2286 -2658
rect 2280 -2670 2286 -2664
rect 2280 -2676 2286 -2670
rect 2280 -2682 2286 -2676
rect 2280 -2688 2286 -2682
rect 2280 -2694 2286 -2688
rect 2280 -2700 2286 -2694
rect 2280 -2706 2286 -2700
rect 2280 -2712 2286 -2706
rect 2280 -2718 2286 -2712
rect 2280 -2724 2286 -2718
rect 2280 -2730 2286 -2724
rect 2280 -2736 2286 -2730
rect 2280 -2742 2286 -2736
rect 2280 -2748 2286 -2742
rect 2280 -2754 2286 -2748
rect 2280 -2760 2286 -2754
rect 2280 -2766 2286 -2760
rect 2280 -2772 2286 -2766
rect 2280 -2778 2286 -2772
rect 2280 -2784 2286 -2778
rect 2280 -2790 2286 -2784
rect 2280 -2796 2286 -2790
rect 2280 -2802 2286 -2796
rect 2280 -2808 2286 -2802
rect 2280 -2814 2286 -2808
rect 2280 -2820 2286 -2814
rect 2280 -2826 2286 -2820
rect 2280 -2832 2286 -2826
rect 2280 -2838 2286 -2832
rect 2280 -2844 2286 -2838
rect 2280 -2850 2286 -2844
rect 2280 -2856 2286 -2850
rect 2280 -2862 2286 -2856
rect 2280 -2868 2286 -2862
rect 2280 -2874 2286 -2868
rect 2280 -2880 2286 -2874
rect 2280 -2886 2286 -2880
rect 2280 -2892 2286 -2886
rect 2280 -2898 2286 -2892
rect 2280 -2904 2286 -2898
rect 2280 -2910 2286 -2904
rect 2280 -2916 2286 -2910
rect 2280 -2922 2286 -2916
rect 2280 -2928 2286 -2922
rect 2280 -2934 2286 -2928
rect 2280 -2940 2286 -2934
rect 2280 -2946 2286 -2940
rect 2280 -2952 2286 -2946
rect 2280 -2958 2286 -2952
rect 2286 -90 2292 -84
rect 2286 -96 2292 -90
rect 2286 -102 2292 -96
rect 2286 -108 2292 -102
rect 2286 -114 2292 -108
rect 2286 -120 2292 -114
rect 2286 -126 2292 -120
rect 2286 -132 2292 -126
rect 2286 -138 2292 -132
rect 2286 -144 2292 -138
rect 2286 -150 2292 -144
rect 2286 -156 2292 -150
rect 2286 -162 2292 -156
rect 2286 -168 2292 -162
rect 2286 -174 2292 -168
rect 2286 -180 2292 -174
rect 2286 -186 2292 -180
rect 2286 -192 2292 -186
rect 2286 -198 2292 -192
rect 2286 -204 2292 -198
rect 2286 -210 2292 -204
rect 2286 -216 2292 -210
rect 2286 -222 2292 -216
rect 2286 -228 2292 -222
rect 2286 -234 2292 -228
rect 2286 -240 2292 -234
rect 2286 -246 2292 -240
rect 2286 -252 2292 -246
rect 2286 -258 2292 -252
rect 2286 -264 2292 -258
rect 2286 -270 2292 -264
rect 2286 -276 2292 -270
rect 2286 -282 2292 -276
rect 2286 -288 2292 -282
rect 2286 -294 2292 -288
rect 2286 -300 2292 -294
rect 2286 -306 2292 -300
rect 2286 -312 2292 -306
rect 2286 -318 2292 -312
rect 2286 -324 2292 -318
rect 2286 -330 2292 -324
rect 2286 -336 2292 -330
rect 2286 -342 2292 -336
rect 2286 -348 2292 -342
rect 2286 -354 2292 -348
rect 2286 -360 2292 -354
rect 2286 -366 2292 -360
rect 2286 -372 2292 -366
rect 2286 -378 2292 -372
rect 2286 -384 2292 -378
rect 2286 -390 2292 -384
rect 2286 -396 2292 -390
rect 2286 -402 2292 -396
rect 2286 -408 2292 -402
rect 2286 -414 2292 -408
rect 2286 -420 2292 -414
rect 2286 -426 2292 -420
rect 2286 -432 2292 -426
rect 2286 -438 2292 -432
rect 2286 -444 2292 -438
rect 2286 -450 2292 -444
rect 2286 -456 2292 -450
rect 2286 -462 2292 -456
rect 2286 -468 2292 -462
rect 2286 -474 2292 -468
rect 2286 -480 2292 -474
rect 2286 -486 2292 -480
rect 2286 -492 2292 -486
rect 2286 -498 2292 -492
rect 2286 -504 2292 -498
rect 2286 -510 2292 -504
rect 2286 -516 2292 -510
rect 2286 -522 2292 -516
rect 2286 -528 2292 -522
rect 2286 -534 2292 -528
rect 2286 -540 2292 -534
rect 2286 -546 2292 -540
rect 2286 -552 2292 -546
rect 2286 -558 2292 -552
rect 2286 -564 2292 -558
rect 2286 -570 2292 -564
rect 2286 -576 2292 -570
rect 2286 -582 2292 -576
rect 2286 -588 2292 -582
rect 2286 -594 2292 -588
rect 2286 -600 2292 -594
rect 2286 -606 2292 -600
rect 2286 -612 2292 -606
rect 2286 -618 2292 -612
rect 2286 -624 2292 -618
rect 2286 -630 2292 -624
rect 2286 -636 2292 -630
rect 2286 -642 2292 -636
rect 2286 -648 2292 -642
rect 2286 -654 2292 -648
rect 2286 -660 2292 -654
rect 2286 -666 2292 -660
rect 2286 -672 2292 -666
rect 2286 -678 2292 -672
rect 2286 -684 2292 -678
rect 2286 -690 2292 -684
rect 2286 -696 2292 -690
rect 2286 -702 2292 -696
rect 2286 -708 2292 -702
rect 2286 -714 2292 -708
rect 2286 -720 2292 -714
rect 2286 -726 2292 -720
rect 2286 -732 2292 -726
rect 2286 -738 2292 -732
rect 2286 -744 2292 -738
rect 2286 -750 2292 -744
rect 2286 -756 2292 -750
rect 2286 -762 2292 -756
rect 2286 -768 2292 -762
rect 2286 -774 2292 -768
rect 2286 -780 2292 -774
rect 2286 -786 2292 -780
rect 2286 -792 2292 -786
rect 2286 -798 2292 -792
rect 2286 -804 2292 -798
rect 2286 -810 2292 -804
rect 2286 -816 2292 -810
rect 2286 -822 2292 -816
rect 2286 -828 2292 -822
rect 2286 -834 2292 -828
rect 2286 -840 2292 -834
rect 2286 -846 2292 -840
rect 2286 -852 2292 -846
rect 2286 -858 2292 -852
rect 2286 -864 2292 -858
rect 2286 -870 2292 -864
rect 2286 -876 2292 -870
rect 2286 -882 2292 -876
rect 2286 -888 2292 -882
rect 2286 -894 2292 -888
rect 2286 -900 2292 -894
rect 2286 -906 2292 -900
rect 2286 -912 2292 -906
rect 2286 -918 2292 -912
rect 2286 -924 2292 -918
rect 2286 -930 2292 -924
rect 2286 -936 2292 -930
rect 2286 -942 2292 -936
rect 2286 -948 2292 -942
rect 2286 -954 2292 -948
rect 2286 -960 2292 -954
rect 2286 -966 2292 -960
rect 2286 -972 2292 -966
rect 2286 -978 2292 -972
rect 2286 -984 2292 -978
rect 2286 -990 2292 -984
rect 2286 -996 2292 -990
rect 2286 -1002 2292 -996
rect 2286 -1008 2292 -1002
rect 2286 -1014 2292 -1008
rect 2286 -1020 2292 -1014
rect 2286 -1026 2292 -1020
rect 2286 -1482 2292 -1476
rect 2286 -1488 2292 -1482
rect 2286 -1494 2292 -1488
rect 2286 -1500 2292 -1494
rect 2286 -1506 2292 -1500
rect 2286 -1512 2292 -1506
rect 2286 -1518 2292 -1512
rect 2286 -1524 2292 -1518
rect 2286 -1530 2292 -1524
rect 2286 -1536 2292 -1530
rect 2286 -1542 2292 -1536
rect 2286 -1548 2292 -1542
rect 2286 -1554 2292 -1548
rect 2286 -1560 2292 -1554
rect 2286 -1566 2292 -1560
rect 2286 -1572 2292 -1566
rect 2286 -1578 2292 -1572
rect 2286 -1584 2292 -1578
rect 2286 -1590 2292 -1584
rect 2286 -1596 2292 -1590
rect 2286 -1602 2292 -1596
rect 2286 -1608 2292 -1602
rect 2286 -1614 2292 -1608
rect 2286 -1620 2292 -1614
rect 2286 -1626 2292 -1620
rect 2286 -1632 2292 -1626
rect 2286 -1638 2292 -1632
rect 2286 -1644 2292 -1638
rect 2286 -1650 2292 -1644
rect 2286 -1656 2292 -1650
rect 2286 -1662 2292 -1656
rect 2286 -1668 2292 -1662
rect 2286 -1674 2292 -1668
rect 2286 -1680 2292 -1674
rect 2286 -1686 2292 -1680
rect 2286 -1692 2292 -1686
rect 2286 -1698 2292 -1692
rect 2286 -1704 2292 -1698
rect 2286 -1710 2292 -1704
rect 2286 -1716 2292 -1710
rect 2286 -1722 2292 -1716
rect 2286 -1728 2292 -1722
rect 2286 -1734 2292 -1728
rect 2286 -1740 2292 -1734
rect 2286 -1746 2292 -1740
rect 2286 -1752 2292 -1746
rect 2286 -1758 2292 -1752
rect 2286 -1764 2292 -1758
rect 2286 -1770 2292 -1764
rect 2286 -1776 2292 -1770
rect 2286 -1782 2292 -1776
rect 2286 -1788 2292 -1782
rect 2286 -1794 2292 -1788
rect 2286 -1800 2292 -1794
rect 2286 -1806 2292 -1800
rect 2286 -1812 2292 -1806
rect 2286 -1818 2292 -1812
rect 2286 -1824 2292 -1818
rect 2286 -1830 2292 -1824
rect 2286 -1836 2292 -1830
rect 2286 -1842 2292 -1836
rect 2286 -1848 2292 -1842
rect 2286 -1854 2292 -1848
rect 2286 -1860 2292 -1854
rect 2286 -1866 2292 -1860
rect 2286 -1872 2292 -1866
rect 2286 -1878 2292 -1872
rect 2286 -1884 2292 -1878
rect 2286 -1890 2292 -1884
rect 2286 -1896 2292 -1890
rect 2286 -1902 2292 -1896
rect 2286 -1908 2292 -1902
rect 2286 -1914 2292 -1908
rect 2286 -1920 2292 -1914
rect 2286 -1926 2292 -1920
rect 2286 -1932 2292 -1926
rect 2286 -1938 2292 -1932
rect 2286 -1944 2292 -1938
rect 2286 -1950 2292 -1944
rect 2286 -1956 2292 -1950
rect 2286 -1962 2292 -1956
rect 2286 -1968 2292 -1962
rect 2286 -1974 2292 -1968
rect 2286 -1980 2292 -1974
rect 2286 -1986 2292 -1980
rect 2286 -1992 2292 -1986
rect 2286 -1998 2292 -1992
rect 2286 -2004 2292 -1998
rect 2286 -2010 2292 -2004
rect 2286 -2016 2292 -2010
rect 2286 -2022 2292 -2016
rect 2286 -2028 2292 -2022
rect 2286 -2034 2292 -2028
rect 2286 -2040 2292 -2034
rect 2286 -2046 2292 -2040
rect 2286 -2052 2292 -2046
rect 2286 -2058 2292 -2052
rect 2286 -2064 2292 -2058
rect 2286 -2070 2292 -2064
rect 2286 -2076 2292 -2070
rect 2286 -2082 2292 -2076
rect 2286 -2088 2292 -2082
rect 2286 -2094 2292 -2088
rect 2286 -2100 2292 -2094
rect 2286 -2106 2292 -2100
rect 2286 -2112 2292 -2106
rect 2286 -2118 2292 -2112
rect 2286 -2124 2292 -2118
rect 2286 -2130 2292 -2124
rect 2286 -2136 2292 -2130
rect 2286 -2142 2292 -2136
rect 2286 -2148 2292 -2142
rect 2286 -2154 2292 -2148
rect 2286 -2160 2292 -2154
rect 2286 -2166 2292 -2160
rect 2286 -2172 2292 -2166
rect 2286 -2178 2292 -2172
rect 2286 -2184 2292 -2178
rect 2286 -2190 2292 -2184
rect 2286 -2196 2292 -2190
rect 2286 -2202 2292 -2196
rect 2286 -2208 2292 -2202
rect 2286 -2214 2292 -2208
rect 2286 -2220 2292 -2214
rect 2286 -2226 2292 -2220
rect 2286 -2232 2292 -2226
rect 2286 -2238 2292 -2232
rect 2286 -2310 2292 -2304
rect 2286 -2316 2292 -2310
rect 2286 -2322 2292 -2316
rect 2286 -2328 2292 -2322
rect 2286 -2334 2292 -2328
rect 2286 -2340 2292 -2334
rect 2286 -2346 2292 -2340
rect 2286 -2352 2292 -2346
rect 2286 -2358 2292 -2352
rect 2286 -2364 2292 -2358
rect 2286 -2370 2292 -2364
rect 2286 -2376 2292 -2370
rect 2286 -2382 2292 -2376
rect 2286 -2388 2292 -2382
rect 2286 -2394 2292 -2388
rect 2286 -2400 2292 -2394
rect 2286 -2406 2292 -2400
rect 2286 -2412 2292 -2406
rect 2286 -2418 2292 -2412
rect 2286 -2424 2292 -2418
rect 2286 -2430 2292 -2424
rect 2286 -2436 2292 -2430
rect 2286 -2442 2292 -2436
rect 2286 -2448 2292 -2442
rect 2286 -2508 2292 -2502
rect 2286 -2514 2292 -2508
rect 2286 -2520 2292 -2514
rect 2286 -2526 2292 -2520
rect 2286 -2532 2292 -2526
rect 2286 -2538 2292 -2532
rect 2286 -2544 2292 -2538
rect 2286 -2550 2292 -2544
rect 2286 -2556 2292 -2550
rect 2286 -2562 2292 -2556
rect 2286 -2568 2292 -2562
rect 2286 -2574 2292 -2568
rect 2286 -2580 2292 -2574
rect 2286 -2586 2292 -2580
rect 2286 -2592 2292 -2586
rect 2286 -2598 2292 -2592
rect 2286 -2604 2292 -2598
rect 2286 -2610 2292 -2604
rect 2286 -2616 2292 -2610
rect 2286 -2622 2292 -2616
rect 2286 -2628 2292 -2622
rect 2286 -2634 2292 -2628
rect 2286 -2640 2292 -2634
rect 2286 -2646 2292 -2640
rect 2286 -2652 2292 -2646
rect 2286 -2658 2292 -2652
rect 2286 -2664 2292 -2658
rect 2286 -2670 2292 -2664
rect 2286 -2676 2292 -2670
rect 2286 -2682 2292 -2676
rect 2286 -2688 2292 -2682
rect 2286 -2694 2292 -2688
rect 2286 -2700 2292 -2694
rect 2286 -2706 2292 -2700
rect 2286 -2712 2292 -2706
rect 2286 -2718 2292 -2712
rect 2286 -2724 2292 -2718
rect 2286 -2730 2292 -2724
rect 2286 -2736 2292 -2730
rect 2286 -2742 2292 -2736
rect 2286 -2748 2292 -2742
rect 2286 -2754 2292 -2748
rect 2286 -2760 2292 -2754
rect 2286 -2766 2292 -2760
rect 2286 -2772 2292 -2766
rect 2286 -2778 2292 -2772
rect 2286 -2784 2292 -2778
rect 2286 -2790 2292 -2784
rect 2286 -2796 2292 -2790
rect 2286 -2802 2292 -2796
rect 2286 -2808 2292 -2802
rect 2286 -2814 2292 -2808
rect 2286 -2820 2292 -2814
rect 2286 -2826 2292 -2820
rect 2286 -2832 2292 -2826
rect 2286 -2838 2292 -2832
rect 2286 -2844 2292 -2838
rect 2286 -2850 2292 -2844
rect 2286 -2856 2292 -2850
rect 2286 -2862 2292 -2856
rect 2286 -2868 2292 -2862
rect 2286 -2874 2292 -2868
rect 2286 -2880 2292 -2874
rect 2286 -2886 2292 -2880
rect 2286 -2892 2292 -2886
rect 2286 -2898 2292 -2892
rect 2286 -2904 2292 -2898
rect 2286 -2910 2292 -2904
rect 2286 -2916 2292 -2910
rect 2286 -2922 2292 -2916
rect 2286 -2928 2292 -2922
rect 2286 -2934 2292 -2928
rect 2286 -2940 2292 -2934
rect 2286 -2946 2292 -2940
rect 2286 -2952 2292 -2946
rect 2292 -84 2298 -78
rect 2292 -90 2298 -84
rect 2292 -96 2298 -90
rect 2292 -102 2298 -96
rect 2292 -108 2298 -102
rect 2292 -114 2298 -108
rect 2292 -120 2298 -114
rect 2292 -126 2298 -120
rect 2292 -132 2298 -126
rect 2292 -138 2298 -132
rect 2292 -144 2298 -138
rect 2292 -150 2298 -144
rect 2292 -156 2298 -150
rect 2292 -162 2298 -156
rect 2292 -168 2298 -162
rect 2292 -174 2298 -168
rect 2292 -180 2298 -174
rect 2292 -186 2298 -180
rect 2292 -192 2298 -186
rect 2292 -198 2298 -192
rect 2292 -204 2298 -198
rect 2292 -210 2298 -204
rect 2292 -216 2298 -210
rect 2292 -222 2298 -216
rect 2292 -228 2298 -222
rect 2292 -234 2298 -228
rect 2292 -240 2298 -234
rect 2292 -246 2298 -240
rect 2292 -252 2298 -246
rect 2292 -258 2298 -252
rect 2292 -264 2298 -258
rect 2292 -270 2298 -264
rect 2292 -276 2298 -270
rect 2292 -282 2298 -276
rect 2292 -288 2298 -282
rect 2292 -294 2298 -288
rect 2292 -300 2298 -294
rect 2292 -306 2298 -300
rect 2292 -312 2298 -306
rect 2292 -318 2298 -312
rect 2292 -324 2298 -318
rect 2292 -330 2298 -324
rect 2292 -336 2298 -330
rect 2292 -342 2298 -336
rect 2292 -348 2298 -342
rect 2292 -354 2298 -348
rect 2292 -360 2298 -354
rect 2292 -366 2298 -360
rect 2292 -372 2298 -366
rect 2292 -378 2298 -372
rect 2292 -384 2298 -378
rect 2292 -390 2298 -384
rect 2292 -396 2298 -390
rect 2292 -402 2298 -396
rect 2292 -408 2298 -402
rect 2292 -414 2298 -408
rect 2292 -420 2298 -414
rect 2292 -426 2298 -420
rect 2292 -432 2298 -426
rect 2292 -438 2298 -432
rect 2292 -444 2298 -438
rect 2292 -450 2298 -444
rect 2292 -456 2298 -450
rect 2292 -462 2298 -456
rect 2292 -468 2298 -462
rect 2292 -474 2298 -468
rect 2292 -480 2298 -474
rect 2292 -486 2298 -480
rect 2292 -492 2298 -486
rect 2292 -498 2298 -492
rect 2292 -504 2298 -498
rect 2292 -510 2298 -504
rect 2292 -516 2298 -510
rect 2292 -522 2298 -516
rect 2292 -528 2298 -522
rect 2292 -534 2298 -528
rect 2292 -540 2298 -534
rect 2292 -546 2298 -540
rect 2292 -552 2298 -546
rect 2292 -558 2298 -552
rect 2292 -564 2298 -558
rect 2292 -570 2298 -564
rect 2292 -576 2298 -570
rect 2292 -582 2298 -576
rect 2292 -588 2298 -582
rect 2292 -594 2298 -588
rect 2292 -600 2298 -594
rect 2292 -606 2298 -600
rect 2292 -612 2298 -606
rect 2292 -618 2298 -612
rect 2292 -624 2298 -618
rect 2292 -630 2298 -624
rect 2292 -636 2298 -630
rect 2292 -642 2298 -636
rect 2292 -648 2298 -642
rect 2292 -654 2298 -648
rect 2292 -660 2298 -654
rect 2292 -666 2298 -660
rect 2292 -672 2298 -666
rect 2292 -678 2298 -672
rect 2292 -684 2298 -678
rect 2292 -690 2298 -684
rect 2292 -696 2298 -690
rect 2292 -702 2298 -696
rect 2292 -708 2298 -702
rect 2292 -714 2298 -708
rect 2292 -720 2298 -714
rect 2292 -726 2298 -720
rect 2292 -732 2298 -726
rect 2292 -738 2298 -732
rect 2292 -744 2298 -738
rect 2292 -750 2298 -744
rect 2292 -756 2298 -750
rect 2292 -762 2298 -756
rect 2292 -768 2298 -762
rect 2292 -774 2298 -768
rect 2292 -780 2298 -774
rect 2292 -786 2298 -780
rect 2292 -792 2298 -786
rect 2292 -798 2298 -792
rect 2292 -804 2298 -798
rect 2292 -810 2298 -804
rect 2292 -816 2298 -810
rect 2292 -822 2298 -816
rect 2292 -828 2298 -822
rect 2292 -834 2298 -828
rect 2292 -840 2298 -834
rect 2292 -846 2298 -840
rect 2292 -852 2298 -846
rect 2292 -858 2298 -852
rect 2292 -864 2298 -858
rect 2292 -870 2298 -864
rect 2292 -876 2298 -870
rect 2292 -882 2298 -876
rect 2292 -888 2298 -882
rect 2292 -894 2298 -888
rect 2292 -900 2298 -894
rect 2292 -906 2298 -900
rect 2292 -912 2298 -906
rect 2292 -918 2298 -912
rect 2292 -924 2298 -918
rect 2292 -930 2298 -924
rect 2292 -936 2298 -930
rect 2292 -942 2298 -936
rect 2292 -948 2298 -942
rect 2292 -954 2298 -948
rect 2292 -960 2298 -954
rect 2292 -966 2298 -960
rect 2292 -972 2298 -966
rect 2292 -978 2298 -972
rect 2292 -984 2298 -978
rect 2292 -990 2298 -984
rect 2292 -996 2298 -990
rect 2292 -1002 2298 -996
rect 2292 -1008 2298 -1002
rect 2292 -1014 2298 -1008
rect 2292 -1476 2298 -1470
rect 2292 -1482 2298 -1476
rect 2292 -1488 2298 -1482
rect 2292 -1494 2298 -1488
rect 2292 -1500 2298 -1494
rect 2292 -1506 2298 -1500
rect 2292 -1512 2298 -1506
rect 2292 -1518 2298 -1512
rect 2292 -1524 2298 -1518
rect 2292 -1530 2298 -1524
rect 2292 -1536 2298 -1530
rect 2292 -1542 2298 -1536
rect 2292 -1548 2298 -1542
rect 2292 -1554 2298 -1548
rect 2292 -1560 2298 -1554
rect 2292 -1566 2298 -1560
rect 2292 -1572 2298 -1566
rect 2292 -1578 2298 -1572
rect 2292 -1584 2298 -1578
rect 2292 -1590 2298 -1584
rect 2292 -1596 2298 -1590
rect 2292 -1602 2298 -1596
rect 2292 -1608 2298 -1602
rect 2292 -1614 2298 -1608
rect 2292 -1620 2298 -1614
rect 2292 -1626 2298 -1620
rect 2292 -1632 2298 -1626
rect 2292 -1638 2298 -1632
rect 2292 -1644 2298 -1638
rect 2292 -1650 2298 -1644
rect 2292 -1656 2298 -1650
rect 2292 -1662 2298 -1656
rect 2292 -1668 2298 -1662
rect 2292 -1674 2298 -1668
rect 2292 -1680 2298 -1674
rect 2292 -1686 2298 -1680
rect 2292 -1692 2298 -1686
rect 2292 -1698 2298 -1692
rect 2292 -1704 2298 -1698
rect 2292 -1710 2298 -1704
rect 2292 -1716 2298 -1710
rect 2292 -1722 2298 -1716
rect 2292 -1728 2298 -1722
rect 2292 -1734 2298 -1728
rect 2292 -1740 2298 -1734
rect 2292 -1746 2298 -1740
rect 2292 -1752 2298 -1746
rect 2292 -1758 2298 -1752
rect 2292 -1764 2298 -1758
rect 2292 -1770 2298 -1764
rect 2292 -1776 2298 -1770
rect 2292 -1782 2298 -1776
rect 2292 -1788 2298 -1782
rect 2292 -1794 2298 -1788
rect 2292 -1800 2298 -1794
rect 2292 -1806 2298 -1800
rect 2292 -1812 2298 -1806
rect 2292 -1818 2298 -1812
rect 2292 -1824 2298 -1818
rect 2292 -1830 2298 -1824
rect 2292 -1836 2298 -1830
rect 2292 -1842 2298 -1836
rect 2292 -1848 2298 -1842
rect 2292 -1854 2298 -1848
rect 2292 -1860 2298 -1854
rect 2292 -1866 2298 -1860
rect 2292 -1872 2298 -1866
rect 2292 -1878 2298 -1872
rect 2292 -1884 2298 -1878
rect 2292 -1890 2298 -1884
rect 2292 -1896 2298 -1890
rect 2292 -1902 2298 -1896
rect 2292 -1908 2298 -1902
rect 2292 -1914 2298 -1908
rect 2292 -1920 2298 -1914
rect 2292 -1926 2298 -1920
rect 2292 -1932 2298 -1926
rect 2292 -1938 2298 -1932
rect 2292 -1944 2298 -1938
rect 2292 -1950 2298 -1944
rect 2292 -1956 2298 -1950
rect 2292 -1962 2298 -1956
rect 2292 -1968 2298 -1962
rect 2292 -1974 2298 -1968
rect 2292 -1980 2298 -1974
rect 2292 -1986 2298 -1980
rect 2292 -1992 2298 -1986
rect 2292 -1998 2298 -1992
rect 2292 -2004 2298 -1998
rect 2292 -2010 2298 -2004
rect 2292 -2016 2298 -2010
rect 2292 -2022 2298 -2016
rect 2292 -2028 2298 -2022
rect 2292 -2034 2298 -2028
rect 2292 -2040 2298 -2034
rect 2292 -2046 2298 -2040
rect 2292 -2052 2298 -2046
rect 2292 -2058 2298 -2052
rect 2292 -2064 2298 -2058
rect 2292 -2070 2298 -2064
rect 2292 -2076 2298 -2070
rect 2292 -2082 2298 -2076
rect 2292 -2088 2298 -2082
rect 2292 -2094 2298 -2088
rect 2292 -2100 2298 -2094
rect 2292 -2106 2298 -2100
rect 2292 -2112 2298 -2106
rect 2292 -2118 2298 -2112
rect 2292 -2124 2298 -2118
rect 2292 -2130 2298 -2124
rect 2292 -2136 2298 -2130
rect 2292 -2142 2298 -2136
rect 2292 -2148 2298 -2142
rect 2292 -2154 2298 -2148
rect 2292 -2160 2298 -2154
rect 2292 -2166 2298 -2160
rect 2292 -2172 2298 -2166
rect 2292 -2178 2298 -2172
rect 2292 -2184 2298 -2178
rect 2292 -2190 2298 -2184
rect 2292 -2196 2298 -2190
rect 2292 -2202 2298 -2196
rect 2292 -2208 2298 -2202
rect 2292 -2214 2298 -2208
rect 2292 -2220 2298 -2214
rect 2292 -2226 2298 -2220
rect 2292 -2232 2298 -2226
rect 2292 -2304 2298 -2298
rect 2292 -2310 2298 -2304
rect 2292 -2316 2298 -2310
rect 2292 -2322 2298 -2316
rect 2292 -2328 2298 -2322
rect 2292 -2334 2298 -2328
rect 2292 -2340 2298 -2334
rect 2292 -2346 2298 -2340
rect 2292 -2352 2298 -2346
rect 2292 -2358 2298 -2352
rect 2292 -2364 2298 -2358
rect 2292 -2370 2298 -2364
rect 2292 -2376 2298 -2370
rect 2292 -2382 2298 -2376
rect 2292 -2388 2298 -2382
rect 2292 -2394 2298 -2388
rect 2292 -2400 2298 -2394
rect 2292 -2406 2298 -2400
rect 2292 -2412 2298 -2406
rect 2292 -2418 2298 -2412
rect 2292 -2424 2298 -2418
rect 2292 -2430 2298 -2424
rect 2292 -2436 2298 -2430
rect 2292 -2442 2298 -2436
rect 2292 -2448 2298 -2442
rect 2292 -2508 2298 -2502
rect 2292 -2514 2298 -2508
rect 2292 -2520 2298 -2514
rect 2292 -2526 2298 -2520
rect 2292 -2532 2298 -2526
rect 2292 -2538 2298 -2532
rect 2292 -2544 2298 -2538
rect 2292 -2550 2298 -2544
rect 2292 -2556 2298 -2550
rect 2292 -2562 2298 -2556
rect 2292 -2568 2298 -2562
rect 2292 -2574 2298 -2568
rect 2292 -2580 2298 -2574
rect 2292 -2586 2298 -2580
rect 2292 -2592 2298 -2586
rect 2292 -2598 2298 -2592
rect 2292 -2604 2298 -2598
rect 2292 -2610 2298 -2604
rect 2292 -2616 2298 -2610
rect 2292 -2622 2298 -2616
rect 2292 -2628 2298 -2622
rect 2292 -2634 2298 -2628
rect 2292 -2640 2298 -2634
rect 2292 -2646 2298 -2640
rect 2292 -2652 2298 -2646
rect 2292 -2658 2298 -2652
rect 2292 -2664 2298 -2658
rect 2292 -2670 2298 -2664
rect 2292 -2676 2298 -2670
rect 2292 -2682 2298 -2676
rect 2292 -2688 2298 -2682
rect 2292 -2694 2298 -2688
rect 2292 -2700 2298 -2694
rect 2292 -2706 2298 -2700
rect 2292 -2712 2298 -2706
rect 2292 -2718 2298 -2712
rect 2292 -2724 2298 -2718
rect 2292 -2730 2298 -2724
rect 2292 -2736 2298 -2730
rect 2292 -2742 2298 -2736
rect 2292 -2748 2298 -2742
rect 2292 -2754 2298 -2748
rect 2292 -2760 2298 -2754
rect 2292 -2766 2298 -2760
rect 2292 -2772 2298 -2766
rect 2292 -2778 2298 -2772
rect 2292 -2784 2298 -2778
rect 2292 -2790 2298 -2784
rect 2292 -2796 2298 -2790
rect 2292 -2802 2298 -2796
rect 2292 -2808 2298 -2802
rect 2292 -2814 2298 -2808
rect 2292 -2820 2298 -2814
rect 2292 -2826 2298 -2820
rect 2292 -2832 2298 -2826
rect 2292 -2838 2298 -2832
rect 2292 -2844 2298 -2838
rect 2292 -2850 2298 -2844
rect 2292 -2856 2298 -2850
rect 2292 -2862 2298 -2856
rect 2292 -2868 2298 -2862
rect 2292 -2874 2298 -2868
rect 2292 -2880 2298 -2874
rect 2292 -2886 2298 -2880
rect 2292 -2892 2298 -2886
rect 2292 -2898 2298 -2892
rect 2292 -2904 2298 -2898
rect 2292 -2910 2298 -2904
rect 2292 -2916 2298 -2910
rect 2292 -2922 2298 -2916
rect 2292 -2928 2298 -2922
rect 2292 -2934 2298 -2928
rect 2292 -2940 2298 -2934
rect 2292 -2946 2298 -2940
rect 2292 -2952 2298 -2946
rect 2298 -78 2304 -72
rect 2298 -84 2304 -78
rect 2298 -90 2304 -84
rect 2298 -96 2304 -90
rect 2298 -102 2304 -96
rect 2298 -108 2304 -102
rect 2298 -114 2304 -108
rect 2298 -120 2304 -114
rect 2298 -126 2304 -120
rect 2298 -132 2304 -126
rect 2298 -138 2304 -132
rect 2298 -144 2304 -138
rect 2298 -150 2304 -144
rect 2298 -156 2304 -150
rect 2298 -162 2304 -156
rect 2298 -168 2304 -162
rect 2298 -174 2304 -168
rect 2298 -180 2304 -174
rect 2298 -186 2304 -180
rect 2298 -192 2304 -186
rect 2298 -198 2304 -192
rect 2298 -204 2304 -198
rect 2298 -210 2304 -204
rect 2298 -216 2304 -210
rect 2298 -222 2304 -216
rect 2298 -228 2304 -222
rect 2298 -234 2304 -228
rect 2298 -240 2304 -234
rect 2298 -246 2304 -240
rect 2298 -252 2304 -246
rect 2298 -258 2304 -252
rect 2298 -264 2304 -258
rect 2298 -270 2304 -264
rect 2298 -276 2304 -270
rect 2298 -282 2304 -276
rect 2298 -288 2304 -282
rect 2298 -294 2304 -288
rect 2298 -300 2304 -294
rect 2298 -306 2304 -300
rect 2298 -312 2304 -306
rect 2298 -318 2304 -312
rect 2298 -324 2304 -318
rect 2298 -330 2304 -324
rect 2298 -336 2304 -330
rect 2298 -342 2304 -336
rect 2298 -348 2304 -342
rect 2298 -354 2304 -348
rect 2298 -360 2304 -354
rect 2298 -366 2304 -360
rect 2298 -372 2304 -366
rect 2298 -378 2304 -372
rect 2298 -384 2304 -378
rect 2298 -390 2304 -384
rect 2298 -396 2304 -390
rect 2298 -402 2304 -396
rect 2298 -408 2304 -402
rect 2298 -414 2304 -408
rect 2298 -420 2304 -414
rect 2298 -426 2304 -420
rect 2298 -432 2304 -426
rect 2298 -438 2304 -432
rect 2298 -444 2304 -438
rect 2298 -450 2304 -444
rect 2298 -456 2304 -450
rect 2298 -462 2304 -456
rect 2298 -468 2304 -462
rect 2298 -474 2304 -468
rect 2298 -480 2304 -474
rect 2298 -486 2304 -480
rect 2298 -492 2304 -486
rect 2298 -498 2304 -492
rect 2298 -504 2304 -498
rect 2298 -510 2304 -504
rect 2298 -516 2304 -510
rect 2298 -522 2304 -516
rect 2298 -528 2304 -522
rect 2298 -534 2304 -528
rect 2298 -540 2304 -534
rect 2298 -546 2304 -540
rect 2298 -552 2304 -546
rect 2298 -558 2304 -552
rect 2298 -564 2304 -558
rect 2298 -570 2304 -564
rect 2298 -576 2304 -570
rect 2298 -582 2304 -576
rect 2298 -588 2304 -582
rect 2298 -594 2304 -588
rect 2298 -600 2304 -594
rect 2298 -606 2304 -600
rect 2298 -612 2304 -606
rect 2298 -618 2304 -612
rect 2298 -624 2304 -618
rect 2298 -630 2304 -624
rect 2298 -636 2304 -630
rect 2298 -642 2304 -636
rect 2298 -648 2304 -642
rect 2298 -654 2304 -648
rect 2298 -660 2304 -654
rect 2298 -666 2304 -660
rect 2298 -672 2304 -666
rect 2298 -678 2304 -672
rect 2298 -684 2304 -678
rect 2298 -690 2304 -684
rect 2298 -696 2304 -690
rect 2298 -702 2304 -696
rect 2298 -708 2304 -702
rect 2298 -714 2304 -708
rect 2298 -720 2304 -714
rect 2298 -726 2304 -720
rect 2298 -732 2304 -726
rect 2298 -738 2304 -732
rect 2298 -744 2304 -738
rect 2298 -750 2304 -744
rect 2298 -756 2304 -750
rect 2298 -762 2304 -756
rect 2298 -768 2304 -762
rect 2298 -774 2304 -768
rect 2298 -780 2304 -774
rect 2298 -786 2304 -780
rect 2298 -792 2304 -786
rect 2298 -798 2304 -792
rect 2298 -804 2304 -798
rect 2298 -810 2304 -804
rect 2298 -816 2304 -810
rect 2298 -822 2304 -816
rect 2298 -828 2304 -822
rect 2298 -834 2304 -828
rect 2298 -840 2304 -834
rect 2298 -846 2304 -840
rect 2298 -852 2304 -846
rect 2298 -858 2304 -852
rect 2298 -864 2304 -858
rect 2298 -870 2304 -864
rect 2298 -876 2304 -870
rect 2298 -882 2304 -876
rect 2298 -888 2304 -882
rect 2298 -894 2304 -888
rect 2298 -900 2304 -894
rect 2298 -906 2304 -900
rect 2298 -912 2304 -906
rect 2298 -918 2304 -912
rect 2298 -924 2304 -918
rect 2298 -930 2304 -924
rect 2298 -936 2304 -930
rect 2298 -942 2304 -936
rect 2298 -948 2304 -942
rect 2298 -954 2304 -948
rect 2298 -960 2304 -954
rect 2298 -966 2304 -960
rect 2298 -972 2304 -966
rect 2298 -978 2304 -972
rect 2298 -984 2304 -978
rect 2298 -990 2304 -984
rect 2298 -996 2304 -990
rect 2298 -1470 2304 -1464
rect 2298 -1476 2304 -1470
rect 2298 -1482 2304 -1476
rect 2298 -1488 2304 -1482
rect 2298 -1494 2304 -1488
rect 2298 -1500 2304 -1494
rect 2298 -1506 2304 -1500
rect 2298 -1512 2304 -1506
rect 2298 -1518 2304 -1512
rect 2298 -1524 2304 -1518
rect 2298 -1530 2304 -1524
rect 2298 -1536 2304 -1530
rect 2298 -1542 2304 -1536
rect 2298 -1548 2304 -1542
rect 2298 -1554 2304 -1548
rect 2298 -1560 2304 -1554
rect 2298 -1566 2304 -1560
rect 2298 -1572 2304 -1566
rect 2298 -1578 2304 -1572
rect 2298 -1584 2304 -1578
rect 2298 -1590 2304 -1584
rect 2298 -1596 2304 -1590
rect 2298 -1602 2304 -1596
rect 2298 -1608 2304 -1602
rect 2298 -1614 2304 -1608
rect 2298 -1620 2304 -1614
rect 2298 -1626 2304 -1620
rect 2298 -1632 2304 -1626
rect 2298 -1638 2304 -1632
rect 2298 -1644 2304 -1638
rect 2298 -1650 2304 -1644
rect 2298 -1656 2304 -1650
rect 2298 -1662 2304 -1656
rect 2298 -1668 2304 -1662
rect 2298 -1674 2304 -1668
rect 2298 -1680 2304 -1674
rect 2298 -1686 2304 -1680
rect 2298 -1692 2304 -1686
rect 2298 -1698 2304 -1692
rect 2298 -1704 2304 -1698
rect 2298 -1710 2304 -1704
rect 2298 -1716 2304 -1710
rect 2298 -1722 2304 -1716
rect 2298 -1728 2304 -1722
rect 2298 -1734 2304 -1728
rect 2298 -1740 2304 -1734
rect 2298 -1746 2304 -1740
rect 2298 -1752 2304 -1746
rect 2298 -1758 2304 -1752
rect 2298 -1764 2304 -1758
rect 2298 -1770 2304 -1764
rect 2298 -1776 2304 -1770
rect 2298 -1782 2304 -1776
rect 2298 -1788 2304 -1782
rect 2298 -1794 2304 -1788
rect 2298 -1800 2304 -1794
rect 2298 -1806 2304 -1800
rect 2298 -1812 2304 -1806
rect 2298 -1818 2304 -1812
rect 2298 -1824 2304 -1818
rect 2298 -1830 2304 -1824
rect 2298 -1836 2304 -1830
rect 2298 -1842 2304 -1836
rect 2298 -1848 2304 -1842
rect 2298 -1854 2304 -1848
rect 2298 -1860 2304 -1854
rect 2298 -1866 2304 -1860
rect 2298 -1872 2304 -1866
rect 2298 -1878 2304 -1872
rect 2298 -1884 2304 -1878
rect 2298 -1890 2304 -1884
rect 2298 -1896 2304 -1890
rect 2298 -1902 2304 -1896
rect 2298 -1908 2304 -1902
rect 2298 -1914 2304 -1908
rect 2298 -1920 2304 -1914
rect 2298 -1926 2304 -1920
rect 2298 -1932 2304 -1926
rect 2298 -1938 2304 -1932
rect 2298 -1944 2304 -1938
rect 2298 -1950 2304 -1944
rect 2298 -1956 2304 -1950
rect 2298 -1962 2304 -1956
rect 2298 -1968 2304 -1962
rect 2298 -1974 2304 -1968
rect 2298 -1980 2304 -1974
rect 2298 -1986 2304 -1980
rect 2298 -1992 2304 -1986
rect 2298 -1998 2304 -1992
rect 2298 -2004 2304 -1998
rect 2298 -2010 2304 -2004
rect 2298 -2016 2304 -2010
rect 2298 -2022 2304 -2016
rect 2298 -2028 2304 -2022
rect 2298 -2034 2304 -2028
rect 2298 -2040 2304 -2034
rect 2298 -2046 2304 -2040
rect 2298 -2052 2304 -2046
rect 2298 -2058 2304 -2052
rect 2298 -2064 2304 -2058
rect 2298 -2070 2304 -2064
rect 2298 -2076 2304 -2070
rect 2298 -2082 2304 -2076
rect 2298 -2088 2304 -2082
rect 2298 -2094 2304 -2088
rect 2298 -2100 2304 -2094
rect 2298 -2106 2304 -2100
rect 2298 -2112 2304 -2106
rect 2298 -2118 2304 -2112
rect 2298 -2124 2304 -2118
rect 2298 -2130 2304 -2124
rect 2298 -2136 2304 -2130
rect 2298 -2142 2304 -2136
rect 2298 -2148 2304 -2142
rect 2298 -2154 2304 -2148
rect 2298 -2160 2304 -2154
rect 2298 -2166 2304 -2160
rect 2298 -2172 2304 -2166
rect 2298 -2178 2304 -2172
rect 2298 -2184 2304 -2178
rect 2298 -2190 2304 -2184
rect 2298 -2196 2304 -2190
rect 2298 -2202 2304 -2196
rect 2298 -2208 2304 -2202
rect 2298 -2214 2304 -2208
rect 2298 -2220 2304 -2214
rect 2298 -2298 2304 -2292
rect 2298 -2304 2304 -2298
rect 2298 -2310 2304 -2304
rect 2298 -2316 2304 -2310
rect 2298 -2322 2304 -2316
rect 2298 -2328 2304 -2322
rect 2298 -2334 2304 -2328
rect 2298 -2340 2304 -2334
rect 2298 -2346 2304 -2340
rect 2298 -2352 2304 -2346
rect 2298 -2358 2304 -2352
rect 2298 -2364 2304 -2358
rect 2298 -2370 2304 -2364
rect 2298 -2376 2304 -2370
rect 2298 -2382 2304 -2376
rect 2298 -2388 2304 -2382
rect 2298 -2394 2304 -2388
rect 2298 -2400 2304 -2394
rect 2298 -2406 2304 -2400
rect 2298 -2412 2304 -2406
rect 2298 -2418 2304 -2412
rect 2298 -2424 2304 -2418
rect 2298 -2430 2304 -2424
rect 2298 -2436 2304 -2430
rect 2298 -2442 2304 -2436
rect 2298 -2508 2304 -2502
rect 2298 -2514 2304 -2508
rect 2298 -2520 2304 -2514
rect 2298 -2526 2304 -2520
rect 2298 -2532 2304 -2526
rect 2298 -2538 2304 -2532
rect 2298 -2544 2304 -2538
rect 2298 -2550 2304 -2544
rect 2298 -2556 2304 -2550
rect 2298 -2562 2304 -2556
rect 2298 -2568 2304 -2562
rect 2298 -2574 2304 -2568
rect 2298 -2580 2304 -2574
rect 2298 -2586 2304 -2580
rect 2298 -2592 2304 -2586
rect 2298 -2598 2304 -2592
rect 2298 -2604 2304 -2598
rect 2298 -2610 2304 -2604
rect 2298 -2616 2304 -2610
rect 2298 -2622 2304 -2616
rect 2298 -2628 2304 -2622
rect 2298 -2634 2304 -2628
rect 2298 -2640 2304 -2634
rect 2298 -2646 2304 -2640
rect 2298 -2652 2304 -2646
rect 2298 -2658 2304 -2652
rect 2298 -2664 2304 -2658
rect 2298 -2670 2304 -2664
rect 2298 -2676 2304 -2670
rect 2298 -2682 2304 -2676
rect 2298 -2688 2304 -2682
rect 2298 -2694 2304 -2688
rect 2298 -2700 2304 -2694
rect 2298 -2706 2304 -2700
rect 2298 -2712 2304 -2706
rect 2298 -2718 2304 -2712
rect 2298 -2724 2304 -2718
rect 2298 -2730 2304 -2724
rect 2298 -2736 2304 -2730
rect 2298 -2742 2304 -2736
rect 2298 -2748 2304 -2742
rect 2298 -2754 2304 -2748
rect 2298 -2760 2304 -2754
rect 2298 -2766 2304 -2760
rect 2298 -2772 2304 -2766
rect 2298 -2778 2304 -2772
rect 2298 -2784 2304 -2778
rect 2298 -2790 2304 -2784
rect 2298 -2796 2304 -2790
rect 2298 -2802 2304 -2796
rect 2298 -2808 2304 -2802
rect 2298 -2814 2304 -2808
rect 2298 -2820 2304 -2814
rect 2298 -2826 2304 -2820
rect 2298 -2832 2304 -2826
rect 2298 -2838 2304 -2832
rect 2298 -2844 2304 -2838
rect 2298 -2850 2304 -2844
rect 2298 -2856 2304 -2850
rect 2298 -2862 2304 -2856
rect 2298 -2868 2304 -2862
rect 2298 -2874 2304 -2868
rect 2298 -2880 2304 -2874
rect 2298 -2886 2304 -2880
rect 2298 -2892 2304 -2886
rect 2298 -2898 2304 -2892
rect 2298 -2904 2304 -2898
rect 2298 -2910 2304 -2904
rect 2298 -2916 2304 -2910
rect 2298 -2922 2304 -2916
rect 2298 -2928 2304 -2922
rect 2298 -2934 2304 -2928
rect 2298 -2940 2304 -2934
rect 2298 -2946 2304 -2940
rect 2304 -72 2310 -66
rect 2304 -78 2310 -72
rect 2304 -84 2310 -78
rect 2304 -90 2310 -84
rect 2304 -96 2310 -90
rect 2304 -102 2310 -96
rect 2304 -108 2310 -102
rect 2304 -114 2310 -108
rect 2304 -120 2310 -114
rect 2304 -126 2310 -120
rect 2304 -132 2310 -126
rect 2304 -138 2310 -132
rect 2304 -144 2310 -138
rect 2304 -150 2310 -144
rect 2304 -156 2310 -150
rect 2304 -162 2310 -156
rect 2304 -168 2310 -162
rect 2304 -174 2310 -168
rect 2304 -180 2310 -174
rect 2304 -186 2310 -180
rect 2304 -192 2310 -186
rect 2304 -198 2310 -192
rect 2304 -204 2310 -198
rect 2304 -210 2310 -204
rect 2304 -216 2310 -210
rect 2304 -222 2310 -216
rect 2304 -228 2310 -222
rect 2304 -234 2310 -228
rect 2304 -240 2310 -234
rect 2304 -246 2310 -240
rect 2304 -252 2310 -246
rect 2304 -258 2310 -252
rect 2304 -264 2310 -258
rect 2304 -270 2310 -264
rect 2304 -276 2310 -270
rect 2304 -282 2310 -276
rect 2304 -288 2310 -282
rect 2304 -294 2310 -288
rect 2304 -300 2310 -294
rect 2304 -306 2310 -300
rect 2304 -312 2310 -306
rect 2304 -318 2310 -312
rect 2304 -324 2310 -318
rect 2304 -330 2310 -324
rect 2304 -336 2310 -330
rect 2304 -342 2310 -336
rect 2304 -348 2310 -342
rect 2304 -354 2310 -348
rect 2304 -360 2310 -354
rect 2304 -366 2310 -360
rect 2304 -372 2310 -366
rect 2304 -378 2310 -372
rect 2304 -384 2310 -378
rect 2304 -390 2310 -384
rect 2304 -396 2310 -390
rect 2304 -402 2310 -396
rect 2304 -408 2310 -402
rect 2304 -414 2310 -408
rect 2304 -420 2310 -414
rect 2304 -426 2310 -420
rect 2304 -432 2310 -426
rect 2304 -438 2310 -432
rect 2304 -444 2310 -438
rect 2304 -450 2310 -444
rect 2304 -456 2310 -450
rect 2304 -462 2310 -456
rect 2304 -468 2310 -462
rect 2304 -474 2310 -468
rect 2304 -480 2310 -474
rect 2304 -486 2310 -480
rect 2304 -492 2310 -486
rect 2304 -498 2310 -492
rect 2304 -504 2310 -498
rect 2304 -510 2310 -504
rect 2304 -516 2310 -510
rect 2304 -522 2310 -516
rect 2304 -528 2310 -522
rect 2304 -534 2310 -528
rect 2304 -540 2310 -534
rect 2304 -546 2310 -540
rect 2304 -552 2310 -546
rect 2304 -558 2310 -552
rect 2304 -564 2310 -558
rect 2304 -570 2310 -564
rect 2304 -576 2310 -570
rect 2304 -582 2310 -576
rect 2304 -588 2310 -582
rect 2304 -594 2310 -588
rect 2304 -600 2310 -594
rect 2304 -606 2310 -600
rect 2304 -612 2310 -606
rect 2304 -618 2310 -612
rect 2304 -624 2310 -618
rect 2304 -630 2310 -624
rect 2304 -636 2310 -630
rect 2304 -642 2310 -636
rect 2304 -648 2310 -642
rect 2304 -654 2310 -648
rect 2304 -660 2310 -654
rect 2304 -666 2310 -660
rect 2304 -672 2310 -666
rect 2304 -678 2310 -672
rect 2304 -684 2310 -678
rect 2304 -690 2310 -684
rect 2304 -696 2310 -690
rect 2304 -702 2310 -696
rect 2304 -708 2310 -702
rect 2304 -714 2310 -708
rect 2304 -720 2310 -714
rect 2304 -726 2310 -720
rect 2304 -732 2310 -726
rect 2304 -738 2310 -732
rect 2304 -744 2310 -738
rect 2304 -750 2310 -744
rect 2304 -756 2310 -750
rect 2304 -762 2310 -756
rect 2304 -768 2310 -762
rect 2304 -774 2310 -768
rect 2304 -780 2310 -774
rect 2304 -786 2310 -780
rect 2304 -792 2310 -786
rect 2304 -798 2310 -792
rect 2304 -804 2310 -798
rect 2304 -810 2310 -804
rect 2304 -816 2310 -810
rect 2304 -822 2310 -816
rect 2304 -828 2310 -822
rect 2304 -834 2310 -828
rect 2304 -840 2310 -834
rect 2304 -846 2310 -840
rect 2304 -852 2310 -846
rect 2304 -858 2310 -852
rect 2304 -864 2310 -858
rect 2304 -870 2310 -864
rect 2304 -876 2310 -870
rect 2304 -882 2310 -876
rect 2304 -888 2310 -882
rect 2304 -894 2310 -888
rect 2304 -900 2310 -894
rect 2304 -906 2310 -900
rect 2304 -912 2310 -906
rect 2304 -918 2310 -912
rect 2304 -924 2310 -918
rect 2304 -930 2310 -924
rect 2304 -936 2310 -930
rect 2304 -942 2310 -936
rect 2304 -948 2310 -942
rect 2304 -954 2310 -948
rect 2304 -960 2310 -954
rect 2304 -966 2310 -960
rect 2304 -972 2310 -966
rect 2304 -978 2310 -972
rect 2304 -1464 2310 -1458
rect 2304 -1470 2310 -1464
rect 2304 -1476 2310 -1470
rect 2304 -1482 2310 -1476
rect 2304 -1488 2310 -1482
rect 2304 -1494 2310 -1488
rect 2304 -1500 2310 -1494
rect 2304 -1506 2310 -1500
rect 2304 -1512 2310 -1506
rect 2304 -1518 2310 -1512
rect 2304 -1524 2310 -1518
rect 2304 -1530 2310 -1524
rect 2304 -1536 2310 -1530
rect 2304 -1542 2310 -1536
rect 2304 -1548 2310 -1542
rect 2304 -1554 2310 -1548
rect 2304 -1560 2310 -1554
rect 2304 -1566 2310 -1560
rect 2304 -1572 2310 -1566
rect 2304 -1578 2310 -1572
rect 2304 -1584 2310 -1578
rect 2304 -1590 2310 -1584
rect 2304 -1596 2310 -1590
rect 2304 -1602 2310 -1596
rect 2304 -1608 2310 -1602
rect 2304 -1614 2310 -1608
rect 2304 -1620 2310 -1614
rect 2304 -1626 2310 -1620
rect 2304 -1632 2310 -1626
rect 2304 -1638 2310 -1632
rect 2304 -1644 2310 -1638
rect 2304 -1650 2310 -1644
rect 2304 -1656 2310 -1650
rect 2304 -1662 2310 -1656
rect 2304 -1668 2310 -1662
rect 2304 -1674 2310 -1668
rect 2304 -1680 2310 -1674
rect 2304 -1686 2310 -1680
rect 2304 -1692 2310 -1686
rect 2304 -1698 2310 -1692
rect 2304 -1704 2310 -1698
rect 2304 -1710 2310 -1704
rect 2304 -1716 2310 -1710
rect 2304 -1722 2310 -1716
rect 2304 -1728 2310 -1722
rect 2304 -1734 2310 -1728
rect 2304 -1740 2310 -1734
rect 2304 -1746 2310 -1740
rect 2304 -1752 2310 -1746
rect 2304 -1758 2310 -1752
rect 2304 -1764 2310 -1758
rect 2304 -1770 2310 -1764
rect 2304 -1776 2310 -1770
rect 2304 -1782 2310 -1776
rect 2304 -1788 2310 -1782
rect 2304 -1794 2310 -1788
rect 2304 -1800 2310 -1794
rect 2304 -1806 2310 -1800
rect 2304 -1812 2310 -1806
rect 2304 -1818 2310 -1812
rect 2304 -1824 2310 -1818
rect 2304 -1830 2310 -1824
rect 2304 -1836 2310 -1830
rect 2304 -1842 2310 -1836
rect 2304 -1848 2310 -1842
rect 2304 -1854 2310 -1848
rect 2304 -1860 2310 -1854
rect 2304 -1866 2310 -1860
rect 2304 -1872 2310 -1866
rect 2304 -1878 2310 -1872
rect 2304 -1884 2310 -1878
rect 2304 -1890 2310 -1884
rect 2304 -1896 2310 -1890
rect 2304 -1902 2310 -1896
rect 2304 -1908 2310 -1902
rect 2304 -1914 2310 -1908
rect 2304 -1920 2310 -1914
rect 2304 -1926 2310 -1920
rect 2304 -1932 2310 -1926
rect 2304 -1938 2310 -1932
rect 2304 -1944 2310 -1938
rect 2304 -1950 2310 -1944
rect 2304 -1956 2310 -1950
rect 2304 -1962 2310 -1956
rect 2304 -1968 2310 -1962
rect 2304 -1974 2310 -1968
rect 2304 -1980 2310 -1974
rect 2304 -1986 2310 -1980
rect 2304 -1992 2310 -1986
rect 2304 -1998 2310 -1992
rect 2304 -2004 2310 -1998
rect 2304 -2010 2310 -2004
rect 2304 -2016 2310 -2010
rect 2304 -2022 2310 -2016
rect 2304 -2028 2310 -2022
rect 2304 -2034 2310 -2028
rect 2304 -2040 2310 -2034
rect 2304 -2046 2310 -2040
rect 2304 -2052 2310 -2046
rect 2304 -2058 2310 -2052
rect 2304 -2064 2310 -2058
rect 2304 -2070 2310 -2064
rect 2304 -2076 2310 -2070
rect 2304 -2082 2310 -2076
rect 2304 -2088 2310 -2082
rect 2304 -2094 2310 -2088
rect 2304 -2100 2310 -2094
rect 2304 -2106 2310 -2100
rect 2304 -2112 2310 -2106
rect 2304 -2118 2310 -2112
rect 2304 -2124 2310 -2118
rect 2304 -2130 2310 -2124
rect 2304 -2136 2310 -2130
rect 2304 -2142 2310 -2136
rect 2304 -2148 2310 -2142
rect 2304 -2154 2310 -2148
rect 2304 -2160 2310 -2154
rect 2304 -2166 2310 -2160
rect 2304 -2172 2310 -2166
rect 2304 -2178 2310 -2172
rect 2304 -2184 2310 -2178
rect 2304 -2190 2310 -2184
rect 2304 -2196 2310 -2190
rect 2304 -2202 2310 -2196
rect 2304 -2208 2310 -2202
rect 2304 -2214 2310 -2208
rect 2304 -2286 2310 -2280
rect 2304 -2292 2310 -2286
rect 2304 -2298 2310 -2292
rect 2304 -2304 2310 -2298
rect 2304 -2310 2310 -2304
rect 2304 -2316 2310 -2310
rect 2304 -2322 2310 -2316
rect 2304 -2328 2310 -2322
rect 2304 -2334 2310 -2328
rect 2304 -2340 2310 -2334
rect 2304 -2346 2310 -2340
rect 2304 -2352 2310 -2346
rect 2304 -2358 2310 -2352
rect 2304 -2364 2310 -2358
rect 2304 -2370 2310 -2364
rect 2304 -2376 2310 -2370
rect 2304 -2382 2310 -2376
rect 2304 -2388 2310 -2382
rect 2304 -2394 2310 -2388
rect 2304 -2400 2310 -2394
rect 2304 -2406 2310 -2400
rect 2304 -2412 2310 -2406
rect 2304 -2418 2310 -2412
rect 2304 -2424 2310 -2418
rect 2304 -2430 2310 -2424
rect 2304 -2436 2310 -2430
rect 2304 -2442 2310 -2436
rect 2304 -2508 2310 -2502
rect 2304 -2514 2310 -2508
rect 2304 -2520 2310 -2514
rect 2304 -2526 2310 -2520
rect 2304 -2532 2310 -2526
rect 2304 -2538 2310 -2532
rect 2304 -2544 2310 -2538
rect 2304 -2550 2310 -2544
rect 2304 -2556 2310 -2550
rect 2304 -2562 2310 -2556
rect 2304 -2568 2310 -2562
rect 2304 -2574 2310 -2568
rect 2304 -2580 2310 -2574
rect 2304 -2586 2310 -2580
rect 2304 -2592 2310 -2586
rect 2304 -2598 2310 -2592
rect 2304 -2604 2310 -2598
rect 2304 -2610 2310 -2604
rect 2304 -2616 2310 -2610
rect 2304 -2622 2310 -2616
rect 2304 -2628 2310 -2622
rect 2304 -2634 2310 -2628
rect 2304 -2640 2310 -2634
rect 2304 -2646 2310 -2640
rect 2304 -2652 2310 -2646
rect 2304 -2658 2310 -2652
rect 2304 -2664 2310 -2658
rect 2304 -2670 2310 -2664
rect 2304 -2676 2310 -2670
rect 2304 -2682 2310 -2676
rect 2304 -2688 2310 -2682
rect 2304 -2694 2310 -2688
rect 2304 -2700 2310 -2694
rect 2304 -2706 2310 -2700
rect 2304 -2712 2310 -2706
rect 2304 -2718 2310 -2712
rect 2304 -2724 2310 -2718
rect 2304 -2730 2310 -2724
rect 2304 -2736 2310 -2730
rect 2304 -2742 2310 -2736
rect 2304 -2748 2310 -2742
rect 2304 -2754 2310 -2748
rect 2304 -2760 2310 -2754
rect 2304 -2766 2310 -2760
rect 2304 -2772 2310 -2766
rect 2304 -2778 2310 -2772
rect 2304 -2784 2310 -2778
rect 2304 -2790 2310 -2784
rect 2304 -2796 2310 -2790
rect 2304 -2802 2310 -2796
rect 2304 -2808 2310 -2802
rect 2304 -2814 2310 -2808
rect 2304 -2820 2310 -2814
rect 2304 -2826 2310 -2820
rect 2304 -2832 2310 -2826
rect 2304 -2838 2310 -2832
rect 2304 -2844 2310 -2838
rect 2304 -2850 2310 -2844
rect 2304 -2856 2310 -2850
rect 2304 -2862 2310 -2856
rect 2304 -2868 2310 -2862
rect 2304 -2874 2310 -2868
rect 2304 -2880 2310 -2874
rect 2304 -2886 2310 -2880
rect 2304 -2892 2310 -2886
rect 2304 -2898 2310 -2892
rect 2304 -2904 2310 -2898
rect 2304 -2910 2310 -2904
rect 2304 -2916 2310 -2910
rect 2304 -2922 2310 -2916
rect 2304 -2928 2310 -2922
rect 2304 -2934 2310 -2928
rect 2304 -2940 2310 -2934
rect 2304 -2946 2310 -2940
rect 2310 -60 2316 -54
rect 2310 -66 2316 -60
rect 2310 -72 2316 -66
rect 2310 -78 2316 -72
rect 2310 -84 2316 -78
rect 2310 -90 2316 -84
rect 2310 -96 2316 -90
rect 2310 -102 2316 -96
rect 2310 -108 2316 -102
rect 2310 -114 2316 -108
rect 2310 -120 2316 -114
rect 2310 -126 2316 -120
rect 2310 -132 2316 -126
rect 2310 -138 2316 -132
rect 2310 -144 2316 -138
rect 2310 -150 2316 -144
rect 2310 -156 2316 -150
rect 2310 -162 2316 -156
rect 2310 -168 2316 -162
rect 2310 -174 2316 -168
rect 2310 -180 2316 -174
rect 2310 -186 2316 -180
rect 2310 -192 2316 -186
rect 2310 -198 2316 -192
rect 2310 -204 2316 -198
rect 2310 -210 2316 -204
rect 2310 -216 2316 -210
rect 2310 -222 2316 -216
rect 2310 -228 2316 -222
rect 2310 -234 2316 -228
rect 2310 -240 2316 -234
rect 2310 -246 2316 -240
rect 2310 -252 2316 -246
rect 2310 -258 2316 -252
rect 2310 -264 2316 -258
rect 2310 -270 2316 -264
rect 2310 -276 2316 -270
rect 2310 -282 2316 -276
rect 2310 -288 2316 -282
rect 2310 -294 2316 -288
rect 2310 -300 2316 -294
rect 2310 -306 2316 -300
rect 2310 -312 2316 -306
rect 2310 -318 2316 -312
rect 2310 -324 2316 -318
rect 2310 -330 2316 -324
rect 2310 -336 2316 -330
rect 2310 -342 2316 -336
rect 2310 -348 2316 -342
rect 2310 -354 2316 -348
rect 2310 -360 2316 -354
rect 2310 -366 2316 -360
rect 2310 -372 2316 -366
rect 2310 -378 2316 -372
rect 2310 -384 2316 -378
rect 2310 -390 2316 -384
rect 2310 -396 2316 -390
rect 2310 -402 2316 -396
rect 2310 -408 2316 -402
rect 2310 -414 2316 -408
rect 2310 -420 2316 -414
rect 2310 -426 2316 -420
rect 2310 -432 2316 -426
rect 2310 -438 2316 -432
rect 2310 -444 2316 -438
rect 2310 -450 2316 -444
rect 2310 -456 2316 -450
rect 2310 -462 2316 -456
rect 2310 -468 2316 -462
rect 2310 -474 2316 -468
rect 2310 -480 2316 -474
rect 2310 -486 2316 -480
rect 2310 -492 2316 -486
rect 2310 -498 2316 -492
rect 2310 -504 2316 -498
rect 2310 -510 2316 -504
rect 2310 -516 2316 -510
rect 2310 -522 2316 -516
rect 2310 -528 2316 -522
rect 2310 -534 2316 -528
rect 2310 -540 2316 -534
rect 2310 -546 2316 -540
rect 2310 -552 2316 -546
rect 2310 -558 2316 -552
rect 2310 -564 2316 -558
rect 2310 -570 2316 -564
rect 2310 -576 2316 -570
rect 2310 -582 2316 -576
rect 2310 -588 2316 -582
rect 2310 -594 2316 -588
rect 2310 -600 2316 -594
rect 2310 -606 2316 -600
rect 2310 -612 2316 -606
rect 2310 -618 2316 -612
rect 2310 -624 2316 -618
rect 2310 -630 2316 -624
rect 2310 -636 2316 -630
rect 2310 -642 2316 -636
rect 2310 -648 2316 -642
rect 2310 -654 2316 -648
rect 2310 -660 2316 -654
rect 2310 -666 2316 -660
rect 2310 -672 2316 -666
rect 2310 -678 2316 -672
rect 2310 -684 2316 -678
rect 2310 -690 2316 -684
rect 2310 -696 2316 -690
rect 2310 -702 2316 -696
rect 2310 -708 2316 -702
rect 2310 -714 2316 -708
rect 2310 -720 2316 -714
rect 2310 -726 2316 -720
rect 2310 -732 2316 -726
rect 2310 -738 2316 -732
rect 2310 -744 2316 -738
rect 2310 -750 2316 -744
rect 2310 -756 2316 -750
rect 2310 -762 2316 -756
rect 2310 -768 2316 -762
rect 2310 -774 2316 -768
rect 2310 -780 2316 -774
rect 2310 -786 2316 -780
rect 2310 -792 2316 -786
rect 2310 -798 2316 -792
rect 2310 -804 2316 -798
rect 2310 -810 2316 -804
rect 2310 -816 2316 -810
rect 2310 -822 2316 -816
rect 2310 -828 2316 -822
rect 2310 -834 2316 -828
rect 2310 -840 2316 -834
rect 2310 -846 2316 -840
rect 2310 -852 2316 -846
rect 2310 -858 2316 -852
rect 2310 -864 2316 -858
rect 2310 -870 2316 -864
rect 2310 -876 2316 -870
rect 2310 -882 2316 -876
rect 2310 -888 2316 -882
rect 2310 -894 2316 -888
rect 2310 -900 2316 -894
rect 2310 -906 2316 -900
rect 2310 -912 2316 -906
rect 2310 -918 2316 -912
rect 2310 -924 2316 -918
rect 2310 -930 2316 -924
rect 2310 -936 2316 -930
rect 2310 -942 2316 -936
rect 2310 -948 2316 -942
rect 2310 -954 2316 -948
rect 2310 -960 2316 -954
rect 2310 -966 2316 -960
rect 2310 -1458 2316 -1452
rect 2310 -1464 2316 -1458
rect 2310 -1470 2316 -1464
rect 2310 -1476 2316 -1470
rect 2310 -1482 2316 -1476
rect 2310 -1488 2316 -1482
rect 2310 -1494 2316 -1488
rect 2310 -1500 2316 -1494
rect 2310 -1506 2316 -1500
rect 2310 -1512 2316 -1506
rect 2310 -1518 2316 -1512
rect 2310 -1524 2316 -1518
rect 2310 -1530 2316 -1524
rect 2310 -1536 2316 -1530
rect 2310 -1542 2316 -1536
rect 2310 -1548 2316 -1542
rect 2310 -1554 2316 -1548
rect 2310 -1560 2316 -1554
rect 2310 -1566 2316 -1560
rect 2310 -1572 2316 -1566
rect 2310 -1578 2316 -1572
rect 2310 -1584 2316 -1578
rect 2310 -1590 2316 -1584
rect 2310 -1596 2316 -1590
rect 2310 -1602 2316 -1596
rect 2310 -1608 2316 -1602
rect 2310 -1614 2316 -1608
rect 2310 -1620 2316 -1614
rect 2310 -1626 2316 -1620
rect 2310 -1632 2316 -1626
rect 2310 -1638 2316 -1632
rect 2310 -1644 2316 -1638
rect 2310 -1650 2316 -1644
rect 2310 -1656 2316 -1650
rect 2310 -1662 2316 -1656
rect 2310 -1668 2316 -1662
rect 2310 -1674 2316 -1668
rect 2310 -1680 2316 -1674
rect 2310 -1686 2316 -1680
rect 2310 -1692 2316 -1686
rect 2310 -1698 2316 -1692
rect 2310 -1704 2316 -1698
rect 2310 -1710 2316 -1704
rect 2310 -1716 2316 -1710
rect 2310 -1722 2316 -1716
rect 2310 -1728 2316 -1722
rect 2310 -1734 2316 -1728
rect 2310 -1740 2316 -1734
rect 2310 -1746 2316 -1740
rect 2310 -1752 2316 -1746
rect 2310 -1758 2316 -1752
rect 2310 -1764 2316 -1758
rect 2310 -1770 2316 -1764
rect 2310 -1776 2316 -1770
rect 2310 -1782 2316 -1776
rect 2310 -1788 2316 -1782
rect 2310 -1794 2316 -1788
rect 2310 -1800 2316 -1794
rect 2310 -1806 2316 -1800
rect 2310 -1812 2316 -1806
rect 2310 -1818 2316 -1812
rect 2310 -1824 2316 -1818
rect 2310 -1830 2316 -1824
rect 2310 -1836 2316 -1830
rect 2310 -1842 2316 -1836
rect 2310 -1848 2316 -1842
rect 2310 -1854 2316 -1848
rect 2310 -1860 2316 -1854
rect 2310 -1866 2316 -1860
rect 2310 -1872 2316 -1866
rect 2310 -1878 2316 -1872
rect 2310 -1884 2316 -1878
rect 2310 -1890 2316 -1884
rect 2310 -1896 2316 -1890
rect 2310 -1902 2316 -1896
rect 2310 -1908 2316 -1902
rect 2310 -1914 2316 -1908
rect 2310 -1920 2316 -1914
rect 2310 -1926 2316 -1920
rect 2310 -1932 2316 -1926
rect 2310 -1938 2316 -1932
rect 2310 -1944 2316 -1938
rect 2310 -1950 2316 -1944
rect 2310 -1956 2316 -1950
rect 2310 -1962 2316 -1956
rect 2310 -1968 2316 -1962
rect 2310 -1974 2316 -1968
rect 2310 -1980 2316 -1974
rect 2310 -1986 2316 -1980
rect 2310 -1992 2316 -1986
rect 2310 -1998 2316 -1992
rect 2310 -2004 2316 -1998
rect 2310 -2010 2316 -2004
rect 2310 -2016 2316 -2010
rect 2310 -2022 2316 -2016
rect 2310 -2028 2316 -2022
rect 2310 -2034 2316 -2028
rect 2310 -2040 2316 -2034
rect 2310 -2046 2316 -2040
rect 2310 -2052 2316 -2046
rect 2310 -2058 2316 -2052
rect 2310 -2064 2316 -2058
rect 2310 -2070 2316 -2064
rect 2310 -2076 2316 -2070
rect 2310 -2082 2316 -2076
rect 2310 -2088 2316 -2082
rect 2310 -2094 2316 -2088
rect 2310 -2100 2316 -2094
rect 2310 -2106 2316 -2100
rect 2310 -2112 2316 -2106
rect 2310 -2118 2316 -2112
rect 2310 -2124 2316 -2118
rect 2310 -2130 2316 -2124
rect 2310 -2136 2316 -2130
rect 2310 -2142 2316 -2136
rect 2310 -2148 2316 -2142
rect 2310 -2154 2316 -2148
rect 2310 -2160 2316 -2154
rect 2310 -2166 2316 -2160
rect 2310 -2172 2316 -2166
rect 2310 -2178 2316 -2172
rect 2310 -2184 2316 -2178
rect 2310 -2190 2316 -2184
rect 2310 -2196 2316 -2190
rect 2310 -2202 2316 -2196
rect 2310 -2208 2316 -2202
rect 2310 -2280 2316 -2274
rect 2310 -2286 2316 -2280
rect 2310 -2292 2316 -2286
rect 2310 -2298 2316 -2292
rect 2310 -2304 2316 -2298
rect 2310 -2310 2316 -2304
rect 2310 -2316 2316 -2310
rect 2310 -2322 2316 -2316
rect 2310 -2328 2316 -2322
rect 2310 -2334 2316 -2328
rect 2310 -2340 2316 -2334
rect 2310 -2346 2316 -2340
rect 2310 -2352 2316 -2346
rect 2310 -2358 2316 -2352
rect 2310 -2364 2316 -2358
rect 2310 -2370 2316 -2364
rect 2310 -2376 2316 -2370
rect 2310 -2382 2316 -2376
rect 2310 -2388 2316 -2382
rect 2310 -2394 2316 -2388
rect 2310 -2400 2316 -2394
rect 2310 -2406 2316 -2400
rect 2310 -2412 2316 -2406
rect 2310 -2418 2316 -2412
rect 2310 -2424 2316 -2418
rect 2310 -2430 2316 -2424
rect 2310 -2436 2316 -2430
rect 2310 -2442 2316 -2436
rect 2310 -2502 2316 -2496
rect 2310 -2508 2316 -2502
rect 2310 -2514 2316 -2508
rect 2310 -2520 2316 -2514
rect 2310 -2526 2316 -2520
rect 2310 -2532 2316 -2526
rect 2310 -2538 2316 -2532
rect 2310 -2544 2316 -2538
rect 2310 -2550 2316 -2544
rect 2310 -2556 2316 -2550
rect 2310 -2562 2316 -2556
rect 2310 -2568 2316 -2562
rect 2310 -2574 2316 -2568
rect 2310 -2580 2316 -2574
rect 2310 -2586 2316 -2580
rect 2310 -2592 2316 -2586
rect 2310 -2598 2316 -2592
rect 2310 -2604 2316 -2598
rect 2310 -2610 2316 -2604
rect 2310 -2616 2316 -2610
rect 2310 -2622 2316 -2616
rect 2310 -2628 2316 -2622
rect 2310 -2634 2316 -2628
rect 2310 -2640 2316 -2634
rect 2310 -2646 2316 -2640
rect 2310 -2652 2316 -2646
rect 2310 -2658 2316 -2652
rect 2310 -2664 2316 -2658
rect 2310 -2670 2316 -2664
rect 2310 -2676 2316 -2670
rect 2310 -2682 2316 -2676
rect 2310 -2688 2316 -2682
rect 2310 -2694 2316 -2688
rect 2310 -2700 2316 -2694
rect 2310 -2706 2316 -2700
rect 2310 -2712 2316 -2706
rect 2310 -2718 2316 -2712
rect 2310 -2724 2316 -2718
rect 2310 -2730 2316 -2724
rect 2310 -2736 2316 -2730
rect 2310 -2742 2316 -2736
rect 2310 -2748 2316 -2742
rect 2310 -2754 2316 -2748
rect 2310 -2760 2316 -2754
rect 2310 -2766 2316 -2760
rect 2310 -2772 2316 -2766
rect 2310 -2778 2316 -2772
rect 2310 -2784 2316 -2778
rect 2310 -2790 2316 -2784
rect 2310 -2796 2316 -2790
rect 2310 -2802 2316 -2796
rect 2310 -2808 2316 -2802
rect 2310 -2814 2316 -2808
rect 2310 -2820 2316 -2814
rect 2310 -2826 2316 -2820
rect 2310 -2832 2316 -2826
rect 2310 -2838 2316 -2832
rect 2310 -2844 2316 -2838
rect 2310 -2850 2316 -2844
rect 2310 -2856 2316 -2850
rect 2310 -2862 2316 -2856
rect 2310 -2868 2316 -2862
rect 2310 -2874 2316 -2868
rect 2310 -2880 2316 -2874
rect 2310 -2886 2316 -2880
rect 2310 -2892 2316 -2886
rect 2310 -2898 2316 -2892
rect 2310 -2904 2316 -2898
rect 2310 -2910 2316 -2904
rect 2310 -2916 2316 -2910
rect 2310 -2922 2316 -2916
rect 2310 -2928 2316 -2922
rect 2310 -2934 2316 -2928
rect 2310 -2940 2316 -2934
rect 2316 -54 2322 -48
rect 2316 -60 2322 -54
rect 2316 -66 2322 -60
rect 2316 -72 2322 -66
rect 2316 -78 2322 -72
rect 2316 -84 2322 -78
rect 2316 -90 2322 -84
rect 2316 -96 2322 -90
rect 2316 -102 2322 -96
rect 2316 -108 2322 -102
rect 2316 -114 2322 -108
rect 2316 -120 2322 -114
rect 2316 -126 2322 -120
rect 2316 -132 2322 -126
rect 2316 -138 2322 -132
rect 2316 -144 2322 -138
rect 2316 -150 2322 -144
rect 2316 -156 2322 -150
rect 2316 -162 2322 -156
rect 2316 -168 2322 -162
rect 2316 -174 2322 -168
rect 2316 -180 2322 -174
rect 2316 -186 2322 -180
rect 2316 -192 2322 -186
rect 2316 -198 2322 -192
rect 2316 -204 2322 -198
rect 2316 -210 2322 -204
rect 2316 -216 2322 -210
rect 2316 -222 2322 -216
rect 2316 -228 2322 -222
rect 2316 -234 2322 -228
rect 2316 -240 2322 -234
rect 2316 -246 2322 -240
rect 2316 -252 2322 -246
rect 2316 -258 2322 -252
rect 2316 -264 2322 -258
rect 2316 -270 2322 -264
rect 2316 -276 2322 -270
rect 2316 -282 2322 -276
rect 2316 -288 2322 -282
rect 2316 -294 2322 -288
rect 2316 -300 2322 -294
rect 2316 -306 2322 -300
rect 2316 -312 2322 -306
rect 2316 -318 2322 -312
rect 2316 -324 2322 -318
rect 2316 -330 2322 -324
rect 2316 -336 2322 -330
rect 2316 -342 2322 -336
rect 2316 -348 2322 -342
rect 2316 -354 2322 -348
rect 2316 -360 2322 -354
rect 2316 -366 2322 -360
rect 2316 -372 2322 -366
rect 2316 -378 2322 -372
rect 2316 -384 2322 -378
rect 2316 -390 2322 -384
rect 2316 -396 2322 -390
rect 2316 -402 2322 -396
rect 2316 -408 2322 -402
rect 2316 -414 2322 -408
rect 2316 -420 2322 -414
rect 2316 -426 2322 -420
rect 2316 -432 2322 -426
rect 2316 -438 2322 -432
rect 2316 -444 2322 -438
rect 2316 -450 2322 -444
rect 2316 -456 2322 -450
rect 2316 -462 2322 -456
rect 2316 -468 2322 -462
rect 2316 -474 2322 -468
rect 2316 -480 2322 -474
rect 2316 -486 2322 -480
rect 2316 -492 2322 -486
rect 2316 -498 2322 -492
rect 2316 -504 2322 -498
rect 2316 -510 2322 -504
rect 2316 -516 2322 -510
rect 2316 -522 2322 -516
rect 2316 -528 2322 -522
rect 2316 -534 2322 -528
rect 2316 -540 2322 -534
rect 2316 -546 2322 -540
rect 2316 -552 2322 -546
rect 2316 -558 2322 -552
rect 2316 -564 2322 -558
rect 2316 -570 2322 -564
rect 2316 -576 2322 -570
rect 2316 -582 2322 -576
rect 2316 -588 2322 -582
rect 2316 -594 2322 -588
rect 2316 -600 2322 -594
rect 2316 -606 2322 -600
rect 2316 -612 2322 -606
rect 2316 -618 2322 -612
rect 2316 -624 2322 -618
rect 2316 -630 2322 -624
rect 2316 -636 2322 -630
rect 2316 -642 2322 -636
rect 2316 -648 2322 -642
rect 2316 -654 2322 -648
rect 2316 -660 2322 -654
rect 2316 -666 2322 -660
rect 2316 -672 2322 -666
rect 2316 -678 2322 -672
rect 2316 -684 2322 -678
rect 2316 -690 2322 -684
rect 2316 -696 2322 -690
rect 2316 -702 2322 -696
rect 2316 -708 2322 -702
rect 2316 -714 2322 -708
rect 2316 -720 2322 -714
rect 2316 -726 2322 -720
rect 2316 -732 2322 -726
rect 2316 -738 2322 -732
rect 2316 -744 2322 -738
rect 2316 -750 2322 -744
rect 2316 -756 2322 -750
rect 2316 -762 2322 -756
rect 2316 -768 2322 -762
rect 2316 -774 2322 -768
rect 2316 -780 2322 -774
rect 2316 -786 2322 -780
rect 2316 -792 2322 -786
rect 2316 -798 2322 -792
rect 2316 -804 2322 -798
rect 2316 -810 2322 -804
rect 2316 -816 2322 -810
rect 2316 -822 2322 -816
rect 2316 -828 2322 -822
rect 2316 -834 2322 -828
rect 2316 -840 2322 -834
rect 2316 -846 2322 -840
rect 2316 -852 2322 -846
rect 2316 -858 2322 -852
rect 2316 -864 2322 -858
rect 2316 -870 2322 -864
rect 2316 -876 2322 -870
rect 2316 -882 2322 -876
rect 2316 -888 2322 -882
rect 2316 -894 2322 -888
rect 2316 -900 2322 -894
rect 2316 -906 2322 -900
rect 2316 -912 2322 -906
rect 2316 -918 2322 -912
rect 2316 -924 2322 -918
rect 2316 -930 2322 -924
rect 2316 -936 2322 -930
rect 2316 -942 2322 -936
rect 2316 -948 2322 -942
rect 2316 -1452 2322 -1446
rect 2316 -1458 2322 -1452
rect 2316 -1464 2322 -1458
rect 2316 -1470 2322 -1464
rect 2316 -1476 2322 -1470
rect 2316 -1482 2322 -1476
rect 2316 -1488 2322 -1482
rect 2316 -1494 2322 -1488
rect 2316 -1500 2322 -1494
rect 2316 -1506 2322 -1500
rect 2316 -1512 2322 -1506
rect 2316 -1518 2322 -1512
rect 2316 -1524 2322 -1518
rect 2316 -1530 2322 -1524
rect 2316 -1536 2322 -1530
rect 2316 -1542 2322 -1536
rect 2316 -1548 2322 -1542
rect 2316 -1554 2322 -1548
rect 2316 -1560 2322 -1554
rect 2316 -1566 2322 -1560
rect 2316 -1572 2322 -1566
rect 2316 -1578 2322 -1572
rect 2316 -1584 2322 -1578
rect 2316 -1590 2322 -1584
rect 2316 -1596 2322 -1590
rect 2316 -1602 2322 -1596
rect 2316 -1608 2322 -1602
rect 2316 -1614 2322 -1608
rect 2316 -1620 2322 -1614
rect 2316 -1626 2322 -1620
rect 2316 -1632 2322 -1626
rect 2316 -1638 2322 -1632
rect 2316 -1644 2322 -1638
rect 2316 -1650 2322 -1644
rect 2316 -1656 2322 -1650
rect 2316 -1662 2322 -1656
rect 2316 -1668 2322 -1662
rect 2316 -1674 2322 -1668
rect 2316 -1680 2322 -1674
rect 2316 -1686 2322 -1680
rect 2316 -1692 2322 -1686
rect 2316 -1698 2322 -1692
rect 2316 -1704 2322 -1698
rect 2316 -1710 2322 -1704
rect 2316 -1716 2322 -1710
rect 2316 -1722 2322 -1716
rect 2316 -1728 2322 -1722
rect 2316 -1734 2322 -1728
rect 2316 -1740 2322 -1734
rect 2316 -1746 2322 -1740
rect 2316 -1752 2322 -1746
rect 2316 -1758 2322 -1752
rect 2316 -1764 2322 -1758
rect 2316 -1770 2322 -1764
rect 2316 -1776 2322 -1770
rect 2316 -1782 2322 -1776
rect 2316 -1788 2322 -1782
rect 2316 -1794 2322 -1788
rect 2316 -1800 2322 -1794
rect 2316 -1806 2322 -1800
rect 2316 -1812 2322 -1806
rect 2316 -1818 2322 -1812
rect 2316 -1824 2322 -1818
rect 2316 -1830 2322 -1824
rect 2316 -1836 2322 -1830
rect 2316 -1842 2322 -1836
rect 2316 -1848 2322 -1842
rect 2316 -1854 2322 -1848
rect 2316 -1860 2322 -1854
rect 2316 -1866 2322 -1860
rect 2316 -1872 2322 -1866
rect 2316 -1878 2322 -1872
rect 2316 -1884 2322 -1878
rect 2316 -1890 2322 -1884
rect 2316 -1896 2322 -1890
rect 2316 -1902 2322 -1896
rect 2316 -1908 2322 -1902
rect 2316 -1914 2322 -1908
rect 2316 -1920 2322 -1914
rect 2316 -1926 2322 -1920
rect 2316 -1932 2322 -1926
rect 2316 -1938 2322 -1932
rect 2316 -1944 2322 -1938
rect 2316 -1950 2322 -1944
rect 2316 -1956 2322 -1950
rect 2316 -1962 2322 -1956
rect 2316 -1968 2322 -1962
rect 2316 -1974 2322 -1968
rect 2316 -1980 2322 -1974
rect 2316 -1986 2322 -1980
rect 2316 -1992 2322 -1986
rect 2316 -1998 2322 -1992
rect 2316 -2004 2322 -1998
rect 2316 -2010 2322 -2004
rect 2316 -2016 2322 -2010
rect 2316 -2022 2322 -2016
rect 2316 -2028 2322 -2022
rect 2316 -2034 2322 -2028
rect 2316 -2040 2322 -2034
rect 2316 -2046 2322 -2040
rect 2316 -2052 2322 -2046
rect 2316 -2058 2322 -2052
rect 2316 -2064 2322 -2058
rect 2316 -2070 2322 -2064
rect 2316 -2076 2322 -2070
rect 2316 -2082 2322 -2076
rect 2316 -2088 2322 -2082
rect 2316 -2094 2322 -2088
rect 2316 -2100 2322 -2094
rect 2316 -2106 2322 -2100
rect 2316 -2112 2322 -2106
rect 2316 -2118 2322 -2112
rect 2316 -2124 2322 -2118
rect 2316 -2130 2322 -2124
rect 2316 -2136 2322 -2130
rect 2316 -2142 2322 -2136
rect 2316 -2148 2322 -2142
rect 2316 -2154 2322 -2148
rect 2316 -2160 2322 -2154
rect 2316 -2166 2322 -2160
rect 2316 -2172 2322 -2166
rect 2316 -2178 2322 -2172
rect 2316 -2184 2322 -2178
rect 2316 -2190 2322 -2184
rect 2316 -2196 2322 -2190
rect 2316 -2202 2322 -2196
rect 2316 -2274 2322 -2268
rect 2316 -2280 2322 -2274
rect 2316 -2286 2322 -2280
rect 2316 -2292 2322 -2286
rect 2316 -2298 2322 -2292
rect 2316 -2304 2322 -2298
rect 2316 -2310 2322 -2304
rect 2316 -2316 2322 -2310
rect 2316 -2322 2322 -2316
rect 2316 -2328 2322 -2322
rect 2316 -2334 2322 -2328
rect 2316 -2340 2322 -2334
rect 2316 -2346 2322 -2340
rect 2316 -2352 2322 -2346
rect 2316 -2358 2322 -2352
rect 2316 -2364 2322 -2358
rect 2316 -2370 2322 -2364
rect 2316 -2376 2322 -2370
rect 2316 -2382 2322 -2376
rect 2316 -2388 2322 -2382
rect 2316 -2394 2322 -2388
rect 2316 -2400 2322 -2394
rect 2316 -2406 2322 -2400
rect 2316 -2412 2322 -2406
rect 2316 -2418 2322 -2412
rect 2316 -2424 2322 -2418
rect 2316 -2430 2322 -2424
rect 2316 -2436 2322 -2430
rect 2316 -2502 2322 -2496
rect 2316 -2508 2322 -2502
rect 2316 -2514 2322 -2508
rect 2316 -2520 2322 -2514
rect 2316 -2526 2322 -2520
rect 2316 -2532 2322 -2526
rect 2316 -2538 2322 -2532
rect 2316 -2544 2322 -2538
rect 2316 -2550 2322 -2544
rect 2316 -2556 2322 -2550
rect 2316 -2562 2322 -2556
rect 2316 -2568 2322 -2562
rect 2316 -2574 2322 -2568
rect 2316 -2580 2322 -2574
rect 2316 -2586 2322 -2580
rect 2316 -2592 2322 -2586
rect 2316 -2598 2322 -2592
rect 2316 -2604 2322 -2598
rect 2316 -2610 2322 -2604
rect 2316 -2616 2322 -2610
rect 2316 -2622 2322 -2616
rect 2316 -2628 2322 -2622
rect 2316 -2634 2322 -2628
rect 2316 -2640 2322 -2634
rect 2316 -2646 2322 -2640
rect 2316 -2652 2322 -2646
rect 2316 -2658 2322 -2652
rect 2316 -2664 2322 -2658
rect 2316 -2670 2322 -2664
rect 2316 -2676 2322 -2670
rect 2316 -2682 2322 -2676
rect 2316 -2688 2322 -2682
rect 2316 -2694 2322 -2688
rect 2316 -2700 2322 -2694
rect 2316 -2706 2322 -2700
rect 2316 -2712 2322 -2706
rect 2316 -2718 2322 -2712
rect 2316 -2724 2322 -2718
rect 2316 -2730 2322 -2724
rect 2316 -2736 2322 -2730
rect 2316 -2742 2322 -2736
rect 2316 -2748 2322 -2742
rect 2316 -2754 2322 -2748
rect 2316 -2760 2322 -2754
rect 2316 -2766 2322 -2760
rect 2316 -2772 2322 -2766
rect 2316 -2778 2322 -2772
rect 2316 -2784 2322 -2778
rect 2316 -2790 2322 -2784
rect 2316 -2796 2322 -2790
rect 2316 -2802 2322 -2796
rect 2316 -2808 2322 -2802
rect 2316 -2814 2322 -2808
rect 2316 -2820 2322 -2814
rect 2316 -2826 2322 -2820
rect 2316 -2832 2322 -2826
rect 2316 -2838 2322 -2832
rect 2316 -2844 2322 -2838
rect 2316 -2850 2322 -2844
rect 2316 -2856 2322 -2850
rect 2316 -2862 2322 -2856
rect 2316 -2868 2322 -2862
rect 2316 -2874 2322 -2868
rect 2316 -2880 2322 -2874
rect 2316 -2886 2322 -2880
rect 2316 -2892 2322 -2886
rect 2316 -2898 2322 -2892
rect 2316 -2904 2322 -2898
rect 2316 -2910 2322 -2904
rect 2316 -2916 2322 -2910
rect 2316 -2922 2322 -2916
rect 2316 -2928 2322 -2922
rect 2316 -2934 2322 -2928
rect 2322 -48 2328 -42
rect 2322 -54 2328 -48
rect 2322 -60 2328 -54
rect 2322 -66 2328 -60
rect 2322 -72 2328 -66
rect 2322 -78 2328 -72
rect 2322 -84 2328 -78
rect 2322 -90 2328 -84
rect 2322 -96 2328 -90
rect 2322 -102 2328 -96
rect 2322 -108 2328 -102
rect 2322 -114 2328 -108
rect 2322 -120 2328 -114
rect 2322 -126 2328 -120
rect 2322 -132 2328 -126
rect 2322 -138 2328 -132
rect 2322 -144 2328 -138
rect 2322 -150 2328 -144
rect 2322 -156 2328 -150
rect 2322 -162 2328 -156
rect 2322 -168 2328 -162
rect 2322 -174 2328 -168
rect 2322 -180 2328 -174
rect 2322 -186 2328 -180
rect 2322 -192 2328 -186
rect 2322 -198 2328 -192
rect 2322 -204 2328 -198
rect 2322 -210 2328 -204
rect 2322 -216 2328 -210
rect 2322 -222 2328 -216
rect 2322 -228 2328 -222
rect 2322 -234 2328 -228
rect 2322 -240 2328 -234
rect 2322 -246 2328 -240
rect 2322 -252 2328 -246
rect 2322 -258 2328 -252
rect 2322 -264 2328 -258
rect 2322 -270 2328 -264
rect 2322 -276 2328 -270
rect 2322 -282 2328 -276
rect 2322 -288 2328 -282
rect 2322 -294 2328 -288
rect 2322 -300 2328 -294
rect 2322 -306 2328 -300
rect 2322 -312 2328 -306
rect 2322 -318 2328 -312
rect 2322 -324 2328 -318
rect 2322 -330 2328 -324
rect 2322 -336 2328 -330
rect 2322 -342 2328 -336
rect 2322 -348 2328 -342
rect 2322 -354 2328 -348
rect 2322 -360 2328 -354
rect 2322 -366 2328 -360
rect 2322 -372 2328 -366
rect 2322 -378 2328 -372
rect 2322 -384 2328 -378
rect 2322 -390 2328 -384
rect 2322 -396 2328 -390
rect 2322 -402 2328 -396
rect 2322 -408 2328 -402
rect 2322 -414 2328 -408
rect 2322 -420 2328 -414
rect 2322 -426 2328 -420
rect 2322 -432 2328 -426
rect 2322 -438 2328 -432
rect 2322 -444 2328 -438
rect 2322 -450 2328 -444
rect 2322 -456 2328 -450
rect 2322 -462 2328 -456
rect 2322 -468 2328 -462
rect 2322 -474 2328 -468
rect 2322 -480 2328 -474
rect 2322 -486 2328 -480
rect 2322 -492 2328 -486
rect 2322 -498 2328 -492
rect 2322 -504 2328 -498
rect 2322 -510 2328 -504
rect 2322 -516 2328 -510
rect 2322 -522 2328 -516
rect 2322 -528 2328 -522
rect 2322 -534 2328 -528
rect 2322 -540 2328 -534
rect 2322 -546 2328 -540
rect 2322 -552 2328 -546
rect 2322 -558 2328 -552
rect 2322 -564 2328 -558
rect 2322 -570 2328 -564
rect 2322 -576 2328 -570
rect 2322 -582 2328 -576
rect 2322 -588 2328 -582
rect 2322 -594 2328 -588
rect 2322 -600 2328 -594
rect 2322 -606 2328 -600
rect 2322 -612 2328 -606
rect 2322 -618 2328 -612
rect 2322 -624 2328 -618
rect 2322 -630 2328 -624
rect 2322 -636 2328 -630
rect 2322 -642 2328 -636
rect 2322 -648 2328 -642
rect 2322 -654 2328 -648
rect 2322 -660 2328 -654
rect 2322 -666 2328 -660
rect 2322 -672 2328 -666
rect 2322 -678 2328 -672
rect 2322 -684 2328 -678
rect 2322 -690 2328 -684
rect 2322 -696 2328 -690
rect 2322 -702 2328 -696
rect 2322 -708 2328 -702
rect 2322 -714 2328 -708
rect 2322 -720 2328 -714
rect 2322 -726 2328 -720
rect 2322 -732 2328 -726
rect 2322 -738 2328 -732
rect 2322 -744 2328 -738
rect 2322 -750 2328 -744
rect 2322 -756 2328 -750
rect 2322 -762 2328 -756
rect 2322 -768 2328 -762
rect 2322 -774 2328 -768
rect 2322 -780 2328 -774
rect 2322 -786 2328 -780
rect 2322 -792 2328 -786
rect 2322 -798 2328 -792
rect 2322 -804 2328 -798
rect 2322 -810 2328 -804
rect 2322 -816 2328 -810
rect 2322 -822 2328 -816
rect 2322 -828 2328 -822
rect 2322 -834 2328 -828
rect 2322 -840 2328 -834
rect 2322 -846 2328 -840
rect 2322 -852 2328 -846
rect 2322 -858 2328 -852
rect 2322 -864 2328 -858
rect 2322 -870 2328 -864
rect 2322 -876 2328 -870
rect 2322 -882 2328 -876
rect 2322 -888 2328 -882
rect 2322 -894 2328 -888
rect 2322 -900 2328 -894
rect 2322 -906 2328 -900
rect 2322 -912 2328 -906
rect 2322 -918 2328 -912
rect 2322 -924 2328 -918
rect 2322 -930 2328 -924
rect 2322 -1452 2328 -1446
rect 2322 -1458 2328 -1452
rect 2322 -1464 2328 -1458
rect 2322 -1470 2328 -1464
rect 2322 -1476 2328 -1470
rect 2322 -1482 2328 -1476
rect 2322 -1488 2328 -1482
rect 2322 -1494 2328 -1488
rect 2322 -1500 2328 -1494
rect 2322 -1506 2328 -1500
rect 2322 -1512 2328 -1506
rect 2322 -1518 2328 -1512
rect 2322 -1524 2328 -1518
rect 2322 -1530 2328 -1524
rect 2322 -1536 2328 -1530
rect 2322 -1542 2328 -1536
rect 2322 -1548 2328 -1542
rect 2322 -1554 2328 -1548
rect 2322 -1560 2328 -1554
rect 2322 -1566 2328 -1560
rect 2322 -1572 2328 -1566
rect 2322 -1578 2328 -1572
rect 2322 -1584 2328 -1578
rect 2322 -1590 2328 -1584
rect 2322 -1596 2328 -1590
rect 2322 -1602 2328 -1596
rect 2322 -1608 2328 -1602
rect 2322 -1614 2328 -1608
rect 2322 -1620 2328 -1614
rect 2322 -1626 2328 -1620
rect 2322 -1632 2328 -1626
rect 2322 -1638 2328 -1632
rect 2322 -1644 2328 -1638
rect 2322 -1650 2328 -1644
rect 2322 -1656 2328 -1650
rect 2322 -1662 2328 -1656
rect 2322 -1668 2328 -1662
rect 2322 -1674 2328 -1668
rect 2322 -1680 2328 -1674
rect 2322 -1686 2328 -1680
rect 2322 -1692 2328 -1686
rect 2322 -1698 2328 -1692
rect 2322 -1704 2328 -1698
rect 2322 -1710 2328 -1704
rect 2322 -1716 2328 -1710
rect 2322 -1722 2328 -1716
rect 2322 -1728 2328 -1722
rect 2322 -1734 2328 -1728
rect 2322 -1740 2328 -1734
rect 2322 -1746 2328 -1740
rect 2322 -1752 2328 -1746
rect 2322 -1758 2328 -1752
rect 2322 -1764 2328 -1758
rect 2322 -1770 2328 -1764
rect 2322 -1776 2328 -1770
rect 2322 -1782 2328 -1776
rect 2322 -1788 2328 -1782
rect 2322 -1794 2328 -1788
rect 2322 -1800 2328 -1794
rect 2322 -1806 2328 -1800
rect 2322 -1812 2328 -1806
rect 2322 -1818 2328 -1812
rect 2322 -1824 2328 -1818
rect 2322 -1830 2328 -1824
rect 2322 -1836 2328 -1830
rect 2322 -1842 2328 -1836
rect 2322 -1848 2328 -1842
rect 2322 -1854 2328 -1848
rect 2322 -1860 2328 -1854
rect 2322 -1866 2328 -1860
rect 2322 -1872 2328 -1866
rect 2322 -1878 2328 -1872
rect 2322 -1884 2328 -1878
rect 2322 -1890 2328 -1884
rect 2322 -1896 2328 -1890
rect 2322 -1902 2328 -1896
rect 2322 -1908 2328 -1902
rect 2322 -1914 2328 -1908
rect 2322 -1920 2328 -1914
rect 2322 -1926 2328 -1920
rect 2322 -1932 2328 -1926
rect 2322 -1938 2328 -1932
rect 2322 -1944 2328 -1938
rect 2322 -1950 2328 -1944
rect 2322 -1956 2328 -1950
rect 2322 -1962 2328 -1956
rect 2322 -1968 2328 -1962
rect 2322 -1974 2328 -1968
rect 2322 -1980 2328 -1974
rect 2322 -1986 2328 -1980
rect 2322 -1992 2328 -1986
rect 2322 -1998 2328 -1992
rect 2322 -2004 2328 -1998
rect 2322 -2010 2328 -2004
rect 2322 -2016 2328 -2010
rect 2322 -2022 2328 -2016
rect 2322 -2028 2328 -2022
rect 2322 -2034 2328 -2028
rect 2322 -2040 2328 -2034
rect 2322 -2046 2328 -2040
rect 2322 -2052 2328 -2046
rect 2322 -2058 2328 -2052
rect 2322 -2064 2328 -2058
rect 2322 -2070 2328 -2064
rect 2322 -2076 2328 -2070
rect 2322 -2082 2328 -2076
rect 2322 -2088 2328 -2082
rect 2322 -2094 2328 -2088
rect 2322 -2100 2328 -2094
rect 2322 -2106 2328 -2100
rect 2322 -2112 2328 -2106
rect 2322 -2118 2328 -2112
rect 2322 -2124 2328 -2118
rect 2322 -2130 2328 -2124
rect 2322 -2136 2328 -2130
rect 2322 -2142 2328 -2136
rect 2322 -2148 2328 -2142
rect 2322 -2154 2328 -2148
rect 2322 -2160 2328 -2154
rect 2322 -2166 2328 -2160
rect 2322 -2172 2328 -2166
rect 2322 -2178 2328 -2172
rect 2322 -2184 2328 -2178
rect 2322 -2190 2328 -2184
rect 2322 -2196 2328 -2190
rect 2322 -2268 2328 -2262
rect 2322 -2274 2328 -2268
rect 2322 -2280 2328 -2274
rect 2322 -2286 2328 -2280
rect 2322 -2292 2328 -2286
rect 2322 -2298 2328 -2292
rect 2322 -2304 2328 -2298
rect 2322 -2310 2328 -2304
rect 2322 -2316 2328 -2310
rect 2322 -2322 2328 -2316
rect 2322 -2328 2328 -2322
rect 2322 -2334 2328 -2328
rect 2322 -2340 2328 -2334
rect 2322 -2346 2328 -2340
rect 2322 -2352 2328 -2346
rect 2322 -2358 2328 -2352
rect 2322 -2364 2328 -2358
rect 2322 -2370 2328 -2364
rect 2322 -2376 2328 -2370
rect 2322 -2382 2328 -2376
rect 2322 -2388 2328 -2382
rect 2322 -2394 2328 -2388
rect 2322 -2400 2328 -2394
rect 2322 -2406 2328 -2400
rect 2322 -2412 2328 -2406
rect 2322 -2418 2328 -2412
rect 2322 -2424 2328 -2418
rect 2322 -2430 2328 -2424
rect 2322 -2436 2328 -2430
rect 2322 -2502 2328 -2496
rect 2322 -2508 2328 -2502
rect 2322 -2514 2328 -2508
rect 2322 -2520 2328 -2514
rect 2322 -2526 2328 -2520
rect 2322 -2532 2328 -2526
rect 2322 -2538 2328 -2532
rect 2322 -2544 2328 -2538
rect 2322 -2550 2328 -2544
rect 2322 -2556 2328 -2550
rect 2322 -2562 2328 -2556
rect 2322 -2568 2328 -2562
rect 2322 -2574 2328 -2568
rect 2322 -2580 2328 -2574
rect 2322 -2586 2328 -2580
rect 2322 -2592 2328 -2586
rect 2322 -2598 2328 -2592
rect 2322 -2604 2328 -2598
rect 2322 -2610 2328 -2604
rect 2322 -2616 2328 -2610
rect 2322 -2622 2328 -2616
rect 2322 -2628 2328 -2622
rect 2322 -2634 2328 -2628
rect 2322 -2640 2328 -2634
rect 2322 -2646 2328 -2640
rect 2322 -2652 2328 -2646
rect 2322 -2658 2328 -2652
rect 2322 -2664 2328 -2658
rect 2322 -2670 2328 -2664
rect 2322 -2676 2328 -2670
rect 2322 -2682 2328 -2676
rect 2322 -2688 2328 -2682
rect 2322 -2694 2328 -2688
rect 2322 -2700 2328 -2694
rect 2322 -2706 2328 -2700
rect 2322 -2712 2328 -2706
rect 2322 -2718 2328 -2712
rect 2322 -2724 2328 -2718
rect 2322 -2730 2328 -2724
rect 2322 -2736 2328 -2730
rect 2322 -2742 2328 -2736
rect 2322 -2748 2328 -2742
rect 2322 -2754 2328 -2748
rect 2322 -2760 2328 -2754
rect 2322 -2766 2328 -2760
rect 2322 -2772 2328 -2766
rect 2322 -2778 2328 -2772
rect 2322 -2784 2328 -2778
rect 2322 -2790 2328 -2784
rect 2322 -2796 2328 -2790
rect 2322 -2802 2328 -2796
rect 2322 -2808 2328 -2802
rect 2322 -2814 2328 -2808
rect 2322 -2820 2328 -2814
rect 2322 -2826 2328 -2820
rect 2322 -2832 2328 -2826
rect 2322 -2838 2328 -2832
rect 2322 -2844 2328 -2838
rect 2322 -2850 2328 -2844
rect 2322 -2856 2328 -2850
rect 2322 -2862 2328 -2856
rect 2322 -2868 2328 -2862
rect 2322 -2874 2328 -2868
rect 2322 -2880 2328 -2874
rect 2322 -2886 2328 -2880
rect 2322 -2892 2328 -2886
rect 2322 -2898 2328 -2892
rect 2322 -2904 2328 -2898
rect 2322 -2910 2328 -2904
rect 2322 -2916 2328 -2910
rect 2322 -2922 2328 -2916
rect 2322 -2928 2328 -2922
rect 2322 -2934 2328 -2928
rect 2328 -42 2334 -36
rect 2328 -48 2334 -42
rect 2328 -54 2334 -48
rect 2328 -60 2334 -54
rect 2328 -66 2334 -60
rect 2328 -72 2334 -66
rect 2328 -78 2334 -72
rect 2328 -84 2334 -78
rect 2328 -90 2334 -84
rect 2328 -96 2334 -90
rect 2328 -102 2334 -96
rect 2328 -108 2334 -102
rect 2328 -114 2334 -108
rect 2328 -120 2334 -114
rect 2328 -126 2334 -120
rect 2328 -132 2334 -126
rect 2328 -138 2334 -132
rect 2328 -144 2334 -138
rect 2328 -150 2334 -144
rect 2328 -156 2334 -150
rect 2328 -162 2334 -156
rect 2328 -168 2334 -162
rect 2328 -174 2334 -168
rect 2328 -180 2334 -174
rect 2328 -186 2334 -180
rect 2328 -192 2334 -186
rect 2328 -198 2334 -192
rect 2328 -204 2334 -198
rect 2328 -210 2334 -204
rect 2328 -216 2334 -210
rect 2328 -222 2334 -216
rect 2328 -228 2334 -222
rect 2328 -234 2334 -228
rect 2328 -240 2334 -234
rect 2328 -246 2334 -240
rect 2328 -252 2334 -246
rect 2328 -258 2334 -252
rect 2328 -264 2334 -258
rect 2328 -270 2334 -264
rect 2328 -276 2334 -270
rect 2328 -282 2334 -276
rect 2328 -288 2334 -282
rect 2328 -294 2334 -288
rect 2328 -300 2334 -294
rect 2328 -306 2334 -300
rect 2328 -312 2334 -306
rect 2328 -318 2334 -312
rect 2328 -324 2334 -318
rect 2328 -330 2334 -324
rect 2328 -336 2334 -330
rect 2328 -342 2334 -336
rect 2328 -348 2334 -342
rect 2328 -354 2334 -348
rect 2328 -360 2334 -354
rect 2328 -366 2334 -360
rect 2328 -372 2334 -366
rect 2328 -378 2334 -372
rect 2328 -384 2334 -378
rect 2328 -390 2334 -384
rect 2328 -396 2334 -390
rect 2328 -402 2334 -396
rect 2328 -408 2334 -402
rect 2328 -414 2334 -408
rect 2328 -420 2334 -414
rect 2328 -426 2334 -420
rect 2328 -432 2334 -426
rect 2328 -438 2334 -432
rect 2328 -444 2334 -438
rect 2328 -450 2334 -444
rect 2328 -456 2334 -450
rect 2328 -462 2334 -456
rect 2328 -468 2334 -462
rect 2328 -474 2334 -468
rect 2328 -480 2334 -474
rect 2328 -486 2334 -480
rect 2328 -492 2334 -486
rect 2328 -498 2334 -492
rect 2328 -504 2334 -498
rect 2328 -510 2334 -504
rect 2328 -516 2334 -510
rect 2328 -522 2334 -516
rect 2328 -528 2334 -522
rect 2328 -534 2334 -528
rect 2328 -540 2334 -534
rect 2328 -546 2334 -540
rect 2328 -552 2334 -546
rect 2328 -558 2334 -552
rect 2328 -564 2334 -558
rect 2328 -570 2334 -564
rect 2328 -576 2334 -570
rect 2328 -582 2334 -576
rect 2328 -588 2334 -582
rect 2328 -594 2334 -588
rect 2328 -600 2334 -594
rect 2328 -606 2334 -600
rect 2328 -612 2334 -606
rect 2328 -618 2334 -612
rect 2328 -624 2334 -618
rect 2328 -630 2334 -624
rect 2328 -636 2334 -630
rect 2328 -642 2334 -636
rect 2328 -648 2334 -642
rect 2328 -654 2334 -648
rect 2328 -660 2334 -654
rect 2328 -666 2334 -660
rect 2328 -672 2334 -666
rect 2328 -678 2334 -672
rect 2328 -684 2334 -678
rect 2328 -690 2334 -684
rect 2328 -696 2334 -690
rect 2328 -702 2334 -696
rect 2328 -708 2334 -702
rect 2328 -714 2334 -708
rect 2328 -720 2334 -714
rect 2328 -726 2334 -720
rect 2328 -732 2334 -726
rect 2328 -738 2334 -732
rect 2328 -744 2334 -738
rect 2328 -750 2334 -744
rect 2328 -756 2334 -750
rect 2328 -762 2334 -756
rect 2328 -768 2334 -762
rect 2328 -774 2334 -768
rect 2328 -780 2334 -774
rect 2328 -786 2334 -780
rect 2328 -792 2334 -786
rect 2328 -798 2334 -792
rect 2328 -804 2334 -798
rect 2328 -810 2334 -804
rect 2328 -816 2334 -810
rect 2328 -822 2334 -816
rect 2328 -828 2334 -822
rect 2328 -834 2334 -828
rect 2328 -840 2334 -834
rect 2328 -846 2334 -840
rect 2328 -852 2334 -846
rect 2328 -858 2334 -852
rect 2328 -864 2334 -858
rect 2328 -870 2334 -864
rect 2328 -876 2334 -870
rect 2328 -882 2334 -876
rect 2328 -888 2334 -882
rect 2328 -894 2334 -888
rect 2328 -900 2334 -894
rect 2328 -906 2334 -900
rect 2328 -912 2334 -906
rect 2328 -918 2334 -912
rect 2328 -1446 2334 -1440
rect 2328 -1452 2334 -1446
rect 2328 -1458 2334 -1452
rect 2328 -1464 2334 -1458
rect 2328 -1470 2334 -1464
rect 2328 -1476 2334 -1470
rect 2328 -1482 2334 -1476
rect 2328 -1488 2334 -1482
rect 2328 -1494 2334 -1488
rect 2328 -1500 2334 -1494
rect 2328 -1506 2334 -1500
rect 2328 -1512 2334 -1506
rect 2328 -1518 2334 -1512
rect 2328 -1524 2334 -1518
rect 2328 -1530 2334 -1524
rect 2328 -1536 2334 -1530
rect 2328 -1542 2334 -1536
rect 2328 -1548 2334 -1542
rect 2328 -1554 2334 -1548
rect 2328 -1560 2334 -1554
rect 2328 -1566 2334 -1560
rect 2328 -1572 2334 -1566
rect 2328 -1578 2334 -1572
rect 2328 -1584 2334 -1578
rect 2328 -1590 2334 -1584
rect 2328 -1596 2334 -1590
rect 2328 -1602 2334 -1596
rect 2328 -1608 2334 -1602
rect 2328 -1614 2334 -1608
rect 2328 -1620 2334 -1614
rect 2328 -1626 2334 -1620
rect 2328 -1632 2334 -1626
rect 2328 -1638 2334 -1632
rect 2328 -1644 2334 -1638
rect 2328 -1650 2334 -1644
rect 2328 -1656 2334 -1650
rect 2328 -1662 2334 -1656
rect 2328 -1668 2334 -1662
rect 2328 -1674 2334 -1668
rect 2328 -1680 2334 -1674
rect 2328 -1686 2334 -1680
rect 2328 -1692 2334 -1686
rect 2328 -1698 2334 -1692
rect 2328 -1704 2334 -1698
rect 2328 -1710 2334 -1704
rect 2328 -1716 2334 -1710
rect 2328 -1722 2334 -1716
rect 2328 -1728 2334 -1722
rect 2328 -1734 2334 -1728
rect 2328 -1740 2334 -1734
rect 2328 -1746 2334 -1740
rect 2328 -1752 2334 -1746
rect 2328 -1758 2334 -1752
rect 2328 -1764 2334 -1758
rect 2328 -1770 2334 -1764
rect 2328 -1776 2334 -1770
rect 2328 -1782 2334 -1776
rect 2328 -1788 2334 -1782
rect 2328 -1794 2334 -1788
rect 2328 -1800 2334 -1794
rect 2328 -1806 2334 -1800
rect 2328 -1812 2334 -1806
rect 2328 -1818 2334 -1812
rect 2328 -1824 2334 -1818
rect 2328 -1830 2334 -1824
rect 2328 -1836 2334 -1830
rect 2328 -1842 2334 -1836
rect 2328 -1848 2334 -1842
rect 2328 -1854 2334 -1848
rect 2328 -1860 2334 -1854
rect 2328 -1866 2334 -1860
rect 2328 -1872 2334 -1866
rect 2328 -1878 2334 -1872
rect 2328 -1884 2334 -1878
rect 2328 -1890 2334 -1884
rect 2328 -1896 2334 -1890
rect 2328 -1902 2334 -1896
rect 2328 -1908 2334 -1902
rect 2328 -1914 2334 -1908
rect 2328 -1920 2334 -1914
rect 2328 -1926 2334 -1920
rect 2328 -1932 2334 -1926
rect 2328 -1938 2334 -1932
rect 2328 -1944 2334 -1938
rect 2328 -1950 2334 -1944
rect 2328 -1956 2334 -1950
rect 2328 -1962 2334 -1956
rect 2328 -1968 2334 -1962
rect 2328 -1974 2334 -1968
rect 2328 -1980 2334 -1974
rect 2328 -1986 2334 -1980
rect 2328 -1992 2334 -1986
rect 2328 -1998 2334 -1992
rect 2328 -2004 2334 -1998
rect 2328 -2010 2334 -2004
rect 2328 -2016 2334 -2010
rect 2328 -2022 2334 -2016
rect 2328 -2028 2334 -2022
rect 2328 -2034 2334 -2028
rect 2328 -2040 2334 -2034
rect 2328 -2046 2334 -2040
rect 2328 -2052 2334 -2046
rect 2328 -2058 2334 -2052
rect 2328 -2064 2334 -2058
rect 2328 -2070 2334 -2064
rect 2328 -2076 2334 -2070
rect 2328 -2082 2334 -2076
rect 2328 -2088 2334 -2082
rect 2328 -2094 2334 -2088
rect 2328 -2100 2334 -2094
rect 2328 -2106 2334 -2100
rect 2328 -2112 2334 -2106
rect 2328 -2118 2334 -2112
rect 2328 -2124 2334 -2118
rect 2328 -2130 2334 -2124
rect 2328 -2136 2334 -2130
rect 2328 -2142 2334 -2136
rect 2328 -2148 2334 -2142
rect 2328 -2154 2334 -2148
rect 2328 -2160 2334 -2154
rect 2328 -2166 2334 -2160
rect 2328 -2172 2334 -2166
rect 2328 -2178 2334 -2172
rect 2328 -2184 2334 -2178
rect 2328 -2262 2334 -2256
rect 2328 -2268 2334 -2262
rect 2328 -2274 2334 -2268
rect 2328 -2280 2334 -2274
rect 2328 -2286 2334 -2280
rect 2328 -2292 2334 -2286
rect 2328 -2298 2334 -2292
rect 2328 -2304 2334 -2298
rect 2328 -2310 2334 -2304
rect 2328 -2316 2334 -2310
rect 2328 -2322 2334 -2316
rect 2328 -2328 2334 -2322
rect 2328 -2334 2334 -2328
rect 2328 -2340 2334 -2334
rect 2328 -2346 2334 -2340
rect 2328 -2352 2334 -2346
rect 2328 -2358 2334 -2352
rect 2328 -2364 2334 -2358
rect 2328 -2370 2334 -2364
rect 2328 -2376 2334 -2370
rect 2328 -2382 2334 -2376
rect 2328 -2388 2334 -2382
rect 2328 -2394 2334 -2388
rect 2328 -2400 2334 -2394
rect 2328 -2406 2334 -2400
rect 2328 -2412 2334 -2406
rect 2328 -2418 2334 -2412
rect 2328 -2424 2334 -2418
rect 2328 -2430 2334 -2424
rect 2328 -2436 2334 -2430
rect 2328 -2496 2334 -2490
rect 2328 -2502 2334 -2496
rect 2328 -2508 2334 -2502
rect 2328 -2514 2334 -2508
rect 2328 -2520 2334 -2514
rect 2328 -2526 2334 -2520
rect 2328 -2532 2334 -2526
rect 2328 -2538 2334 -2532
rect 2328 -2544 2334 -2538
rect 2328 -2550 2334 -2544
rect 2328 -2556 2334 -2550
rect 2328 -2562 2334 -2556
rect 2328 -2568 2334 -2562
rect 2328 -2574 2334 -2568
rect 2328 -2580 2334 -2574
rect 2328 -2586 2334 -2580
rect 2328 -2592 2334 -2586
rect 2328 -2598 2334 -2592
rect 2328 -2604 2334 -2598
rect 2328 -2610 2334 -2604
rect 2328 -2616 2334 -2610
rect 2328 -2622 2334 -2616
rect 2328 -2628 2334 -2622
rect 2328 -2634 2334 -2628
rect 2328 -2640 2334 -2634
rect 2328 -2646 2334 -2640
rect 2328 -2652 2334 -2646
rect 2328 -2658 2334 -2652
rect 2328 -2664 2334 -2658
rect 2328 -2670 2334 -2664
rect 2328 -2676 2334 -2670
rect 2328 -2682 2334 -2676
rect 2328 -2688 2334 -2682
rect 2328 -2694 2334 -2688
rect 2328 -2700 2334 -2694
rect 2328 -2706 2334 -2700
rect 2328 -2712 2334 -2706
rect 2328 -2718 2334 -2712
rect 2328 -2724 2334 -2718
rect 2328 -2730 2334 -2724
rect 2328 -2736 2334 -2730
rect 2328 -2742 2334 -2736
rect 2328 -2748 2334 -2742
rect 2328 -2754 2334 -2748
rect 2328 -2760 2334 -2754
rect 2328 -2766 2334 -2760
rect 2328 -2772 2334 -2766
rect 2328 -2778 2334 -2772
rect 2328 -2784 2334 -2778
rect 2328 -2790 2334 -2784
rect 2328 -2796 2334 -2790
rect 2328 -2802 2334 -2796
rect 2328 -2808 2334 -2802
rect 2328 -2814 2334 -2808
rect 2328 -2820 2334 -2814
rect 2328 -2826 2334 -2820
rect 2328 -2832 2334 -2826
rect 2328 -2838 2334 -2832
rect 2328 -2844 2334 -2838
rect 2328 -2850 2334 -2844
rect 2328 -2856 2334 -2850
rect 2328 -2862 2334 -2856
rect 2328 -2868 2334 -2862
rect 2328 -2874 2334 -2868
rect 2328 -2880 2334 -2874
rect 2328 -2886 2334 -2880
rect 2328 -2892 2334 -2886
rect 2328 -2898 2334 -2892
rect 2328 -2904 2334 -2898
rect 2328 -2910 2334 -2904
rect 2328 -2916 2334 -2910
rect 2328 -2922 2334 -2916
rect 2328 -2928 2334 -2922
rect 2334 -36 2340 -30
rect 2334 -42 2340 -36
rect 2334 -48 2340 -42
rect 2334 -54 2340 -48
rect 2334 -60 2340 -54
rect 2334 -66 2340 -60
rect 2334 -72 2340 -66
rect 2334 -78 2340 -72
rect 2334 -84 2340 -78
rect 2334 -90 2340 -84
rect 2334 -96 2340 -90
rect 2334 -102 2340 -96
rect 2334 -108 2340 -102
rect 2334 -114 2340 -108
rect 2334 -120 2340 -114
rect 2334 -126 2340 -120
rect 2334 -132 2340 -126
rect 2334 -138 2340 -132
rect 2334 -144 2340 -138
rect 2334 -150 2340 -144
rect 2334 -156 2340 -150
rect 2334 -162 2340 -156
rect 2334 -168 2340 -162
rect 2334 -174 2340 -168
rect 2334 -180 2340 -174
rect 2334 -186 2340 -180
rect 2334 -192 2340 -186
rect 2334 -198 2340 -192
rect 2334 -204 2340 -198
rect 2334 -210 2340 -204
rect 2334 -216 2340 -210
rect 2334 -222 2340 -216
rect 2334 -228 2340 -222
rect 2334 -234 2340 -228
rect 2334 -240 2340 -234
rect 2334 -246 2340 -240
rect 2334 -252 2340 -246
rect 2334 -258 2340 -252
rect 2334 -264 2340 -258
rect 2334 -270 2340 -264
rect 2334 -276 2340 -270
rect 2334 -282 2340 -276
rect 2334 -288 2340 -282
rect 2334 -294 2340 -288
rect 2334 -300 2340 -294
rect 2334 -306 2340 -300
rect 2334 -312 2340 -306
rect 2334 -318 2340 -312
rect 2334 -324 2340 -318
rect 2334 -330 2340 -324
rect 2334 -336 2340 -330
rect 2334 -342 2340 -336
rect 2334 -348 2340 -342
rect 2334 -354 2340 -348
rect 2334 -360 2340 -354
rect 2334 -366 2340 -360
rect 2334 -372 2340 -366
rect 2334 -378 2340 -372
rect 2334 -384 2340 -378
rect 2334 -390 2340 -384
rect 2334 -396 2340 -390
rect 2334 -402 2340 -396
rect 2334 -408 2340 -402
rect 2334 -414 2340 -408
rect 2334 -420 2340 -414
rect 2334 -426 2340 -420
rect 2334 -432 2340 -426
rect 2334 -438 2340 -432
rect 2334 -444 2340 -438
rect 2334 -450 2340 -444
rect 2334 -456 2340 -450
rect 2334 -462 2340 -456
rect 2334 -468 2340 -462
rect 2334 -474 2340 -468
rect 2334 -480 2340 -474
rect 2334 -486 2340 -480
rect 2334 -492 2340 -486
rect 2334 -498 2340 -492
rect 2334 -504 2340 -498
rect 2334 -510 2340 -504
rect 2334 -516 2340 -510
rect 2334 -522 2340 -516
rect 2334 -528 2340 -522
rect 2334 -534 2340 -528
rect 2334 -540 2340 -534
rect 2334 -546 2340 -540
rect 2334 -552 2340 -546
rect 2334 -558 2340 -552
rect 2334 -564 2340 -558
rect 2334 -570 2340 -564
rect 2334 -576 2340 -570
rect 2334 -582 2340 -576
rect 2334 -588 2340 -582
rect 2334 -594 2340 -588
rect 2334 -600 2340 -594
rect 2334 -606 2340 -600
rect 2334 -612 2340 -606
rect 2334 -618 2340 -612
rect 2334 -624 2340 -618
rect 2334 -630 2340 -624
rect 2334 -636 2340 -630
rect 2334 -642 2340 -636
rect 2334 -648 2340 -642
rect 2334 -654 2340 -648
rect 2334 -660 2340 -654
rect 2334 -666 2340 -660
rect 2334 -672 2340 -666
rect 2334 -678 2340 -672
rect 2334 -684 2340 -678
rect 2334 -690 2340 -684
rect 2334 -696 2340 -690
rect 2334 -702 2340 -696
rect 2334 -708 2340 -702
rect 2334 -714 2340 -708
rect 2334 -720 2340 -714
rect 2334 -726 2340 -720
rect 2334 -732 2340 -726
rect 2334 -738 2340 -732
rect 2334 -744 2340 -738
rect 2334 -750 2340 -744
rect 2334 -756 2340 -750
rect 2334 -762 2340 -756
rect 2334 -768 2340 -762
rect 2334 -774 2340 -768
rect 2334 -780 2340 -774
rect 2334 -786 2340 -780
rect 2334 -792 2340 -786
rect 2334 -798 2340 -792
rect 2334 -804 2340 -798
rect 2334 -810 2340 -804
rect 2334 -816 2340 -810
rect 2334 -822 2340 -816
rect 2334 -828 2340 -822
rect 2334 -834 2340 -828
rect 2334 -840 2340 -834
rect 2334 -846 2340 -840
rect 2334 -852 2340 -846
rect 2334 -858 2340 -852
rect 2334 -864 2340 -858
rect 2334 -870 2340 -864
rect 2334 -876 2340 -870
rect 2334 -882 2340 -876
rect 2334 -888 2340 -882
rect 2334 -894 2340 -888
rect 2334 -900 2340 -894
rect 2334 -1440 2340 -1434
rect 2334 -1446 2340 -1440
rect 2334 -1452 2340 -1446
rect 2334 -1458 2340 -1452
rect 2334 -1464 2340 -1458
rect 2334 -1470 2340 -1464
rect 2334 -1476 2340 -1470
rect 2334 -1482 2340 -1476
rect 2334 -1488 2340 -1482
rect 2334 -1494 2340 -1488
rect 2334 -1500 2340 -1494
rect 2334 -1506 2340 -1500
rect 2334 -1512 2340 -1506
rect 2334 -1518 2340 -1512
rect 2334 -1524 2340 -1518
rect 2334 -1530 2340 -1524
rect 2334 -1536 2340 -1530
rect 2334 -1542 2340 -1536
rect 2334 -1548 2340 -1542
rect 2334 -1554 2340 -1548
rect 2334 -1560 2340 -1554
rect 2334 -1566 2340 -1560
rect 2334 -1572 2340 -1566
rect 2334 -1578 2340 -1572
rect 2334 -1584 2340 -1578
rect 2334 -1590 2340 -1584
rect 2334 -1596 2340 -1590
rect 2334 -1602 2340 -1596
rect 2334 -1608 2340 -1602
rect 2334 -1614 2340 -1608
rect 2334 -1620 2340 -1614
rect 2334 -1626 2340 -1620
rect 2334 -1632 2340 -1626
rect 2334 -1638 2340 -1632
rect 2334 -1644 2340 -1638
rect 2334 -1650 2340 -1644
rect 2334 -1656 2340 -1650
rect 2334 -1662 2340 -1656
rect 2334 -1668 2340 -1662
rect 2334 -1674 2340 -1668
rect 2334 -1680 2340 -1674
rect 2334 -1686 2340 -1680
rect 2334 -1692 2340 -1686
rect 2334 -1698 2340 -1692
rect 2334 -1704 2340 -1698
rect 2334 -1710 2340 -1704
rect 2334 -1716 2340 -1710
rect 2334 -1722 2340 -1716
rect 2334 -1728 2340 -1722
rect 2334 -1734 2340 -1728
rect 2334 -1740 2340 -1734
rect 2334 -1746 2340 -1740
rect 2334 -1752 2340 -1746
rect 2334 -1758 2340 -1752
rect 2334 -1764 2340 -1758
rect 2334 -1770 2340 -1764
rect 2334 -1776 2340 -1770
rect 2334 -1782 2340 -1776
rect 2334 -1788 2340 -1782
rect 2334 -1794 2340 -1788
rect 2334 -1800 2340 -1794
rect 2334 -1806 2340 -1800
rect 2334 -1812 2340 -1806
rect 2334 -1818 2340 -1812
rect 2334 -1824 2340 -1818
rect 2334 -1830 2340 -1824
rect 2334 -1836 2340 -1830
rect 2334 -1842 2340 -1836
rect 2334 -1848 2340 -1842
rect 2334 -1854 2340 -1848
rect 2334 -1860 2340 -1854
rect 2334 -1866 2340 -1860
rect 2334 -1872 2340 -1866
rect 2334 -1878 2340 -1872
rect 2334 -1884 2340 -1878
rect 2334 -1890 2340 -1884
rect 2334 -1896 2340 -1890
rect 2334 -1902 2340 -1896
rect 2334 -1908 2340 -1902
rect 2334 -1914 2340 -1908
rect 2334 -1920 2340 -1914
rect 2334 -1926 2340 -1920
rect 2334 -1932 2340 -1926
rect 2334 -1938 2340 -1932
rect 2334 -1944 2340 -1938
rect 2334 -1950 2340 -1944
rect 2334 -1956 2340 -1950
rect 2334 -1962 2340 -1956
rect 2334 -1968 2340 -1962
rect 2334 -1974 2340 -1968
rect 2334 -1980 2340 -1974
rect 2334 -1986 2340 -1980
rect 2334 -1992 2340 -1986
rect 2334 -1998 2340 -1992
rect 2334 -2004 2340 -1998
rect 2334 -2010 2340 -2004
rect 2334 -2016 2340 -2010
rect 2334 -2022 2340 -2016
rect 2334 -2028 2340 -2022
rect 2334 -2034 2340 -2028
rect 2334 -2040 2340 -2034
rect 2334 -2046 2340 -2040
rect 2334 -2052 2340 -2046
rect 2334 -2058 2340 -2052
rect 2334 -2064 2340 -2058
rect 2334 -2070 2340 -2064
rect 2334 -2076 2340 -2070
rect 2334 -2082 2340 -2076
rect 2334 -2088 2340 -2082
rect 2334 -2094 2340 -2088
rect 2334 -2100 2340 -2094
rect 2334 -2106 2340 -2100
rect 2334 -2112 2340 -2106
rect 2334 -2118 2340 -2112
rect 2334 -2124 2340 -2118
rect 2334 -2130 2340 -2124
rect 2334 -2136 2340 -2130
rect 2334 -2142 2340 -2136
rect 2334 -2148 2340 -2142
rect 2334 -2154 2340 -2148
rect 2334 -2160 2340 -2154
rect 2334 -2166 2340 -2160
rect 2334 -2172 2340 -2166
rect 2334 -2178 2340 -2172
rect 2334 -2256 2340 -2250
rect 2334 -2262 2340 -2256
rect 2334 -2268 2340 -2262
rect 2334 -2274 2340 -2268
rect 2334 -2280 2340 -2274
rect 2334 -2286 2340 -2280
rect 2334 -2292 2340 -2286
rect 2334 -2298 2340 -2292
rect 2334 -2304 2340 -2298
rect 2334 -2310 2340 -2304
rect 2334 -2316 2340 -2310
rect 2334 -2322 2340 -2316
rect 2334 -2328 2340 -2322
rect 2334 -2334 2340 -2328
rect 2334 -2340 2340 -2334
rect 2334 -2346 2340 -2340
rect 2334 -2352 2340 -2346
rect 2334 -2358 2340 -2352
rect 2334 -2364 2340 -2358
rect 2334 -2370 2340 -2364
rect 2334 -2376 2340 -2370
rect 2334 -2382 2340 -2376
rect 2334 -2388 2340 -2382
rect 2334 -2394 2340 -2388
rect 2334 -2400 2340 -2394
rect 2334 -2406 2340 -2400
rect 2334 -2412 2340 -2406
rect 2334 -2418 2340 -2412
rect 2334 -2424 2340 -2418
rect 2334 -2430 2340 -2424
rect 2334 -2496 2340 -2490
rect 2334 -2502 2340 -2496
rect 2334 -2508 2340 -2502
rect 2334 -2514 2340 -2508
rect 2334 -2520 2340 -2514
rect 2334 -2526 2340 -2520
rect 2334 -2532 2340 -2526
rect 2334 -2538 2340 -2532
rect 2334 -2544 2340 -2538
rect 2334 -2550 2340 -2544
rect 2334 -2556 2340 -2550
rect 2334 -2562 2340 -2556
rect 2334 -2568 2340 -2562
rect 2334 -2574 2340 -2568
rect 2334 -2580 2340 -2574
rect 2334 -2586 2340 -2580
rect 2334 -2592 2340 -2586
rect 2334 -2598 2340 -2592
rect 2334 -2604 2340 -2598
rect 2334 -2610 2340 -2604
rect 2334 -2616 2340 -2610
rect 2334 -2622 2340 -2616
rect 2334 -2628 2340 -2622
rect 2334 -2634 2340 -2628
rect 2334 -2640 2340 -2634
rect 2334 -2646 2340 -2640
rect 2334 -2652 2340 -2646
rect 2334 -2658 2340 -2652
rect 2334 -2664 2340 -2658
rect 2334 -2670 2340 -2664
rect 2334 -2676 2340 -2670
rect 2334 -2682 2340 -2676
rect 2334 -2688 2340 -2682
rect 2334 -2694 2340 -2688
rect 2334 -2700 2340 -2694
rect 2334 -2706 2340 -2700
rect 2334 -2712 2340 -2706
rect 2334 -2718 2340 -2712
rect 2334 -2724 2340 -2718
rect 2334 -2730 2340 -2724
rect 2334 -2736 2340 -2730
rect 2334 -2742 2340 -2736
rect 2334 -2748 2340 -2742
rect 2334 -2754 2340 -2748
rect 2334 -2760 2340 -2754
rect 2334 -2766 2340 -2760
rect 2334 -2772 2340 -2766
rect 2334 -2778 2340 -2772
rect 2334 -2784 2340 -2778
rect 2334 -2790 2340 -2784
rect 2334 -2796 2340 -2790
rect 2334 -2802 2340 -2796
rect 2334 -2808 2340 -2802
rect 2334 -2814 2340 -2808
rect 2334 -2820 2340 -2814
rect 2334 -2826 2340 -2820
rect 2334 -2832 2340 -2826
rect 2334 -2838 2340 -2832
rect 2334 -2844 2340 -2838
rect 2334 -2850 2340 -2844
rect 2334 -2856 2340 -2850
rect 2334 -2862 2340 -2856
rect 2334 -2868 2340 -2862
rect 2334 -2874 2340 -2868
rect 2334 -2880 2340 -2874
rect 2334 -2886 2340 -2880
rect 2334 -2892 2340 -2886
rect 2334 -2898 2340 -2892
rect 2334 -2904 2340 -2898
rect 2334 -2910 2340 -2904
rect 2334 -2916 2340 -2910
rect 2334 -2922 2340 -2916
rect 2334 -2928 2340 -2922
rect 2340 -24 2346 -18
rect 2340 -30 2346 -24
rect 2340 -36 2346 -30
rect 2340 -42 2346 -36
rect 2340 -48 2346 -42
rect 2340 -54 2346 -48
rect 2340 -60 2346 -54
rect 2340 -66 2346 -60
rect 2340 -72 2346 -66
rect 2340 -78 2346 -72
rect 2340 -84 2346 -78
rect 2340 -90 2346 -84
rect 2340 -96 2346 -90
rect 2340 -102 2346 -96
rect 2340 -108 2346 -102
rect 2340 -114 2346 -108
rect 2340 -120 2346 -114
rect 2340 -126 2346 -120
rect 2340 -132 2346 -126
rect 2340 -138 2346 -132
rect 2340 -144 2346 -138
rect 2340 -150 2346 -144
rect 2340 -156 2346 -150
rect 2340 -162 2346 -156
rect 2340 -168 2346 -162
rect 2340 -174 2346 -168
rect 2340 -180 2346 -174
rect 2340 -186 2346 -180
rect 2340 -192 2346 -186
rect 2340 -198 2346 -192
rect 2340 -204 2346 -198
rect 2340 -210 2346 -204
rect 2340 -216 2346 -210
rect 2340 -222 2346 -216
rect 2340 -228 2346 -222
rect 2340 -234 2346 -228
rect 2340 -240 2346 -234
rect 2340 -246 2346 -240
rect 2340 -252 2346 -246
rect 2340 -258 2346 -252
rect 2340 -264 2346 -258
rect 2340 -270 2346 -264
rect 2340 -276 2346 -270
rect 2340 -282 2346 -276
rect 2340 -288 2346 -282
rect 2340 -294 2346 -288
rect 2340 -300 2346 -294
rect 2340 -306 2346 -300
rect 2340 -312 2346 -306
rect 2340 -318 2346 -312
rect 2340 -324 2346 -318
rect 2340 -330 2346 -324
rect 2340 -336 2346 -330
rect 2340 -342 2346 -336
rect 2340 -348 2346 -342
rect 2340 -354 2346 -348
rect 2340 -360 2346 -354
rect 2340 -366 2346 -360
rect 2340 -372 2346 -366
rect 2340 -378 2346 -372
rect 2340 -384 2346 -378
rect 2340 -390 2346 -384
rect 2340 -396 2346 -390
rect 2340 -402 2346 -396
rect 2340 -408 2346 -402
rect 2340 -414 2346 -408
rect 2340 -420 2346 -414
rect 2340 -426 2346 -420
rect 2340 -432 2346 -426
rect 2340 -438 2346 -432
rect 2340 -444 2346 -438
rect 2340 -450 2346 -444
rect 2340 -456 2346 -450
rect 2340 -462 2346 -456
rect 2340 -468 2346 -462
rect 2340 -474 2346 -468
rect 2340 -480 2346 -474
rect 2340 -486 2346 -480
rect 2340 -492 2346 -486
rect 2340 -498 2346 -492
rect 2340 -504 2346 -498
rect 2340 -510 2346 -504
rect 2340 -516 2346 -510
rect 2340 -522 2346 -516
rect 2340 -528 2346 -522
rect 2340 -534 2346 -528
rect 2340 -540 2346 -534
rect 2340 -546 2346 -540
rect 2340 -552 2346 -546
rect 2340 -558 2346 -552
rect 2340 -564 2346 -558
rect 2340 -570 2346 -564
rect 2340 -576 2346 -570
rect 2340 -582 2346 -576
rect 2340 -588 2346 -582
rect 2340 -594 2346 -588
rect 2340 -600 2346 -594
rect 2340 -606 2346 -600
rect 2340 -612 2346 -606
rect 2340 -618 2346 -612
rect 2340 -624 2346 -618
rect 2340 -630 2346 -624
rect 2340 -636 2346 -630
rect 2340 -642 2346 -636
rect 2340 -648 2346 -642
rect 2340 -654 2346 -648
rect 2340 -660 2346 -654
rect 2340 -666 2346 -660
rect 2340 -672 2346 -666
rect 2340 -678 2346 -672
rect 2340 -684 2346 -678
rect 2340 -690 2346 -684
rect 2340 -696 2346 -690
rect 2340 -702 2346 -696
rect 2340 -708 2346 -702
rect 2340 -714 2346 -708
rect 2340 -720 2346 -714
rect 2340 -726 2346 -720
rect 2340 -732 2346 -726
rect 2340 -738 2346 -732
rect 2340 -744 2346 -738
rect 2340 -750 2346 -744
rect 2340 -756 2346 -750
rect 2340 -762 2346 -756
rect 2340 -768 2346 -762
rect 2340 -774 2346 -768
rect 2340 -780 2346 -774
rect 2340 -786 2346 -780
rect 2340 -792 2346 -786
rect 2340 -798 2346 -792
rect 2340 -804 2346 -798
rect 2340 -810 2346 -804
rect 2340 -816 2346 -810
rect 2340 -822 2346 -816
rect 2340 -828 2346 -822
rect 2340 -834 2346 -828
rect 2340 -840 2346 -834
rect 2340 -846 2346 -840
rect 2340 -852 2346 -846
rect 2340 -858 2346 -852
rect 2340 -864 2346 -858
rect 2340 -870 2346 -864
rect 2340 -876 2346 -870
rect 2340 -882 2346 -876
rect 2340 -1434 2346 -1428
rect 2340 -1440 2346 -1434
rect 2340 -1446 2346 -1440
rect 2340 -1452 2346 -1446
rect 2340 -1458 2346 -1452
rect 2340 -1464 2346 -1458
rect 2340 -1470 2346 -1464
rect 2340 -1476 2346 -1470
rect 2340 -1482 2346 -1476
rect 2340 -1488 2346 -1482
rect 2340 -1494 2346 -1488
rect 2340 -1500 2346 -1494
rect 2340 -1506 2346 -1500
rect 2340 -1512 2346 -1506
rect 2340 -1518 2346 -1512
rect 2340 -1524 2346 -1518
rect 2340 -1530 2346 -1524
rect 2340 -1536 2346 -1530
rect 2340 -1542 2346 -1536
rect 2340 -1548 2346 -1542
rect 2340 -1554 2346 -1548
rect 2340 -1560 2346 -1554
rect 2340 -1566 2346 -1560
rect 2340 -1572 2346 -1566
rect 2340 -1578 2346 -1572
rect 2340 -1584 2346 -1578
rect 2340 -1590 2346 -1584
rect 2340 -1596 2346 -1590
rect 2340 -1602 2346 -1596
rect 2340 -1608 2346 -1602
rect 2340 -1614 2346 -1608
rect 2340 -1620 2346 -1614
rect 2340 -1626 2346 -1620
rect 2340 -1632 2346 -1626
rect 2340 -1638 2346 -1632
rect 2340 -1644 2346 -1638
rect 2340 -1650 2346 -1644
rect 2340 -1656 2346 -1650
rect 2340 -1662 2346 -1656
rect 2340 -1668 2346 -1662
rect 2340 -1674 2346 -1668
rect 2340 -1680 2346 -1674
rect 2340 -1686 2346 -1680
rect 2340 -1692 2346 -1686
rect 2340 -1698 2346 -1692
rect 2340 -1704 2346 -1698
rect 2340 -1710 2346 -1704
rect 2340 -1716 2346 -1710
rect 2340 -1722 2346 -1716
rect 2340 -1728 2346 -1722
rect 2340 -1734 2346 -1728
rect 2340 -1740 2346 -1734
rect 2340 -1746 2346 -1740
rect 2340 -1752 2346 -1746
rect 2340 -1758 2346 -1752
rect 2340 -1764 2346 -1758
rect 2340 -1770 2346 -1764
rect 2340 -1776 2346 -1770
rect 2340 -1782 2346 -1776
rect 2340 -1788 2346 -1782
rect 2340 -1794 2346 -1788
rect 2340 -1800 2346 -1794
rect 2340 -1806 2346 -1800
rect 2340 -1812 2346 -1806
rect 2340 -1818 2346 -1812
rect 2340 -1824 2346 -1818
rect 2340 -1830 2346 -1824
rect 2340 -1836 2346 -1830
rect 2340 -1842 2346 -1836
rect 2340 -1848 2346 -1842
rect 2340 -1854 2346 -1848
rect 2340 -1860 2346 -1854
rect 2340 -1866 2346 -1860
rect 2340 -1872 2346 -1866
rect 2340 -1878 2346 -1872
rect 2340 -1884 2346 -1878
rect 2340 -1890 2346 -1884
rect 2340 -1896 2346 -1890
rect 2340 -1902 2346 -1896
rect 2340 -1908 2346 -1902
rect 2340 -1914 2346 -1908
rect 2340 -1920 2346 -1914
rect 2340 -1926 2346 -1920
rect 2340 -1932 2346 -1926
rect 2340 -1938 2346 -1932
rect 2340 -1944 2346 -1938
rect 2340 -1950 2346 -1944
rect 2340 -1956 2346 -1950
rect 2340 -1962 2346 -1956
rect 2340 -1968 2346 -1962
rect 2340 -1974 2346 -1968
rect 2340 -1980 2346 -1974
rect 2340 -1986 2346 -1980
rect 2340 -1992 2346 -1986
rect 2340 -1998 2346 -1992
rect 2340 -2004 2346 -1998
rect 2340 -2010 2346 -2004
rect 2340 -2016 2346 -2010
rect 2340 -2022 2346 -2016
rect 2340 -2028 2346 -2022
rect 2340 -2034 2346 -2028
rect 2340 -2040 2346 -2034
rect 2340 -2046 2346 -2040
rect 2340 -2052 2346 -2046
rect 2340 -2058 2346 -2052
rect 2340 -2064 2346 -2058
rect 2340 -2070 2346 -2064
rect 2340 -2076 2346 -2070
rect 2340 -2082 2346 -2076
rect 2340 -2088 2346 -2082
rect 2340 -2094 2346 -2088
rect 2340 -2100 2346 -2094
rect 2340 -2106 2346 -2100
rect 2340 -2112 2346 -2106
rect 2340 -2118 2346 -2112
rect 2340 -2124 2346 -2118
rect 2340 -2130 2346 -2124
rect 2340 -2136 2346 -2130
rect 2340 -2142 2346 -2136
rect 2340 -2148 2346 -2142
rect 2340 -2154 2346 -2148
rect 2340 -2160 2346 -2154
rect 2340 -2166 2346 -2160
rect 2340 -2172 2346 -2166
rect 2340 -2250 2346 -2244
rect 2340 -2256 2346 -2250
rect 2340 -2262 2346 -2256
rect 2340 -2268 2346 -2262
rect 2340 -2274 2346 -2268
rect 2340 -2280 2346 -2274
rect 2340 -2286 2346 -2280
rect 2340 -2292 2346 -2286
rect 2340 -2298 2346 -2292
rect 2340 -2304 2346 -2298
rect 2340 -2310 2346 -2304
rect 2340 -2316 2346 -2310
rect 2340 -2322 2346 -2316
rect 2340 -2328 2346 -2322
rect 2340 -2334 2346 -2328
rect 2340 -2340 2346 -2334
rect 2340 -2346 2346 -2340
rect 2340 -2352 2346 -2346
rect 2340 -2358 2346 -2352
rect 2340 -2364 2346 -2358
rect 2340 -2370 2346 -2364
rect 2340 -2376 2346 -2370
rect 2340 -2382 2346 -2376
rect 2340 -2388 2346 -2382
rect 2340 -2394 2346 -2388
rect 2340 -2400 2346 -2394
rect 2340 -2406 2346 -2400
rect 2340 -2412 2346 -2406
rect 2340 -2418 2346 -2412
rect 2340 -2424 2346 -2418
rect 2340 -2430 2346 -2424
rect 2340 -2496 2346 -2490
rect 2340 -2502 2346 -2496
rect 2340 -2508 2346 -2502
rect 2340 -2514 2346 -2508
rect 2340 -2520 2346 -2514
rect 2340 -2526 2346 -2520
rect 2340 -2532 2346 -2526
rect 2340 -2538 2346 -2532
rect 2340 -2544 2346 -2538
rect 2340 -2550 2346 -2544
rect 2340 -2556 2346 -2550
rect 2340 -2562 2346 -2556
rect 2340 -2568 2346 -2562
rect 2340 -2574 2346 -2568
rect 2340 -2580 2346 -2574
rect 2340 -2586 2346 -2580
rect 2340 -2592 2346 -2586
rect 2340 -2598 2346 -2592
rect 2340 -2604 2346 -2598
rect 2340 -2610 2346 -2604
rect 2340 -2616 2346 -2610
rect 2340 -2622 2346 -2616
rect 2340 -2628 2346 -2622
rect 2340 -2634 2346 -2628
rect 2340 -2640 2346 -2634
rect 2340 -2646 2346 -2640
rect 2340 -2652 2346 -2646
rect 2340 -2658 2346 -2652
rect 2340 -2664 2346 -2658
rect 2340 -2670 2346 -2664
rect 2340 -2676 2346 -2670
rect 2340 -2682 2346 -2676
rect 2340 -2688 2346 -2682
rect 2340 -2694 2346 -2688
rect 2340 -2700 2346 -2694
rect 2340 -2706 2346 -2700
rect 2340 -2712 2346 -2706
rect 2340 -2718 2346 -2712
rect 2340 -2724 2346 -2718
rect 2340 -2730 2346 -2724
rect 2340 -2736 2346 -2730
rect 2340 -2742 2346 -2736
rect 2340 -2748 2346 -2742
rect 2340 -2754 2346 -2748
rect 2340 -2760 2346 -2754
rect 2340 -2766 2346 -2760
rect 2340 -2772 2346 -2766
rect 2340 -2778 2346 -2772
rect 2340 -2784 2346 -2778
rect 2340 -2790 2346 -2784
rect 2340 -2796 2346 -2790
rect 2340 -2802 2346 -2796
rect 2340 -2808 2346 -2802
rect 2340 -2814 2346 -2808
rect 2340 -2820 2346 -2814
rect 2340 -2826 2346 -2820
rect 2340 -2832 2346 -2826
rect 2340 -2838 2346 -2832
rect 2340 -2844 2346 -2838
rect 2340 -2850 2346 -2844
rect 2340 -2856 2346 -2850
rect 2340 -2862 2346 -2856
rect 2340 -2868 2346 -2862
rect 2340 -2874 2346 -2868
rect 2340 -2880 2346 -2874
rect 2340 -2886 2346 -2880
rect 2340 -2892 2346 -2886
rect 2340 -2898 2346 -2892
rect 2340 -2904 2346 -2898
rect 2340 -2910 2346 -2904
rect 2340 -2916 2346 -2910
rect 2340 -2922 2346 -2916
rect 2346 -18 2352 -12
rect 2346 -24 2352 -18
rect 2346 -30 2352 -24
rect 2346 -36 2352 -30
rect 2346 -42 2352 -36
rect 2346 -48 2352 -42
rect 2346 -54 2352 -48
rect 2346 -60 2352 -54
rect 2346 -66 2352 -60
rect 2346 -72 2352 -66
rect 2346 -78 2352 -72
rect 2346 -84 2352 -78
rect 2346 -90 2352 -84
rect 2346 -96 2352 -90
rect 2346 -102 2352 -96
rect 2346 -108 2352 -102
rect 2346 -114 2352 -108
rect 2346 -120 2352 -114
rect 2346 -126 2352 -120
rect 2346 -132 2352 -126
rect 2346 -138 2352 -132
rect 2346 -144 2352 -138
rect 2346 -150 2352 -144
rect 2346 -156 2352 -150
rect 2346 -162 2352 -156
rect 2346 -168 2352 -162
rect 2346 -174 2352 -168
rect 2346 -180 2352 -174
rect 2346 -186 2352 -180
rect 2346 -192 2352 -186
rect 2346 -198 2352 -192
rect 2346 -204 2352 -198
rect 2346 -210 2352 -204
rect 2346 -216 2352 -210
rect 2346 -222 2352 -216
rect 2346 -228 2352 -222
rect 2346 -234 2352 -228
rect 2346 -240 2352 -234
rect 2346 -246 2352 -240
rect 2346 -252 2352 -246
rect 2346 -258 2352 -252
rect 2346 -264 2352 -258
rect 2346 -270 2352 -264
rect 2346 -276 2352 -270
rect 2346 -282 2352 -276
rect 2346 -288 2352 -282
rect 2346 -294 2352 -288
rect 2346 -300 2352 -294
rect 2346 -306 2352 -300
rect 2346 -312 2352 -306
rect 2346 -318 2352 -312
rect 2346 -324 2352 -318
rect 2346 -330 2352 -324
rect 2346 -336 2352 -330
rect 2346 -342 2352 -336
rect 2346 -348 2352 -342
rect 2346 -354 2352 -348
rect 2346 -360 2352 -354
rect 2346 -366 2352 -360
rect 2346 -372 2352 -366
rect 2346 -378 2352 -372
rect 2346 -384 2352 -378
rect 2346 -390 2352 -384
rect 2346 -396 2352 -390
rect 2346 -402 2352 -396
rect 2346 -408 2352 -402
rect 2346 -414 2352 -408
rect 2346 -420 2352 -414
rect 2346 -426 2352 -420
rect 2346 -432 2352 -426
rect 2346 -438 2352 -432
rect 2346 -444 2352 -438
rect 2346 -450 2352 -444
rect 2346 -456 2352 -450
rect 2346 -462 2352 -456
rect 2346 -468 2352 -462
rect 2346 -474 2352 -468
rect 2346 -480 2352 -474
rect 2346 -486 2352 -480
rect 2346 -492 2352 -486
rect 2346 -498 2352 -492
rect 2346 -504 2352 -498
rect 2346 -510 2352 -504
rect 2346 -516 2352 -510
rect 2346 -522 2352 -516
rect 2346 -528 2352 -522
rect 2346 -534 2352 -528
rect 2346 -540 2352 -534
rect 2346 -546 2352 -540
rect 2346 -552 2352 -546
rect 2346 -558 2352 -552
rect 2346 -564 2352 -558
rect 2346 -570 2352 -564
rect 2346 -576 2352 -570
rect 2346 -582 2352 -576
rect 2346 -588 2352 -582
rect 2346 -594 2352 -588
rect 2346 -600 2352 -594
rect 2346 -606 2352 -600
rect 2346 -612 2352 -606
rect 2346 -618 2352 -612
rect 2346 -624 2352 -618
rect 2346 -630 2352 -624
rect 2346 -636 2352 -630
rect 2346 -642 2352 -636
rect 2346 -648 2352 -642
rect 2346 -654 2352 -648
rect 2346 -660 2352 -654
rect 2346 -666 2352 -660
rect 2346 -672 2352 -666
rect 2346 -678 2352 -672
rect 2346 -684 2352 -678
rect 2346 -690 2352 -684
rect 2346 -696 2352 -690
rect 2346 -702 2352 -696
rect 2346 -708 2352 -702
rect 2346 -714 2352 -708
rect 2346 -720 2352 -714
rect 2346 -726 2352 -720
rect 2346 -732 2352 -726
rect 2346 -738 2352 -732
rect 2346 -744 2352 -738
rect 2346 -750 2352 -744
rect 2346 -756 2352 -750
rect 2346 -762 2352 -756
rect 2346 -768 2352 -762
rect 2346 -774 2352 -768
rect 2346 -780 2352 -774
rect 2346 -786 2352 -780
rect 2346 -792 2352 -786
rect 2346 -798 2352 -792
rect 2346 -804 2352 -798
rect 2346 -810 2352 -804
rect 2346 -816 2352 -810
rect 2346 -822 2352 -816
rect 2346 -828 2352 -822
rect 2346 -834 2352 -828
rect 2346 -840 2352 -834
rect 2346 -846 2352 -840
rect 2346 -852 2352 -846
rect 2346 -858 2352 -852
rect 2346 -864 2352 -858
rect 2346 -1428 2352 -1422
rect 2346 -1434 2352 -1428
rect 2346 -1440 2352 -1434
rect 2346 -1446 2352 -1440
rect 2346 -1452 2352 -1446
rect 2346 -1458 2352 -1452
rect 2346 -1464 2352 -1458
rect 2346 -1470 2352 -1464
rect 2346 -1476 2352 -1470
rect 2346 -1482 2352 -1476
rect 2346 -1488 2352 -1482
rect 2346 -1494 2352 -1488
rect 2346 -1500 2352 -1494
rect 2346 -1506 2352 -1500
rect 2346 -1512 2352 -1506
rect 2346 -1518 2352 -1512
rect 2346 -1524 2352 -1518
rect 2346 -1530 2352 -1524
rect 2346 -1536 2352 -1530
rect 2346 -1542 2352 -1536
rect 2346 -1548 2352 -1542
rect 2346 -1554 2352 -1548
rect 2346 -1560 2352 -1554
rect 2346 -1566 2352 -1560
rect 2346 -1572 2352 -1566
rect 2346 -1578 2352 -1572
rect 2346 -1584 2352 -1578
rect 2346 -1590 2352 -1584
rect 2346 -1596 2352 -1590
rect 2346 -1602 2352 -1596
rect 2346 -1608 2352 -1602
rect 2346 -1614 2352 -1608
rect 2346 -1620 2352 -1614
rect 2346 -1626 2352 -1620
rect 2346 -1632 2352 -1626
rect 2346 -1638 2352 -1632
rect 2346 -1644 2352 -1638
rect 2346 -1650 2352 -1644
rect 2346 -1656 2352 -1650
rect 2346 -1662 2352 -1656
rect 2346 -1668 2352 -1662
rect 2346 -1674 2352 -1668
rect 2346 -1680 2352 -1674
rect 2346 -1686 2352 -1680
rect 2346 -1692 2352 -1686
rect 2346 -1698 2352 -1692
rect 2346 -1704 2352 -1698
rect 2346 -1710 2352 -1704
rect 2346 -1716 2352 -1710
rect 2346 -1722 2352 -1716
rect 2346 -1728 2352 -1722
rect 2346 -1734 2352 -1728
rect 2346 -1740 2352 -1734
rect 2346 -1746 2352 -1740
rect 2346 -1752 2352 -1746
rect 2346 -1758 2352 -1752
rect 2346 -1764 2352 -1758
rect 2346 -1770 2352 -1764
rect 2346 -1776 2352 -1770
rect 2346 -1782 2352 -1776
rect 2346 -1788 2352 -1782
rect 2346 -1794 2352 -1788
rect 2346 -1800 2352 -1794
rect 2346 -1806 2352 -1800
rect 2346 -1812 2352 -1806
rect 2346 -1818 2352 -1812
rect 2346 -1824 2352 -1818
rect 2346 -1830 2352 -1824
rect 2346 -1836 2352 -1830
rect 2346 -1842 2352 -1836
rect 2346 -1848 2352 -1842
rect 2346 -1854 2352 -1848
rect 2346 -1860 2352 -1854
rect 2346 -1866 2352 -1860
rect 2346 -1872 2352 -1866
rect 2346 -1878 2352 -1872
rect 2346 -1884 2352 -1878
rect 2346 -1890 2352 -1884
rect 2346 -1896 2352 -1890
rect 2346 -1902 2352 -1896
rect 2346 -1908 2352 -1902
rect 2346 -1914 2352 -1908
rect 2346 -1920 2352 -1914
rect 2346 -1926 2352 -1920
rect 2346 -1932 2352 -1926
rect 2346 -1938 2352 -1932
rect 2346 -1944 2352 -1938
rect 2346 -1950 2352 -1944
rect 2346 -1956 2352 -1950
rect 2346 -1962 2352 -1956
rect 2346 -1968 2352 -1962
rect 2346 -1974 2352 -1968
rect 2346 -1980 2352 -1974
rect 2346 -1986 2352 -1980
rect 2346 -1992 2352 -1986
rect 2346 -1998 2352 -1992
rect 2346 -2004 2352 -1998
rect 2346 -2010 2352 -2004
rect 2346 -2016 2352 -2010
rect 2346 -2022 2352 -2016
rect 2346 -2028 2352 -2022
rect 2346 -2034 2352 -2028
rect 2346 -2040 2352 -2034
rect 2346 -2046 2352 -2040
rect 2346 -2052 2352 -2046
rect 2346 -2058 2352 -2052
rect 2346 -2064 2352 -2058
rect 2346 -2070 2352 -2064
rect 2346 -2076 2352 -2070
rect 2346 -2082 2352 -2076
rect 2346 -2088 2352 -2082
rect 2346 -2094 2352 -2088
rect 2346 -2100 2352 -2094
rect 2346 -2106 2352 -2100
rect 2346 -2112 2352 -2106
rect 2346 -2118 2352 -2112
rect 2346 -2124 2352 -2118
rect 2346 -2130 2352 -2124
rect 2346 -2136 2352 -2130
rect 2346 -2142 2352 -2136
rect 2346 -2148 2352 -2142
rect 2346 -2154 2352 -2148
rect 2346 -2160 2352 -2154
rect 2346 -2166 2352 -2160
rect 2346 -2238 2352 -2232
rect 2346 -2244 2352 -2238
rect 2346 -2250 2352 -2244
rect 2346 -2256 2352 -2250
rect 2346 -2262 2352 -2256
rect 2346 -2268 2352 -2262
rect 2346 -2274 2352 -2268
rect 2346 -2280 2352 -2274
rect 2346 -2286 2352 -2280
rect 2346 -2292 2352 -2286
rect 2346 -2298 2352 -2292
rect 2346 -2304 2352 -2298
rect 2346 -2310 2352 -2304
rect 2346 -2316 2352 -2310
rect 2346 -2322 2352 -2316
rect 2346 -2328 2352 -2322
rect 2346 -2334 2352 -2328
rect 2346 -2340 2352 -2334
rect 2346 -2346 2352 -2340
rect 2346 -2352 2352 -2346
rect 2346 -2358 2352 -2352
rect 2346 -2364 2352 -2358
rect 2346 -2370 2352 -2364
rect 2346 -2376 2352 -2370
rect 2346 -2382 2352 -2376
rect 2346 -2388 2352 -2382
rect 2346 -2394 2352 -2388
rect 2346 -2400 2352 -2394
rect 2346 -2406 2352 -2400
rect 2346 -2412 2352 -2406
rect 2346 -2418 2352 -2412
rect 2346 -2424 2352 -2418
rect 2346 -2496 2352 -2490
rect 2346 -2502 2352 -2496
rect 2346 -2508 2352 -2502
rect 2346 -2514 2352 -2508
rect 2346 -2520 2352 -2514
rect 2346 -2526 2352 -2520
rect 2346 -2532 2352 -2526
rect 2346 -2538 2352 -2532
rect 2346 -2544 2352 -2538
rect 2346 -2550 2352 -2544
rect 2346 -2556 2352 -2550
rect 2346 -2562 2352 -2556
rect 2346 -2568 2352 -2562
rect 2346 -2574 2352 -2568
rect 2346 -2580 2352 -2574
rect 2346 -2586 2352 -2580
rect 2346 -2592 2352 -2586
rect 2346 -2598 2352 -2592
rect 2346 -2604 2352 -2598
rect 2346 -2610 2352 -2604
rect 2346 -2616 2352 -2610
rect 2346 -2622 2352 -2616
rect 2346 -2628 2352 -2622
rect 2346 -2634 2352 -2628
rect 2346 -2640 2352 -2634
rect 2346 -2646 2352 -2640
rect 2346 -2652 2352 -2646
rect 2346 -2658 2352 -2652
rect 2346 -2664 2352 -2658
rect 2346 -2670 2352 -2664
rect 2346 -2676 2352 -2670
rect 2346 -2682 2352 -2676
rect 2346 -2688 2352 -2682
rect 2346 -2694 2352 -2688
rect 2346 -2700 2352 -2694
rect 2346 -2706 2352 -2700
rect 2346 -2712 2352 -2706
rect 2346 -2718 2352 -2712
rect 2346 -2724 2352 -2718
rect 2346 -2730 2352 -2724
rect 2346 -2736 2352 -2730
rect 2346 -2742 2352 -2736
rect 2346 -2748 2352 -2742
rect 2346 -2754 2352 -2748
rect 2346 -2760 2352 -2754
rect 2346 -2766 2352 -2760
rect 2346 -2772 2352 -2766
rect 2346 -2778 2352 -2772
rect 2346 -2784 2352 -2778
rect 2346 -2790 2352 -2784
rect 2346 -2796 2352 -2790
rect 2346 -2802 2352 -2796
rect 2346 -2808 2352 -2802
rect 2346 -2814 2352 -2808
rect 2346 -2820 2352 -2814
rect 2346 -2826 2352 -2820
rect 2346 -2832 2352 -2826
rect 2346 -2838 2352 -2832
rect 2346 -2844 2352 -2838
rect 2346 -2850 2352 -2844
rect 2346 -2856 2352 -2850
rect 2346 -2862 2352 -2856
rect 2346 -2868 2352 -2862
rect 2346 -2874 2352 -2868
rect 2346 -2880 2352 -2874
rect 2346 -2886 2352 -2880
rect 2346 -2892 2352 -2886
rect 2346 -2898 2352 -2892
rect 2346 -2904 2352 -2898
rect 2346 -2910 2352 -2904
rect 2346 -2916 2352 -2910
rect 2352 -12 2358 -6
rect 2352 -18 2358 -12
rect 2352 -24 2358 -18
rect 2352 -30 2358 -24
rect 2352 -36 2358 -30
rect 2352 -42 2358 -36
rect 2352 -48 2358 -42
rect 2352 -54 2358 -48
rect 2352 -60 2358 -54
rect 2352 -66 2358 -60
rect 2352 -72 2358 -66
rect 2352 -78 2358 -72
rect 2352 -84 2358 -78
rect 2352 -90 2358 -84
rect 2352 -96 2358 -90
rect 2352 -102 2358 -96
rect 2352 -108 2358 -102
rect 2352 -114 2358 -108
rect 2352 -120 2358 -114
rect 2352 -126 2358 -120
rect 2352 -132 2358 -126
rect 2352 -138 2358 -132
rect 2352 -144 2358 -138
rect 2352 -150 2358 -144
rect 2352 -156 2358 -150
rect 2352 -162 2358 -156
rect 2352 -168 2358 -162
rect 2352 -174 2358 -168
rect 2352 -180 2358 -174
rect 2352 -186 2358 -180
rect 2352 -192 2358 -186
rect 2352 -198 2358 -192
rect 2352 -204 2358 -198
rect 2352 -210 2358 -204
rect 2352 -216 2358 -210
rect 2352 -222 2358 -216
rect 2352 -228 2358 -222
rect 2352 -234 2358 -228
rect 2352 -240 2358 -234
rect 2352 -246 2358 -240
rect 2352 -252 2358 -246
rect 2352 -258 2358 -252
rect 2352 -264 2358 -258
rect 2352 -270 2358 -264
rect 2352 -276 2358 -270
rect 2352 -282 2358 -276
rect 2352 -288 2358 -282
rect 2352 -294 2358 -288
rect 2352 -300 2358 -294
rect 2352 -306 2358 -300
rect 2352 -312 2358 -306
rect 2352 -318 2358 -312
rect 2352 -324 2358 -318
rect 2352 -330 2358 -324
rect 2352 -336 2358 -330
rect 2352 -342 2358 -336
rect 2352 -348 2358 -342
rect 2352 -354 2358 -348
rect 2352 -360 2358 -354
rect 2352 -366 2358 -360
rect 2352 -372 2358 -366
rect 2352 -378 2358 -372
rect 2352 -384 2358 -378
rect 2352 -390 2358 -384
rect 2352 -396 2358 -390
rect 2352 -402 2358 -396
rect 2352 -408 2358 -402
rect 2352 -414 2358 -408
rect 2352 -420 2358 -414
rect 2352 -426 2358 -420
rect 2352 -432 2358 -426
rect 2352 -438 2358 -432
rect 2352 -444 2358 -438
rect 2352 -450 2358 -444
rect 2352 -456 2358 -450
rect 2352 -462 2358 -456
rect 2352 -468 2358 -462
rect 2352 -474 2358 -468
rect 2352 -480 2358 -474
rect 2352 -486 2358 -480
rect 2352 -492 2358 -486
rect 2352 -498 2358 -492
rect 2352 -504 2358 -498
rect 2352 -510 2358 -504
rect 2352 -516 2358 -510
rect 2352 -522 2358 -516
rect 2352 -528 2358 -522
rect 2352 -534 2358 -528
rect 2352 -540 2358 -534
rect 2352 -546 2358 -540
rect 2352 -552 2358 -546
rect 2352 -558 2358 -552
rect 2352 -564 2358 -558
rect 2352 -570 2358 -564
rect 2352 -576 2358 -570
rect 2352 -582 2358 -576
rect 2352 -588 2358 -582
rect 2352 -594 2358 -588
rect 2352 -600 2358 -594
rect 2352 -606 2358 -600
rect 2352 -612 2358 -606
rect 2352 -618 2358 -612
rect 2352 -624 2358 -618
rect 2352 -630 2358 -624
rect 2352 -636 2358 -630
rect 2352 -642 2358 -636
rect 2352 -648 2358 -642
rect 2352 -654 2358 -648
rect 2352 -660 2358 -654
rect 2352 -666 2358 -660
rect 2352 -672 2358 -666
rect 2352 -678 2358 -672
rect 2352 -684 2358 -678
rect 2352 -690 2358 -684
rect 2352 -696 2358 -690
rect 2352 -702 2358 -696
rect 2352 -708 2358 -702
rect 2352 -714 2358 -708
rect 2352 -720 2358 -714
rect 2352 -726 2358 -720
rect 2352 -732 2358 -726
rect 2352 -738 2358 -732
rect 2352 -744 2358 -738
rect 2352 -750 2358 -744
rect 2352 -756 2358 -750
rect 2352 -762 2358 -756
rect 2352 -768 2358 -762
rect 2352 -774 2358 -768
rect 2352 -780 2358 -774
rect 2352 -786 2358 -780
rect 2352 -792 2358 -786
rect 2352 -798 2358 -792
rect 2352 -804 2358 -798
rect 2352 -810 2358 -804
rect 2352 -816 2358 -810
rect 2352 -822 2358 -816
rect 2352 -828 2358 -822
rect 2352 -834 2358 -828
rect 2352 -840 2358 -834
rect 2352 -846 2358 -840
rect 2352 -1428 2358 -1422
rect 2352 -1434 2358 -1428
rect 2352 -1440 2358 -1434
rect 2352 -1446 2358 -1440
rect 2352 -1452 2358 -1446
rect 2352 -1458 2358 -1452
rect 2352 -1464 2358 -1458
rect 2352 -1470 2358 -1464
rect 2352 -1476 2358 -1470
rect 2352 -1482 2358 -1476
rect 2352 -1488 2358 -1482
rect 2352 -1494 2358 -1488
rect 2352 -1500 2358 -1494
rect 2352 -1506 2358 -1500
rect 2352 -1512 2358 -1506
rect 2352 -1518 2358 -1512
rect 2352 -1524 2358 -1518
rect 2352 -1530 2358 -1524
rect 2352 -1536 2358 -1530
rect 2352 -1542 2358 -1536
rect 2352 -1548 2358 -1542
rect 2352 -1554 2358 -1548
rect 2352 -1560 2358 -1554
rect 2352 -1566 2358 -1560
rect 2352 -1572 2358 -1566
rect 2352 -1578 2358 -1572
rect 2352 -1584 2358 -1578
rect 2352 -1590 2358 -1584
rect 2352 -1596 2358 -1590
rect 2352 -1602 2358 -1596
rect 2352 -1608 2358 -1602
rect 2352 -1614 2358 -1608
rect 2352 -1620 2358 -1614
rect 2352 -1626 2358 -1620
rect 2352 -1632 2358 -1626
rect 2352 -1638 2358 -1632
rect 2352 -1644 2358 -1638
rect 2352 -1650 2358 -1644
rect 2352 -1656 2358 -1650
rect 2352 -1662 2358 -1656
rect 2352 -1668 2358 -1662
rect 2352 -1674 2358 -1668
rect 2352 -1680 2358 -1674
rect 2352 -1686 2358 -1680
rect 2352 -1692 2358 -1686
rect 2352 -1698 2358 -1692
rect 2352 -1704 2358 -1698
rect 2352 -1710 2358 -1704
rect 2352 -1716 2358 -1710
rect 2352 -1722 2358 -1716
rect 2352 -1728 2358 -1722
rect 2352 -1734 2358 -1728
rect 2352 -1740 2358 -1734
rect 2352 -1746 2358 -1740
rect 2352 -1752 2358 -1746
rect 2352 -1758 2358 -1752
rect 2352 -1764 2358 -1758
rect 2352 -1770 2358 -1764
rect 2352 -1776 2358 -1770
rect 2352 -1782 2358 -1776
rect 2352 -1788 2358 -1782
rect 2352 -1794 2358 -1788
rect 2352 -1800 2358 -1794
rect 2352 -1806 2358 -1800
rect 2352 -1812 2358 -1806
rect 2352 -1818 2358 -1812
rect 2352 -1824 2358 -1818
rect 2352 -1830 2358 -1824
rect 2352 -1836 2358 -1830
rect 2352 -1842 2358 -1836
rect 2352 -1848 2358 -1842
rect 2352 -1854 2358 -1848
rect 2352 -1860 2358 -1854
rect 2352 -1866 2358 -1860
rect 2352 -1872 2358 -1866
rect 2352 -1878 2358 -1872
rect 2352 -1884 2358 -1878
rect 2352 -1890 2358 -1884
rect 2352 -1896 2358 -1890
rect 2352 -1902 2358 -1896
rect 2352 -1908 2358 -1902
rect 2352 -1914 2358 -1908
rect 2352 -1920 2358 -1914
rect 2352 -1926 2358 -1920
rect 2352 -1932 2358 -1926
rect 2352 -1938 2358 -1932
rect 2352 -1944 2358 -1938
rect 2352 -1950 2358 -1944
rect 2352 -1956 2358 -1950
rect 2352 -1962 2358 -1956
rect 2352 -1968 2358 -1962
rect 2352 -1974 2358 -1968
rect 2352 -1980 2358 -1974
rect 2352 -1986 2358 -1980
rect 2352 -1992 2358 -1986
rect 2352 -1998 2358 -1992
rect 2352 -2004 2358 -1998
rect 2352 -2010 2358 -2004
rect 2352 -2016 2358 -2010
rect 2352 -2022 2358 -2016
rect 2352 -2028 2358 -2022
rect 2352 -2034 2358 -2028
rect 2352 -2040 2358 -2034
rect 2352 -2046 2358 -2040
rect 2352 -2052 2358 -2046
rect 2352 -2058 2358 -2052
rect 2352 -2064 2358 -2058
rect 2352 -2070 2358 -2064
rect 2352 -2076 2358 -2070
rect 2352 -2082 2358 -2076
rect 2352 -2088 2358 -2082
rect 2352 -2094 2358 -2088
rect 2352 -2100 2358 -2094
rect 2352 -2106 2358 -2100
rect 2352 -2112 2358 -2106
rect 2352 -2118 2358 -2112
rect 2352 -2124 2358 -2118
rect 2352 -2130 2358 -2124
rect 2352 -2136 2358 -2130
rect 2352 -2142 2358 -2136
rect 2352 -2148 2358 -2142
rect 2352 -2154 2358 -2148
rect 2352 -2232 2358 -2226
rect 2352 -2238 2358 -2232
rect 2352 -2244 2358 -2238
rect 2352 -2250 2358 -2244
rect 2352 -2256 2358 -2250
rect 2352 -2262 2358 -2256
rect 2352 -2268 2358 -2262
rect 2352 -2274 2358 -2268
rect 2352 -2280 2358 -2274
rect 2352 -2286 2358 -2280
rect 2352 -2292 2358 -2286
rect 2352 -2298 2358 -2292
rect 2352 -2304 2358 -2298
rect 2352 -2310 2358 -2304
rect 2352 -2316 2358 -2310
rect 2352 -2322 2358 -2316
rect 2352 -2328 2358 -2322
rect 2352 -2334 2358 -2328
rect 2352 -2340 2358 -2334
rect 2352 -2346 2358 -2340
rect 2352 -2352 2358 -2346
rect 2352 -2358 2358 -2352
rect 2352 -2364 2358 -2358
rect 2352 -2370 2358 -2364
rect 2352 -2376 2358 -2370
rect 2352 -2382 2358 -2376
rect 2352 -2388 2358 -2382
rect 2352 -2394 2358 -2388
rect 2352 -2400 2358 -2394
rect 2352 -2406 2358 -2400
rect 2352 -2412 2358 -2406
rect 2352 -2418 2358 -2412
rect 2352 -2424 2358 -2418
rect 2352 -2490 2358 -2484
rect 2352 -2496 2358 -2490
rect 2352 -2502 2358 -2496
rect 2352 -2508 2358 -2502
rect 2352 -2514 2358 -2508
rect 2352 -2520 2358 -2514
rect 2352 -2526 2358 -2520
rect 2352 -2532 2358 -2526
rect 2352 -2538 2358 -2532
rect 2352 -2544 2358 -2538
rect 2352 -2550 2358 -2544
rect 2352 -2556 2358 -2550
rect 2352 -2562 2358 -2556
rect 2352 -2568 2358 -2562
rect 2352 -2574 2358 -2568
rect 2352 -2580 2358 -2574
rect 2352 -2586 2358 -2580
rect 2352 -2592 2358 -2586
rect 2352 -2598 2358 -2592
rect 2352 -2604 2358 -2598
rect 2352 -2610 2358 -2604
rect 2352 -2616 2358 -2610
rect 2352 -2622 2358 -2616
rect 2352 -2628 2358 -2622
rect 2352 -2634 2358 -2628
rect 2352 -2640 2358 -2634
rect 2352 -2646 2358 -2640
rect 2352 -2652 2358 -2646
rect 2352 -2658 2358 -2652
rect 2352 -2664 2358 -2658
rect 2352 -2670 2358 -2664
rect 2352 -2676 2358 -2670
rect 2352 -2682 2358 -2676
rect 2352 -2688 2358 -2682
rect 2352 -2694 2358 -2688
rect 2352 -2700 2358 -2694
rect 2352 -2706 2358 -2700
rect 2352 -2712 2358 -2706
rect 2352 -2718 2358 -2712
rect 2352 -2724 2358 -2718
rect 2352 -2730 2358 -2724
rect 2352 -2736 2358 -2730
rect 2352 -2742 2358 -2736
rect 2352 -2748 2358 -2742
rect 2352 -2754 2358 -2748
rect 2352 -2760 2358 -2754
rect 2352 -2766 2358 -2760
rect 2352 -2772 2358 -2766
rect 2352 -2778 2358 -2772
rect 2352 -2784 2358 -2778
rect 2352 -2790 2358 -2784
rect 2352 -2796 2358 -2790
rect 2352 -2802 2358 -2796
rect 2352 -2808 2358 -2802
rect 2352 -2814 2358 -2808
rect 2352 -2820 2358 -2814
rect 2352 -2826 2358 -2820
rect 2352 -2832 2358 -2826
rect 2352 -2838 2358 -2832
rect 2352 -2844 2358 -2838
rect 2352 -2850 2358 -2844
rect 2352 -2856 2358 -2850
rect 2352 -2862 2358 -2856
rect 2352 -2868 2358 -2862
rect 2352 -2874 2358 -2868
rect 2352 -2880 2358 -2874
rect 2352 -2886 2358 -2880
rect 2352 -2892 2358 -2886
rect 2352 -2898 2358 -2892
rect 2352 -2904 2358 -2898
rect 2352 -2910 2358 -2904
rect 2352 -2916 2358 -2910
rect 2358 -12 2364 -6
rect 2358 -18 2364 -12
rect 2358 -24 2364 -18
rect 2358 -30 2364 -24
rect 2358 -36 2364 -30
rect 2358 -42 2364 -36
rect 2358 -48 2364 -42
rect 2358 -54 2364 -48
rect 2358 -60 2364 -54
rect 2358 -66 2364 -60
rect 2358 -72 2364 -66
rect 2358 -78 2364 -72
rect 2358 -84 2364 -78
rect 2358 -90 2364 -84
rect 2358 -96 2364 -90
rect 2358 -102 2364 -96
rect 2358 -108 2364 -102
rect 2358 -114 2364 -108
rect 2358 -120 2364 -114
rect 2358 -126 2364 -120
rect 2358 -132 2364 -126
rect 2358 -138 2364 -132
rect 2358 -144 2364 -138
rect 2358 -150 2364 -144
rect 2358 -156 2364 -150
rect 2358 -162 2364 -156
rect 2358 -168 2364 -162
rect 2358 -174 2364 -168
rect 2358 -180 2364 -174
rect 2358 -186 2364 -180
rect 2358 -192 2364 -186
rect 2358 -198 2364 -192
rect 2358 -204 2364 -198
rect 2358 -210 2364 -204
rect 2358 -216 2364 -210
rect 2358 -222 2364 -216
rect 2358 -228 2364 -222
rect 2358 -234 2364 -228
rect 2358 -240 2364 -234
rect 2358 -246 2364 -240
rect 2358 -252 2364 -246
rect 2358 -258 2364 -252
rect 2358 -264 2364 -258
rect 2358 -270 2364 -264
rect 2358 -276 2364 -270
rect 2358 -282 2364 -276
rect 2358 -288 2364 -282
rect 2358 -294 2364 -288
rect 2358 -300 2364 -294
rect 2358 -306 2364 -300
rect 2358 -312 2364 -306
rect 2358 -318 2364 -312
rect 2358 -324 2364 -318
rect 2358 -330 2364 -324
rect 2358 -336 2364 -330
rect 2358 -342 2364 -336
rect 2358 -348 2364 -342
rect 2358 -354 2364 -348
rect 2358 -360 2364 -354
rect 2358 -366 2364 -360
rect 2358 -372 2364 -366
rect 2358 -378 2364 -372
rect 2358 -384 2364 -378
rect 2358 -390 2364 -384
rect 2358 -396 2364 -390
rect 2358 -402 2364 -396
rect 2358 -408 2364 -402
rect 2358 -414 2364 -408
rect 2358 -420 2364 -414
rect 2358 -426 2364 -420
rect 2358 -432 2364 -426
rect 2358 -438 2364 -432
rect 2358 -444 2364 -438
rect 2358 -450 2364 -444
rect 2358 -456 2364 -450
rect 2358 -462 2364 -456
rect 2358 -468 2364 -462
rect 2358 -474 2364 -468
rect 2358 -480 2364 -474
rect 2358 -486 2364 -480
rect 2358 -492 2364 -486
rect 2358 -498 2364 -492
rect 2358 -504 2364 -498
rect 2358 -510 2364 -504
rect 2358 -516 2364 -510
rect 2358 -522 2364 -516
rect 2358 -528 2364 -522
rect 2358 -534 2364 -528
rect 2358 -540 2364 -534
rect 2358 -546 2364 -540
rect 2358 -552 2364 -546
rect 2358 -558 2364 -552
rect 2358 -564 2364 -558
rect 2358 -570 2364 -564
rect 2358 -576 2364 -570
rect 2358 -582 2364 -576
rect 2358 -588 2364 -582
rect 2358 -594 2364 -588
rect 2358 -600 2364 -594
rect 2358 -606 2364 -600
rect 2358 -612 2364 -606
rect 2358 -618 2364 -612
rect 2358 -624 2364 -618
rect 2358 -630 2364 -624
rect 2358 -636 2364 -630
rect 2358 -642 2364 -636
rect 2358 -648 2364 -642
rect 2358 -654 2364 -648
rect 2358 -660 2364 -654
rect 2358 -666 2364 -660
rect 2358 -672 2364 -666
rect 2358 -678 2364 -672
rect 2358 -684 2364 -678
rect 2358 -690 2364 -684
rect 2358 -696 2364 -690
rect 2358 -702 2364 -696
rect 2358 -708 2364 -702
rect 2358 -714 2364 -708
rect 2358 -720 2364 -714
rect 2358 -726 2364 -720
rect 2358 -732 2364 -726
rect 2358 -738 2364 -732
rect 2358 -744 2364 -738
rect 2358 -750 2364 -744
rect 2358 -756 2364 -750
rect 2358 -762 2364 -756
rect 2358 -768 2364 -762
rect 2358 -774 2364 -768
rect 2358 -780 2364 -774
rect 2358 -786 2364 -780
rect 2358 -792 2364 -786
rect 2358 -798 2364 -792
rect 2358 -804 2364 -798
rect 2358 -810 2364 -804
rect 2358 -816 2364 -810
rect 2358 -822 2364 -816
rect 2358 -828 2364 -822
rect 2358 -1422 2364 -1416
rect 2358 -1428 2364 -1422
rect 2358 -1434 2364 -1428
rect 2358 -1440 2364 -1434
rect 2358 -1446 2364 -1440
rect 2358 -1452 2364 -1446
rect 2358 -1458 2364 -1452
rect 2358 -1464 2364 -1458
rect 2358 -1470 2364 -1464
rect 2358 -1476 2364 -1470
rect 2358 -1482 2364 -1476
rect 2358 -1488 2364 -1482
rect 2358 -1494 2364 -1488
rect 2358 -1500 2364 -1494
rect 2358 -1506 2364 -1500
rect 2358 -1512 2364 -1506
rect 2358 -1518 2364 -1512
rect 2358 -1524 2364 -1518
rect 2358 -1530 2364 -1524
rect 2358 -1536 2364 -1530
rect 2358 -1542 2364 -1536
rect 2358 -1548 2364 -1542
rect 2358 -1554 2364 -1548
rect 2358 -1560 2364 -1554
rect 2358 -1566 2364 -1560
rect 2358 -1572 2364 -1566
rect 2358 -1578 2364 -1572
rect 2358 -1584 2364 -1578
rect 2358 -1590 2364 -1584
rect 2358 -1596 2364 -1590
rect 2358 -1602 2364 -1596
rect 2358 -1608 2364 -1602
rect 2358 -1614 2364 -1608
rect 2358 -1620 2364 -1614
rect 2358 -1626 2364 -1620
rect 2358 -1632 2364 -1626
rect 2358 -1638 2364 -1632
rect 2358 -1644 2364 -1638
rect 2358 -1650 2364 -1644
rect 2358 -1656 2364 -1650
rect 2358 -1662 2364 -1656
rect 2358 -1668 2364 -1662
rect 2358 -1674 2364 -1668
rect 2358 -1680 2364 -1674
rect 2358 -1686 2364 -1680
rect 2358 -1692 2364 -1686
rect 2358 -1698 2364 -1692
rect 2358 -1704 2364 -1698
rect 2358 -1710 2364 -1704
rect 2358 -1716 2364 -1710
rect 2358 -1722 2364 -1716
rect 2358 -1728 2364 -1722
rect 2358 -1734 2364 -1728
rect 2358 -1740 2364 -1734
rect 2358 -1746 2364 -1740
rect 2358 -1752 2364 -1746
rect 2358 -1758 2364 -1752
rect 2358 -1764 2364 -1758
rect 2358 -1770 2364 -1764
rect 2358 -1776 2364 -1770
rect 2358 -1782 2364 -1776
rect 2358 -1788 2364 -1782
rect 2358 -1794 2364 -1788
rect 2358 -1800 2364 -1794
rect 2358 -1806 2364 -1800
rect 2358 -1812 2364 -1806
rect 2358 -1818 2364 -1812
rect 2358 -1824 2364 -1818
rect 2358 -1830 2364 -1824
rect 2358 -1836 2364 -1830
rect 2358 -1842 2364 -1836
rect 2358 -1848 2364 -1842
rect 2358 -1854 2364 -1848
rect 2358 -1860 2364 -1854
rect 2358 -1866 2364 -1860
rect 2358 -1872 2364 -1866
rect 2358 -1878 2364 -1872
rect 2358 -1884 2364 -1878
rect 2358 -1890 2364 -1884
rect 2358 -1896 2364 -1890
rect 2358 -1902 2364 -1896
rect 2358 -1908 2364 -1902
rect 2358 -1914 2364 -1908
rect 2358 -1920 2364 -1914
rect 2358 -1926 2364 -1920
rect 2358 -1932 2364 -1926
rect 2358 -1938 2364 -1932
rect 2358 -1944 2364 -1938
rect 2358 -1950 2364 -1944
rect 2358 -1956 2364 -1950
rect 2358 -1962 2364 -1956
rect 2358 -1968 2364 -1962
rect 2358 -1974 2364 -1968
rect 2358 -1980 2364 -1974
rect 2358 -1986 2364 -1980
rect 2358 -1992 2364 -1986
rect 2358 -1998 2364 -1992
rect 2358 -2004 2364 -1998
rect 2358 -2010 2364 -2004
rect 2358 -2016 2364 -2010
rect 2358 -2022 2364 -2016
rect 2358 -2028 2364 -2022
rect 2358 -2034 2364 -2028
rect 2358 -2040 2364 -2034
rect 2358 -2046 2364 -2040
rect 2358 -2052 2364 -2046
rect 2358 -2058 2364 -2052
rect 2358 -2064 2364 -2058
rect 2358 -2070 2364 -2064
rect 2358 -2076 2364 -2070
rect 2358 -2082 2364 -2076
rect 2358 -2088 2364 -2082
rect 2358 -2094 2364 -2088
rect 2358 -2100 2364 -2094
rect 2358 -2106 2364 -2100
rect 2358 -2112 2364 -2106
rect 2358 -2118 2364 -2112
rect 2358 -2124 2364 -2118
rect 2358 -2130 2364 -2124
rect 2358 -2136 2364 -2130
rect 2358 -2142 2364 -2136
rect 2358 -2148 2364 -2142
rect 2358 -2226 2364 -2220
rect 2358 -2232 2364 -2226
rect 2358 -2238 2364 -2232
rect 2358 -2244 2364 -2238
rect 2358 -2250 2364 -2244
rect 2358 -2256 2364 -2250
rect 2358 -2262 2364 -2256
rect 2358 -2268 2364 -2262
rect 2358 -2274 2364 -2268
rect 2358 -2280 2364 -2274
rect 2358 -2286 2364 -2280
rect 2358 -2292 2364 -2286
rect 2358 -2298 2364 -2292
rect 2358 -2304 2364 -2298
rect 2358 -2310 2364 -2304
rect 2358 -2316 2364 -2310
rect 2358 -2322 2364 -2316
rect 2358 -2328 2364 -2322
rect 2358 -2334 2364 -2328
rect 2358 -2340 2364 -2334
rect 2358 -2346 2364 -2340
rect 2358 -2352 2364 -2346
rect 2358 -2358 2364 -2352
rect 2358 -2364 2364 -2358
rect 2358 -2370 2364 -2364
rect 2358 -2376 2364 -2370
rect 2358 -2382 2364 -2376
rect 2358 -2388 2364 -2382
rect 2358 -2394 2364 -2388
rect 2358 -2400 2364 -2394
rect 2358 -2406 2364 -2400
rect 2358 -2412 2364 -2406
rect 2358 -2418 2364 -2412
rect 2358 -2424 2364 -2418
rect 2358 -2490 2364 -2484
rect 2358 -2496 2364 -2490
rect 2358 -2502 2364 -2496
rect 2358 -2508 2364 -2502
rect 2358 -2514 2364 -2508
rect 2358 -2520 2364 -2514
rect 2358 -2526 2364 -2520
rect 2358 -2532 2364 -2526
rect 2358 -2538 2364 -2532
rect 2358 -2544 2364 -2538
rect 2358 -2550 2364 -2544
rect 2358 -2556 2364 -2550
rect 2358 -2562 2364 -2556
rect 2358 -2568 2364 -2562
rect 2358 -2574 2364 -2568
rect 2358 -2580 2364 -2574
rect 2358 -2586 2364 -2580
rect 2358 -2592 2364 -2586
rect 2358 -2598 2364 -2592
rect 2358 -2604 2364 -2598
rect 2358 -2610 2364 -2604
rect 2358 -2616 2364 -2610
rect 2358 -2622 2364 -2616
rect 2358 -2628 2364 -2622
rect 2358 -2634 2364 -2628
rect 2358 -2640 2364 -2634
rect 2358 -2646 2364 -2640
rect 2358 -2652 2364 -2646
rect 2358 -2658 2364 -2652
rect 2358 -2664 2364 -2658
rect 2358 -2670 2364 -2664
rect 2358 -2676 2364 -2670
rect 2358 -2682 2364 -2676
rect 2358 -2688 2364 -2682
rect 2358 -2694 2364 -2688
rect 2358 -2700 2364 -2694
rect 2358 -2706 2364 -2700
rect 2358 -2712 2364 -2706
rect 2358 -2718 2364 -2712
rect 2358 -2724 2364 -2718
rect 2358 -2730 2364 -2724
rect 2358 -2736 2364 -2730
rect 2358 -2742 2364 -2736
rect 2358 -2748 2364 -2742
rect 2358 -2754 2364 -2748
rect 2358 -2760 2364 -2754
rect 2358 -2766 2364 -2760
rect 2358 -2772 2364 -2766
rect 2358 -2778 2364 -2772
rect 2358 -2784 2364 -2778
rect 2358 -2790 2364 -2784
rect 2358 -2796 2364 -2790
rect 2358 -2802 2364 -2796
rect 2358 -2808 2364 -2802
rect 2358 -2814 2364 -2808
rect 2358 -2820 2364 -2814
rect 2358 -2826 2364 -2820
rect 2358 -2832 2364 -2826
rect 2358 -2838 2364 -2832
rect 2358 -2844 2364 -2838
rect 2358 -2850 2364 -2844
rect 2358 -2856 2364 -2850
rect 2358 -2862 2364 -2856
rect 2358 -2868 2364 -2862
rect 2358 -2874 2364 -2868
rect 2358 -2880 2364 -2874
rect 2358 -2886 2364 -2880
rect 2358 -2892 2364 -2886
rect 2358 -2898 2364 -2892
rect 2358 -2904 2364 -2898
rect 2358 -2910 2364 -2904
rect 2364 -36 2370 -30
rect 2364 -42 2370 -36
rect 2364 -48 2370 -42
rect 2364 -54 2370 -48
rect 2364 -60 2370 -54
rect 2364 -66 2370 -60
rect 2364 -72 2370 -66
rect 2364 -78 2370 -72
rect 2364 -84 2370 -78
rect 2364 -90 2370 -84
rect 2364 -96 2370 -90
rect 2364 -102 2370 -96
rect 2364 -108 2370 -102
rect 2364 -114 2370 -108
rect 2364 -120 2370 -114
rect 2364 -126 2370 -120
rect 2364 -132 2370 -126
rect 2364 -138 2370 -132
rect 2364 -144 2370 -138
rect 2364 -150 2370 -144
rect 2364 -156 2370 -150
rect 2364 -162 2370 -156
rect 2364 -168 2370 -162
rect 2364 -174 2370 -168
rect 2364 -180 2370 -174
rect 2364 -186 2370 -180
rect 2364 -192 2370 -186
rect 2364 -198 2370 -192
rect 2364 -204 2370 -198
rect 2364 -210 2370 -204
rect 2364 -216 2370 -210
rect 2364 -222 2370 -216
rect 2364 -228 2370 -222
rect 2364 -234 2370 -228
rect 2364 -240 2370 -234
rect 2364 -246 2370 -240
rect 2364 -252 2370 -246
rect 2364 -258 2370 -252
rect 2364 -264 2370 -258
rect 2364 -270 2370 -264
rect 2364 -276 2370 -270
rect 2364 -282 2370 -276
rect 2364 -288 2370 -282
rect 2364 -294 2370 -288
rect 2364 -300 2370 -294
rect 2364 -306 2370 -300
rect 2364 -312 2370 -306
rect 2364 -318 2370 -312
rect 2364 -324 2370 -318
rect 2364 -330 2370 -324
rect 2364 -336 2370 -330
rect 2364 -342 2370 -336
rect 2364 -348 2370 -342
rect 2364 -354 2370 -348
rect 2364 -360 2370 -354
rect 2364 -366 2370 -360
rect 2364 -372 2370 -366
rect 2364 -378 2370 -372
rect 2364 -384 2370 -378
rect 2364 -390 2370 -384
rect 2364 -396 2370 -390
rect 2364 -402 2370 -396
rect 2364 -408 2370 -402
rect 2364 -414 2370 -408
rect 2364 -420 2370 -414
rect 2364 -426 2370 -420
rect 2364 -432 2370 -426
rect 2364 -438 2370 -432
rect 2364 -444 2370 -438
rect 2364 -450 2370 -444
rect 2364 -456 2370 -450
rect 2364 -462 2370 -456
rect 2364 -468 2370 -462
rect 2364 -474 2370 -468
rect 2364 -480 2370 -474
rect 2364 -486 2370 -480
rect 2364 -492 2370 -486
rect 2364 -498 2370 -492
rect 2364 -504 2370 -498
rect 2364 -510 2370 -504
rect 2364 -516 2370 -510
rect 2364 -522 2370 -516
rect 2364 -528 2370 -522
rect 2364 -534 2370 -528
rect 2364 -540 2370 -534
rect 2364 -546 2370 -540
rect 2364 -552 2370 -546
rect 2364 -558 2370 -552
rect 2364 -564 2370 -558
rect 2364 -570 2370 -564
rect 2364 -576 2370 -570
rect 2364 -582 2370 -576
rect 2364 -588 2370 -582
rect 2364 -594 2370 -588
rect 2364 -600 2370 -594
rect 2364 -606 2370 -600
rect 2364 -612 2370 -606
rect 2364 -618 2370 -612
rect 2364 -624 2370 -618
rect 2364 -630 2370 -624
rect 2364 -636 2370 -630
rect 2364 -642 2370 -636
rect 2364 -648 2370 -642
rect 2364 -654 2370 -648
rect 2364 -660 2370 -654
rect 2364 -666 2370 -660
rect 2364 -672 2370 -666
rect 2364 -678 2370 -672
rect 2364 -684 2370 -678
rect 2364 -690 2370 -684
rect 2364 -696 2370 -690
rect 2364 -702 2370 -696
rect 2364 -708 2370 -702
rect 2364 -714 2370 -708
rect 2364 -720 2370 -714
rect 2364 -726 2370 -720
rect 2364 -732 2370 -726
rect 2364 -738 2370 -732
rect 2364 -744 2370 -738
rect 2364 -750 2370 -744
rect 2364 -756 2370 -750
rect 2364 -762 2370 -756
rect 2364 -768 2370 -762
rect 2364 -774 2370 -768
rect 2364 -780 2370 -774
rect 2364 -786 2370 -780
rect 2364 -792 2370 -786
rect 2364 -798 2370 -792
rect 2364 -804 2370 -798
rect 2364 -810 2370 -804
rect 2364 -1416 2370 -1410
rect 2364 -1422 2370 -1416
rect 2364 -1428 2370 -1422
rect 2364 -1434 2370 -1428
rect 2364 -1440 2370 -1434
rect 2364 -1446 2370 -1440
rect 2364 -1452 2370 -1446
rect 2364 -1458 2370 -1452
rect 2364 -1464 2370 -1458
rect 2364 -1470 2370 -1464
rect 2364 -1476 2370 -1470
rect 2364 -1482 2370 -1476
rect 2364 -1488 2370 -1482
rect 2364 -1494 2370 -1488
rect 2364 -1500 2370 -1494
rect 2364 -1506 2370 -1500
rect 2364 -1512 2370 -1506
rect 2364 -1518 2370 -1512
rect 2364 -1524 2370 -1518
rect 2364 -1530 2370 -1524
rect 2364 -1536 2370 -1530
rect 2364 -1542 2370 -1536
rect 2364 -1548 2370 -1542
rect 2364 -1554 2370 -1548
rect 2364 -1560 2370 -1554
rect 2364 -1566 2370 -1560
rect 2364 -1572 2370 -1566
rect 2364 -1578 2370 -1572
rect 2364 -1584 2370 -1578
rect 2364 -1590 2370 -1584
rect 2364 -1596 2370 -1590
rect 2364 -1602 2370 -1596
rect 2364 -1608 2370 -1602
rect 2364 -1614 2370 -1608
rect 2364 -1620 2370 -1614
rect 2364 -1626 2370 -1620
rect 2364 -1632 2370 -1626
rect 2364 -1638 2370 -1632
rect 2364 -1644 2370 -1638
rect 2364 -1650 2370 -1644
rect 2364 -1656 2370 -1650
rect 2364 -1662 2370 -1656
rect 2364 -1668 2370 -1662
rect 2364 -1674 2370 -1668
rect 2364 -1680 2370 -1674
rect 2364 -1686 2370 -1680
rect 2364 -1692 2370 -1686
rect 2364 -1698 2370 -1692
rect 2364 -1704 2370 -1698
rect 2364 -1710 2370 -1704
rect 2364 -1716 2370 -1710
rect 2364 -1722 2370 -1716
rect 2364 -1728 2370 -1722
rect 2364 -1734 2370 -1728
rect 2364 -1740 2370 -1734
rect 2364 -1746 2370 -1740
rect 2364 -1752 2370 -1746
rect 2364 -1758 2370 -1752
rect 2364 -1764 2370 -1758
rect 2364 -1770 2370 -1764
rect 2364 -1776 2370 -1770
rect 2364 -1782 2370 -1776
rect 2364 -1788 2370 -1782
rect 2364 -1794 2370 -1788
rect 2364 -1800 2370 -1794
rect 2364 -1806 2370 -1800
rect 2364 -1812 2370 -1806
rect 2364 -1818 2370 -1812
rect 2364 -1824 2370 -1818
rect 2364 -1830 2370 -1824
rect 2364 -1836 2370 -1830
rect 2364 -1842 2370 -1836
rect 2364 -1848 2370 -1842
rect 2364 -1854 2370 -1848
rect 2364 -1860 2370 -1854
rect 2364 -1866 2370 -1860
rect 2364 -1872 2370 -1866
rect 2364 -1878 2370 -1872
rect 2364 -1884 2370 -1878
rect 2364 -1890 2370 -1884
rect 2364 -1896 2370 -1890
rect 2364 -1902 2370 -1896
rect 2364 -1908 2370 -1902
rect 2364 -1914 2370 -1908
rect 2364 -1920 2370 -1914
rect 2364 -1926 2370 -1920
rect 2364 -1932 2370 -1926
rect 2364 -1938 2370 -1932
rect 2364 -1944 2370 -1938
rect 2364 -1950 2370 -1944
rect 2364 -1956 2370 -1950
rect 2364 -1962 2370 -1956
rect 2364 -1968 2370 -1962
rect 2364 -1974 2370 -1968
rect 2364 -1980 2370 -1974
rect 2364 -1986 2370 -1980
rect 2364 -1992 2370 -1986
rect 2364 -1998 2370 -1992
rect 2364 -2004 2370 -1998
rect 2364 -2010 2370 -2004
rect 2364 -2016 2370 -2010
rect 2364 -2022 2370 -2016
rect 2364 -2028 2370 -2022
rect 2364 -2034 2370 -2028
rect 2364 -2040 2370 -2034
rect 2364 -2046 2370 -2040
rect 2364 -2052 2370 -2046
rect 2364 -2058 2370 -2052
rect 2364 -2064 2370 -2058
rect 2364 -2070 2370 -2064
rect 2364 -2076 2370 -2070
rect 2364 -2082 2370 -2076
rect 2364 -2088 2370 -2082
rect 2364 -2094 2370 -2088
rect 2364 -2100 2370 -2094
rect 2364 -2106 2370 -2100
rect 2364 -2112 2370 -2106
rect 2364 -2118 2370 -2112
rect 2364 -2124 2370 -2118
rect 2364 -2130 2370 -2124
rect 2364 -2136 2370 -2130
rect 2364 -2142 2370 -2136
rect 2364 -2220 2370 -2214
rect 2364 -2226 2370 -2220
rect 2364 -2232 2370 -2226
rect 2364 -2238 2370 -2232
rect 2364 -2244 2370 -2238
rect 2364 -2250 2370 -2244
rect 2364 -2256 2370 -2250
rect 2364 -2262 2370 -2256
rect 2364 -2268 2370 -2262
rect 2364 -2274 2370 -2268
rect 2364 -2280 2370 -2274
rect 2364 -2286 2370 -2280
rect 2364 -2292 2370 -2286
rect 2364 -2298 2370 -2292
rect 2364 -2304 2370 -2298
rect 2364 -2310 2370 -2304
rect 2364 -2316 2370 -2310
rect 2364 -2322 2370 -2316
rect 2364 -2328 2370 -2322
rect 2364 -2334 2370 -2328
rect 2364 -2340 2370 -2334
rect 2364 -2346 2370 -2340
rect 2364 -2352 2370 -2346
rect 2364 -2358 2370 -2352
rect 2364 -2364 2370 -2358
rect 2364 -2370 2370 -2364
rect 2364 -2376 2370 -2370
rect 2364 -2382 2370 -2376
rect 2364 -2388 2370 -2382
rect 2364 -2394 2370 -2388
rect 2364 -2400 2370 -2394
rect 2364 -2406 2370 -2400
rect 2364 -2412 2370 -2406
rect 2364 -2418 2370 -2412
rect 2364 -2490 2370 -2484
rect 2364 -2496 2370 -2490
rect 2364 -2502 2370 -2496
rect 2364 -2508 2370 -2502
rect 2364 -2514 2370 -2508
rect 2364 -2520 2370 -2514
rect 2364 -2526 2370 -2520
rect 2364 -2532 2370 -2526
rect 2364 -2538 2370 -2532
rect 2364 -2544 2370 -2538
rect 2364 -2550 2370 -2544
rect 2364 -2556 2370 -2550
rect 2364 -2562 2370 -2556
rect 2364 -2568 2370 -2562
rect 2364 -2574 2370 -2568
rect 2364 -2580 2370 -2574
rect 2364 -2586 2370 -2580
rect 2364 -2592 2370 -2586
rect 2364 -2598 2370 -2592
rect 2364 -2604 2370 -2598
rect 2364 -2610 2370 -2604
rect 2364 -2616 2370 -2610
rect 2364 -2622 2370 -2616
rect 2364 -2628 2370 -2622
rect 2364 -2634 2370 -2628
rect 2364 -2640 2370 -2634
rect 2364 -2646 2370 -2640
rect 2364 -2652 2370 -2646
rect 2364 -2658 2370 -2652
rect 2364 -2664 2370 -2658
rect 2364 -2670 2370 -2664
rect 2364 -2676 2370 -2670
rect 2364 -2682 2370 -2676
rect 2364 -2688 2370 -2682
rect 2364 -2694 2370 -2688
rect 2364 -2700 2370 -2694
rect 2364 -2706 2370 -2700
rect 2364 -2712 2370 -2706
rect 2364 -2718 2370 -2712
rect 2364 -2724 2370 -2718
rect 2364 -2730 2370 -2724
rect 2364 -2736 2370 -2730
rect 2364 -2742 2370 -2736
rect 2364 -2748 2370 -2742
rect 2364 -2754 2370 -2748
rect 2364 -2760 2370 -2754
rect 2364 -2766 2370 -2760
rect 2364 -2772 2370 -2766
rect 2364 -2778 2370 -2772
rect 2364 -2784 2370 -2778
rect 2364 -2790 2370 -2784
rect 2364 -2796 2370 -2790
rect 2364 -2802 2370 -2796
rect 2364 -2808 2370 -2802
rect 2364 -2814 2370 -2808
rect 2364 -2820 2370 -2814
rect 2364 -2826 2370 -2820
rect 2364 -2832 2370 -2826
rect 2364 -2838 2370 -2832
rect 2364 -2844 2370 -2838
rect 2364 -2850 2370 -2844
rect 2364 -2856 2370 -2850
rect 2364 -2862 2370 -2856
rect 2364 -2868 2370 -2862
rect 2364 -2874 2370 -2868
rect 2364 -2880 2370 -2874
rect 2364 -2886 2370 -2880
rect 2364 -2892 2370 -2886
rect 2364 -2898 2370 -2892
rect 2364 -2904 2370 -2898
rect 2364 -2910 2370 -2904
rect 2370 -60 2376 -54
rect 2370 -66 2376 -60
rect 2370 -72 2376 -66
rect 2370 -78 2376 -72
rect 2370 -84 2376 -78
rect 2370 -90 2376 -84
rect 2370 -96 2376 -90
rect 2370 -102 2376 -96
rect 2370 -108 2376 -102
rect 2370 -114 2376 -108
rect 2370 -120 2376 -114
rect 2370 -126 2376 -120
rect 2370 -132 2376 -126
rect 2370 -138 2376 -132
rect 2370 -144 2376 -138
rect 2370 -150 2376 -144
rect 2370 -156 2376 -150
rect 2370 -162 2376 -156
rect 2370 -168 2376 -162
rect 2370 -174 2376 -168
rect 2370 -180 2376 -174
rect 2370 -186 2376 -180
rect 2370 -192 2376 -186
rect 2370 -198 2376 -192
rect 2370 -204 2376 -198
rect 2370 -210 2376 -204
rect 2370 -216 2376 -210
rect 2370 -222 2376 -216
rect 2370 -228 2376 -222
rect 2370 -234 2376 -228
rect 2370 -240 2376 -234
rect 2370 -246 2376 -240
rect 2370 -252 2376 -246
rect 2370 -258 2376 -252
rect 2370 -264 2376 -258
rect 2370 -270 2376 -264
rect 2370 -276 2376 -270
rect 2370 -282 2376 -276
rect 2370 -288 2376 -282
rect 2370 -294 2376 -288
rect 2370 -300 2376 -294
rect 2370 -306 2376 -300
rect 2370 -312 2376 -306
rect 2370 -318 2376 -312
rect 2370 -324 2376 -318
rect 2370 -330 2376 -324
rect 2370 -336 2376 -330
rect 2370 -342 2376 -336
rect 2370 -348 2376 -342
rect 2370 -354 2376 -348
rect 2370 -360 2376 -354
rect 2370 -366 2376 -360
rect 2370 -372 2376 -366
rect 2370 -378 2376 -372
rect 2370 -384 2376 -378
rect 2370 -390 2376 -384
rect 2370 -396 2376 -390
rect 2370 -402 2376 -396
rect 2370 -408 2376 -402
rect 2370 -414 2376 -408
rect 2370 -420 2376 -414
rect 2370 -426 2376 -420
rect 2370 -432 2376 -426
rect 2370 -438 2376 -432
rect 2370 -444 2376 -438
rect 2370 -450 2376 -444
rect 2370 -456 2376 -450
rect 2370 -462 2376 -456
rect 2370 -468 2376 -462
rect 2370 -474 2376 -468
rect 2370 -480 2376 -474
rect 2370 -486 2376 -480
rect 2370 -492 2376 -486
rect 2370 -498 2376 -492
rect 2370 -504 2376 -498
rect 2370 -510 2376 -504
rect 2370 -516 2376 -510
rect 2370 -522 2376 -516
rect 2370 -528 2376 -522
rect 2370 -534 2376 -528
rect 2370 -540 2376 -534
rect 2370 -546 2376 -540
rect 2370 -552 2376 -546
rect 2370 -558 2376 -552
rect 2370 -564 2376 -558
rect 2370 -570 2376 -564
rect 2370 -576 2376 -570
rect 2370 -582 2376 -576
rect 2370 -588 2376 -582
rect 2370 -594 2376 -588
rect 2370 -600 2376 -594
rect 2370 -606 2376 -600
rect 2370 -612 2376 -606
rect 2370 -618 2376 -612
rect 2370 -624 2376 -618
rect 2370 -630 2376 -624
rect 2370 -636 2376 -630
rect 2370 -642 2376 -636
rect 2370 -648 2376 -642
rect 2370 -654 2376 -648
rect 2370 -660 2376 -654
rect 2370 -666 2376 -660
rect 2370 -672 2376 -666
rect 2370 -678 2376 -672
rect 2370 -684 2376 -678
rect 2370 -690 2376 -684
rect 2370 -696 2376 -690
rect 2370 -702 2376 -696
rect 2370 -708 2376 -702
rect 2370 -714 2376 -708
rect 2370 -720 2376 -714
rect 2370 -726 2376 -720
rect 2370 -732 2376 -726
rect 2370 -738 2376 -732
rect 2370 -744 2376 -738
rect 2370 -750 2376 -744
rect 2370 -756 2376 -750
rect 2370 -762 2376 -756
rect 2370 -768 2376 -762
rect 2370 -774 2376 -768
rect 2370 -780 2376 -774
rect 2370 -786 2376 -780
rect 2370 -792 2376 -786
rect 2370 -1410 2376 -1404
rect 2370 -1416 2376 -1410
rect 2370 -1422 2376 -1416
rect 2370 -1428 2376 -1422
rect 2370 -1434 2376 -1428
rect 2370 -1440 2376 -1434
rect 2370 -1446 2376 -1440
rect 2370 -1452 2376 -1446
rect 2370 -1458 2376 -1452
rect 2370 -1464 2376 -1458
rect 2370 -1470 2376 -1464
rect 2370 -1476 2376 -1470
rect 2370 -1482 2376 -1476
rect 2370 -1488 2376 -1482
rect 2370 -1494 2376 -1488
rect 2370 -1500 2376 -1494
rect 2370 -1506 2376 -1500
rect 2370 -1512 2376 -1506
rect 2370 -1518 2376 -1512
rect 2370 -1524 2376 -1518
rect 2370 -1530 2376 -1524
rect 2370 -1536 2376 -1530
rect 2370 -1542 2376 -1536
rect 2370 -1548 2376 -1542
rect 2370 -1554 2376 -1548
rect 2370 -1560 2376 -1554
rect 2370 -1566 2376 -1560
rect 2370 -1572 2376 -1566
rect 2370 -1578 2376 -1572
rect 2370 -1584 2376 -1578
rect 2370 -1590 2376 -1584
rect 2370 -1596 2376 -1590
rect 2370 -1602 2376 -1596
rect 2370 -1608 2376 -1602
rect 2370 -1614 2376 -1608
rect 2370 -1620 2376 -1614
rect 2370 -1626 2376 -1620
rect 2370 -1632 2376 -1626
rect 2370 -1638 2376 -1632
rect 2370 -1644 2376 -1638
rect 2370 -1650 2376 -1644
rect 2370 -1656 2376 -1650
rect 2370 -1662 2376 -1656
rect 2370 -1668 2376 -1662
rect 2370 -1674 2376 -1668
rect 2370 -1680 2376 -1674
rect 2370 -1686 2376 -1680
rect 2370 -1692 2376 -1686
rect 2370 -1698 2376 -1692
rect 2370 -1704 2376 -1698
rect 2370 -1710 2376 -1704
rect 2370 -1716 2376 -1710
rect 2370 -1722 2376 -1716
rect 2370 -1728 2376 -1722
rect 2370 -1734 2376 -1728
rect 2370 -1740 2376 -1734
rect 2370 -1746 2376 -1740
rect 2370 -1752 2376 -1746
rect 2370 -1758 2376 -1752
rect 2370 -1764 2376 -1758
rect 2370 -1770 2376 -1764
rect 2370 -1776 2376 -1770
rect 2370 -1782 2376 -1776
rect 2370 -1788 2376 -1782
rect 2370 -1794 2376 -1788
rect 2370 -1800 2376 -1794
rect 2370 -1806 2376 -1800
rect 2370 -1812 2376 -1806
rect 2370 -1818 2376 -1812
rect 2370 -1824 2376 -1818
rect 2370 -1830 2376 -1824
rect 2370 -1836 2376 -1830
rect 2370 -1842 2376 -1836
rect 2370 -1848 2376 -1842
rect 2370 -1854 2376 -1848
rect 2370 -1860 2376 -1854
rect 2370 -1866 2376 -1860
rect 2370 -1872 2376 -1866
rect 2370 -1878 2376 -1872
rect 2370 -1884 2376 -1878
rect 2370 -1890 2376 -1884
rect 2370 -1896 2376 -1890
rect 2370 -1902 2376 -1896
rect 2370 -1908 2376 -1902
rect 2370 -1914 2376 -1908
rect 2370 -1920 2376 -1914
rect 2370 -1926 2376 -1920
rect 2370 -1932 2376 -1926
rect 2370 -1938 2376 -1932
rect 2370 -1944 2376 -1938
rect 2370 -1950 2376 -1944
rect 2370 -1956 2376 -1950
rect 2370 -1962 2376 -1956
rect 2370 -1968 2376 -1962
rect 2370 -1974 2376 -1968
rect 2370 -1980 2376 -1974
rect 2370 -1986 2376 -1980
rect 2370 -1992 2376 -1986
rect 2370 -1998 2376 -1992
rect 2370 -2004 2376 -1998
rect 2370 -2010 2376 -2004
rect 2370 -2016 2376 -2010
rect 2370 -2022 2376 -2016
rect 2370 -2028 2376 -2022
rect 2370 -2034 2376 -2028
rect 2370 -2040 2376 -2034
rect 2370 -2046 2376 -2040
rect 2370 -2052 2376 -2046
rect 2370 -2058 2376 -2052
rect 2370 -2064 2376 -2058
rect 2370 -2070 2376 -2064
rect 2370 -2076 2376 -2070
rect 2370 -2082 2376 -2076
rect 2370 -2088 2376 -2082
rect 2370 -2094 2376 -2088
rect 2370 -2100 2376 -2094
rect 2370 -2106 2376 -2100
rect 2370 -2112 2376 -2106
rect 2370 -2118 2376 -2112
rect 2370 -2124 2376 -2118
rect 2370 -2130 2376 -2124
rect 2370 -2136 2376 -2130
rect 2370 -2214 2376 -2208
rect 2370 -2220 2376 -2214
rect 2370 -2226 2376 -2220
rect 2370 -2232 2376 -2226
rect 2370 -2238 2376 -2232
rect 2370 -2244 2376 -2238
rect 2370 -2250 2376 -2244
rect 2370 -2256 2376 -2250
rect 2370 -2262 2376 -2256
rect 2370 -2268 2376 -2262
rect 2370 -2274 2376 -2268
rect 2370 -2280 2376 -2274
rect 2370 -2286 2376 -2280
rect 2370 -2292 2376 -2286
rect 2370 -2298 2376 -2292
rect 2370 -2304 2376 -2298
rect 2370 -2310 2376 -2304
rect 2370 -2316 2376 -2310
rect 2370 -2322 2376 -2316
rect 2370 -2328 2376 -2322
rect 2370 -2334 2376 -2328
rect 2370 -2340 2376 -2334
rect 2370 -2346 2376 -2340
rect 2370 -2352 2376 -2346
rect 2370 -2358 2376 -2352
rect 2370 -2364 2376 -2358
rect 2370 -2370 2376 -2364
rect 2370 -2376 2376 -2370
rect 2370 -2382 2376 -2376
rect 2370 -2388 2376 -2382
rect 2370 -2394 2376 -2388
rect 2370 -2400 2376 -2394
rect 2370 -2406 2376 -2400
rect 2370 -2412 2376 -2406
rect 2370 -2418 2376 -2412
rect 2370 -2484 2376 -2478
rect 2370 -2490 2376 -2484
rect 2370 -2496 2376 -2490
rect 2370 -2502 2376 -2496
rect 2370 -2508 2376 -2502
rect 2370 -2514 2376 -2508
rect 2370 -2520 2376 -2514
rect 2370 -2526 2376 -2520
rect 2370 -2532 2376 -2526
rect 2370 -2538 2376 -2532
rect 2370 -2544 2376 -2538
rect 2370 -2550 2376 -2544
rect 2370 -2556 2376 -2550
rect 2370 -2562 2376 -2556
rect 2370 -2568 2376 -2562
rect 2370 -2574 2376 -2568
rect 2370 -2580 2376 -2574
rect 2370 -2586 2376 -2580
rect 2370 -2592 2376 -2586
rect 2370 -2598 2376 -2592
rect 2370 -2604 2376 -2598
rect 2370 -2610 2376 -2604
rect 2370 -2616 2376 -2610
rect 2370 -2622 2376 -2616
rect 2370 -2628 2376 -2622
rect 2370 -2634 2376 -2628
rect 2370 -2640 2376 -2634
rect 2370 -2646 2376 -2640
rect 2370 -2652 2376 -2646
rect 2370 -2658 2376 -2652
rect 2370 -2664 2376 -2658
rect 2370 -2670 2376 -2664
rect 2370 -2676 2376 -2670
rect 2370 -2682 2376 -2676
rect 2370 -2688 2376 -2682
rect 2370 -2694 2376 -2688
rect 2370 -2700 2376 -2694
rect 2370 -2706 2376 -2700
rect 2370 -2712 2376 -2706
rect 2370 -2718 2376 -2712
rect 2370 -2724 2376 -2718
rect 2370 -2730 2376 -2724
rect 2370 -2736 2376 -2730
rect 2370 -2742 2376 -2736
rect 2370 -2748 2376 -2742
rect 2370 -2754 2376 -2748
rect 2370 -2760 2376 -2754
rect 2370 -2766 2376 -2760
rect 2370 -2772 2376 -2766
rect 2370 -2778 2376 -2772
rect 2370 -2784 2376 -2778
rect 2370 -2790 2376 -2784
rect 2370 -2796 2376 -2790
rect 2370 -2802 2376 -2796
rect 2370 -2808 2376 -2802
rect 2370 -2814 2376 -2808
rect 2370 -2820 2376 -2814
rect 2370 -2826 2376 -2820
rect 2370 -2832 2376 -2826
rect 2370 -2838 2376 -2832
rect 2370 -2844 2376 -2838
rect 2370 -2850 2376 -2844
rect 2370 -2856 2376 -2850
rect 2370 -2862 2376 -2856
rect 2370 -2868 2376 -2862
rect 2370 -2874 2376 -2868
rect 2370 -2880 2376 -2874
rect 2370 -2886 2376 -2880
rect 2370 -2892 2376 -2886
rect 2370 -2898 2376 -2892
rect 2370 -2904 2376 -2898
rect 2376 -78 2382 -72
rect 2376 -84 2382 -78
rect 2376 -90 2382 -84
rect 2376 -96 2382 -90
rect 2376 -102 2382 -96
rect 2376 -108 2382 -102
rect 2376 -114 2382 -108
rect 2376 -120 2382 -114
rect 2376 -126 2382 -120
rect 2376 -132 2382 -126
rect 2376 -138 2382 -132
rect 2376 -144 2382 -138
rect 2376 -150 2382 -144
rect 2376 -156 2382 -150
rect 2376 -162 2382 -156
rect 2376 -168 2382 -162
rect 2376 -174 2382 -168
rect 2376 -180 2382 -174
rect 2376 -186 2382 -180
rect 2376 -192 2382 -186
rect 2376 -198 2382 -192
rect 2376 -204 2382 -198
rect 2376 -210 2382 -204
rect 2376 -216 2382 -210
rect 2376 -222 2382 -216
rect 2376 -228 2382 -222
rect 2376 -234 2382 -228
rect 2376 -240 2382 -234
rect 2376 -246 2382 -240
rect 2376 -252 2382 -246
rect 2376 -258 2382 -252
rect 2376 -264 2382 -258
rect 2376 -270 2382 -264
rect 2376 -276 2382 -270
rect 2376 -282 2382 -276
rect 2376 -288 2382 -282
rect 2376 -294 2382 -288
rect 2376 -300 2382 -294
rect 2376 -306 2382 -300
rect 2376 -312 2382 -306
rect 2376 -318 2382 -312
rect 2376 -324 2382 -318
rect 2376 -330 2382 -324
rect 2376 -336 2382 -330
rect 2376 -342 2382 -336
rect 2376 -348 2382 -342
rect 2376 -354 2382 -348
rect 2376 -360 2382 -354
rect 2376 -366 2382 -360
rect 2376 -372 2382 -366
rect 2376 -378 2382 -372
rect 2376 -384 2382 -378
rect 2376 -390 2382 -384
rect 2376 -396 2382 -390
rect 2376 -402 2382 -396
rect 2376 -408 2382 -402
rect 2376 -414 2382 -408
rect 2376 -420 2382 -414
rect 2376 -426 2382 -420
rect 2376 -432 2382 -426
rect 2376 -438 2382 -432
rect 2376 -444 2382 -438
rect 2376 -450 2382 -444
rect 2376 -456 2382 -450
rect 2376 -462 2382 -456
rect 2376 -468 2382 -462
rect 2376 -474 2382 -468
rect 2376 -480 2382 -474
rect 2376 -486 2382 -480
rect 2376 -492 2382 -486
rect 2376 -498 2382 -492
rect 2376 -504 2382 -498
rect 2376 -510 2382 -504
rect 2376 -516 2382 -510
rect 2376 -522 2382 -516
rect 2376 -528 2382 -522
rect 2376 -534 2382 -528
rect 2376 -540 2382 -534
rect 2376 -546 2382 -540
rect 2376 -552 2382 -546
rect 2376 -558 2382 -552
rect 2376 -564 2382 -558
rect 2376 -570 2382 -564
rect 2376 -576 2382 -570
rect 2376 -582 2382 -576
rect 2376 -588 2382 -582
rect 2376 -594 2382 -588
rect 2376 -600 2382 -594
rect 2376 -606 2382 -600
rect 2376 -612 2382 -606
rect 2376 -618 2382 -612
rect 2376 -624 2382 -618
rect 2376 -630 2382 -624
rect 2376 -636 2382 -630
rect 2376 -642 2382 -636
rect 2376 -648 2382 -642
rect 2376 -654 2382 -648
rect 2376 -660 2382 -654
rect 2376 -666 2382 -660
rect 2376 -672 2382 -666
rect 2376 -678 2382 -672
rect 2376 -684 2382 -678
rect 2376 -690 2382 -684
rect 2376 -696 2382 -690
rect 2376 -702 2382 -696
rect 2376 -708 2382 -702
rect 2376 -714 2382 -708
rect 2376 -720 2382 -714
rect 2376 -726 2382 -720
rect 2376 -732 2382 -726
rect 2376 -738 2382 -732
rect 2376 -744 2382 -738
rect 2376 -750 2382 -744
rect 2376 -756 2382 -750
rect 2376 -762 2382 -756
rect 2376 -768 2382 -762
rect 2376 -774 2382 -768
rect 2376 -1404 2382 -1398
rect 2376 -1410 2382 -1404
rect 2376 -1416 2382 -1410
rect 2376 -1422 2382 -1416
rect 2376 -1428 2382 -1422
rect 2376 -1434 2382 -1428
rect 2376 -1440 2382 -1434
rect 2376 -1446 2382 -1440
rect 2376 -1452 2382 -1446
rect 2376 -1458 2382 -1452
rect 2376 -1464 2382 -1458
rect 2376 -1470 2382 -1464
rect 2376 -1476 2382 -1470
rect 2376 -1482 2382 -1476
rect 2376 -1488 2382 -1482
rect 2376 -1494 2382 -1488
rect 2376 -1500 2382 -1494
rect 2376 -1506 2382 -1500
rect 2376 -1512 2382 -1506
rect 2376 -1518 2382 -1512
rect 2376 -1524 2382 -1518
rect 2376 -1530 2382 -1524
rect 2376 -1536 2382 -1530
rect 2376 -1542 2382 -1536
rect 2376 -1548 2382 -1542
rect 2376 -1554 2382 -1548
rect 2376 -1560 2382 -1554
rect 2376 -1566 2382 -1560
rect 2376 -1572 2382 -1566
rect 2376 -1578 2382 -1572
rect 2376 -1584 2382 -1578
rect 2376 -1590 2382 -1584
rect 2376 -1596 2382 -1590
rect 2376 -1602 2382 -1596
rect 2376 -1608 2382 -1602
rect 2376 -1614 2382 -1608
rect 2376 -1620 2382 -1614
rect 2376 -1626 2382 -1620
rect 2376 -1632 2382 -1626
rect 2376 -1638 2382 -1632
rect 2376 -1644 2382 -1638
rect 2376 -1650 2382 -1644
rect 2376 -1656 2382 -1650
rect 2376 -1662 2382 -1656
rect 2376 -1668 2382 -1662
rect 2376 -1674 2382 -1668
rect 2376 -1680 2382 -1674
rect 2376 -1686 2382 -1680
rect 2376 -1692 2382 -1686
rect 2376 -1698 2382 -1692
rect 2376 -1704 2382 -1698
rect 2376 -1710 2382 -1704
rect 2376 -1716 2382 -1710
rect 2376 -1722 2382 -1716
rect 2376 -1728 2382 -1722
rect 2376 -1734 2382 -1728
rect 2376 -1740 2382 -1734
rect 2376 -1746 2382 -1740
rect 2376 -1752 2382 -1746
rect 2376 -1758 2382 -1752
rect 2376 -1764 2382 -1758
rect 2376 -1770 2382 -1764
rect 2376 -1776 2382 -1770
rect 2376 -1782 2382 -1776
rect 2376 -1788 2382 -1782
rect 2376 -1794 2382 -1788
rect 2376 -1800 2382 -1794
rect 2376 -1806 2382 -1800
rect 2376 -1812 2382 -1806
rect 2376 -1818 2382 -1812
rect 2376 -1824 2382 -1818
rect 2376 -1830 2382 -1824
rect 2376 -1836 2382 -1830
rect 2376 -1842 2382 -1836
rect 2376 -1848 2382 -1842
rect 2376 -1854 2382 -1848
rect 2376 -1860 2382 -1854
rect 2376 -1866 2382 -1860
rect 2376 -1872 2382 -1866
rect 2376 -1878 2382 -1872
rect 2376 -1884 2382 -1878
rect 2376 -1890 2382 -1884
rect 2376 -1896 2382 -1890
rect 2376 -1902 2382 -1896
rect 2376 -1908 2382 -1902
rect 2376 -1914 2382 -1908
rect 2376 -1920 2382 -1914
rect 2376 -1926 2382 -1920
rect 2376 -1932 2382 -1926
rect 2376 -1938 2382 -1932
rect 2376 -1944 2382 -1938
rect 2376 -1950 2382 -1944
rect 2376 -1956 2382 -1950
rect 2376 -1962 2382 -1956
rect 2376 -1968 2382 -1962
rect 2376 -1974 2382 -1968
rect 2376 -1980 2382 -1974
rect 2376 -1986 2382 -1980
rect 2376 -1992 2382 -1986
rect 2376 -1998 2382 -1992
rect 2376 -2004 2382 -1998
rect 2376 -2010 2382 -2004
rect 2376 -2016 2382 -2010
rect 2376 -2022 2382 -2016
rect 2376 -2028 2382 -2022
rect 2376 -2034 2382 -2028
rect 2376 -2040 2382 -2034
rect 2376 -2046 2382 -2040
rect 2376 -2052 2382 -2046
rect 2376 -2058 2382 -2052
rect 2376 -2064 2382 -2058
rect 2376 -2070 2382 -2064
rect 2376 -2076 2382 -2070
rect 2376 -2082 2382 -2076
rect 2376 -2088 2382 -2082
rect 2376 -2094 2382 -2088
rect 2376 -2100 2382 -2094
rect 2376 -2106 2382 -2100
rect 2376 -2112 2382 -2106
rect 2376 -2118 2382 -2112
rect 2376 -2124 2382 -2118
rect 2376 -2130 2382 -2124
rect 2376 -2208 2382 -2202
rect 2376 -2214 2382 -2208
rect 2376 -2220 2382 -2214
rect 2376 -2226 2382 -2220
rect 2376 -2232 2382 -2226
rect 2376 -2238 2382 -2232
rect 2376 -2244 2382 -2238
rect 2376 -2250 2382 -2244
rect 2376 -2256 2382 -2250
rect 2376 -2262 2382 -2256
rect 2376 -2268 2382 -2262
rect 2376 -2274 2382 -2268
rect 2376 -2280 2382 -2274
rect 2376 -2286 2382 -2280
rect 2376 -2292 2382 -2286
rect 2376 -2298 2382 -2292
rect 2376 -2304 2382 -2298
rect 2376 -2310 2382 -2304
rect 2376 -2316 2382 -2310
rect 2376 -2322 2382 -2316
rect 2376 -2328 2382 -2322
rect 2376 -2334 2382 -2328
rect 2376 -2340 2382 -2334
rect 2376 -2346 2382 -2340
rect 2376 -2352 2382 -2346
rect 2376 -2358 2382 -2352
rect 2376 -2364 2382 -2358
rect 2376 -2370 2382 -2364
rect 2376 -2376 2382 -2370
rect 2376 -2382 2382 -2376
rect 2376 -2388 2382 -2382
rect 2376 -2394 2382 -2388
rect 2376 -2400 2382 -2394
rect 2376 -2406 2382 -2400
rect 2376 -2412 2382 -2406
rect 2376 -2418 2382 -2412
rect 2376 -2484 2382 -2478
rect 2376 -2490 2382 -2484
rect 2376 -2496 2382 -2490
rect 2376 -2502 2382 -2496
rect 2376 -2508 2382 -2502
rect 2376 -2514 2382 -2508
rect 2376 -2520 2382 -2514
rect 2376 -2526 2382 -2520
rect 2376 -2532 2382 -2526
rect 2376 -2538 2382 -2532
rect 2376 -2544 2382 -2538
rect 2376 -2550 2382 -2544
rect 2376 -2556 2382 -2550
rect 2376 -2562 2382 -2556
rect 2376 -2568 2382 -2562
rect 2376 -2574 2382 -2568
rect 2376 -2580 2382 -2574
rect 2376 -2586 2382 -2580
rect 2376 -2592 2382 -2586
rect 2376 -2598 2382 -2592
rect 2376 -2604 2382 -2598
rect 2376 -2610 2382 -2604
rect 2376 -2616 2382 -2610
rect 2376 -2622 2382 -2616
rect 2376 -2628 2382 -2622
rect 2376 -2634 2382 -2628
rect 2376 -2640 2382 -2634
rect 2376 -2646 2382 -2640
rect 2376 -2652 2382 -2646
rect 2376 -2658 2382 -2652
rect 2376 -2664 2382 -2658
rect 2376 -2670 2382 -2664
rect 2376 -2676 2382 -2670
rect 2376 -2682 2382 -2676
rect 2376 -2688 2382 -2682
rect 2376 -2694 2382 -2688
rect 2376 -2700 2382 -2694
rect 2376 -2706 2382 -2700
rect 2376 -2712 2382 -2706
rect 2376 -2718 2382 -2712
rect 2376 -2724 2382 -2718
rect 2376 -2730 2382 -2724
rect 2376 -2736 2382 -2730
rect 2376 -2742 2382 -2736
rect 2376 -2748 2382 -2742
rect 2376 -2754 2382 -2748
rect 2376 -2760 2382 -2754
rect 2376 -2766 2382 -2760
rect 2376 -2772 2382 -2766
rect 2376 -2778 2382 -2772
rect 2376 -2784 2382 -2778
rect 2376 -2790 2382 -2784
rect 2376 -2796 2382 -2790
rect 2376 -2802 2382 -2796
rect 2376 -2808 2382 -2802
rect 2376 -2814 2382 -2808
rect 2376 -2820 2382 -2814
rect 2376 -2826 2382 -2820
rect 2376 -2832 2382 -2826
rect 2376 -2838 2382 -2832
rect 2376 -2844 2382 -2838
rect 2376 -2850 2382 -2844
rect 2376 -2856 2382 -2850
rect 2376 -2862 2382 -2856
rect 2376 -2868 2382 -2862
rect 2376 -2874 2382 -2868
rect 2376 -2880 2382 -2874
rect 2376 -2886 2382 -2880
rect 2376 -2892 2382 -2886
rect 2376 -2898 2382 -2892
rect 2382 -102 2388 -96
rect 2382 -108 2388 -102
rect 2382 -114 2388 -108
rect 2382 -120 2388 -114
rect 2382 -126 2388 -120
rect 2382 -132 2388 -126
rect 2382 -138 2388 -132
rect 2382 -144 2388 -138
rect 2382 -150 2388 -144
rect 2382 -156 2388 -150
rect 2382 -162 2388 -156
rect 2382 -168 2388 -162
rect 2382 -174 2388 -168
rect 2382 -180 2388 -174
rect 2382 -186 2388 -180
rect 2382 -192 2388 -186
rect 2382 -198 2388 -192
rect 2382 -204 2388 -198
rect 2382 -210 2388 -204
rect 2382 -216 2388 -210
rect 2382 -222 2388 -216
rect 2382 -228 2388 -222
rect 2382 -234 2388 -228
rect 2382 -240 2388 -234
rect 2382 -246 2388 -240
rect 2382 -252 2388 -246
rect 2382 -258 2388 -252
rect 2382 -264 2388 -258
rect 2382 -270 2388 -264
rect 2382 -276 2388 -270
rect 2382 -282 2388 -276
rect 2382 -288 2388 -282
rect 2382 -294 2388 -288
rect 2382 -300 2388 -294
rect 2382 -306 2388 -300
rect 2382 -312 2388 -306
rect 2382 -318 2388 -312
rect 2382 -324 2388 -318
rect 2382 -330 2388 -324
rect 2382 -336 2388 -330
rect 2382 -342 2388 -336
rect 2382 -348 2388 -342
rect 2382 -354 2388 -348
rect 2382 -360 2388 -354
rect 2382 -366 2388 -360
rect 2382 -372 2388 -366
rect 2382 -378 2388 -372
rect 2382 -384 2388 -378
rect 2382 -390 2388 -384
rect 2382 -396 2388 -390
rect 2382 -402 2388 -396
rect 2382 -408 2388 -402
rect 2382 -414 2388 -408
rect 2382 -420 2388 -414
rect 2382 -426 2388 -420
rect 2382 -432 2388 -426
rect 2382 -438 2388 -432
rect 2382 -444 2388 -438
rect 2382 -450 2388 -444
rect 2382 -456 2388 -450
rect 2382 -462 2388 -456
rect 2382 -468 2388 -462
rect 2382 -474 2388 -468
rect 2382 -480 2388 -474
rect 2382 -486 2388 -480
rect 2382 -492 2388 -486
rect 2382 -498 2388 -492
rect 2382 -504 2388 -498
rect 2382 -510 2388 -504
rect 2382 -516 2388 -510
rect 2382 -522 2388 -516
rect 2382 -528 2388 -522
rect 2382 -534 2388 -528
rect 2382 -540 2388 -534
rect 2382 -546 2388 -540
rect 2382 -552 2388 -546
rect 2382 -558 2388 -552
rect 2382 -564 2388 -558
rect 2382 -570 2388 -564
rect 2382 -576 2388 -570
rect 2382 -582 2388 -576
rect 2382 -588 2388 -582
rect 2382 -594 2388 -588
rect 2382 -600 2388 -594
rect 2382 -606 2388 -600
rect 2382 -612 2388 -606
rect 2382 -618 2388 -612
rect 2382 -624 2388 -618
rect 2382 -630 2388 -624
rect 2382 -636 2388 -630
rect 2382 -642 2388 -636
rect 2382 -648 2388 -642
rect 2382 -654 2388 -648
rect 2382 -660 2388 -654
rect 2382 -666 2388 -660
rect 2382 -672 2388 -666
rect 2382 -678 2388 -672
rect 2382 -684 2388 -678
rect 2382 -690 2388 -684
rect 2382 -696 2388 -690
rect 2382 -702 2388 -696
rect 2382 -708 2388 -702
rect 2382 -714 2388 -708
rect 2382 -720 2388 -714
rect 2382 -726 2388 -720
rect 2382 -732 2388 -726
rect 2382 -738 2388 -732
rect 2382 -744 2388 -738
rect 2382 -750 2388 -744
rect 2382 -756 2388 -750
rect 2382 -1404 2388 -1398
rect 2382 -1410 2388 -1404
rect 2382 -1416 2388 -1410
rect 2382 -1422 2388 -1416
rect 2382 -1428 2388 -1422
rect 2382 -1434 2388 -1428
rect 2382 -1440 2388 -1434
rect 2382 -1446 2388 -1440
rect 2382 -1452 2388 -1446
rect 2382 -1458 2388 -1452
rect 2382 -1464 2388 -1458
rect 2382 -1470 2388 -1464
rect 2382 -1476 2388 -1470
rect 2382 -1482 2388 -1476
rect 2382 -1488 2388 -1482
rect 2382 -1494 2388 -1488
rect 2382 -1500 2388 -1494
rect 2382 -1506 2388 -1500
rect 2382 -1512 2388 -1506
rect 2382 -1518 2388 -1512
rect 2382 -1524 2388 -1518
rect 2382 -1530 2388 -1524
rect 2382 -1536 2388 -1530
rect 2382 -1542 2388 -1536
rect 2382 -1548 2388 -1542
rect 2382 -1554 2388 -1548
rect 2382 -1560 2388 -1554
rect 2382 -1566 2388 -1560
rect 2382 -1572 2388 -1566
rect 2382 -1578 2388 -1572
rect 2382 -1584 2388 -1578
rect 2382 -1590 2388 -1584
rect 2382 -1596 2388 -1590
rect 2382 -1602 2388 -1596
rect 2382 -1608 2388 -1602
rect 2382 -1614 2388 -1608
rect 2382 -1620 2388 -1614
rect 2382 -1626 2388 -1620
rect 2382 -1632 2388 -1626
rect 2382 -1638 2388 -1632
rect 2382 -1644 2388 -1638
rect 2382 -1650 2388 -1644
rect 2382 -1656 2388 -1650
rect 2382 -1662 2388 -1656
rect 2382 -1668 2388 -1662
rect 2382 -1674 2388 -1668
rect 2382 -1680 2388 -1674
rect 2382 -1686 2388 -1680
rect 2382 -1692 2388 -1686
rect 2382 -1698 2388 -1692
rect 2382 -1704 2388 -1698
rect 2382 -1710 2388 -1704
rect 2382 -1716 2388 -1710
rect 2382 -1722 2388 -1716
rect 2382 -1728 2388 -1722
rect 2382 -1734 2388 -1728
rect 2382 -1740 2388 -1734
rect 2382 -1746 2388 -1740
rect 2382 -1752 2388 -1746
rect 2382 -1758 2388 -1752
rect 2382 -1764 2388 -1758
rect 2382 -1770 2388 -1764
rect 2382 -1776 2388 -1770
rect 2382 -1782 2388 -1776
rect 2382 -1788 2388 -1782
rect 2382 -1794 2388 -1788
rect 2382 -1800 2388 -1794
rect 2382 -1806 2388 -1800
rect 2382 -1812 2388 -1806
rect 2382 -1818 2388 -1812
rect 2382 -1824 2388 -1818
rect 2382 -1830 2388 -1824
rect 2382 -1836 2388 -1830
rect 2382 -1842 2388 -1836
rect 2382 -1848 2388 -1842
rect 2382 -1854 2388 -1848
rect 2382 -1860 2388 -1854
rect 2382 -1866 2388 -1860
rect 2382 -1872 2388 -1866
rect 2382 -1878 2388 -1872
rect 2382 -1884 2388 -1878
rect 2382 -1890 2388 -1884
rect 2382 -1896 2388 -1890
rect 2382 -1902 2388 -1896
rect 2382 -1908 2388 -1902
rect 2382 -1914 2388 -1908
rect 2382 -1920 2388 -1914
rect 2382 -1926 2388 -1920
rect 2382 -1932 2388 -1926
rect 2382 -1938 2388 -1932
rect 2382 -1944 2388 -1938
rect 2382 -1950 2388 -1944
rect 2382 -1956 2388 -1950
rect 2382 -1962 2388 -1956
rect 2382 -1968 2388 -1962
rect 2382 -1974 2388 -1968
rect 2382 -1980 2388 -1974
rect 2382 -1986 2388 -1980
rect 2382 -1992 2388 -1986
rect 2382 -1998 2388 -1992
rect 2382 -2004 2388 -1998
rect 2382 -2010 2388 -2004
rect 2382 -2016 2388 -2010
rect 2382 -2022 2388 -2016
rect 2382 -2028 2388 -2022
rect 2382 -2034 2388 -2028
rect 2382 -2040 2388 -2034
rect 2382 -2046 2388 -2040
rect 2382 -2052 2388 -2046
rect 2382 -2058 2388 -2052
rect 2382 -2064 2388 -2058
rect 2382 -2070 2388 -2064
rect 2382 -2076 2388 -2070
rect 2382 -2082 2388 -2076
rect 2382 -2088 2388 -2082
rect 2382 -2094 2388 -2088
rect 2382 -2100 2388 -2094
rect 2382 -2106 2388 -2100
rect 2382 -2112 2388 -2106
rect 2382 -2118 2388 -2112
rect 2382 -2196 2388 -2190
rect 2382 -2202 2388 -2196
rect 2382 -2208 2388 -2202
rect 2382 -2214 2388 -2208
rect 2382 -2220 2388 -2214
rect 2382 -2226 2388 -2220
rect 2382 -2232 2388 -2226
rect 2382 -2238 2388 -2232
rect 2382 -2244 2388 -2238
rect 2382 -2250 2388 -2244
rect 2382 -2256 2388 -2250
rect 2382 -2262 2388 -2256
rect 2382 -2268 2388 -2262
rect 2382 -2274 2388 -2268
rect 2382 -2280 2388 -2274
rect 2382 -2286 2388 -2280
rect 2382 -2292 2388 -2286
rect 2382 -2298 2388 -2292
rect 2382 -2304 2388 -2298
rect 2382 -2310 2388 -2304
rect 2382 -2316 2388 -2310
rect 2382 -2322 2388 -2316
rect 2382 -2328 2388 -2322
rect 2382 -2334 2388 -2328
rect 2382 -2340 2388 -2334
rect 2382 -2346 2388 -2340
rect 2382 -2352 2388 -2346
rect 2382 -2358 2388 -2352
rect 2382 -2364 2388 -2358
rect 2382 -2370 2388 -2364
rect 2382 -2376 2388 -2370
rect 2382 -2382 2388 -2376
rect 2382 -2388 2388 -2382
rect 2382 -2394 2388 -2388
rect 2382 -2400 2388 -2394
rect 2382 -2406 2388 -2400
rect 2382 -2412 2388 -2406
rect 2382 -2484 2388 -2478
rect 2382 -2490 2388 -2484
rect 2382 -2496 2388 -2490
rect 2382 -2502 2388 -2496
rect 2382 -2508 2388 -2502
rect 2382 -2514 2388 -2508
rect 2382 -2520 2388 -2514
rect 2382 -2526 2388 -2520
rect 2382 -2532 2388 -2526
rect 2382 -2538 2388 -2532
rect 2382 -2544 2388 -2538
rect 2382 -2550 2388 -2544
rect 2382 -2556 2388 -2550
rect 2382 -2562 2388 -2556
rect 2382 -2568 2388 -2562
rect 2382 -2574 2388 -2568
rect 2382 -2580 2388 -2574
rect 2382 -2586 2388 -2580
rect 2382 -2592 2388 -2586
rect 2382 -2598 2388 -2592
rect 2382 -2604 2388 -2598
rect 2382 -2610 2388 -2604
rect 2382 -2616 2388 -2610
rect 2382 -2622 2388 -2616
rect 2382 -2628 2388 -2622
rect 2382 -2634 2388 -2628
rect 2382 -2640 2388 -2634
rect 2382 -2646 2388 -2640
rect 2382 -2652 2388 -2646
rect 2382 -2658 2388 -2652
rect 2382 -2664 2388 -2658
rect 2382 -2670 2388 -2664
rect 2382 -2676 2388 -2670
rect 2382 -2682 2388 -2676
rect 2382 -2688 2388 -2682
rect 2382 -2694 2388 -2688
rect 2382 -2700 2388 -2694
rect 2382 -2706 2388 -2700
rect 2382 -2712 2388 -2706
rect 2382 -2718 2388 -2712
rect 2382 -2724 2388 -2718
rect 2382 -2730 2388 -2724
rect 2382 -2736 2388 -2730
rect 2382 -2742 2388 -2736
rect 2382 -2748 2388 -2742
rect 2382 -2754 2388 -2748
rect 2382 -2760 2388 -2754
rect 2382 -2766 2388 -2760
rect 2382 -2772 2388 -2766
rect 2382 -2778 2388 -2772
rect 2382 -2784 2388 -2778
rect 2382 -2790 2388 -2784
rect 2382 -2796 2388 -2790
rect 2382 -2802 2388 -2796
rect 2382 -2808 2388 -2802
rect 2382 -2814 2388 -2808
rect 2382 -2820 2388 -2814
rect 2382 -2826 2388 -2820
rect 2382 -2832 2388 -2826
rect 2382 -2838 2388 -2832
rect 2382 -2844 2388 -2838
rect 2382 -2850 2388 -2844
rect 2382 -2856 2388 -2850
rect 2382 -2862 2388 -2856
rect 2382 -2868 2388 -2862
rect 2382 -2874 2388 -2868
rect 2382 -2880 2388 -2874
rect 2382 -2886 2388 -2880
rect 2382 -2892 2388 -2886
rect 2382 -2898 2388 -2892
rect 2388 -126 2394 -120
rect 2388 -132 2394 -126
rect 2388 -138 2394 -132
rect 2388 -144 2394 -138
rect 2388 -150 2394 -144
rect 2388 -156 2394 -150
rect 2388 -162 2394 -156
rect 2388 -168 2394 -162
rect 2388 -174 2394 -168
rect 2388 -180 2394 -174
rect 2388 -186 2394 -180
rect 2388 -192 2394 -186
rect 2388 -198 2394 -192
rect 2388 -204 2394 -198
rect 2388 -210 2394 -204
rect 2388 -216 2394 -210
rect 2388 -222 2394 -216
rect 2388 -228 2394 -222
rect 2388 -234 2394 -228
rect 2388 -240 2394 -234
rect 2388 -246 2394 -240
rect 2388 -252 2394 -246
rect 2388 -258 2394 -252
rect 2388 -264 2394 -258
rect 2388 -270 2394 -264
rect 2388 -276 2394 -270
rect 2388 -282 2394 -276
rect 2388 -288 2394 -282
rect 2388 -294 2394 -288
rect 2388 -300 2394 -294
rect 2388 -306 2394 -300
rect 2388 -312 2394 -306
rect 2388 -318 2394 -312
rect 2388 -324 2394 -318
rect 2388 -330 2394 -324
rect 2388 -336 2394 -330
rect 2388 -342 2394 -336
rect 2388 -348 2394 -342
rect 2388 -354 2394 -348
rect 2388 -360 2394 -354
rect 2388 -366 2394 -360
rect 2388 -372 2394 -366
rect 2388 -378 2394 -372
rect 2388 -384 2394 -378
rect 2388 -390 2394 -384
rect 2388 -396 2394 -390
rect 2388 -402 2394 -396
rect 2388 -408 2394 -402
rect 2388 -414 2394 -408
rect 2388 -420 2394 -414
rect 2388 -426 2394 -420
rect 2388 -432 2394 -426
rect 2388 -438 2394 -432
rect 2388 -444 2394 -438
rect 2388 -450 2394 -444
rect 2388 -456 2394 -450
rect 2388 -462 2394 -456
rect 2388 -468 2394 -462
rect 2388 -474 2394 -468
rect 2388 -480 2394 -474
rect 2388 -486 2394 -480
rect 2388 -492 2394 -486
rect 2388 -498 2394 -492
rect 2388 -504 2394 -498
rect 2388 -510 2394 -504
rect 2388 -516 2394 -510
rect 2388 -522 2394 -516
rect 2388 -528 2394 -522
rect 2388 -534 2394 -528
rect 2388 -540 2394 -534
rect 2388 -546 2394 -540
rect 2388 -552 2394 -546
rect 2388 -558 2394 -552
rect 2388 -564 2394 -558
rect 2388 -570 2394 -564
rect 2388 -576 2394 -570
rect 2388 -582 2394 -576
rect 2388 -588 2394 -582
rect 2388 -594 2394 -588
rect 2388 -600 2394 -594
rect 2388 -606 2394 -600
rect 2388 -612 2394 -606
rect 2388 -618 2394 -612
rect 2388 -624 2394 -618
rect 2388 -630 2394 -624
rect 2388 -636 2394 -630
rect 2388 -642 2394 -636
rect 2388 -648 2394 -642
rect 2388 -654 2394 -648
rect 2388 -660 2394 -654
rect 2388 -666 2394 -660
rect 2388 -672 2394 -666
rect 2388 -678 2394 -672
rect 2388 -684 2394 -678
rect 2388 -690 2394 -684
rect 2388 -696 2394 -690
rect 2388 -702 2394 -696
rect 2388 -708 2394 -702
rect 2388 -714 2394 -708
rect 2388 -720 2394 -714
rect 2388 -726 2394 -720
rect 2388 -732 2394 -726
rect 2388 -1398 2394 -1392
rect 2388 -1404 2394 -1398
rect 2388 -1410 2394 -1404
rect 2388 -1416 2394 -1410
rect 2388 -1422 2394 -1416
rect 2388 -1428 2394 -1422
rect 2388 -1434 2394 -1428
rect 2388 -1440 2394 -1434
rect 2388 -1446 2394 -1440
rect 2388 -1452 2394 -1446
rect 2388 -1458 2394 -1452
rect 2388 -1464 2394 -1458
rect 2388 -1470 2394 -1464
rect 2388 -1476 2394 -1470
rect 2388 -1482 2394 -1476
rect 2388 -1488 2394 -1482
rect 2388 -1494 2394 -1488
rect 2388 -1500 2394 -1494
rect 2388 -1506 2394 -1500
rect 2388 -1512 2394 -1506
rect 2388 -1518 2394 -1512
rect 2388 -1524 2394 -1518
rect 2388 -1530 2394 -1524
rect 2388 -1536 2394 -1530
rect 2388 -1542 2394 -1536
rect 2388 -1548 2394 -1542
rect 2388 -1554 2394 -1548
rect 2388 -1560 2394 -1554
rect 2388 -1566 2394 -1560
rect 2388 -1572 2394 -1566
rect 2388 -1578 2394 -1572
rect 2388 -1584 2394 -1578
rect 2388 -1590 2394 -1584
rect 2388 -1596 2394 -1590
rect 2388 -1602 2394 -1596
rect 2388 -1608 2394 -1602
rect 2388 -1614 2394 -1608
rect 2388 -1620 2394 -1614
rect 2388 -1626 2394 -1620
rect 2388 -1632 2394 -1626
rect 2388 -1638 2394 -1632
rect 2388 -1644 2394 -1638
rect 2388 -1650 2394 -1644
rect 2388 -1656 2394 -1650
rect 2388 -1662 2394 -1656
rect 2388 -1668 2394 -1662
rect 2388 -1674 2394 -1668
rect 2388 -1680 2394 -1674
rect 2388 -1686 2394 -1680
rect 2388 -1692 2394 -1686
rect 2388 -1698 2394 -1692
rect 2388 -1704 2394 -1698
rect 2388 -1710 2394 -1704
rect 2388 -1716 2394 -1710
rect 2388 -1722 2394 -1716
rect 2388 -1728 2394 -1722
rect 2388 -1734 2394 -1728
rect 2388 -1740 2394 -1734
rect 2388 -1746 2394 -1740
rect 2388 -1752 2394 -1746
rect 2388 -1758 2394 -1752
rect 2388 -1764 2394 -1758
rect 2388 -1770 2394 -1764
rect 2388 -1776 2394 -1770
rect 2388 -1782 2394 -1776
rect 2388 -1788 2394 -1782
rect 2388 -1794 2394 -1788
rect 2388 -1800 2394 -1794
rect 2388 -1806 2394 -1800
rect 2388 -1812 2394 -1806
rect 2388 -1818 2394 -1812
rect 2388 -1824 2394 -1818
rect 2388 -1830 2394 -1824
rect 2388 -1836 2394 -1830
rect 2388 -1842 2394 -1836
rect 2388 -1848 2394 -1842
rect 2388 -1854 2394 -1848
rect 2388 -1860 2394 -1854
rect 2388 -1866 2394 -1860
rect 2388 -1872 2394 -1866
rect 2388 -1878 2394 -1872
rect 2388 -1884 2394 -1878
rect 2388 -1890 2394 -1884
rect 2388 -1896 2394 -1890
rect 2388 -1902 2394 -1896
rect 2388 -1908 2394 -1902
rect 2388 -1914 2394 -1908
rect 2388 -1920 2394 -1914
rect 2388 -1926 2394 -1920
rect 2388 -1932 2394 -1926
rect 2388 -1938 2394 -1932
rect 2388 -1944 2394 -1938
rect 2388 -1950 2394 -1944
rect 2388 -1956 2394 -1950
rect 2388 -1962 2394 -1956
rect 2388 -1968 2394 -1962
rect 2388 -1974 2394 -1968
rect 2388 -1980 2394 -1974
rect 2388 -1986 2394 -1980
rect 2388 -1992 2394 -1986
rect 2388 -1998 2394 -1992
rect 2388 -2004 2394 -1998
rect 2388 -2010 2394 -2004
rect 2388 -2016 2394 -2010
rect 2388 -2022 2394 -2016
rect 2388 -2028 2394 -2022
rect 2388 -2034 2394 -2028
rect 2388 -2040 2394 -2034
rect 2388 -2046 2394 -2040
rect 2388 -2052 2394 -2046
rect 2388 -2058 2394 -2052
rect 2388 -2064 2394 -2058
rect 2388 -2070 2394 -2064
rect 2388 -2076 2394 -2070
rect 2388 -2082 2394 -2076
rect 2388 -2088 2394 -2082
rect 2388 -2094 2394 -2088
rect 2388 -2100 2394 -2094
rect 2388 -2106 2394 -2100
rect 2388 -2112 2394 -2106
rect 2388 -2190 2394 -2184
rect 2388 -2196 2394 -2190
rect 2388 -2202 2394 -2196
rect 2388 -2208 2394 -2202
rect 2388 -2214 2394 -2208
rect 2388 -2220 2394 -2214
rect 2388 -2226 2394 -2220
rect 2388 -2232 2394 -2226
rect 2388 -2238 2394 -2232
rect 2388 -2244 2394 -2238
rect 2388 -2250 2394 -2244
rect 2388 -2256 2394 -2250
rect 2388 -2262 2394 -2256
rect 2388 -2268 2394 -2262
rect 2388 -2274 2394 -2268
rect 2388 -2280 2394 -2274
rect 2388 -2286 2394 -2280
rect 2388 -2292 2394 -2286
rect 2388 -2298 2394 -2292
rect 2388 -2304 2394 -2298
rect 2388 -2310 2394 -2304
rect 2388 -2316 2394 -2310
rect 2388 -2322 2394 -2316
rect 2388 -2328 2394 -2322
rect 2388 -2334 2394 -2328
rect 2388 -2340 2394 -2334
rect 2388 -2346 2394 -2340
rect 2388 -2352 2394 -2346
rect 2388 -2358 2394 -2352
rect 2388 -2364 2394 -2358
rect 2388 -2370 2394 -2364
rect 2388 -2376 2394 -2370
rect 2388 -2382 2394 -2376
rect 2388 -2388 2394 -2382
rect 2388 -2394 2394 -2388
rect 2388 -2400 2394 -2394
rect 2388 -2406 2394 -2400
rect 2388 -2412 2394 -2406
rect 2388 -2484 2394 -2478
rect 2388 -2490 2394 -2484
rect 2388 -2496 2394 -2490
rect 2388 -2502 2394 -2496
rect 2388 -2508 2394 -2502
rect 2388 -2514 2394 -2508
rect 2388 -2520 2394 -2514
rect 2388 -2526 2394 -2520
rect 2388 -2532 2394 -2526
rect 2388 -2538 2394 -2532
rect 2388 -2544 2394 -2538
rect 2388 -2550 2394 -2544
rect 2388 -2556 2394 -2550
rect 2388 -2562 2394 -2556
rect 2388 -2568 2394 -2562
rect 2388 -2574 2394 -2568
rect 2388 -2580 2394 -2574
rect 2388 -2586 2394 -2580
rect 2388 -2592 2394 -2586
rect 2388 -2598 2394 -2592
rect 2388 -2604 2394 -2598
rect 2388 -2610 2394 -2604
rect 2388 -2616 2394 -2610
rect 2388 -2622 2394 -2616
rect 2388 -2628 2394 -2622
rect 2388 -2634 2394 -2628
rect 2388 -2640 2394 -2634
rect 2388 -2646 2394 -2640
rect 2388 -2652 2394 -2646
rect 2388 -2658 2394 -2652
rect 2388 -2664 2394 -2658
rect 2388 -2670 2394 -2664
rect 2388 -2676 2394 -2670
rect 2388 -2682 2394 -2676
rect 2388 -2688 2394 -2682
rect 2388 -2694 2394 -2688
rect 2388 -2700 2394 -2694
rect 2388 -2706 2394 -2700
rect 2388 -2712 2394 -2706
rect 2388 -2718 2394 -2712
rect 2388 -2724 2394 -2718
rect 2388 -2730 2394 -2724
rect 2388 -2736 2394 -2730
rect 2388 -2742 2394 -2736
rect 2388 -2748 2394 -2742
rect 2388 -2754 2394 -2748
rect 2388 -2760 2394 -2754
rect 2388 -2766 2394 -2760
rect 2388 -2772 2394 -2766
rect 2388 -2778 2394 -2772
rect 2388 -2784 2394 -2778
rect 2388 -2790 2394 -2784
rect 2388 -2796 2394 -2790
rect 2388 -2802 2394 -2796
rect 2388 -2808 2394 -2802
rect 2388 -2814 2394 -2808
rect 2388 -2820 2394 -2814
rect 2388 -2826 2394 -2820
rect 2388 -2832 2394 -2826
rect 2388 -2838 2394 -2832
rect 2388 -2844 2394 -2838
rect 2388 -2850 2394 -2844
rect 2388 -2856 2394 -2850
rect 2388 -2862 2394 -2856
rect 2388 -2868 2394 -2862
rect 2388 -2874 2394 -2868
rect 2388 -2880 2394 -2874
rect 2388 -2886 2394 -2880
rect 2388 -2892 2394 -2886
rect 2394 -150 2400 -144
rect 2394 -156 2400 -150
rect 2394 -162 2400 -156
rect 2394 -168 2400 -162
rect 2394 -174 2400 -168
rect 2394 -180 2400 -174
rect 2394 -186 2400 -180
rect 2394 -192 2400 -186
rect 2394 -198 2400 -192
rect 2394 -204 2400 -198
rect 2394 -210 2400 -204
rect 2394 -216 2400 -210
rect 2394 -222 2400 -216
rect 2394 -228 2400 -222
rect 2394 -234 2400 -228
rect 2394 -240 2400 -234
rect 2394 -246 2400 -240
rect 2394 -252 2400 -246
rect 2394 -258 2400 -252
rect 2394 -264 2400 -258
rect 2394 -270 2400 -264
rect 2394 -276 2400 -270
rect 2394 -282 2400 -276
rect 2394 -288 2400 -282
rect 2394 -294 2400 -288
rect 2394 -300 2400 -294
rect 2394 -306 2400 -300
rect 2394 -312 2400 -306
rect 2394 -318 2400 -312
rect 2394 -324 2400 -318
rect 2394 -330 2400 -324
rect 2394 -336 2400 -330
rect 2394 -342 2400 -336
rect 2394 -348 2400 -342
rect 2394 -354 2400 -348
rect 2394 -360 2400 -354
rect 2394 -366 2400 -360
rect 2394 -372 2400 -366
rect 2394 -378 2400 -372
rect 2394 -384 2400 -378
rect 2394 -390 2400 -384
rect 2394 -396 2400 -390
rect 2394 -402 2400 -396
rect 2394 -408 2400 -402
rect 2394 -414 2400 -408
rect 2394 -420 2400 -414
rect 2394 -426 2400 -420
rect 2394 -432 2400 -426
rect 2394 -438 2400 -432
rect 2394 -444 2400 -438
rect 2394 -450 2400 -444
rect 2394 -456 2400 -450
rect 2394 -462 2400 -456
rect 2394 -468 2400 -462
rect 2394 -474 2400 -468
rect 2394 -480 2400 -474
rect 2394 -486 2400 -480
rect 2394 -492 2400 -486
rect 2394 -498 2400 -492
rect 2394 -504 2400 -498
rect 2394 -510 2400 -504
rect 2394 -516 2400 -510
rect 2394 -522 2400 -516
rect 2394 -528 2400 -522
rect 2394 -534 2400 -528
rect 2394 -540 2400 -534
rect 2394 -546 2400 -540
rect 2394 -552 2400 -546
rect 2394 -558 2400 -552
rect 2394 -564 2400 -558
rect 2394 -570 2400 -564
rect 2394 -576 2400 -570
rect 2394 -582 2400 -576
rect 2394 -588 2400 -582
rect 2394 -594 2400 -588
rect 2394 -600 2400 -594
rect 2394 -606 2400 -600
rect 2394 -612 2400 -606
rect 2394 -618 2400 -612
rect 2394 -624 2400 -618
rect 2394 -630 2400 -624
rect 2394 -636 2400 -630
rect 2394 -642 2400 -636
rect 2394 -648 2400 -642
rect 2394 -654 2400 -648
rect 2394 -660 2400 -654
rect 2394 -666 2400 -660
rect 2394 -672 2400 -666
rect 2394 -678 2400 -672
rect 2394 -684 2400 -678
rect 2394 -690 2400 -684
rect 2394 -696 2400 -690
rect 2394 -702 2400 -696
rect 2394 -708 2400 -702
rect 2394 -714 2400 -708
rect 2394 -1392 2400 -1386
rect 2394 -1398 2400 -1392
rect 2394 -1404 2400 -1398
rect 2394 -1410 2400 -1404
rect 2394 -1416 2400 -1410
rect 2394 -1422 2400 -1416
rect 2394 -1428 2400 -1422
rect 2394 -1434 2400 -1428
rect 2394 -1440 2400 -1434
rect 2394 -1446 2400 -1440
rect 2394 -1452 2400 -1446
rect 2394 -1458 2400 -1452
rect 2394 -1464 2400 -1458
rect 2394 -1470 2400 -1464
rect 2394 -1476 2400 -1470
rect 2394 -1482 2400 -1476
rect 2394 -1488 2400 -1482
rect 2394 -1494 2400 -1488
rect 2394 -1500 2400 -1494
rect 2394 -1506 2400 -1500
rect 2394 -1512 2400 -1506
rect 2394 -1518 2400 -1512
rect 2394 -1524 2400 -1518
rect 2394 -1530 2400 -1524
rect 2394 -1536 2400 -1530
rect 2394 -1542 2400 -1536
rect 2394 -1548 2400 -1542
rect 2394 -1554 2400 -1548
rect 2394 -1560 2400 -1554
rect 2394 -1566 2400 -1560
rect 2394 -1572 2400 -1566
rect 2394 -1578 2400 -1572
rect 2394 -1584 2400 -1578
rect 2394 -1590 2400 -1584
rect 2394 -1596 2400 -1590
rect 2394 -1602 2400 -1596
rect 2394 -1608 2400 -1602
rect 2394 -1614 2400 -1608
rect 2394 -1620 2400 -1614
rect 2394 -1626 2400 -1620
rect 2394 -1632 2400 -1626
rect 2394 -1638 2400 -1632
rect 2394 -1644 2400 -1638
rect 2394 -1650 2400 -1644
rect 2394 -1656 2400 -1650
rect 2394 -1662 2400 -1656
rect 2394 -1668 2400 -1662
rect 2394 -1674 2400 -1668
rect 2394 -1680 2400 -1674
rect 2394 -1686 2400 -1680
rect 2394 -1692 2400 -1686
rect 2394 -1698 2400 -1692
rect 2394 -1704 2400 -1698
rect 2394 -1710 2400 -1704
rect 2394 -1716 2400 -1710
rect 2394 -1722 2400 -1716
rect 2394 -1728 2400 -1722
rect 2394 -1734 2400 -1728
rect 2394 -1740 2400 -1734
rect 2394 -1746 2400 -1740
rect 2394 -1752 2400 -1746
rect 2394 -1758 2400 -1752
rect 2394 -1764 2400 -1758
rect 2394 -1770 2400 -1764
rect 2394 -1776 2400 -1770
rect 2394 -1782 2400 -1776
rect 2394 -1788 2400 -1782
rect 2394 -1794 2400 -1788
rect 2394 -1800 2400 -1794
rect 2394 -1806 2400 -1800
rect 2394 -1812 2400 -1806
rect 2394 -1818 2400 -1812
rect 2394 -1824 2400 -1818
rect 2394 -1830 2400 -1824
rect 2394 -1836 2400 -1830
rect 2394 -1842 2400 -1836
rect 2394 -1848 2400 -1842
rect 2394 -1854 2400 -1848
rect 2394 -1860 2400 -1854
rect 2394 -1866 2400 -1860
rect 2394 -1872 2400 -1866
rect 2394 -1878 2400 -1872
rect 2394 -1884 2400 -1878
rect 2394 -1890 2400 -1884
rect 2394 -1896 2400 -1890
rect 2394 -1902 2400 -1896
rect 2394 -1908 2400 -1902
rect 2394 -1914 2400 -1908
rect 2394 -1920 2400 -1914
rect 2394 -1926 2400 -1920
rect 2394 -1932 2400 -1926
rect 2394 -1938 2400 -1932
rect 2394 -1944 2400 -1938
rect 2394 -1950 2400 -1944
rect 2394 -1956 2400 -1950
rect 2394 -1962 2400 -1956
rect 2394 -1968 2400 -1962
rect 2394 -1974 2400 -1968
rect 2394 -1980 2400 -1974
rect 2394 -1986 2400 -1980
rect 2394 -1992 2400 -1986
rect 2394 -1998 2400 -1992
rect 2394 -2004 2400 -1998
rect 2394 -2010 2400 -2004
rect 2394 -2016 2400 -2010
rect 2394 -2022 2400 -2016
rect 2394 -2028 2400 -2022
rect 2394 -2034 2400 -2028
rect 2394 -2040 2400 -2034
rect 2394 -2046 2400 -2040
rect 2394 -2052 2400 -2046
rect 2394 -2058 2400 -2052
rect 2394 -2064 2400 -2058
rect 2394 -2070 2400 -2064
rect 2394 -2076 2400 -2070
rect 2394 -2082 2400 -2076
rect 2394 -2088 2400 -2082
rect 2394 -2094 2400 -2088
rect 2394 -2100 2400 -2094
rect 2394 -2106 2400 -2100
rect 2394 -2184 2400 -2178
rect 2394 -2190 2400 -2184
rect 2394 -2196 2400 -2190
rect 2394 -2202 2400 -2196
rect 2394 -2208 2400 -2202
rect 2394 -2214 2400 -2208
rect 2394 -2220 2400 -2214
rect 2394 -2226 2400 -2220
rect 2394 -2232 2400 -2226
rect 2394 -2238 2400 -2232
rect 2394 -2244 2400 -2238
rect 2394 -2250 2400 -2244
rect 2394 -2256 2400 -2250
rect 2394 -2262 2400 -2256
rect 2394 -2268 2400 -2262
rect 2394 -2274 2400 -2268
rect 2394 -2280 2400 -2274
rect 2394 -2286 2400 -2280
rect 2394 -2292 2400 -2286
rect 2394 -2298 2400 -2292
rect 2394 -2304 2400 -2298
rect 2394 -2310 2400 -2304
rect 2394 -2316 2400 -2310
rect 2394 -2322 2400 -2316
rect 2394 -2328 2400 -2322
rect 2394 -2334 2400 -2328
rect 2394 -2340 2400 -2334
rect 2394 -2346 2400 -2340
rect 2394 -2352 2400 -2346
rect 2394 -2358 2400 -2352
rect 2394 -2364 2400 -2358
rect 2394 -2370 2400 -2364
rect 2394 -2376 2400 -2370
rect 2394 -2382 2400 -2376
rect 2394 -2388 2400 -2382
rect 2394 -2394 2400 -2388
rect 2394 -2400 2400 -2394
rect 2394 -2406 2400 -2400
rect 2394 -2478 2400 -2472
rect 2394 -2484 2400 -2478
rect 2394 -2490 2400 -2484
rect 2394 -2496 2400 -2490
rect 2394 -2502 2400 -2496
rect 2394 -2508 2400 -2502
rect 2394 -2514 2400 -2508
rect 2394 -2520 2400 -2514
rect 2394 -2526 2400 -2520
rect 2394 -2532 2400 -2526
rect 2394 -2538 2400 -2532
rect 2394 -2544 2400 -2538
rect 2394 -2550 2400 -2544
rect 2394 -2556 2400 -2550
rect 2394 -2562 2400 -2556
rect 2394 -2568 2400 -2562
rect 2394 -2574 2400 -2568
rect 2394 -2580 2400 -2574
rect 2394 -2586 2400 -2580
rect 2394 -2592 2400 -2586
rect 2394 -2598 2400 -2592
rect 2394 -2604 2400 -2598
rect 2394 -2610 2400 -2604
rect 2394 -2616 2400 -2610
rect 2394 -2622 2400 -2616
rect 2394 -2628 2400 -2622
rect 2394 -2634 2400 -2628
rect 2394 -2640 2400 -2634
rect 2394 -2646 2400 -2640
rect 2394 -2652 2400 -2646
rect 2394 -2658 2400 -2652
rect 2394 -2664 2400 -2658
rect 2394 -2670 2400 -2664
rect 2394 -2676 2400 -2670
rect 2394 -2682 2400 -2676
rect 2394 -2688 2400 -2682
rect 2394 -2694 2400 -2688
rect 2394 -2700 2400 -2694
rect 2394 -2706 2400 -2700
rect 2394 -2712 2400 -2706
rect 2394 -2718 2400 -2712
rect 2394 -2724 2400 -2718
rect 2394 -2730 2400 -2724
rect 2394 -2736 2400 -2730
rect 2394 -2742 2400 -2736
rect 2394 -2748 2400 -2742
rect 2394 -2754 2400 -2748
rect 2394 -2760 2400 -2754
rect 2394 -2766 2400 -2760
rect 2394 -2772 2400 -2766
rect 2394 -2778 2400 -2772
rect 2394 -2784 2400 -2778
rect 2394 -2790 2400 -2784
rect 2394 -2796 2400 -2790
rect 2394 -2802 2400 -2796
rect 2394 -2808 2400 -2802
rect 2394 -2814 2400 -2808
rect 2394 -2820 2400 -2814
rect 2394 -2826 2400 -2820
rect 2394 -2832 2400 -2826
rect 2394 -2838 2400 -2832
rect 2394 -2844 2400 -2838
rect 2394 -2850 2400 -2844
rect 2394 -2856 2400 -2850
rect 2394 -2862 2400 -2856
rect 2394 -2868 2400 -2862
rect 2394 -2874 2400 -2868
rect 2394 -2880 2400 -2874
rect 2394 -2886 2400 -2880
rect 2394 -2892 2400 -2886
rect 2400 -174 2406 -168
rect 2400 -180 2406 -174
rect 2400 -186 2406 -180
rect 2400 -192 2406 -186
rect 2400 -198 2406 -192
rect 2400 -204 2406 -198
rect 2400 -210 2406 -204
rect 2400 -216 2406 -210
rect 2400 -222 2406 -216
rect 2400 -228 2406 -222
rect 2400 -234 2406 -228
rect 2400 -240 2406 -234
rect 2400 -246 2406 -240
rect 2400 -252 2406 -246
rect 2400 -258 2406 -252
rect 2400 -264 2406 -258
rect 2400 -270 2406 -264
rect 2400 -276 2406 -270
rect 2400 -282 2406 -276
rect 2400 -288 2406 -282
rect 2400 -294 2406 -288
rect 2400 -300 2406 -294
rect 2400 -306 2406 -300
rect 2400 -312 2406 -306
rect 2400 -318 2406 -312
rect 2400 -324 2406 -318
rect 2400 -330 2406 -324
rect 2400 -336 2406 -330
rect 2400 -342 2406 -336
rect 2400 -348 2406 -342
rect 2400 -354 2406 -348
rect 2400 -360 2406 -354
rect 2400 -366 2406 -360
rect 2400 -372 2406 -366
rect 2400 -378 2406 -372
rect 2400 -384 2406 -378
rect 2400 -390 2406 -384
rect 2400 -396 2406 -390
rect 2400 -402 2406 -396
rect 2400 -408 2406 -402
rect 2400 -414 2406 -408
rect 2400 -420 2406 -414
rect 2400 -426 2406 -420
rect 2400 -432 2406 -426
rect 2400 -438 2406 -432
rect 2400 -444 2406 -438
rect 2400 -450 2406 -444
rect 2400 -456 2406 -450
rect 2400 -462 2406 -456
rect 2400 -468 2406 -462
rect 2400 -474 2406 -468
rect 2400 -480 2406 -474
rect 2400 -486 2406 -480
rect 2400 -492 2406 -486
rect 2400 -498 2406 -492
rect 2400 -504 2406 -498
rect 2400 -510 2406 -504
rect 2400 -516 2406 -510
rect 2400 -522 2406 -516
rect 2400 -528 2406 -522
rect 2400 -534 2406 -528
rect 2400 -540 2406 -534
rect 2400 -546 2406 -540
rect 2400 -552 2406 -546
rect 2400 -558 2406 -552
rect 2400 -564 2406 -558
rect 2400 -570 2406 -564
rect 2400 -576 2406 -570
rect 2400 -582 2406 -576
rect 2400 -588 2406 -582
rect 2400 -594 2406 -588
rect 2400 -600 2406 -594
rect 2400 -606 2406 -600
rect 2400 -612 2406 -606
rect 2400 -618 2406 -612
rect 2400 -624 2406 -618
rect 2400 -630 2406 -624
rect 2400 -636 2406 -630
rect 2400 -642 2406 -636
rect 2400 -648 2406 -642
rect 2400 -654 2406 -648
rect 2400 -660 2406 -654
rect 2400 -666 2406 -660
rect 2400 -672 2406 -666
rect 2400 -678 2406 -672
rect 2400 -684 2406 -678
rect 2400 -690 2406 -684
rect 2400 -696 2406 -690
rect 2400 -1386 2406 -1380
rect 2400 -1392 2406 -1386
rect 2400 -1398 2406 -1392
rect 2400 -1404 2406 -1398
rect 2400 -1410 2406 -1404
rect 2400 -1416 2406 -1410
rect 2400 -1422 2406 -1416
rect 2400 -1428 2406 -1422
rect 2400 -1434 2406 -1428
rect 2400 -1440 2406 -1434
rect 2400 -1446 2406 -1440
rect 2400 -1452 2406 -1446
rect 2400 -1458 2406 -1452
rect 2400 -1464 2406 -1458
rect 2400 -1470 2406 -1464
rect 2400 -1476 2406 -1470
rect 2400 -1482 2406 -1476
rect 2400 -1488 2406 -1482
rect 2400 -1494 2406 -1488
rect 2400 -1500 2406 -1494
rect 2400 -1506 2406 -1500
rect 2400 -1512 2406 -1506
rect 2400 -1518 2406 -1512
rect 2400 -1524 2406 -1518
rect 2400 -1530 2406 -1524
rect 2400 -1536 2406 -1530
rect 2400 -1542 2406 -1536
rect 2400 -1548 2406 -1542
rect 2400 -1554 2406 -1548
rect 2400 -1560 2406 -1554
rect 2400 -1566 2406 -1560
rect 2400 -1572 2406 -1566
rect 2400 -1578 2406 -1572
rect 2400 -1584 2406 -1578
rect 2400 -1590 2406 -1584
rect 2400 -1596 2406 -1590
rect 2400 -1602 2406 -1596
rect 2400 -1608 2406 -1602
rect 2400 -1614 2406 -1608
rect 2400 -1620 2406 -1614
rect 2400 -1626 2406 -1620
rect 2400 -1632 2406 -1626
rect 2400 -1638 2406 -1632
rect 2400 -1644 2406 -1638
rect 2400 -1650 2406 -1644
rect 2400 -1656 2406 -1650
rect 2400 -1662 2406 -1656
rect 2400 -1668 2406 -1662
rect 2400 -1674 2406 -1668
rect 2400 -1680 2406 -1674
rect 2400 -1686 2406 -1680
rect 2400 -1692 2406 -1686
rect 2400 -1698 2406 -1692
rect 2400 -1704 2406 -1698
rect 2400 -1710 2406 -1704
rect 2400 -1716 2406 -1710
rect 2400 -1722 2406 -1716
rect 2400 -1728 2406 -1722
rect 2400 -1734 2406 -1728
rect 2400 -1740 2406 -1734
rect 2400 -1746 2406 -1740
rect 2400 -1752 2406 -1746
rect 2400 -1758 2406 -1752
rect 2400 -1764 2406 -1758
rect 2400 -1770 2406 -1764
rect 2400 -1776 2406 -1770
rect 2400 -1782 2406 -1776
rect 2400 -1788 2406 -1782
rect 2400 -1794 2406 -1788
rect 2400 -1800 2406 -1794
rect 2400 -1806 2406 -1800
rect 2400 -1812 2406 -1806
rect 2400 -1818 2406 -1812
rect 2400 -1824 2406 -1818
rect 2400 -1830 2406 -1824
rect 2400 -1836 2406 -1830
rect 2400 -1842 2406 -1836
rect 2400 -1848 2406 -1842
rect 2400 -1854 2406 -1848
rect 2400 -1860 2406 -1854
rect 2400 -1866 2406 -1860
rect 2400 -1872 2406 -1866
rect 2400 -1878 2406 -1872
rect 2400 -1884 2406 -1878
rect 2400 -1890 2406 -1884
rect 2400 -1896 2406 -1890
rect 2400 -1902 2406 -1896
rect 2400 -1908 2406 -1902
rect 2400 -1914 2406 -1908
rect 2400 -1920 2406 -1914
rect 2400 -1926 2406 -1920
rect 2400 -1932 2406 -1926
rect 2400 -1938 2406 -1932
rect 2400 -1944 2406 -1938
rect 2400 -1950 2406 -1944
rect 2400 -1956 2406 -1950
rect 2400 -1962 2406 -1956
rect 2400 -1968 2406 -1962
rect 2400 -1974 2406 -1968
rect 2400 -1980 2406 -1974
rect 2400 -1986 2406 -1980
rect 2400 -1992 2406 -1986
rect 2400 -1998 2406 -1992
rect 2400 -2004 2406 -1998
rect 2400 -2010 2406 -2004
rect 2400 -2016 2406 -2010
rect 2400 -2022 2406 -2016
rect 2400 -2028 2406 -2022
rect 2400 -2034 2406 -2028
rect 2400 -2040 2406 -2034
rect 2400 -2046 2406 -2040
rect 2400 -2052 2406 -2046
rect 2400 -2058 2406 -2052
rect 2400 -2064 2406 -2058
rect 2400 -2070 2406 -2064
rect 2400 -2076 2406 -2070
rect 2400 -2082 2406 -2076
rect 2400 -2088 2406 -2082
rect 2400 -2094 2406 -2088
rect 2400 -2100 2406 -2094
rect 2400 -2178 2406 -2172
rect 2400 -2184 2406 -2178
rect 2400 -2190 2406 -2184
rect 2400 -2196 2406 -2190
rect 2400 -2202 2406 -2196
rect 2400 -2208 2406 -2202
rect 2400 -2214 2406 -2208
rect 2400 -2220 2406 -2214
rect 2400 -2226 2406 -2220
rect 2400 -2232 2406 -2226
rect 2400 -2238 2406 -2232
rect 2400 -2244 2406 -2238
rect 2400 -2250 2406 -2244
rect 2400 -2256 2406 -2250
rect 2400 -2262 2406 -2256
rect 2400 -2268 2406 -2262
rect 2400 -2274 2406 -2268
rect 2400 -2280 2406 -2274
rect 2400 -2286 2406 -2280
rect 2400 -2292 2406 -2286
rect 2400 -2298 2406 -2292
rect 2400 -2304 2406 -2298
rect 2400 -2310 2406 -2304
rect 2400 -2316 2406 -2310
rect 2400 -2322 2406 -2316
rect 2400 -2328 2406 -2322
rect 2400 -2334 2406 -2328
rect 2400 -2340 2406 -2334
rect 2400 -2346 2406 -2340
rect 2400 -2352 2406 -2346
rect 2400 -2358 2406 -2352
rect 2400 -2364 2406 -2358
rect 2400 -2370 2406 -2364
rect 2400 -2376 2406 -2370
rect 2400 -2382 2406 -2376
rect 2400 -2388 2406 -2382
rect 2400 -2394 2406 -2388
rect 2400 -2400 2406 -2394
rect 2400 -2406 2406 -2400
rect 2400 -2478 2406 -2472
rect 2400 -2484 2406 -2478
rect 2400 -2490 2406 -2484
rect 2400 -2496 2406 -2490
rect 2400 -2502 2406 -2496
rect 2400 -2508 2406 -2502
rect 2400 -2514 2406 -2508
rect 2400 -2520 2406 -2514
rect 2400 -2526 2406 -2520
rect 2400 -2532 2406 -2526
rect 2400 -2538 2406 -2532
rect 2400 -2544 2406 -2538
rect 2400 -2550 2406 -2544
rect 2400 -2556 2406 -2550
rect 2400 -2562 2406 -2556
rect 2400 -2568 2406 -2562
rect 2400 -2574 2406 -2568
rect 2400 -2580 2406 -2574
rect 2400 -2586 2406 -2580
rect 2400 -2592 2406 -2586
rect 2400 -2598 2406 -2592
rect 2400 -2604 2406 -2598
rect 2400 -2610 2406 -2604
rect 2400 -2616 2406 -2610
rect 2400 -2622 2406 -2616
rect 2400 -2628 2406 -2622
rect 2400 -2634 2406 -2628
rect 2400 -2640 2406 -2634
rect 2400 -2646 2406 -2640
rect 2400 -2652 2406 -2646
rect 2400 -2658 2406 -2652
rect 2400 -2664 2406 -2658
rect 2400 -2670 2406 -2664
rect 2400 -2676 2406 -2670
rect 2400 -2682 2406 -2676
rect 2400 -2688 2406 -2682
rect 2400 -2694 2406 -2688
rect 2400 -2700 2406 -2694
rect 2400 -2706 2406 -2700
rect 2400 -2712 2406 -2706
rect 2400 -2718 2406 -2712
rect 2400 -2724 2406 -2718
rect 2400 -2730 2406 -2724
rect 2400 -2736 2406 -2730
rect 2400 -2742 2406 -2736
rect 2400 -2748 2406 -2742
rect 2400 -2754 2406 -2748
rect 2400 -2760 2406 -2754
rect 2400 -2766 2406 -2760
rect 2400 -2772 2406 -2766
rect 2400 -2778 2406 -2772
rect 2400 -2784 2406 -2778
rect 2400 -2790 2406 -2784
rect 2400 -2796 2406 -2790
rect 2400 -2802 2406 -2796
rect 2400 -2808 2406 -2802
rect 2400 -2814 2406 -2808
rect 2400 -2820 2406 -2814
rect 2400 -2826 2406 -2820
rect 2400 -2832 2406 -2826
rect 2400 -2838 2406 -2832
rect 2400 -2844 2406 -2838
rect 2400 -2850 2406 -2844
rect 2400 -2856 2406 -2850
rect 2400 -2862 2406 -2856
rect 2400 -2868 2406 -2862
rect 2400 -2874 2406 -2868
rect 2400 -2880 2406 -2874
rect 2400 -2886 2406 -2880
rect 2406 -198 2412 -192
rect 2406 -204 2412 -198
rect 2406 -210 2412 -204
rect 2406 -216 2412 -210
rect 2406 -222 2412 -216
rect 2406 -228 2412 -222
rect 2406 -234 2412 -228
rect 2406 -240 2412 -234
rect 2406 -246 2412 -240
rect 2406 -252 2412 -246
rect 2406 -258 2412 -252
rect 2406 -264 2412 -258
rect 2406 -270 2412 -264
rect 2406 -276 2412 -270
rect 2406 -282 2412 -276
rect 2406 -288 2412 -282
rect 2406 -294 2412 -288
rect 2406 -300 2412 -294
rect 2406 -306 2412 -300
rect 2406 -312 2412 -306
rect 2406 -318 2412 -312
rect 2406 -324 2412 -318
rect 2406 -330 2412 -324
rect 2406 -336 2412 -330
rect 2406 -342 2412 -336
rect 2406 -348 2412 -342
rect 2406 -354 2412 -348
rect 2406 -360 2412 -354
rect 2406 -366 2412 -360
rect 2406 -372 2412 -366
rect 2406 -378 2412 -372
rect 2406 -384 2412 -378
rect 2406 -390 2412 -384
rect 2406 -396 2412 -390
rect 2406 -402 2412 -396
rect 2406 -408 2412 -402
rect 2406 -414 2412 -408
rect 2406 -420 2412 -414
rect 2406 -426 2412 -420
rect 2406 -432 2412 -426
rect 2406 -438 2412 -432
rect 2406 -444 2412 -438
rect 2406 -450 2412 -444
rect 2406 -456 2412 -450
rect 2406 -462 2412 -456
rect 2406 -468 2412 -462
rect 2406 -474 2412 -468
rect 2406 -480 2412 -474
rect 2406 -486 2412 -480
rect 2406 -492 2412 -486
rect 2406 -498 2412 -492
rect 2406 -504 2412 -498
rect 2406 -510 2412 -504
rect 2406 -516 2412 -510
rect 2406 -522 2412 -516
rect 2406 -528 2412 -522
rect 2406 -534 2412 -528
rect 2406 -540 2412 -534
rect 2406 -546 2412 -540
rect 2406 -552 2412 -546
rect 2406 -558 2412 -552
rect 2406 -564 2412 -558
rect 2406 -570 2412 -564
rect 2406 -576 2412 -570
rect 2406 -582 2412 -576
rect 2406 -588 2412 -582
rect 2406 -594 2412 -588
rect 2406 -600 2412 -594
rect 2406 -606 2412 -600
rect 2406 -612 2412 -606
rect 2406 -618 2412 -612
rect 2406 -624 2412 -618
rect 2406 -630 2412 -624
rect 2406 -636 2412 -630
rect 2406 -642 2412 -636
rect 2406 -648 2412 -642
rect 2406 -654 2412 -648
rect 2406 -660 2412 -654
rect 2406 -666 2412 -660
rect 2406 -672 2412 -666
rect 2406 -1380 2412 -1374
rect 2406 -1386 2412 -1380
rect 2406 -1392 2412 -1386
rect 2406 -1398 2412 -1392
rect 2406 -1404 2412 -1398
rect 2406 -1410 2412 -1404
rect 2406 -1416 2412 -1410
rect 2406 -1422 2412 -1416
rect 2406 -1428 2412 -1422
rect 2406 -1434 2412 -1428
rect 2406 -1440 2412 -1434
rect 2406 -1446 2412 -1440
rect 2406 -1452 2412 -1446
rect 2406 -1458 2412 -1452
rect 2406 -1464 2412 -1458
rect 2406 -1470 2412 -1464
rect 2406 -1476 2412 -1470
rect 2406 -1482 2412 -1476
rect 2406 -1488 2412 -1482
rect 2406 -1494 2412 -1488
rect 2406 -1500 2412 -1494
rect 2406 -1506 2412 -1500
rect 2406 -1512 2412 -1506
rect 2406 -1518 2412 -1512
rect 2406 -1524 2412 -1518
rect 2406 -1530 2412 -1524
rect 2406 -1536 2412 -1530
rect 2406 -1542 2412 -1536
rect 2406 -1548 2412 -1542
rect 2406 -1554 2412 -1548
rect 2406 -1560 2412 -1554
rect 2406 -1566 2412 -1560
rect 2406 -1572 2412 -1566
rect 2406 -1578 2412 -1572
rect 2406 -1584 2412 -1578
rect 2406 -1590 2412 -1584
rect 2406 -1596 2412 -1590
rect 2406 -1602 2412 -1596
rect 2406 -1608 2412 -1602
rect 2406 -1614 2412 -1608
rect 2406 -1620 2412 -1614
rect 2406 -1626 2412 -1620
rect 2406 -1632 2412 -1626
rect 2406 -1638 2412 -1632
rect 2406 -1644 2412 -1638
rect 2406 -1650 2412 -1644
rect 2406 -1656 2412 -1650
rect 2406 -1662 2412 -1656
rect 2406 -1668 2412 -1662
rect 2406 -1674 2412 -1668
rect 2406 -1680 2412 -1674
rect 2406 -1686 2412 -1680
rect 2406 -1692 2412 -1686
rect 2406 -1698 2412 -1692
rect 2406 -1704 2412 -1698
rect 2406 -1710 2412 -1704
rect 2406 -1716 2412 -1710
rect 2406 -1722 2412 -1716
rect 2406 -1728 2412 -1722
rect 2406 -1734 2412 -1728
rect 2406 -1740 2412 -1734
rect 2406 -1746 2412 -1740
rect 2406 -1752 2412 -1746
rect 2406 -1758 2412 -1752
rect 2406 -1764 2412 -1758
rect 2406 -1770 2412 -1764
rect 2406 -1776 2412 -1770
rect 2406 -1782 2412 -1776
rect 2406 -1788 2412 -1782
rect 2406 -1794 2412 -1788
rect 2406 -1800 2412 -1794
rect 2406 -1806 2412 -1800
rect 2406 -1812 2412 -1806
rect 2406 -1818 2412 -1812
rect 2406 -1824 2412 -1818
rect 2406 -1830 2412 -1824
rect 2406 -1836 2412 -1830
rect 2406 -1842 2412 -1836
rect 2406 -1848 2412 -1842
rect 2406 -1854 2412 -1848
rect 2406 -1860 2412 -1854
rect 2406 -1866 2412 -1860
rect 2406 -1872 2412 -1866
rect 2406 -1878 2412 -1872
rect 2406 -1884 2412 -1878
rect 2406 -1890 2412 -1884
rect 2406 -1896 2412 -1890
rect 2406 -1902 2412 -1896
rect 2406 -1908 2412 -1902
rect 2406 -1914 2412 -1908
rect 2406 -1920 2412 -1914
rect 2406 -1926 2412 -1920
rect 2406 -1932 2412 -1926
rect 2406 -1938 2412 -1932
rect 2406 -1944 2412 -1938
rect 2406 -1950 2412 -1944
rect 2406 -1956 2412 -1950
rect 2406 -1962 2412 -1956
rect 2406 -1968 2412 -1962
rect 2406 -1974 2412 -1968
rect 2406 -1980 2412 -1974
rect 2406 -1986 2412 -1980
rect 2406 -1992 2412 -1986
rect 2406 -1998 2412 -1992
rect 2406 -2004 2412 -1998
rect 2406 -2010 2412 -2004
rect 2406 -2016 2412 -2010
rect 2406 -2022 2412 -2016
rect 2406 -2028 2412 -2022
rect 2406 -2034 2412 -2028
rect 2406 -2040 2412 -2034
rect 2406 -2046 2412 -2040
rect 2406 -2052 2412 -2046
rect 2406 -2058 2412 -2052
rect 2406 -2064 2412 -2058
rect 2406 -2070 2412 -2064
rect 2406 -2076 2412 -2070
rect 2406 -2082 2412 -2076
rect 2406 -2088 2412 -2082
rect 2406 -2172 2412 -2166
rect 2406 -2178 2412 -2172
rect 2406 -2184 2412 -2178
rect 2406 -2190 2412 -2184
rect 2406 -2196 2412 -2190
rect 2406 -2202 2412 -2196
rect 2406 -2208 2412 -2202
rect 2406 -2214 2412 -2208
rect 2406 -2220 2412 -2214
rect 2406 -2226 2412 -2220
rect 2406 -2232 2412 -2226
rect 2406 -2238 2412 -2232
rect 2406 -2244 2412 -2238
rect 2406 -2250 2412 -2244
rect 2406 -2256 2412 -2250
rect 2406 -2262 2412 -2256
rect 2406 -2268 2412 -2262
rect 2406 -2274 2412 -2268
rect 2406 -2280 2412 -2274
rect 2406 -2286 2412 -2280
rect 2406 -2292 2412 -2286
rect 2406 -2298 2412 -2292
rect 2406 -2304 2412 -2298
rect 2406 -2310 2412 -2304
rect 2406 -2316 2412 -2310
rect 2406 -2322 2412 -2316
rect 2406 -2328 2412 -2322
rect 2406 -2334 2412 -2328
rect 2406 -2340 2412 -2334
rect 2406 -2346 2412 -2340
rect 2406 -2352 2412 -2346
rect 2406 -2358 2412 -2352
rect 2406 -2364 2412 -2358
rect 2406 -2370 2412 -2364
rect 2406 -2376 2412 -2370
rect 2406 -2382 2412 -2376
rect 2406 -2388 2412 -2382
rect 2406 -2394 2412 -2388
rect 2406 -2400 2412 -2394
rect 2406 -2406 2412 -2400
rect 2406 -2478 2412 -2472
rect 2406 -2484 2412 -2478
rect 2406 -2490 2412 -2484
rect 2406 -2496 2412 -2490
rect 2406 -2502 2412 -2496
rect 2406 -2508 2412 -2502
rect 2406 -2514 2412 -2508
rect 2406 -2520 2412 -2514
rect 2406 -2526 2412 -2520
rect 2406 -2532 2412 -2526
rect 2406 -2538 2412 -2532
rect 2406 -2544 2412 -2538
rect 2406 -2550 2412 -2544
rect 2406 -2556 2412 -2550
rect 2406 -2562 2412 -2556
rect 2406 -2568 2412 -2562
rect 2406 -2574 2412 -2568
rect 2406 -2580 2412 -2574
rect 2406 -2586 2412 -2580
rect 2406 -2592 2412 -2586
rect 2406 -2598 2412 -2592
rect 2406 -2604 2412 -2598
rect 2406 -2610 2412 -2604
rect 2406 -2616 2412 -2610
rect 2406 -2622 2412 -2616
rect 2406 -2628 2412 -2622
rect 2406 -2634 2412 -2628
rect 2406 -2640 2412 -2634
rect 2406 -2646 2412 -2640
rect 2406 -2652 2412 -2646
rect 2406 -2658 2412 -2652
rect 2406 -2664 2412 -2658
rect 2406 -2670 2412 -2664
rect 2406 -2676 2412 -2670
rect 2406 -2682 2412 -2676
rect 2406 -2688 2412 -2682
rect 2406 -2694 2412 -2688
rect 2406 -2700 2412 -2694
rect 2406 -2706 2412 -2700
rect 2406 -2712 2412 -2706
rect 2406 -2718 2412 -2712
rect 2406 -2724 2412 -2718
rect 2406 -2730 2412 -2724
rect 2406 -2736 2412 -2730
rect 2406 -2742 2412 -2736
rect 2406 -2748 2412 -2742
rect 2406 -2754 2412 -2748
rect 2406 -2760 2412 -2754
rect 2406 -2766 2412 -2760
rect 2406 -2772 2412 -2766
rect 2406 -2778 2412 -2772
rect 2406 -2784 2412 -2778
rect 2406 -2790 2412 -2784
rect 2406 -2796 2412 -2790
rect 2406 -2802 2412 -2796
rect 2406 -2808 2412 -2802
rect 2406 -2814 2412 -2808
rect 2406 -2820 2412 -2814
rect 2406 -2826 2412 -2820
rect 2406 -2832 2412 -2826
rect 2406 -2838 2412 -2832
rect 2406 -2844 2412 -2838
rect 2406 -2850 2412 -2844
rect 2406 -2856 2412 -2850
rect 2406 -2862 2412 -2856
rect 2406 -2868 2412 -2862
rect 2406 -2874 2412 -2868
rect 2406 -2880 2412 -2874
rect 2412 -222 2418 -216
rect 2412 -228 2418 -222
rect 2412 -234 2418 -228
rect 2412 -240 2418 -234
rect 2412 -246 2418 -240
rect 2412 -252 2418 -246
rect 2412 -258 2418 -252
rect 2412 -264 2418 -258
rect 2412 -270 2418 -264
rect 2412 -276 2418 -270
rect 2412 -282 2418 -276
rect 2412 -288 2418 -282
rect 2412 -294 2418 -288
rect 2412 -300 2418 -294
rect 2412 -306 2418 -300
rect 2412 -312 2418 -306
rect 2412 -318 2418 -312
rect 2412 -324 2418 -318
rect 2412 -330 2418 -324
rect 2412 -336 2418 -330
rect 2412 -342 2418 -336
rect 2412 -348 2418 -342
rect 2412 -354 2418 -348
rect 2412 -360 2418 -354
rect 2412 -366 2418 -360
rect 2412 -372 2418 -366
rect 2412 -378 2418 -372
rect 2412 -384 2418 -378
rect 2412 -390 2418 -384
rect 2412 -396 2418 -390
rect 2412 -402 2418 -396
rect 2412 -408 2418 -402
rect 2412 -414 2418 -408
rect 2412 -420 2418 -414
rect 2412 -426 2418 -420
rect 2412 -432 2418 -426
rect 2412 -438 2418 -432
rect 2412 -444 2418 -438
rect 2412 -450 2418 -444
rect 2412 -456 2418 -450
rect 2412 -462 2418 -456
rect 2412 -468 2418 -462
rect 2412 -474 2418 -468
rect 2412 -480 2418 -474
rect 2412 -486 2418 -480
rect 2412 -492 2418 -486
rect 2412 -498 2418 -492
rect 2412 -504 2418 -498
rect 2412 -510 2418 -504
rect 2412 -516 2418 -510
rect 2412 -522 2418 -516
rect 2412 -528 2418 -522
rect 2412 -534 2418 -528
rect 2412 -540 2418 -534
rect 2412 -546 2418 -540
rect 2412 -552 2418 -546
rect 2412 -558 2418 -552
rect 2412 -564 2418 -558
rect 2412 -570 2418 -564
rect 2412 -576 2418 -570
rect 2412 -582 2418 -576
rect 2412 -588 2418 -582
rect 2412 -594 2418 -588
rect 2412 -600 2418 -594
rect 2412 -606 2418 -600
rect 2412 -612 2418 -606
rect 2412 -618 2418 -612
rect 2412 -624 2418 -618
rect 2412 -630 2418 -624
rect 2412 -636 2418 -630
rect 2412 -642 2418 -636
rect 2412 -648 2418 -642
rect 2412 -1374 2418 -1368
rect 2412 -1380 2418 -1374
rect 2412 -1386 2418 -1380
rect 2412 -1392 2418 -1386
rect 2412 -1398 2418 -1392
rect 2412 -1404 2418 -1398
rect 2412 -1410 2418 -1404
rect 2412 -1416 2418 -1410
rect 2412 -1422 2418 -1416
rect 2412 -1428 2418 -1422
rect 2412 -1434 2418 -1428
rect 2412 -1440 2418 -1434
rect 2412 -1446 2418 -1440
rect 2412 -1452 2418 -1446
rect 2412 -1458 2418 -1452
rect 2412 -1464 2418 -1458
rect 2412 -1470 2418 -1464
rect 2412 -1476 2418 -1470
rect 2412 -1482 2418 -1476
rect 2412 -1488 2418 -1482
rect 2412 -1494 2418 -1488
rect 2412 -1500 2418 -1494
rect 2412 -1506 2418 -1500
rect 2412 -1512 2418 -1506
rect 2412 -1518 2418 -1512
rect 2412 -1524 2418 -1518
rect 2412 -1530 2418 -1524
rect 2412 -1536 2418 -1530
rect 2412 -1542 2418 -1536
rect 2412 -1548 2418 -1542
rect 2412 -1554 2418 -1548
rect 2412 -1560 2418 -1554
rect 2412 -1566 2418 -1560
rect 2412 -1572 2418 -1566
rect 2412 -1578 2418 -1572
rect 2412 -1584 2418 -1578
rect 2412 -1590 2418 -1584
rect 2412 -1596 2418 -1590
rect 2412 -1602 2418 -1596
rect 2412 -1608 2418 -1602
rect 2412 -1614 2418 -1608
rect 2412 -1620 2418 -1614
rect 2412 -1626 2418 -1620
rect 2412 -1632 2418 -1626
rect 2412 -1638 2418 -1632
rect 2412 -1644 2418 -1638
rect 2412 -1650 2418 -1644
rect 2412 -1656 2418 -1650
rect 2412 -1662 2418 -1656
rect 2412 -1668 2418 -1662
rect 2412 -1674 2418 -1668
rect 2412 -1680 2418 -1674
rect 2412 -1686 2418 -1680
rect 2412 -1692 2418 -1686
rect 2412 -1698 2418 -1692
rect 2412 -1704 2418 -1698
rect 2412 -1710 2418 -1704
rect 2412 -1716 2418 -1710
rect 2412 -1722 2418 -1716
rect 2412 -1728 2418 -1722
rect 2412 -1734 2418 -1728
rect 2412 -1740 2418 -1734
rect 2412 -1746 2418 -1740
rect 2412 -1752 2418 -1746
rect 2412 -1758 2418 -1752
rect 2412 -1764 2418 -1758
rect 2412 -1770 2418 -1764
rect 2412 -1776 2418 -1770
rect 2412 -1782 2418 -1776
rect 2412 -1788 2418 -1782
rect 2412 -1794 2418 -1788
rect 2412 -1800 2418 -1794
rect 2412 -1806 2418 -1800
rect 2412 -1812 2418 -1806
rect 2412 -1818 2418 -1812
rect 2412 -1824 2418 -1818
rect 2412 -1830 2418 -1824
rect 2412 -1836 2418 -1830
rect 2412 -1842 2418 -1836
rect 2412 -1848 2418 -1842
rect 2412 -1854 2418 -1848
rect 2412 -1860 2418 -1854
rect 2412 -1866 2418 -1860
rect 2412 -1872 2418 -1866
rect 2412 -1878 2418 -1872
rect 2412 -1884 2418 -1878
rect 2412 -1890 2418 -1884
rect 2412 -1896 2418 -1890
rect 2412 -1902 2418 -1896
rect 2412 -1908 2418 -1902
rect 2412 -1914 2418 -1908
rect 2412 -1920 2418 -1914
rect 2412 -1926 2418 -1920
rect 2412 -1932 2418 -1926
rect 2412 -1938 2418 -1932
rect 2412 -1944 2418 -1938
rect 2412 -1950 2418 -1944
rect 2412 -1956 2418 -1950
rect 2412 -1962 2418 -1956
rect 2412 -1968 2418 -1962
rect 2412 -1974 2418 -1968
rect 2412 -1980 2418 -1974
rect 2412 -1986 2418 -1980
rect 2412 -1992 2418 -1986
rect 2412 -1998 2418 -1992
rect 2412 -2004 2418 -1998
rect 2412 -2010 2418 -2004
rect 2412 -2016 2418 -2010
rect 2412 -2022 2418 -2016
rect 2412 -2028 2418 -2022
rect 2412 -2034 2418 -2028
rect 2412 -2040 2418 -2034
rect 2412 -2046 2418 -2040
rect 2412 -2052 2418 -2046
rect 2412 -2058 2418 -2052
rect 2412 -2064 2418 -2058
rect 2412 -2070 2418 -2064
rect 2412 -2076 2418 -2070
rect 2412 -2082 2418 -2076
rect 2412 -2166 2418 -2160
rect 2412 -2172 2418 -2166
rect 2412 -2178 2418 -2172
rect 2412 -2184 2418 -2178
rect 2412 -2190 2418 -2184
rect 2412 -2196 2418 -2190
rect 2412 -2202 2418 -2196
rect 2412 -2208 2418 -2202
rect 2412 -2214 2418 -2208
rect 2412 -2220 2418 -2214
rect 2412 -2226 2418 -2220
rect 2412 -2232 2418 -2226
rect 2412 -2238 2418 -2232
rect 2412 -2244 2418 -2238
rect 2412 -2250 2418 -2244
rect 2412 -2256 2418 -2250
rect 2412 -2262 2418 -2256
rect 2412 -2268 2418 -2262
rect 2412 -2274 2418 -2268
rect 2412 -2280 2418 -2274
rect 2412 -2286 2418 -2280
rect 2412 -2292 2418 -2286
rect 2412 -2298 2418 -2292
rect 2412 -2304 2418 -2298
rect 2412 -2310 2418 -2304
rect 2412 -2316 2418 -2310
rect 2412 -2322 2418 -2316
rect 2412 -2328 2418 -2322
rect 2412 -2334 2418 -2328
rect 2412 -2340 2418 -2334
rect 2412 -2346 2418 -2340
rect 2412 -2352 2418 -2346
rect 2412 -2358 2418 -2352
rect 2412 -2364 2418 -2358
rect 2412 -2370 2418 -2364
rect 2412 -2376 2418 -2370
rect 2412 -2382 2418 -2376
rect 2412 -2388 2418 -2382
rect 2412 -2394 2418 -2388
rect 2412 -2400 2418 -2394
rect 2412 -2472 2418 -2466
rect 2412 -2478 2418 -2472
rect 2412 -2484 2418 -2478
rect 2412 -2490 2418 -2484
rect 2412 -2496 2418 -2490
rect 2412 -2502 2418 -2496
rect 2412 -2508 2418 -2502
rect 2412 -2514 2418 -2508
rect 2412 -2520 2418 -2514
rect 2412 -2526 2418 -2520
rect 2412 -2532 2418 -2526
rect 2412 -2538 2418 -2532
rect 2412 -2544 2418 -2538
rect 2412 -2550 2418 -2544
rect 2412 -2556 2418 -2550
rect 2412 -2562 2418 -2556
rect 2412 -2568 2418 -2562
rect 2412 -2574 2418 -2568
rect 2412 -2580 2418 -2574
rect 2412 -2586 2418 -2580
rect 2412 -2592 2418 -2586
rect 2412 -2598 2418 -2592
rect 2412 -2604 2418 -2598
rect 2412 -2610 2418 -2604
rect 2412 -2616 2418 -2610
rect 2412 -2622 2418 -2616
rect 2412 -2628 2418 -2622
rect 2412 -2634 2418 -2628
rect 2412 -2640 2418 -2634
rect 2412 -2646 2418 -2640
rect 2412 -2652 2418 -2646
rect 2412 -2658 2418 -2652
rect 2412 -2664 2418 -2658
rect 2412 -2670 2418 -2664
rect 2412 -2676 2418 -2670
rect 2412 -2682 2418 -2676
rect 2412 -2688 2418 -2682
rect 2412 -2694 2418 -2688
rect 2412 -2700 2418 -2694
rect 2412 -2706 2418 -2700
rect 2412 -2712 2418 -2706
rect 2412 -2718 2418 -2712
rect 2412 -2724 2418 -2718
rect 2412 -2730 2418 -2724
rect 2412 -2736 2418 -2730
rect 2412 -2742 2418 -2736
rect 2412 -2748 2418 -2742
rect 2412 -2754 2418 -2748
rect 2412 -2760 2418 -2754
rect 2412 -2766 2418 -2760
rect 2412 -2772 2418 -2766
rect 2412 -2778 2418 -2772
rect 2412 -2784 2418 -2778
rect 2412 -2790 2418 -2784
rect 2412 -2796 2418 -2790
rect 2412 -2802 2418 -2796
rect 2412 -2808 2418 -2802
rect 2412 -2814 2418 -2808
rect 2412 -2820 2418 -2814
rect 2412 -2826 2418 -2820
rect 2412 -2832 2418 -2826
rect 2412 -2838 2418 -2832
rect 2412 -2844 2418 -2838
rect 2412 -2850 2418 -2844
rect 2412 -2856 2418 -2850
rect 2412 -2862 2418 -2856
rect 2412 -2868 2418 -2862
rect 2412 -2874 2418 -2868
rect 2412 -2880 2418 -2874
rect 2418 -252 2424 -246
rect 2418 -258 2424 -252
rect 2418 -264 2424 -258
rect 2418 -270 2424 -264
rect 2418 -276 2424 -270
rect 2418 -282 2424 -276
rect 2418 -288 2424 -282
rect 2418 -294 2424 -288
rect 2418 -300 2424 -294
rect 2418 -306 2424 -300
rect 2418 -312 2424 -306
rect 2418 -318 2424 -312
rect 2418 -324 2424 -318
rect 2418 -330 2424 -324
rect 2418 -336 2424 -330
rect 2418 -342 2424 -336
rect 2418 -348 2424 -342
rect 2418 -354 2424 -348
rect 2418 -360 2424 -354
rect 2418 -366 2424 -360
rect 2418 -372 2424 -366
rect 2418 -378 2424 -372
rect 2418 -384 2424 -378
rect 2418 -390 2424 -384
rect 2418 -396 2424 -390
rect 2418 -402 2424 -396
rect 2418 -408 2424 -402
rect 2418 -414 2424 -408
rect 2418 -420 2424 -414
rect 2418 -426 2424 -420
rect 2418 -432 2424 -426
rect 2418 -438 2424 -432
rect 2418 -444 2424 -438
rect 2418 -450 2424 -444
rect 2418 -456 2424 -450
rect 2418 -462 2424 -456
rect 2418 -468 2424 -462
rect 2418 -474 2424 -468
rect 2418 -480 2424 -474
rect 2418 -486 2424 -480
rect 2418 -492 2424 -486
rect 2418 -498 2424 -492
rect 2418 -504 2424 -498
rect 2418 -510 2424 -504
rect 2418 -516 2424 -510
rect 2418 -522 2424 -516
rect 2418 -528 2424 -522
rect 2418 -534 2424 -528
rect 2418 -540 2424 -534
rect 2418 -546 2424 -540
rect 2418 -552 2424 -546
rect 2418 -558 2424 -552
rect 2418 -564 2424 -558
rect 2418 -570 2424 -564
rect 2418 -576 2424 -570
rect 2418 -582 2424 -576
rect 2418 -588 2424 -582
rect 2418 -594 2424 -588
rect 2418 -600 2424 -594
rect 2418 -606 2424 -600
rect 2418 -612 2424 -606
rect 2418 -618 2424 -612
rect 2418 -624 2424 -618
rect 2418 -1374 2424 -1368
rect 2418 -1380 2424 -1374
rect 2418 -1386 2424 -1380
rect 2418 -1392 2424 -1386
rect 2418 -1398 2424 -1392
rect 2418 -1404 2424 -1398
rect 2418 -1410 2424 -1404
rect 2418 -1416 2424 -1410
rect 2418 -1422 2424 -1416
rect 2418 -1428 2424 -1422
rect 2418 -1434 2424 -1428
rect 2418 -1440 2424 -1434
rect 2418 -1446 2424 -1440
rect 2418 -1452 2424 -1446
rect 2418 -1458 2424 -1452
rect 2418 -1464 2424 -1458
rect 2418 -1470 2424 -1464
rect 2418 -1476 2424 -1470
rect 2418 -1482 2424 -1476
rect 2418 -1488 2424 -1482
rect 2418 -1494 2424 -1488
rect 2418 -1500 2424 -1494
rect 2418 -1506 2424 -1500
rect 2418 -1512 2424 -1506
rect 2418 -1518 2424 -1512
rect 2418 -1524 2424 -1518
rect 2418 -1530 2424 -1524
rect 2418 -1536 2424 -1530
rect 2418 -1542 2424 -1536
rect 2418 -1548 2424 -1542
rect 2418 -1554 2424 -1548
rect 2418 -1560 2424 -1554
rect 2418 -1566 2424 -1560
rect 2418 -1572 2424 -1566
rect 2418 -1578 2424 -1572
rect 2418 -1584 2424 -1578
rect 2418 -1590 2424 -1584
rect 2418 -1596 2424 -1590
rect 2418 -1602 2424 -1596
rect 2418 -1608 2424 -1602
rect 2418 -1614 2424 -1608
rect 2418 -1620 2424 -1614
rect 2418 -1626 2424 -1620
rect 2418 -1632 2424 -1626
rect 2418 -1638 2424 -1632
rect 2418 -1644 2424 -1638
rect 2418 -1650 2424 -1644
rect 2418 -1656 2424 -1650
rect 2418 -1662 2424 -1656
rect 2418 -1668 2424 -1662
rect 2418 -1674 2424 -1668
rect 2418 -1680 2424 -1674
rect 2418 -1686 2424 -1680
rect 2418 -1692 2424 -1686
rect 2418 -1698 2424 -1692
rect 2418 -1704 2424 -1698
rect 2418 -1710 2424 -1704
rect 2418 -1716 2424 -1710
rect 2418 -1722 2424 -1716
rect 2418 -1728 2424 -1722
rect 2418 -1734 2424 -1728
rect 2418 -1740 2424 -1734
rect 2418 -1746 2424 -1740
rect 2418 -1752 2424 -1746
rect 2418 -1758 2424 -1752
rect 2418 -1764 2424 -1758
rect 2418 -1770 2424 -1764
rect 2418 -1776 2424 -1770
rect 2418 -1782 2424 -1776
rect 2418 -1788 2424 -1782
rect 2418 -1794 2424 -1788
rect 2418 -1800 2424 -1794
rect 2418 -1806 2424 -1800
rect 2418 -1812 2424 -1806
rect 2418 -1818 2424 -1812
rect 2418 -1824 2424 -1818
rect 2418 -1830 2424 -1824
rect 2418 -1836 2424 -1830
rect 2418 -1842 2424 -1836
rect 2418 -1848 2424 -1842
rect 2418 -1854 2424 -1848
rect 2418 -1860 2424 -1854
rect 2418 -1866 2424 -1860
rect 2418 -1872 2424 -1866
rect 2418 -1878 2424 -1872
rect 2418 -1884 2424 -1878
rect 2418 -1890 2424 -1884
rect 2418 -1896 2424 -1890
rect 2418 -1902 2424 -1896
rect 2418 -1908 2424 -1902
rect 2418 -1914 2424 -1908
rect 2418 -1920 2424 -1914
rect 2418 -1926 2424 -1920
rect 2418 -1932 2424 -1926
rect 2418 -1938 2424 -1932
rect 2418 -1944 2424 -1938
rect 2418 -1950 2424 -1944
rect 2418 -1956 2424 -1950
rect 2418 -1962 2424 -1956
rect 2418 -1968 2424 -1962
rect 2418 -1974 2424 -1968
rect 2418 -1980 2424 -1974
rect 2418 -1986 2424 -1980
rect 2418 -1992 2424 -1986
rect 2418 -1998 2424 -1992
rect 2418 -2004 2424 -1998
rect 2418 -2010 2424 -2004
rect 2418 -2016 2424 -2010
rect 2418 -2022 2424 -2016
rect 2418 -2028 2424 -2022
rect 2418 -2034 2424 -2028
rect 2418 -2040 2424 -2034
rect 2418 -2046 2424 -2040
rect 2418 -2052 2424 -2046
rect 2418 -2058 2424 -2052
rect 2418 -2064 2424 -2058
rect 2418 -2070 2424 -2064
rect 2418 -2076 2424 -2070
rect 2418 -2178 2424 -2172
rect 2418 -2184 2424 -2178
rect 2418 -2190 2424 -2184
rect 2418 -2196 2424 -2190
rect 2418 -2202 2424 -2196
rect 2418 -2208 2424 -2202
rect 2418 -2214 2424 -2208
rect 2418 -2220 2424 -2214
rect 2418 -2226 2424 -2220
rect 2418 -2232 2424 -2226
rect 2418 -2238 2424 -2232
rect 2418 -2244 2424 -2238
rect 2418 -2250 2424 -2244
rect 2418 -2256 2424 -2250
rect 2418 -2262 2424 -2256
rect 2418 -2268 2424 -2262
rect 2418 -2274 2424 -2268
rect 2418 -2280 2424 -2274
rect 2418 -2286 2424 -2280
rect 2418 -2292 2424 -2286
rect 2418 -2298 2424 -2292
rect 2418 -2304 2424 -2298
rect 2418 -2310 2424 -2304
rect 2418 -2316 2424 -2310
rect 2418 -2322 2424 -2316
rect 2418 -2328 2424 -2322
rect 2418 -2334 2424 -2328
rect 2418 -2340 2424 -2334
rect 2418 -2346 2424 -2340
rect 2418 -2352 2424 -2346
rect 2418 -2358 2424 -2352
rect 2418 -2364 2424 -2358
rect 2418 -2370 2424 -2364
rect 2418 -2376 2424 -2370
rect 2418 -2382 2424 -2376
rect 2418 -2388 2424 -2382
rect 2418 -2394 2424 -2388
rect 2418 -2400 2424 -2394
rect 2418 -2472 2424 -2466
rect 2418 -2478 2424 -2472
rect 2418 -2484 2424 -2478
rect 2418 -2490 2424 -2484
rect 2418 -2496 2424 -2490
rect 2418 -2502 2424 -2496
rect 2418 -2508 2424 -2502
rect 2418 -2514 2424 -2508
rect 2418 -2520 2424 -2514
rect 2418 -2526 2424 -2520
rect 2418 -2532 2424 -2526
rect 2418 -2538 2424 -2532
rect 2418 -2544 2424 -2538
rect 2418 -2550 2424 -2544
rect 2418 -2556 2424 -2550
rect 2418 -2562 2424 -2556
rect 2418 -2568 2424 -2562
rect 2418 -2574 2424 -2568
rect 2418 -2580 2424 -2574
rect 2418 -2586 2424 -2580
rect 2418 -2592 2424 -2586
rect 2418 -2598 2424 -2592
rect 2418 -2604 2424 -2598
rect 2418 -2610 2424 -2604
rect 2418 -2616 2424 -2610
rect 2418 -2622 2424 -2616
rect 2418 -2628 2424 -2622
rect 2418 -2634 2424 -2628
rect 2418 -2640 2424 -2634
rect 2418 -2646 2424 -2640
rect 2418 -2652 2424 -2646
rect 2418 -2658 2424 -2652
rect 2418 -2664 2424 -2658
rect 2418 -2670 2424 -2664
rect 2418 -2676 2424 -2670
rect 2418 -2682 2424 -2676
rect 2418 -2688 2424 -2682
rect 2418 -2694 2424 -2688
rect 2418 -2700 2424 -2694
rect 2418 -2706 2424 -2700
rect 2418 -2712 2424 -2706
rect 2418 -2718 2424 -2712
rect 2418 -2724 2424 -2718
rect 2418 -2730 2424 -2724
rect 2418 -2736 2424 -2730
rect 2418 -2742 2424 -2736
rect 2418 -2748 2424 -2742
rect 2418 -2754 2424 -2748
rect 2418 -2760 2424 -2754
rect 2418 -2766 2424 -2760
rect 2418 -2772 2424 -2766
rect 2418 -2778 2424 -2772
rect 2418 -2784 2424 -2778
rect 2418 -2790 2424 -2784
rect 2418 -2796 2424 -2790
rect 2418 -2802 2424 -2796
rect 2418 -2808 2424 -2802
rect 2418 -2814 2424 -2808
rect 2418 -2820 2424 -2814
rect 2418 -2826 2424 -2820
rect 2418 -2832 2424 -2826
rect 2418 -2838 2424 -2832
rect 2418 -2844 2424 -2838
rect 2418 -2850 2424 -2844
rect 2418 -2856 2424 -2850
rect 2418 -2862 2424 -2856
rect 2418 -2868 2424 -2862
rect 2418 -2874 2424 -2868
rect 2424 -282 2430 -276
rect 2424 -288 2430 -282
rect 2424 -294 2430 -288
rect 2424 -300 2430 -294
rect 2424 -306 2430 -300
rect 2424 -312 2430 -306
rect 2424 -318 2430 -312
rect 2424 -324 2430 -318
rect 2424 -330 2430 -324
rect 2424 -336 2430 -330
rect 2424 -342 2430 -336
rect 2424 -348 2430 -342
rect 2424 -354 2430 -348
rect 2424 -360 2430 -354
rect 2424 -366 2430 -360
rect 2424 -372 2430 -366
rect 2424 -378 2430 -372
rect 2424 -384 2430 -378
rect 2424 -390 2430 -384
rect 2424 -396 2430 -390
rect 2424 -402 2430 -396
rect 2424 -408 2430 -402
rect 2424 -414 2430 -408
rect 2424 -420 2430 -414
rect 2424 -426 2430 -420
rect 2424 -432 2430 -426
rect 2424 -438 2430 -432
rect 2424 -444 2430 -438
rect 2424 -450 2430 -444
rect 2424 -456 2430 -450
rect 2424 -462 2430 -456
rect 2424 -468 2430 -462
rect 2424 -474 2430 -468
rect 2424 -480 2430 -474
rect 2424 -486 2430 -480
rect 2424 -492 2430 -486
rect 2424 -498 2430 -492
rect 2424 -504 2430 -498
rect 2424 -510 2430 -504
rect 2424 -516 2430 -510
rect 2424 -522 2430 -516
rect 2424 -528 2430 -522
rect 2424 -534 2430 -528
rect 2424 -540 2430 -534
rect 2424 -546 2430 -540
rect 2424 -552 2430 -546
rect 2424 -558 2430 -552
rect 2424 -564 2430 -558
rect 2424 -570 2430 -564
rect 2424 -576 2430 -570
rect 2424 -582 2430 -576
rect 2424 -588 2430 -582
rect 2424 -594 2430 -588
rect 2424 -600 2430 -594
rect 2424 -1368 2430 -1362
rect 2424 -1374 2430 -1368
rect 2424 -1380 2430 -1374
rect 2424 -1386 2430 -1380
rect 2424 -1392 2430 -1386
rect 2424 -1398 2430 -1392
rect 2424 -1404 2430 -1398
rect 2424 -1410 2430 -1404
rect 2424 -1416 2430 -1410
rect 2424 -1422 2430 -1416
rect 2424 -1428 2430 -1422
rect 2424 -1434 2430 -1428
rect 2424 -1440 2430 -1434
rect 2424 -1446 2430 -1440
rect 2424 -1452 2430 -1446
rect 2424 -1458 2430 -1452
rect 2424 -1464 2430 -1458
rect 2424 -1470 2430 -1464
rect 2424 -1476 2430 -1470
rect 2424 -1482 2430 -1476
rect 2424 -1488 2430 -1482
rect 2424 -1494 2430 -1488
rect 2424 -1500 2430 -1494
rect 2424 -1506 2430 -1500
rect 2424 -1512 2430 -1506
rect 2424 -1518 2430 -1512
rect 2424 -1524 2430 -1518
rect 2424 -1530 2430 -1524
rect 2424 -1536 2430 -1530
rect 2424 -1542 2430 -1536
rect 2424 -1548 2430 -1542
rect 2424 -1554 2430 -1548
rect 2424 -1560 2430 -1554
rect 2424 -1566 2430 -1560
rect 2424 -1572 2430 -1566
rect 2424 -1578 2430 -1572
rect 2424 -1584 2430 -1578
rect 2424 -1590 2430 -1584
rect 2424 -1596 2430 -1590
rect 2424 -1602 2430 -1596
rect 2424 -1608 2430 -1602
rect 2424 -1614 2430 -1608
rect 2424 -1620 2430 -1614
rect 2424 -1626 2430 -1620
rect 2424 -1632 2430 -1626
rect 2424 -1638 2430 -1632
rect 2424 -1644 2430 -1638
rect 2424 -1650 2430 -1644
rect 2424 -1656 2430 -1650
rect 2424 -1662 2430 -1656
rect 2424 -1668 2430 -1662
rect 2424 -1674 2430 -1668
rect 2424 -1680 2430 -1674
rect 2424 -1686 2430 -1680
rect 2424 -1692 2430 -1686
rect 2424 -1698 2430 -1692
rect 2424 -1704 2430 -1698
rect 2424 -1710 2430 -1704
rect 2424 -1716 2430 -1710
rect 2424 -1722 2430 -1716
rect 2424 -1728 2430 -1722
rect 2424 -1734 2430 -1728
rect 2424 -1740 2430 -1734
rect 2424 -1746 2430 -1740
rect 2424 -1752 2430 -1746
rect 2424 -1758 2430 -1752
rect 2424 -1764 2430 -1758
rect 2424 -1770 2430 -1764
rect 2424 -1776 2430 -1770
rect 2424 -1782 2430 -1776
rect 2424 -1788 2430 -1782
rect 2424 -1794 2430 -1788
rect 2424 -1800 2430 -1794
rect 2424 -1806 2430 -1800
rect 2424 -1812 2430 -1806
rect 2424 -1818 2430 -1812
rect 2424 -1824 2430 -1818
rect 2424 -1830 2430 -1824
rect 2424 -1836 2430 -1830
rect 2424 -1842 2430 -1836
rect 2424 -1848 2430 -1842
rect 2424 -1854 2430 -1848
rect 2424 -1860 2430 -1854
rect 2424 -1866 2430 -1860
rect 2424 -1872 2430 -1866
rect 2424 -1878 2430 -1872
rect 2424 -1884 2430 -1878
rect 2424 -1890 2430 -1884
rect 2424 -1896 2430 -1890
rect 2424 -1902 2430 -1896
rect 2424 -1908 2430 -1902
rect 2424 -1914 2430 -1908
rect 2424 -1920 2430 -1914
rect 2424 -1926 2430 -1920
rect 2424 -1932 2430 -1926
rect 2424 -1938 2430 -1932
rect 2424 -1944 2430 -1938
rect 2424 -1950 2430 -1944
rect 2424 -1956 2430 -1950
rect 2424 -1962 2430 -1956
rect 2424 -1968 2430 -1962
rect 2424 -1974 2430 -1968
rect 2424 -1980 2430 -1974
rect 2424 -1986 2430 -1980
rect 2424 -1992 2430 -1986
rect 2424 -1998 2430 -1992
rect 2424 -2004 2430 -1998
rect 2424 -2010 2430 -2004
rect 2424 -2016 2430 -2010
rect 2424 -2022 2430 -2016
rect 2424 -2028 2430 -2022
rect 2424 -2034 2430 -2028
rect 2424 -2040 2430 -2034
rect 2424 -2046 2430 -2040
rect 2424 -2052 2430 -2046
rect 2424 -2058 2430 -2052
rect 2424 -2064 2430 -2058
rect 2424 -2070 2430 -2064
rect 2424 -2214 2430 -2208
rect 2424 -2220 2430 -2214
rect 2424 -2226 2430 -2220
rect 2424 -2232 2430 -2226
rect 2424 -2238 2430 -2232
rect 2424 -2244 2430 -2238
rect 2424 -2250 2430 -2244
rect 2424 -2256 2430 -2250
rect 2424 -2262 2430 -2256
rect 2424 -2268 2430 -2262
rect 2424 -2274 2430 -2268
rect 2424 -2280 2430 -2274
rect 2424 -2286 2430 -2280
rect 2424 -2292 2430 -2286
rect 2424 -2298 2430 -2292
rect 2424 -2304 2430 -2298
rect 2424 -2310 2430 -2304
rect 2424 -2316 2430 -2310
rect 2424 -2322 2430 -2316
rect 2424 -2328 2430 -2322
rect 2424 -2334 2430 -2328
rect 2424 -2340 2430 -2334
rect 2424 -2346 2430 -2340
rect 2424 -2352 2430 -2346
rect 2424 -2358 2430 -2352
rect 2424 -2364 2430 -2358
rect 2424 -2370 2430 -2364
rect 2424 -2376 2430 -2370
rect 2424 -2472 2430 -2466
rect 2424 -2478 2430 -2472
rect 2424 -2484 2430 -2478
rect 2424 -2490 2430 -2484
rect 2424 -2496 2430 -2490
rect 2424 -2502 2430 -2496
rect 2424 -2508 2430 -2502
rect 2424 -2514 2430 -2508
rect 2424 -2520 2430 -2514
rect 2424 -2526 2430 -2520
rect 2424 -2532 2430 -2526
rect 2424 -2538 2430 -2532
rect 2424 -2544 2430 -2538
rect 2424 -2550 2430 -2544
rect 2424 -2556 2430 -2550
rect 2424 -2562 2430 -2556
rect 2424 -2568 2430 -2562
rect 2424 -2574 2430 -2568
rect 2424 -2580 2430 -2574
rect 2424 -2586 2430 -2580
rect 2424 -2592 2430 -2586
rect 2424 -2598 2430 -2592
rect 2424 -2604 2430 -2598
rect 2424 -2610 2430 -2604
rect 2424 -2616 2430 -2610
rect 2424 -2622 2430 -2616
rect 2424 -2628 2430 -2622
rect 2424 -2634 2430 -2628
rect 2424 -2640 2430 -2634
rect 2424 -2646 2430 -2640
rect 2424 -2652 2430 -2646
rect 2424 -2658 2430 -2652
rect 2424 -2664 2430 -2658
rect 2424 -2670 2430 -2664
rect 2424 -2676 2430 -2670
rect 2424 -2682 2430 -2676
rect 2424 -2688 2430 -2682
rect 2424 -2694 2430 -2688
rect 2424 -2700 2430 -2694
rect 2424 -2706 2430 -2700
rect 2424 -2712 2430 -2706
rect 2424 -2718 2430 -2712
rect 2424 -2724 2430 -2718
rect 2424 -2730 2430 -2724
rect 2424 -2736 2430 -2730
rect 2424 -2742 2430 -2736
rect 2424 -2748 2430 -2742
rect 2424 -2754 2430 -2748
rect 2424 -2760 2430 -2754
rect 2424 -2766 2430 -2760
rect 2424 -2772 2430 -2766
rect 2424 -2778 2430 -2772
rect 2424 -2784 2430 -2778
rect 2424 -2790 2430 -2784
rect 2424 -2796 2430 -2790
rect 2424 -2802 2430 -2796
rect 2424 -2808 2430 -2802
rect 2424 -2814 2430 -2808
rect 2424 -2820 2430 -2814
rect 2424 -2826 2430 -2820
rect 2424 -2832 2430 -2826
rect 2424 -2838 2430 -2832
rect 2424 -2844 2430 -2838
rect 2424 -2850 2430 -2844
rect 2424 -2856 2430 -2850
rect 2424 -2862 2430 -2856
rect 2424 -2868 2430 -2862
rect 2424 -2874 2430 -2868
rect 2430 -312 2436 -306
rect 2430 -318 2436 -312
rect 2430 -324 2436 -318
rect 2430 -330 2436 -324
rect 2430 -336 2436 -330
rect 2430 -342 2436 -336
rect 2430 -348 2436 -342
rect 2430 -354 2436 -348
rect 2430 -360 2436 -354
rect 2430 -366 2436 -360
rect 2430 -372 2436 -366
rect 2430 -378 2436 -372
rect 2430 -384 2436 -378
rect 2430 -390 2436 -384
rect 2430 -396 2436 -390
rect 2430 -402 2436 -396
rect 2430 -408 2436 -402
rect 2430 -414 2436 -408
rect 2430 -420 2436 -414
rect 2430 -426 2436 -420
rect 2430 -432 2436 -426
rect 2430 -438 2436 -432
rect 2430 -444 2436 -438
rect 2430 -450 2436 -444
rect 2430 -456 2436 -450
rect 2430 -462 2436 -456
rect 2430 -468 2436 -462
rect 2430 -474 2436 -468
rect 2430 -480 2436 -474
rect 2430 -486 2436 -480
rect 2430 -492 2436 -486
rect 2430 -498 2436 -492
rect 2430 -504 2436 -498
rect 2430 -510 2436 -504
rect 2430 -516 2436 -510
rect 2430 -522 2436 -516
rect 2430 -528 2436 -522
rect 2430 -534 2436 -528
rect 2430 -540 2436 -534
rect 2430 -546 2436 -540
rect 2430 -552 2436 -546
rect 2430 -558 2436 -552
rect 2430 -564 2436 -558
rect 2430 -1362 2436 -1356
rect 2430 -1368 2436 -1362
rect 2430 -1374 2436 -1368
rect 2430 -1380 2436 -1374
rect 2430 -1386 2436 -1380
rect 2430 -1392 2436 -1386
rect 2430 -1398 2436 -1392
rect 2430 -1404 2436 -1398
rect 2430 -1410 2436 -1404
rect 2430 -1416 2436 -1410
rect 2430 -1422 2436 -1416
rect 2430 -1428 2436 -1422
rect 2430 -1434 2436 -1428
rect 2430 -1440 2436 -1434
rect 2430 -1446 2436 -1440
rect 2430 -1452 2436 -1446
rect 2430 -1458 2436 -1452
rect 2430 -1464 2436 -1458
rect 2430 -1470 2436 -1464
rect 2430 -1476 2436 -1470
rect 2430 -1482 2436 -1476
rect 2430 -1488 2436 -1482
rect 2430 -1494 2436 -1488
rect 2430 -1500 2436 -1494
rect 2430 -1506 2436 -1500
rect 2430 -1512 2436 -1506
rect 2430 -1518 2436 -1512
rect 2430 -1524 2436 -1518
rect 2430 -1530 2436 -1524
rect 2430 -1536 2436 -1530
rect 2430 -1542 2436 -1536
rect 2430 -1548 2436 -1542
rect 2430 -1554 2436 -1548
rect 2430 -1560 2436 -1554
rect 2430 -1566 2436 -1560
rect 2430 -1572 2436 -1566
rect 2430 -1578 2436 -1572
rect 2430 -1584 2436 -1578
rect 2430 -1590 2436 -1584
rect 2430 -1596 2436 -1590
rect 2430 -1602 2436 -1596
rect 2430 -1608 2436 -1602
rect 2430 -1614 2436 -1608
rect 2430 -1620 2436 -1614
rect 2430 -1626 2436 -1620
rect 2430 -1632 2436 -1626
rect 2430 -1638 2436 -1632
rect 2430 -1644 2436 -1638
rect 2430 -1650 2436 -1644
rect 2430 -1656 2436 -1650
rect 2430 -1662 2436 -1656
rect 2430 -1668 2436 -1662
rect 2430 -1674 2436 -1668
rect 2430 -1680 2436 -1674
rect 2430 -1686 2436 -1680
rect 2430 -1692 2436 -1686
rect 2430 -1698 2436 -1692
rect 2430 -1704 2436 -1698
rect 2430 -1710 2436 -1704
rect 2430 -1716 2436 -1710
rect 2430 -1722 2436 -1716
rect 2430 -1728 2436 -1722
rect 2430 -1734 2436 -1728
rect 2430 -1740 2436 -1734
rect 2430 -1746 2436 -1740
rect 2430 -1752 2436 -1746
rect 2430 -1758 2436 -1752
rect 2430 -1764 2436 -1758
rect 2430 -1770 2436 -1764
rect 2430 -1776 2436 -1770
rect 2430 -1782 2436 -1776
rect 2430 -1788 2436 -1782
rect 2430 -1794 2436 -1788
rect 2430 -1800 2436 -1794
rect 2430 -1806 2436 -1800
rect 2430 -1812 2436 -1806
rect 2430 -1818 2436 -1812
rect 2430 -1824 2436 -1818
rect 2430 -1830 2436 -1824
rect 2430 -1836 2436 -1830
rect 2430 -1842 2436 -1836
rect 2430 -1848 2436 -1842
rect 2430 -1854 2436 -1848
rect 2430 -1860 2436 -1854
rect 2430 -1866 2436 -1860
rect 2430 -1872 2436 -1866
rect 2430 -1878 2436 -1872
rect 2430 -1884 2436 -1878
rect 2430 -1890 2436 -1884
rect 2430 -1896 2436 -1890
rect 2430 -1902 2436 -1896
rect 2430 -1908 2436 -1902
rect 2430 -1914 2436 -1908
rect 2430 -1920 2436 -1914
rect 2430 -1926 2436 -1920
rect 2430 -1932 2436 -1926
rect 2430 -1938 2436 -1932
rect 2430 -1944 2436 -1938
rect 2430 -1950 2436 -1944
rect 2430 -1956 2436 -1950
rect 2430 -1962 2436 -1956
rect 2430 -1968 2436 -1962
rect 2430 -1974 2436 -1968
rect 2430 -1980 2436 -1974
rect 2430 -1986 2436 -1980
rect 2430 -1992 2436 -1986
rect 2430 -1998 2436 -1992
rect 2430 -2004 2436 -1998
rect 2430 -2010 2436 -2004
rect 2430 -2016 2436 -2010
rect 2430 -2022 2436 -2016
rect 2430 -2028 2436 -2022
rect 2430 -2034 2436 -2028
rect 2430 -2040 2436 -2034
rect 2430 -2046 2436 -2040
rect 2430 -2052 2436 -2046
rect 2430 -2058 2436 -2052
rect 2430 -2472 2436 -2466
rect 2430 -2478 2436 -2472
rect 2430 -2484 2436 -2478
rect 2430 -2490 2436 -2484
rect 2430 -2496 2436 -2490
rect 2430 -2502 2436 -2496
rect 2430 -2508 2436 -2502
rect 2430 -2514 2436 -2508
rect 2430 -2520 2436 -2514
rect 2430 -2526 2436 -2520
rect 2430 -2532 2436 -2526
rect 2430 -2538 2436 -2532
rect 2430 -2544 2436 -2538
rect 2430 -2550 2436 -2544
rect 2430 -2556 2436 -2550
rect 2430 -2562 2436 -2556
rect 2430 -2568 2436 -2562
rect 2430 -2574 2436 -2568
rect 2430 -2580 2436 -2574
rect 2430 -2586 2436 -2580
rect 2430 -2592 2436 -2586
rect 2430 -2598 2436 -2592
rect 2430 -2604 2436 -2598
rect 2430 -2610 2436 -2604
rect 2430 -2616 2436 -2610
rect 2430 -2622 2436 -2616
rect 2430 -2628 2436 -2622
rect 2430 -2634 2436 -2628
rect 2430 -2640 2436 -2634
rect 2430 -2646 2436 -2640
rect 2430 -2652 2436 -2646
rect 2430 -2658 2436 -2652
rect 2430 -2664 2436 -2658
rect 2430 -2670 2436 -2664
rect 2430 -2676 2436 -2670
rect 2430 -2682 2436 -2676
rect 2430 -2688 2436 -2682
rect 2430 -2694 2436 -2688
rect 2430 -2700 2436 -2694
rect 2430 -2706 2436 -2700
rect 2430 -2712 2436 -2706
rect 2430 -2718 2436 -2712
rect 2430 -2724 2436 -2718
rect 2430 -2730 2436 -2724
rect 2430 -2736 2436 -2730
rect 2430 -2742 2436 -2736
rect 2430 -2748 2436 -2742
rect 2430 -2754 2436 -2748
rect 2430 -2760 2436 -2754
rect 2430 -2766 2436 -2760
rect 2430 -2772 2436 -2766
rect 2430 -2778 2436 -2772
rect 2430 -2784 2436 -2778
rect 2430 -2790 2436 -2784
rect 2430 -2796 2436 -2790
rect 2430 -2802 2436 -2796
rect 2430 -2808 2436 -2802
rect 2430 -2814 2436 -2808
rect 2430 -2820 2436 -2814
rect 2430 -2826 2436 -2820
rect 2430 -2832 2436 -2826
rect 2430 -2838 2436 -2832
rect 2430 -2844 2436 -2838
rect 2430 -2850 2436 -2844
rect 2430 -2856 2436 -2850
rect 2430 -2862 2436 -2856
rect 2430 -2868 2436 -2862
rect 2436 -354 2442 -348
rect 2436 -360 2442 -354
rect 2436 -366 2442 -360
rect 2436 -372 2442 -366
rect 2436 -378 2442 -372
rect 2436 -384 2442 -378
rect 2436 -390 2442 -384
rect 2436 -396 2442 -390
rect 2436 -402 2442 -396
rect 2436 -408 2442 -402
rect 2436 -414 2442 -408
rect 2436 -420 2442 -414
rect 2436 -426 2442 -420
rect 2436 -432 2442 -426
rect 2436 -438 2442 -432
rect 2436 -444 2442 -438
rect 2436 -450 2442 -444
rect 2436 -456 2442 -450
rect 2436 -462 2442 -456
rect 2436 -468 2442 -462
rect 2436 -474 2442 -468
rect 2436 -480 2442 -474
rect 2436 -486 2442 -480
rect 2436 -492 2442 -486
rect 2436 -498 2442 -492
rect 2436 -504 2442 -498
rect 2436 -510 2442 -504
rect 2436 -516 2442 -510
rect 2436 -522 2442 -516
rect 2436 -528 2442 -522
rect 2436 -1356 2442 -1350
rect 2436 -1362 2442 -1356
rect 2436 -1368 2442 -1362
rect 2436 -1374 2442 -1368
rect 2436 -1380 2442 -1374
rect 2436 -1386 2442 -1380
rect 2436 -1392 2442 -1386
rect 2436 -1398 2442 -1392
rect 2436 -1404 2442 -1398
rect 2436 -1410 2442 -1404
rect 2436 -1416 2442 -1410
rect 2436 -1422 2442 -1416
rect 2436 -1428 2442 -1422
rect 2436 -1434 2442 -1428
rect 2436 -1440 2442 -1434
rect 2436 -1446 2442 -1440
rect 2436 -1452 2442 -1446
rect 2436 -1458 2442 -1452
rect 2436 -1464 2442 -1458
rect 2436 -1470 2442 -1464
rect 2436 -1476 2442 -1470
rect 2436 -1482 2442 -1476
rect 2436 -1488 2442 -1482
rect 2436 -1494 2442 -1488
rect 2436 -1500 2442 -1494
rect 2436 -1506 2442 -1500
rect 2436 -1512 2442 -1506
rect 2436 -1518 2442 -1512
rect 2436 -1524 2442 -1518
rect 2436 -1530 2442 -1524
rect 2436 -1536 2442 -1530
rect 2436 -1542 2442 -1536
rect 2436 -1548 2442 -1542
rect 2436 -1554 2442 -1548
rect 2436 -1560 2442 -1554
rect 2436 -1566 2442 -1560
rect 2436 -1572 2442 -1566
rect 2436 -1578 2442 -1572
rect 2436 -1584 2442 -1578
rect 2436 -1590 2442 -1584
rect 2436 -1596 2442 -1590
rect 2436 -1602 2442 -1596
rect 2436 -1608 2442 -1602
rect 2436 -1614 2442 -1608
rect 2436 -1620 2442 -1614
rect 2436 -1626 2442 -1620
rect 2436 -1632 2442 -1626
rect 2436 -1638 2442 -1632
rect 2436 -1644 2442 -1638
rect 2436 -1650 2442 -1644
rect 2436 -1656 2442 -1650
rect 2436 -1662 2442 -1656
rect 2436 -1668 2442 -1662
rect 2436 -1674 2442 -1668
rect 2436 -1680 2442 -1674
rect 2436 -1686 2442 -1680
rect 2436 -1692 2442 -1686
rect 2436 -1698 2442 -1692
rect 2436 -1704 2442 -1698
rect 2436 -1710 2442 -1704
rect 2436 -1716 2442 -1710
rect 2436 -1722 2442 -1716
rect 2436 -1728 2442 -1722
rect 2436 -1734 2442 -1728
rect 2436 -1740 2442 -1734
rect 2436 -1746 2442 -1740
rect 2436 -1752 2442 -1746
rect 2436 -1758 2442 -1752
rect 2436 -1764 2442 -1758
rect 2436 -1770 2442 -1764
rect 2436 -1776 2442 -1770
rect 2436 -1782 2442 -1776
rect 2436 -1788 2442 -1782
rect 2436 -1794 2442 -1788
rect 2436 -1800 2442 -1794
rect 2436 -1806 2442 -1800
rect 2436 -1812 2442 -1806
rect 2436 -1818 2442 -1812
rect 2436 -1824 2442 -1818
rect 2436 -1830 2442 -1824
rect 2436 -1836 2442 -1830
rect 2436 -1842 2442 -1836
rect 2436 -1848 2442 -1842
rect 2436 -1854 2442 -1848
rect 2436 -1860 2442 -1854
rect 2436 -1866 2442 -1860
rect 2436 -1872 2442 -1866
rect 2436 -1878 2442 -1872
rect 2436 -1884 2442 -1878
rect 2436 -1890 2442 -1884
rect 2436 -1896 2442 -1890
rect 2436 -1902 2442 -1896
rect 2436 -1908 2442 -1902
rect 2436 -1914 2442 -1908
rect 2436 -1920 2442 -1914
rect 2436 -1926 2442 -1920
rect 2436 -1932 2442 -1926
rect 2436 -1938 2442 -1932
rect 2436 -1944 2442 -1938
rect 2436 -1950 2442 -1944
rect 2436 -1956 2442 -1950
rect 2436 -1962 2442 -1956
rect 2436 -1968 2442 -1962
rect 2436 -1974 2442 -1968
rect 2436 -1980 2442 -1974
rect 2436 -1986 2442 -1980
rect 2436 -1992 2442 -1986
rect 2436 -1998 2442 -1992
rect 2436 -2004 2442 -1998
rect 2436 -2010 2442 -2004
rect 2436 -2016 2442 -2010
rect 2436 -2022 2442 -2016
rect 2436 -2028 2442 -2022
rect 2436 -2034 2442 -2028
rect 2436 -2040 2442 -2034
rect 2436 -2046 2442 -2040
rect 2436 -2052 2442 -2046
rect 2436 -2466 2442 -2460
rect 2436 -2472 2442 -2466
rect 2436 -2478 2442 -2472
rect 2436 -2484 2442 -2478
rect 2436 -2490 2442 -2484
rect 2436 -2496 2442 -2490
rect 2436 -2502 2442 -2496
rect 2436 -2508 2442 -2502
rect 2436 -2514 2442 -2508
rect 2436 -2520 2442 -2514
rect 2436 -2526 2442 -2520
rect 2436 -2532 2442 -2526
rect 2436 -2538 2442 -2532
rect 2436 -2544 2442 -2538
rect 2436 -2550 2442 -2544
rect 2436 -2556 2442 -2550
rect 2436 -2562 2442 -2556
rect 2436 -2568 2442 -2562
rect 2436 -2574 2442 -2568
rect 2436 -2580 2442 -2574
rect 2436 -2586 2442 -2580
rect 2436 -2592 2442 -2586
rect 2436 -2598 2442 -2592
rect 2436 -2604 2442 -2598
rect 2436 -2610 2442 -2604
rect 2436 -2616 2442 -2610
rect 2436 -2622 2442 -2616
rect 2436 -2628 2442 -2622
rect 2436 -2634 2442 -2628
rect 2436 -2640 2442 -2634
rect 2436 -2646 2442 -2640
rect 2436 -2652 2442 -2646
rect 2436 -2658 2442 -2652
rect 2436 -2664 2442 -2658
rect 2436 -2670 2442 -2664
rect 2436 -2676 2442 -2670
rect 2436 -2682 2442 -2676
rect 2436 -2688 2442 -2682
rect 2436 -2694 2442 -2688
rect 2436 -2700 2442 -2694
rect 2436 -2706 2442 -2700
rect 2436 -2712 2442 -2706
rect 2436 -2718 2442 -2712
rect 2436 -2724 2442 -2718
rect 2436 -2730 2442 -2724
rect 2436 -2736 2442 -2730
rect 2436 -2742 2442 -2736
rect 2436 -2748 2442 -2742
rect 2436 -2754 2442 -2748
rect 2436 -2760 2442 -2754
rect 2436 -2766 2442 -2760
rect 2436 -2772 2442 -2766
rect 2436 -2778 2442 -2772
rect 2436 -2784 2442 -2778
rect 2436 -2790 2442 -2784
rect 2436 -2796 2442 -2790
rect 2436 -2802 2442 -2796
rect 2436 -2808 2442 -2802
rect 2436 -2814 2442 -2808
rect 2436 -2820 2442 -2814
rect 2436 -2826 2442 -2820
rect 2436 -2832 2442 -2826
rect 2436 -2838 2442 -2832
rect 2436 -2844 2442 -2838
rect 2436 -2850 2442 -2844
rect 2436 -2856 2442 -2850
rect 2436 -2862 2442 -2856
rect 2442 -432 2448 -426
rect 2442 -438 2448 -432
rect 2442 -444 2448 -438
rect 2442 -450 2448 -444
rect 2442 -456 2448 -450
rect 2442 -1356 2448 -1350
rect 2442 -1362 2448 -1356
rect 2442 -1368 2448 -1362
rect 2442 -1374 2448 -1368
rect 2442 -1380 2448 -1374
rect 2442 -1386 2448 -1380
rect 2442 -1392 2448 -1386
rect 2442 -1398 2448 -1392
rect 2442 -1404 2448 -1398
rect 2442 -1410 2448 -1404
rect 2442 -1416 2448 -1410
rect 2442 -1422 2448 -1416
rect 2442 -1428 2448 -1422
rect 2442 -1434 2448 -1428
rect 2442 -1440 2448 -1434
rect 2442 -1446 2448 -1440
rect 2442 -1452 2448 -1446
rect 2442 -1458 2448 -1452
rect 2442 -1464 2448 -1458
rect 2442 -1470 2448 -1464
rect 2442 -1476 2448 -1470
rect 2442 -1482 2448 -1476
rect 2442 -1488 2448 -1482
rect 2442 -1494 2448 -1488
rect 2442 -1500 2448 -1494
rect 2442 -1506 2448 -1500
rect 2442 -1512 2448 -1506
rect 2442 -1518 2448 -1512
rect 2442 -1524 2448 -1518
rect 2442 -1530 2448 -1524
rect 2442 -1536 2448 -1530
rect 2442 -1542 2448 -1536
rect 2442 -1548 2448 -1542
rect 2442 -1554 2448 -1548
rect 2442 -1560 2448 -1554
rect 2442 -1566 2448 -1560
rect 2442 -1572 2448 -1566
rect 2442 -1578 2448 -1572
rect 2442 -1584 2448 -1578
rect 2442 -1590 2448 -1584
rect 2442 -1596 2448 -1590
rect 2442 -1602 2448 -1596
rect 2442 -1608 2448 -1602
rect 2442 -1614 2448 -1608
rect 2442 -1620 2448 -1614
rect 2442 -1626 2448 -1620
rect 2442 -1632 2448 -1626
rect 2442 -1638 2448 -1632
rect 2442 -1644 2448 -1638
rect 2442 -1650 2448 -1644
rect 2442 -1656 2448 -1650
rect 2442 -1662 2448 -1656
rect 2442 -1668 2448 -1662
rect 2442 -1674 2448 -1668
rect 2442 -1680 2448 -1674
rect 2442 -1686 2448 -1680
rect 2442 -1692 2448 -1686
rect 2442 -1698 2448 -1692
rect 2442 -1704 2448 -1698
rect 2442 -1710 2448 -1704
rect 2442 -1716 2448 -1710
rect 2442 -1722 2448 -1716
rect 2442 -1728 2448 -1722
rect 2442 -1734 2448 -1728
rect 2442 -1740 2448 -1734
rect 2442 -1746 2448 -1740
rect 2442 -1752 2448 -1746
rect 2442 -1758 2448 -1752
rect 2442 -1764 2448 -1758
rect 2442 -1770 2448 -1764
rect 2442 -1776 2448 -1770
rect 2442 -1782 2448 -1776
rect 2442 -1788 2448 -1782
rect 2442 -1794 2448 -1788
rect 2442 -1800 2448 -1794
rect 2442 -1806 2448 -1800
rect 2442 -1812 2448 -1806
rect 2442 -1818 2448 -1812
rect 2442 -1824 2448 -1818
rect 2442 -1830 2448 -1824
rect 2442 -1836 2448 -1830
rect 2442 -1842 2448 -1836
rect 2442 -1848 2448 -1842
rect 2442 -1854 2448 -1848
rect 2442 -1860 2448 -1854
rect 2442 -1866 2448 -1860
rect 2442 -1872 2448 -1866
rect 2442 -1878 2448 -1872
rect 2442 -1884 2448 -1878
rect 2442 -1890 2448 -1884
rect 2442 -1896 2448 -1890
rect 2442 -1902 2448 -1896
rect 2442 -1908 2448 -1902
rect 2442 -1914 2448 -1908
rect 2442 -1920 2448 -1914
rect 2442 -1926 2448 -1920
rect 2442 -1932 2448 -1926
rect 2442 -1938 2448 -1932
rect 2442 -1944 2448 -1938
rect 2442 -1950 2448 -1944
rect 2442 -1956 2448 -1950
rect 2442 -1962 2448 -1956
rect 2442 -1968 2448 -1962
rect 2442 -1974 2448 -1968
rect 2442 -1980 2448 -1974
rect 2442 -1986 2448 -1980
rect 2442 -1992 2448 -1986
rect 2442 -1998 2448 -1992
rect 2442 -2004 2448 -1998
rect 2442 -2010 2448 -2004
rect 2442 -2016 2448 -2010
rect 2442 -2022 2448 -2016
rect 2442 -2028 2448 -2022
rect 2442 -2034 2448 -2028
rect 2442 -2040 2448 -2034
rect 2442 -2046 2448 -2040
rect 2442 -2466 2448 -2460
rect 2442 -2472 2448 -2466
rect 2442 -2478 2448 -2472
rect 2442 -2484 2448 -2478
rect 2442 -2490 2448 -2484
rect 2442 -2496 2448 -2490
rect 2442 -2502 2448 -2496
rect 2442 -2508 2448 -2502
rect 2442 -2514 2448 -2508
rect 2442 -2520 2448 -2514
rect 2442 -2526 2448 -2520
rect 2442 -2532 2448 -2526
rect 2442 -2538 2448 -2532
rect 2442 -2544 2448 -2538
rect 2442 -2550 2448 -2544
rect 2442 -2556 2448 -2550
rect 2442 -2562 2448 -2556
rect 2442 -2568 2448 -2562
rect 2442 -2574 2448 -2568
rect 2442 -2580 2448 -2574
rect 2442 -2586 2448 -2580
rect 2442 -2592 2448 -2586
rect 2442 -2598 2448 -2592
rect 2442 -2604 2448 -2598
rect 2442 -2610 2448 -2604
rect 2442 -2616 2448 -2610
rect 2442 -2622 2448 -2616
rect 2442 -2628 2448 -2622
rect 2442 -2634 2448 -2628
rect 2442 -2640 2448 -2634
rect 2442 -2646 2448 -2640
rect 2442 -2652 2448 -2646
rect 2442 -2658 2448 -2652
rect 2442 -2664 2448 -2658
rect 2442 -2670 2448 -2664
rect 2442 -2676 2448 -2670
rect 2442 -2682 2448 -2676
rect 2442 -2688 2448 -2682
rect 2442 -2694 2448 -2688
rect 2442 -2700 2448 -2694
rect 2442 -2706 2448 -2700
rect 2442 -2712 2448 -2706
rect 2442 -2718 2448 -2712
rect 2442 -2724 2448 -2718
rect 2442 -2730 2448 -2724
rect 2442 -2736 2448 -2730
rect 2442 -2742 2448 -2736
rect 2442 -2748 2448 -2742
rect 2442 -2754 2448 -2748
rect 2442 -2760 2448 -2754
rect 2442 -2766 2448 -2760
rect 2442 -2772 2448 -2766
rect 2442 -2778 2448 -2772
rect 2442 -2784 2448 -2778
rect 2442 -2790 2448 -2784
rect 2442 -2796 2448 -2790
rect 2442 -2802 2448 -2796
rect 2442 -2808 2448 -2802
rect 2442 -2814 2448 -2808
rect 2442 -2820 2448 -2814
rect 2442 -2826 2448 -2820
rect 2442 -2832 2448 -2826
rect 2442 -2838 2448 -2832
rect 2442 -2844 2448 -2838
rect 2442 -2850 2448 -2844
rect 2442 -2856 2448 -2850
rect 2442 -2862 2448 -2856
rect 2448 -1350 2454 -1344
rect 2448 -1356 2454 -1350
rect 2448 -1362 2454 -1356
rect 2448 -1368 2454 -1362
rect 2448 -1374 2454 -1368
rect 2448 -1380 2454 -1374
rect 2448 -1386 2454 -1380
rect 2448 -1392 2454 -1386
rect 2448 -1398 2454 -1392
rect 2448 -1404 2454 -1398
rect 2448 -1410 2454 -1404
rect 2448 -1416 2454 -1410
rect 2448 -1422 2454 -1416
rect 2448 -1428 2454 -1422
rect 2448 -1434 2454 -1428
rect 2448 -1440 2454 -1434
rect 2448 -1446 2454 -1440
rect 2448 -1452 2454 -1446
rect 2448 -1458 2454 -1452
rect 2448 -1464 2454 -1458
rect 2448 -1470 2454 -1464
rect 2448 -1476 2454 -1470
rect 2448 -1482 2454 -1476
rect 2448 -1488 2454 -1482
rect 2448 -1494 2454 -1488
rect 2448 -1500 2454 -1494
rect 2448 -1506 2454 -1500
rect 2448 -1512 2454 -1506
rect 2448 -1518 2454 -1512
rect 2448 -1524 2454 -1518
rect 2448 -1530 2454 -1524
rect 2448 -1536 2454 -1530
rect 2448 -1542 2454 -1536
rect 2448 -1548 2454 -1542
rect 2448 -1554 2454 -1548
rect 2448 -1560 2454 -1554
rect 2448 -1566 2454 -1560
rect 2448 -1572 2454 -1566
rect 2448 -1578 2454 -1572
rect 2448 -1584 2454 -1578
rect 2448 -1590 2454 -1584
rect 2448 -1596 2454 -1590
rect 2448 -1602 2454 -1596
rect 2448 -1608 2454 -1602
rect 2448 -1614 2454 -1608
rect 2448 -1620 2454 -1614
rect 2448 -1626 2454 -1620
rect 2448 -1632 2454 -1626
rect 2448 -1638 2454 -1632
rect 2448 -1644 2454 -1638
rect 2448 -1650 2454 -1644
rect 2448 -1656 2454 -1650
rect 2448 -1662 2454 -1656
rect 2448 -1668 2454 -1662
rect 2448 -1674 2454 -1668
rect 2448 -1680 2454 -1674
rect 2448 -1686 2454 -1680
rect 2448 -1692 2454 -1686
rect 2448 -1698 2454 -1692
rect 2448 -1704 2454 -1698
rect 2448 -1710 2454 -1704
rect 2448 -1716 2454 -1710
rect 2448 -1722 2454 -1716
rect 2448 -1728 2454 -1722
rect 2448 -1734 2454 -1728
rect 2448 -1740 2454 -1734
rect 2448 -1746 2454 -1740
rect 2448 -1752 2454 -1746
rect 2448 -1758 2454 -1752
rect 2448 -1764 2454 -1758
rect 2448 -1770 2454 -1764
rect 2448 -1776 2454 -1770
rect 2448 -1782 2454 -1776
rect 2448 -1788 2454 -1782
rect 2448 -1794 2454 -1788
rect 2448 -1800 2454 -1794
rect 2448 -1806 2454 -1800
rect 2448 -1812 2454 -1806
rect 2448 -1818 2454 -1812
rect 2448 -1824 2454 -1818
rect 2448 -1830 2454 -1824
rect 2448 -1836 2454 -1830
rect 2448 -1842 2454 -1836
rect 2448 -1848 2454 -1842
rect 2448 -1854 2454 -1848
rect 2448 -1860 2454 -1854
rect 2448 -1866 2454 -1860
rect 2448 -1872 2454 -1866
rect 2448 -1878 2454 -1872
rect 2448 -1884 2454 -1878
rect 2448 -1890 2454 -1884
rect 2448 -1896 2454 -1890
rect 2448 -1902 2454 -1896
rect 2448 -1908 2454 -1902
rect 2448 -1914 2454 -1908
rect 2448 -1920 2454 -1914
rect 2448 -1926 2454 -1920
rect 2448 -1932 2454 -1926
rect 2448 -1938 2454 -1932
rect 2448 -1944 2454 -1938
rect 2448 -1950 2454 -1944
rect 2448 -1956 2454 -1950
rect 2448 -1962 2454 -1956
rect 2448 -1968 2454 -1962
rect 2448 -1974 2454 -1968
rect 2448 -1980 2454 -1974
rect 2448 -1986 2454 -1980
rect 2448 -1992 2454 -1986
rect 2448 -1998 2454 -1992
rect 2448 -2004 2454 -1998
rect 2448 -2010 2454 -2004
rect 2448 -2016 2454 -2010
rect 2448 -2022 2454 -2016
rect 2448 -2028 2454 -2022
rect 2448 -2034 2454 -2028
rect 2448 -2040 2454 -2034
rect 2448 -2466 2454 -2460
rect 2448 -2472 2454 -2466
rect 2448 -2478 2454 -2472
rect 2448 -2484 2454 -2478
rect 2448 -2490 2454 -2484
rect 2448 -2496 2454 -2490
rect 2448 -2502 2454 -2496
rect 2448 -2508 2454 -2502
rect 2448 -2514 2454 -2508
rect 2448 -2520 2454 -2514
rect 2448 -2526 2454 -2520
rect 2448 -2532 2454 -2526
rect 2448 -2538 2454 -2532
rect 2448 -2544 2454 -2538
rect 2448 -2550 2454 -2544
rect 2448 -2556 2454 -2550
rect 2448 -2562 2454 -2556
rect 2448 -2568 2454 -2562
rect 2448 -2574 2454 -2568
rect 2448 -2580 2454 -2574
rect 2448 -2586 2454 -2580
rect 2448 -2592 2454 -2586
rect 2448 -2598 2454 -2592
rect 2448 -2604 2454 -2598
rect 2448 -2610 2454 -2604
rect 2448 -2616 2454 -2610
rect 2448 -2622 2454 -2616
rect 2448 -2628 2454 -2622
rect 2448 -2634 2454 -2628
rect 2448 -2640 2454 -2634
rect 2448 -2646 2454 -2640
rect 2448 -2652 2454 -2646
rect 2448 -2658 2454 -2652
rect 2448 -2664 2454 -2658
rect 2448 -2670 2454 -2664
rect 2448 -2676 2454 -2670
rect 2448 -2682 2454 -2676
rect 2448 -2688 2454 -2682
rect 2448 -2694 2454 -2688
rect 2448 -2700 2454 -2694
rect 2448 -2706 2454 -2700
rect 2448 -2712 2454 -2706
rect 2448 -2718 2454 -2712
rect 2448 -2724 2454 -2718
rect 2448 -2730 2454 -2724
rect 2448 -2736 2454 -2730
rect 2448 -2742 2454 -2736
rect 2448 -2748 2454 -2742
rect 2448 -2754 2454 -2748
rect 2448 -2760 2454 -2754
rect 2448 -2766 2454 -2760
rect 2448 -2772 2454 -2766
rect 2448 -2778 2454 -2772
rect 2448 -2784 2454 -2778
rect 2448 -2790 2454 -2784
rect 2448 -2796 2454 -2790
rect 2448 -2802 2454 -2796
rect 2448 -2808 2454 -2802
rect 2448 -2814 2454 -2808
rect 2448 -2820 2454 -2814
rect 2448 -2826 2454 -2820
rect 2448 -2832 2454 -2826
rect 2448 -2838 2454 -2832
rect 2448 -2844 2454 -2838
rect 2448 -2850 2454 -2844
rect 2448 -2856 2454 -2850
rect 2454 -1344 2460 -1338
rect 2454 -1350 2460 -1344
rect 2454 -1356 2460 -1350
rect 2454 -1362 2460 -1356
rect 2454 -1368 2460 -1362
rect 2454 -1374 2460 -1368
rect 2454 -1380 2460 -1374
rect 2454 -1386 2460 -1380
rect 2454 -1392 2460 -1386
rect 2454 -1398 2460 -1392
rect 2454 -1404 2460 -1398
rect 2454 -1410 2460 -1404
rect 2454 -1416 2460 -1410
rect 2454 -1422 2460 -1416
rect 2454 -1428 2460 -1422
rect 2454 -1434 2460 -1428
rect 2454 -1440 2460 -1434
rect 2454 -1446 2460 -1440
rect 2454 -1452 2460 -1446
rect 2454 -1458 2460 -1452
rect 2454 -1464 2460 -1458
rect 2454 -1470 2460 -1464
rect 2454 -1476 2460 -1470
rect 2454 -1482 2460 -1476
rect 2454 -1488 2460 -1482
rect 2454 -1494 2460 -1488
rect 2454 -1500 2460 -1494
rect 2454 -1506 2460 -1500
rect 2454 -1512 2460 -1506
rect 2454 -1518 2460 -1512
rect 2454 -1524 2460 -1518
rect 2454 -1530 2460 -1524
rect 2454 -1536 2460 -1530
rect 2454 -1542 2460 -1536
rect 2454 -1548 2460 -1542
rect 2454 -1554 2460 -1548
rect 2454 -1560 2460 -1554
rect 2454 -1566 2460 -1560
rect 2454 -1572 2460 -1566
rect 2454 -1578 2460 -1572
rect 2454 -1584 2460 -1578
rect 2454 -1590 2460 -1584
rect 2454 -1596 2460 -1590
rect 2454 -1602 2460 -1596
rect 2454 -1608 2460 -1602
rect 2454 -1614 2460 -1608
rect 2454 -1620 2460 -1614
rect 2454 -1626 2460 -1620
rect 2454 -1632 2460 -1626
rect 2454 -1638 2460 -1632
rect 2454 -1644 2460 -1638
rect 2454 -1650 2460 -1644
rect 2454 -1656 2460 -1650
rect 2454 -1662 2460 -1656
rect 2454 -1668 2460 -1662
rect 2454 -1674 2460 -1668
rect 2454 -1680 2460 -1674
rect 2454 -1686 2460 -1680
rect 2454 -1692 2460 -1686
rect 2454 -1698 2460 -1692
rect 2454 -1704 2460 -1698
rect 2454 -1710 2460 -1704
rect 2454 -1716 2460 -1710
rect 2454 -1722 2460 -1716
rect 2454 -1728 2460 -1722
rect 2454 -1734 2460 -1728
rect 2454 -1740 2460 -1734
rect 2454 -1746 2460 -1740
rect 2454 -1752 2460 -1746
rect 2454 -1758 2460 -1752
rect 2454 -1764 2460 -1758
rect 2454 -1770 2460 -1764
rect 2454 -1776 2460 -1770
rect 2454 -1782 2460 -1776
rect 2454 -1788 2460 -1782
rect 2454 -1794 2460 -1788
rect 2454 -1800 2460 -1794
rect 2454 -1806 2460 -1800
rect 2454 -1812 2460 -1806
rect 2454 -1818 2460 -1812
rect 2454 -1824 2460 -1818
rect 2454 -1830 2460 -1824
rect 2454 -1836 2460 -1830
rect 2454 -1842 2460 -1836
rect 2454 -1848 2460 -1842
rect 2454 -1854 2460 -1848
rect 2454 -1860 2460 -1854
rect 2454 -1866 2460 -1860
rect 2454 -1872 2460 -1866
rect 2454 -1878 2460 -1872
rect 2454 -1884 2460 -1878
rect 2454 -1890 2460 -1884
rect 2454 -1896 2460 -1890
rect 2454 -1902 2460 -1896
rect 2454 -1908 2460 -1902
rect 2454 -1914 2460 -1908
rect 2454 -1920 2460 -1914
rect 2454 -1926 2460 -1920
rect 2454 -1932 2460 -1926
rect 2454 -1938 2460 -1932
rect 2454 -1944 2460 -1938
rect 2454 -1950 2460 -1944
rect 2454 -1956 2460 -1950
rect 2454 -1962 2460 -1956
rect 2454 -1968 2460 -1962
rect 2454 -1974 2460 -1968
rect 2454 -1980 2460 -1974
rect 2454 -1986 2460 -1980
rect 2454 -1992 2460 -1986
rect 2454 -1998 2460 -1992
rect 2454 -2004 2460 -1998
rect 2454 -2010 2460 -2004
rect 2454 -2016 2460 -2010
rect 2454 -2022 2460 -2016
rect 2454 -2028 2460 -2022
rect 2454 -2034 2460 -2028
rect 2454 -2460 2460 -2454
rect 2454 -2466 2460 -2460
rect 2454 -2472 2460 -2466
rect 2454 -2478 2460 -2472
rect 2454 -2484 2460 -2478
rect 2454 -2490 2460 -2484
rect 2454 -2496 2460 -2490
rect 2454 -2502 2460 -2496
rect 2454 -2508 2460 -2502
rect 2454 -2514 2460 -2508
rect 2454 -2520 2460 -2514
rect 2454 -2526 2460 -2520
rect 2454 -2532 2460 -2526
rect 2454 -2538 2460 -2532
rect 2454 -2544 2460 -2538
rect 2454 -2550 2460 -2544
rect 2454 -2556 2460 -2550
rect 2454 -2562 2460 -2556
rect 2454 -2568 2460 -2562
rect 2454 -2574 2460 -2568
rect 2454 -2580 2460 -2574
rect 2454 -2586 2460 -2580
rect 2454 -2592 2460 -2586
rect 2454 -2598 2460 -2592
rect 2454 -2604 2460 -2598
rect 2454 -2610 2460 -2604
rect 2454 -2616 2460 -2610
rect 2454 -2622 2460 -2616
rect 2454 -2628 2460 -2622
rect 2454 -2634 2460 -2628
rect 2454 -2640 2460 -2634
rect 2454 -2646 2460 -2640
rect 2454 -2652 2460 -2646
rect 2454 -2658 2460 -2652
rect 2454 -2664 2460 -2658
rect 2454 -2670 2460 -2664
rect 2454 -2676 2460 -2670
rect 2454 -2682 2460 -2676
rect 2454 -2688 2460 -2682
rect 2454 -2694 2460 -2688
rect 2454 -2700 2460 -2694
rect 2454 -2706 2460 -2700
rect 2454 -2712 2460 -2706
rect 2454 -2718 2460 -2712
rect 2454 -2724 2460 -2718
rect 2454 -2730 2460 -2724
rect 2454 -2736 2460 -2730
rect 2454 -2742 2460 -2736
rect 2454 -2748 2460 -2742
rect 2454 -2754 2460 -2748
rect 2454 -2760 2460 -2754
rect 2454 -2766 2460 -2760
rect 2454 -2772 2460 -2766
rect 2454 -2778 2460 -2772
rect 2454 -2784 2460 -2778
rect 2454 -2790 2460 -2784
rect 2454 -2796 2460 -2790
rect 2454 -2802 2460 -2796
rect 2454 -2808 2460 -2802
rect 2454 -2814 2460 -2808
rect 2454 -2820 2460 -2814
rect 2454 -2826 2460 -2820
rect 2454 -2832 2460 -2826
rect 2454 -2838 2460 -2832
rect 2454 -2844 2460 -2838
rect 2454 -2850 2460 -2844
rect 2454 -2856 2460 -2850
rect 2460 -1338 2466 -1332
rect 2460 -1344 2466 -1338
rect 2460 -1350 2466 -1344
rect 2460 -1356 2466 -1350
rect 2460 -1362 2466 -1356
rect 2460 -1368 2466 -1362
rect 2460 -1374 2466 -1368
rect 2460 -1380 2466 -1374
rect 2460 -1386 2466 -1380
rect 2460 -1392 2466 -1386
rect 2460 -1398 2466 -1392
rect 2460 -1404 2466 -1398
rect 2460 -1410 2466 -1404
rect 2460 -1416 2466 -1410
rect 2460 -1422 2466 -1416
rect 2460 -1428 2466 -1422
rect 2460 -1434 2466 -1428
rect 2460 -1440 2466 -1434
rect 2460 -1446 2466 -1440
rect 2460 -1452 2466 -1446
rect 2460 -1458 2466 -1452
rect 2460 -1464 2466 -1458
rect 2460 -1470 2466 -1464
rect 2460 -1476 2466 -1470
rect 2460 -1482 2466 -1476
rect 2460 -1488 2466 -1482
rect 2460 -1494 2466 -1488
rect 2460 -1500 2466 -1494
rect 2460 -1506 2466 -1500
rect 2460 -1512 2466 -1506
rect 2460 -1518 2466 -1512
rect 2460 -1524 2466 -1518
rect 2460 -1530 2466 -1524
rect 2460 -1536 2466 -1530
rect 2460 -1542 2466 -1536
rect 2460 -1548 2466 -1542
rect 2460 -1554 2466 -1548
rect 2460 -1560 2466 -1554
rect 2460 -1566 2466 -1560
rect 2460 -1572 2466 -1566
rect 2460 -1578 2466 -1572
rect 2460 -1584 2466 -1578
rect 2460 -1590 2466 -1584
rect 2460 -1596 2466 -1590
rect 2460 -1602 2466 -1596
rect 2460 -1608 2466 -1602
rect 2460 -1614 2466 -1608
rect 2460 -1620 2466 -1614
rect 2460 -1626 2466 -1620
rect 2460 -1632 2466 -1626
rect 2460 -1638 2466 -1632
rect 2460 -1644 2466 -1638
rect 2460 -1650 2466 -1644
rect 2460 -1656 2466 -1650
rect 2460 -1662 2466 -1656
rect 2460 -1668 2466 -1662
rect 2460 -1674 2466 -1668
rect 2460 -1680 2466 -1674
rect 2460 -1686 2466 -1680
rect 2460 -1692 2466 -1686
rect 2460 -1698 2466 -1692
rect 2460 -1704 2466 -1698
rect 2460 -1710 2466 -1704
rect 2460 -1716 2466 -1710
rect 2460 -1722 2466 -1716
rect 2460 -1728 2466 -1722
rect 2460 -1734 2466 -1728
rect 2460 -1740 2466 -1734
rect 2460 -1746 2466 -1740
rect 2460 -1752 2466 -1746
rect 2460 -1758 2466 -1752
rect 2460 -1764 2466 -1758
rect 2460 -1770 2466 -1764
rect 2460 -1776 2466 -1770
rect 2460 -1782 2466 -1776
rect 2460 -1788 2466 -1782
rect 2460 -1794 2466 -1788
rect 2460 -1800 2466 -1794
rect 2460 -1806 2466 -1800
rect 2460 -1812 2466 -1806
rect 2460 -1818 2466 -1812
rect 2460 -1824 2466 -1818
rect 2460 -1830 2466 -1824
rect 2460 -1836 2466 -1830
rect 2460 -1842 2466 -1836
rect 2460 -1848 2466 -1842
rect 2460 -1854 2466 -1848
rect 2460 -1860 2466 -1854
rect 2460 -1866 2466 -1860
rect 2460 -1872 2466 -1866
rect 2460 -1878 2466 -1872
rect 2460 -1884 2466 -1878
rect 2460 -1890 2466 -1884
rect 2460 -1896 2466 -1890
rect 2460 -1902 2466 -1896
rect 2460 -1908 2466 -1902
rect 2460 -1914 2466 -1908
rect 2460 -1920 2466 -1914
rect 2460 -1926 2466 -1920
rect 2460 -1932 2466 -1926
rect 2460 -1938 2466 -1932
rect 2460 -1944 2466 -1938
rect 2460 -1950 2466 -1944
rect 2460 -1956 2466 -1950
rect 2460 -1962 2466 -1956
rect 2460 -1968 2466 -1962
rect 2460 -1974 2466 -1968
rect 2460 -1980 2466 -1974
rect 2460 -1986 2466 -1980
rect 2460 -1992 2466 -1986
rect 2460 -1998 2466 -1992
rect 2460 -2004 2466 -1998
rect 2460 -2010 2466 -2004
rect 2460 -2016 2466 -2010
rect 2460 -2022 2466 -2016
rect 2460 -2460 2466 -2454
rect 2460 -2466 2466 -2460
rect 2460 -2472 2466 -2466
rect 2460 -2478 2466 -2472
rect 2460 -2484 2466 -2478
rect 2460 -2490 2466 -2484
rect 2460 -2496 2466 -2490
rect 2460 -2502 2466 -2496
rect 2460 -2508 2466 -2502
rect 2460 -2514 2466 -2508
rect 2460 -2520 2466 -2514
rect 2460 -2526 2466 -2520
rect 2460 -2532 2466 -2526
rect 2460 -2538 2466 -2532
rect 2460 -2544 2466 -2538
rect 2460 -2550 2466 -2544
rect 2460 -2556 2466 -2550
rect 2460 -2562 2466 -2556
rect 2460 -2568 2466 -2562
rect 2460 -2574 2466 -2568
rect 2460 -2580 2466 -2574
rect 2460 -2586 2466 -2580
rect 2460 -2592 2466 -2586
rect 2460 -2598 2466 -2592
rect 2460 -2604 2466 -2598
rect 2460 -2610 2466 -2604
rect 2460 -2616 2466 -2610
rect 2460 -2622 2466 -2616
rect 2460 -2628 2466 -2622
rect 2460 -2634 2466 -2628
rect 2460 -2640 2466 -2634
rect 2460 -2646 2466 -2640
rect 2460 -2652 2466 -2646
rect 2460 -2658 2466 -2652
rect 2460 -2664 2466 -2658
rect 2460 -2670 2466 -2664
rect 2460 -2676 2466 -2670
rect 2460 -2682 2466 -2676
rect 2460 -2688 2466 -2682
rect 2460 -2694 2466 -2688
rect 2460 -2700 2466 -2694
rect 2460 -2706 2466 -2700
rect 2460 -2712 2466 -2706
rect 2460 -2718 2466 -2712
rect 2460 -2724 2466 -2718
rect 2460 -2730 2466 -2724
rect 2460 -2736 2466 -2730
rect 2460 -2742 2466 -2736
rect 2460 -2748 2466 -2742
rect 2460 -2754 2466 -2748
rect 2460 -2760 2466 -2754
rect 2460 -2766 2466 -2760
rect 2460 -2772 2466 -2766
rect 2460 -2778 2466 -2772
rect 2460 -2784 2466 -2778
rect 2460 -2790 2466 -2784
rect 2460 -2796 2466 -2790
rect 2460 -2802 2466 -2796
rect 2460 -2808 2466 -2802
rect 2460 -2814 2466 -2808
rect 2460 -2820 2466 -2814
rect 2460 -2826 2466 -2820
rect 2460 -2832 2466 -2826
rect 2460 -2838 2466 -2832
rect 2460 -2844 2466 -2838
rect 2460 -2850 2466 -2844
rect 2466 -1332 2472 -1326
rect 2466 -1338 2472 -1332
rect 2466 -1344 2472 -1338
rect 2466 -1350 2472 -1344
rect 2466 -1356 2472 -1350
rect 2466 -1362 2472 -1356
rect 2466 -1368 2472 -1362
rect 2466 -1374 2472 -1368
rect 2466 -1380 2472 -1374
rect 2466 -1386 2472 -1380
rect 2466 -1392 2472 -1386
rect 2466 -1398 2472 -1392
rect 2466 -1404 2472 -1398
rect 2466 -1410 2472 -1404
rect 2466 -1416 2472 -1410
rect 2466 -1422 2472 -1416
rect 2466 -1428 2472 -1422
rect 2466 -1434 2472 -1428
rect 2466 -1440 2472 -1434
rect 2466 -1446 2472 -1440
rect 2466 -1452 2472 -1446
rect 2466 -1458 2472 -1452
rect 2466 -1464 2472 -1458
rect 2466 -1470 2472 -1464
rect 2466 -1476 2472 -1470
rect 2466 -1482 2472 -1476
rect 2466 -1488 2472 -1482
rect 2466 -1494 2472 -1488
rect 2466 -1500 2472 -1494
rect 2466 -1506 2472 -1500
rect 2466 -1512 2472 -1506
rect 2466 -1518 2472 -1512
rect 2466 -1524 2472 -1518
rect 2466 -1530 2472 -1524
rect 2466 -1536 2472 -1530
rect 2466 -1542 2472 -1536
rect 2466 -1548 2472 -1542
rect 2466 -1554 2472 -1548
rect 2466 -1560 2472 -1554
rect 2466 -1566 2472 -1560
rect 2466 -1572 2472 -1566
rect 2466 -1578 2472 -1572
rect 2466 -1584 2472 -1578
rect 2466 -1590 2472 -1584
rect 2466 -1596 2472 -1590
rect 2466 -1602 2472 -1596
rect 2466 -1608 2472 -1602
rect 2466 -1614 2472 -1608
rect 2466 -1620 2472 -1614
rect 2466 -1626 2472 -1620
rect 2466 -1632 2472 -1626
rect 2466 -1638 2472 -1632
rect 2466 -1644 2472 -1638
rect 2466 -1650 2472 -1644
rect 2466 -1656 2472 -1650
rect 2466 -1662 2472 -1656
rect 2466 -1668 2472 -1662
rect 2466 -1674 2472 -1668
rect 2466 -1680 2472 -1674
rect 2466 -1686 2472 -1680
rect 2466 -1692 2472 -1686
rect 2466 -1698 2472 -1692
rect 2466 -1704 2472 -1698
rect 2466 -1710 2472 -1704
rect 2466 -1716 2472 -1710
rect 2466 -1722 2472 -1716
rect 2466 -1728 2472 -1722
rect 2466 -1734 2472 -1728
rect 2466 -1740 2472 -1734
rect 2466 -1746 2472 -1740
rect 2466 -1752 2472 -1746
rect 2466 -1758 2472 -1752
rect 2466 -1764 2472 -1758
rect 2466 -1770 2472 -1764
rect 2466 -1776 2472 -1770
rect 2466 -1782 2472 -1776
rect 2466 -1788 2472 -1782
rect 2466 -1794 2472 -1788
rect 2466 -1800 2472 -1794
rect 2466 -1806 2472 -1800
rect 2466 -1812 2472 -1806
rect 2466 -1818 2472 -1812
rect 2466 -1824 2472 -1818
rect 2466 -1830 2472 -1824
rect 2466 -1836 2472 -1830
rect 2466 -1842 2472 -1836
rect 2466 -1848 2472 -1842
rect 2466 -1854 2472 -1848
rect 2466 -1860 2472 -1854
rect 2466 -1866 2472 -1860
rect 2466 -1872 2472 -1866
rect 2466 -1878 2472 -1872
rect 2466 -1884 2472 -1878
rect 2466 -1890 2472 -1884
rect 2466 -1896 2472 -1890
rect 2466 -1902 2472 -1896
rect 2466 -1908 2472 -1902
rect 2466 -1914 2472 -1908
rect 2466 -1920 2472 -1914
rect 2466 -1926 2472 -1920
rect 2466 -1932 2472 -1926
rect 2466 -1938 2472 -1932
rect 2466 -1944 2472 -1938
rect 2466 -1950 2472 -1944
rect 2466 -1956 2472 -1950
rect 2466 -1962 2472 -1956
rect 2466 -1968 2472 -1962
rect 2466 -1974 2472 -1968
rect 2466 -1980 2472 -1974
rect 2466 -1986 2472 -1980
rect 2466 -1992 2472 -1986
rect 2466 -1998 2472 -1992
rect 2466 -2004 2472 -1998
rect 2466 -2010 2472 -2004
rect 2466 -2016 2472 -2010
rect 2466 -2460 2472 -2454
rect 2466 -2466 2472 -2460
rect 2466 -2472 2472 -2466
rect 2466 -2478 2472 -2472
rect 2466 -2484 2472 -2478
rect 2466 -2490 2472 -2484
rect 2466 -2496 2472 -2490
rect 2466 -2502 2472 -2496
rect 2466 -2508 2472 -2502
rect 2466 -2514 2472 -2508
rect 2466 -2520 2472 -2514
rect 2466 -2526 2472 -2520
rect 2466 -2532 2472 -2526
rect 2466 -2538 2472 -2532
rect 2466 -2544 2472 -2538
rect 2466 -2550 2472 -2544
rect 2466 -2556 2472 -2550
rect 2466 -2562 2472 -2556
rect 2466 -2568 2472 -2562
rect 2466 -2574 2472 -2568
rect 2466 -2580 2472 -2574
rect 2466 -2586 2472 -2580
rect 2466 -2592 2472 -2586
rect 2466 -2598 2472 -2592
rect 2466 -2604 2472 -2598
rect 2466 -2610 2472 -2604
rect 2466 -2616 2472 -2610
rect 2466 -2622 2472 -2616
rect 2466 -2628 2472 -2622
rect 2466 -2634 2472 -2628
rect 2466 -2640 2472 -2634
rect 2466 -2646 2472 -2640
rect 2466 -2652 2472 -2646
rect 2466 -2658 2472 -2652
rect 2466 -2664 2472 -2658
rect 2466 -2670 2472 -2664
rect 2466 -2676 2472 -2670
rect 2466 -2682 2472 -2676
rect 2466 -2688 2472 -2682
rect 2466 -2694 2472 -2688
rect 2466 -2700 2472 -2694
rect 2466 -2706 2472 -2700
rect 2466 -2712 2472 -2706
rect 2466 -2718 2472 -2712
rect 2466 -2724 2472 -2718
rect 2466 -2730 2472 -2724
rect 2466 -2736 2472 -2730
rect 2466 -2742 2472 -2736
rect 2466 -2748 2472 -2742
rect 2466 -2754 2472 -2748
rect 2466 -2760 2472 -2754
rect 2466 -2766 2472 -2760
rect 2466 -2772 2472 -2766
rect 2466 -2778 2472 -2772
rect 2466 -2784 2472 -2778
rect 2466 -2790 2472 -2784
rect 2466 -2796 2472 -2790
rect 2466 -2802 2472 -2796
rect 2466 -2808 2472 -2802
rect 2466 -2814 2472 -2808
rect 2466 -2820 2472 -2814
rect 2466 -2826 2472 -2820
rect 2466 -2832 2472 -2826
rect 2466 -2838 2472 -2832
rect 2466 -2844 2472 -2838
rect 2472 -1332 2478 -1326
rect 2472 -1338 2478 -1332
rect 2472 -1344 2478 -1338
rect 2472 -1350 2478 -1344
rect 2472 -1356 2478 -1350
rect 2472 -1362 2478 -1356
rect 2472 -1368 2478 -1362
rect 2472 -1374 2478 -1368
rect 2472 -1380 2478 -1374
rect 2472 -1386 2478 -1380
rect 2472 -1392 2478 -1386
rect 2472 -1398 2478 -1392
rect 2472 -1404 2478 -1398
rect 2472 -1410 2478 -1404
rect 2472 -1416 2478 -1410
rect 2472 -1422 2478 -1416
rect 2472 -1428 2478 -1422
rect 2472 -1434 2478 -1428
rect 2472 -1440 2478 -1434
rect 2472 -1446 2478 -1440
rect 2472 -1452 2478 -1446
rect 2472 -1458 2478 -1452
rect 2472 -1464 2478 -1458
rect 2472 -1470 2478 -1464
rect 2472 -1476 2478 -1470
rect 2472 -1482 2478 -1476
rect 2472 -1488 2478 -1482
rect 2472 -1494 2478 -1488
rect 2472 -1500 2478 -1494
rect 2472 -1506 2478 -1500
rect 2472 -1512 2478 -1506
rect 2472 -1518 2478 -1512
rect 2472 -1524 2478 -1518
rect 2472 -1530 2478 -1524
rect 2472 -1536 2478 -1530
rect 2472 -1542 2478 -1536
rect 2472 -1548 2478 -1542
rect 2472 -1554 2478 -1548
rect 2472 -1560 2478 -1554
rect 2472 -1566 2478 -1560
rect 2472 -1572 2478 -1566
rect 2472 -1578 2478 -1572
rect 2472 -1584 2478 -1578
rect 2472 -1590 2478 -1584
rect 2472 -1596 2478 -1590
rect 2472 -1602 2478 -1596
rect 2472 -1608 2478 -1602
rect 2472 -1614 2478 -1608
rect 2472 -1620 2478 -1614
rect 2472 -1626 2478 -1620
rect 2472 -1632 2478 -1626
rect 2472 -1638 2478 -1632
rect 2472 -1644 2478 -1638
rect 2472 -1650 2478 -1644
rect 2472 -1656 2478 -1650
rect 2472 -1662 2478 -1656
rect 2472 -1668 2478 -1662
rect 2472 -1674 2478 -1668
rect 2472 -1680 2478 -1674
rect 2472 -1686 2478 -1680
rect 2472 -1692 2478 -1686
rect 2472 -1698 2478 -1692
rect 2472 -1704 2478 -1698
rect 2472 -1710 2478 -1704
rect 2472 -1716 2478 -1710
rect 2472 -1722 2478 -1716
rect 2472 -1728 2478 -1722
rect 2472 -1734 2478 -1728
rect 2472 -1740 2478 -1734
rect 2472 -1746 2478 -1740
rect 2472 -1752 2478 -1746
rect 2472 -1758 2478 -1752
rect 2472 -1764 2478 -1758
rect 2472 -1770 2478 -1764
rect 2472 -1776 2478 -1770
rect 2472 -1782 2478 -1776
rect 2472 -1788 2478 -1782
rect 2472 -1794 2478 -1788
rect 2472 -1800 2478 -1794
rect 2472 -1806 2478 -1800
rect 2472 -1812 2478 -1806
rect 2472 -1818 2478 -1812
rect 2472 -1824 2478 -1818
rect 2472 -1830 2478 -1824
rect 2472 -1836 2478 -1830
rect 2472 -1842 2478 -1836
rect 2472 -1848 2478 -1842
rect 2472 -1854 2478 -1848
rect 2472 -1860 2478 -1854
rect 2472 -1866 2478 -1860
rect 2472 -1872 2478 -1866
rect 2472 -1878 2478 -1872
rect 2472 -1884 2478 -1878
rect 2472 -1890 2478 -1884
rect 2472 -1896 2478 -1890
rect 2472 -1902 2478 -1896
rect 2472 -1908 2478 -1902
rect 2472 -1914 2478 -1908
rect 2472 -1920 2478 -1914
rect 2472 -1926 2478 -1920
rect 2472 -1932 2478 -1926
rect 2472 -1938 2478 -1932
rect 2472 -1944 2478 -1938
rect 2472 -1950 2478 -1944
rect 2472 -1956 2478 -1950
rect 2472 -1962 2478 -1956
rect 2472 -1968 2478 -1962
rect 2472 -1974 2478 -1968
rect 2472 -1980 2478 -1974
rect 2472 -1986 2478 -1980
rect 2472 -1992 2478 -1986
rect 2472 -1998 2478 -1992
rect 2472 -2004 2478 -1998
rect 2472 -2010 2478 -2004
rect 2472 -2460 2478 -2454
rect 2472 -2466 2478 -2460
rect 2472 -2472 2478 -2466
rect 2472 -2478 2478 -2472
rect 2472 -2484 2478 -2478
rect 2472 -2490 2478 -2484
rect 2472 -2496 2478 -2490
rect 2472 -2502 2478 -2496
rect 2472 -2508 2478 -2502
rect 2472 -2514 2478 -2508
rect 2472 -2520 2478 -2514
rect 2472 -2526 2478 -2520
rect 2472 -2532 2478 -2526
rect 2472 -2538 2478 -2532
rect 2472 -2544 2478 -2538
rect 2472 -2550 2478 -2544
rect 2472 -2556 2478 -2550
rect 2472 -2562 2478 -2556
rect 2472 -2568 2478 -2562
rect 2472 -2574 2478 -2568
rect 2472 -2580 2478 -2574
rect 2472 -2586 2478 -2580
rect 2472 -2592 2478 -2586
rect 2472 -2598 2478 -2592
rect 2472 -2604 2478 -2598
rect 2472 -2610 2478 -2604
rect 2472 -2616 2478 -2610
rect 2472 -2622 2478 -2616
rect 2472 -2628 2478 -2622
rect 2472 -2634 2478 -2628
rect 2472 -2640 2478 -2634
rect 2472 -2646 2478 -2640
rect 2472 -2652 2478 -2646
rect 2472 -2658 2478 -2652
rect 2472 -2664 2478 -2658
rect 2472 -2670 2478 -2664
rect 2472 -2676 2478 -2670
rect 2472 -2682 2478 -2676
rect 2472 -2688 2478 -2682
rect 2472 -2694 2478 -2688
rect 2472 -2700 2478 -2694
rect 2472 -2706 2478 -2700
rect 2472 -2712 2478 -2706
rect 2472 -2718 2478 -2712
rect 2472 -2724 2478 -2718
rect 2472 -2730 2478 -2724
rect 2472 -2736 2478 -2730
rect 2472 -2742 2478 -2736
rect 2472 -2748 2478 -2742
rect 2472 -2754 2478 -2748
rect 2472 -2760 2478 -2754
rect 2472 -2766 2478 -2760
rect 2472 -2772 2478 -2766
rect 2472 -2778 2478 -2772
rect 2472 -2784 2478 -2778
rect 2472 -2790 2478 -2784
rect 2472 -2796 2478 -2790
rect 2472 -2802 2478 -2796
rect 2472 -2808 2478 -2802
rect 2472 -2814 2478 -2808
rect 2472 -2820 2478 -2814
rect 2472 -2826 2478 -2820
rect 2472 -2832 2478 -2826
rect 2472 -2838 2478 -2832
rect 2472 -2844 2478 -2838
rect 2478 -1326 2484 -1320
rect 2478 -1332 2484 -1326
rect 2478 -1338 2484 -1332
rect 2478 -1344 2484 -1338
rect 2478 -1350 2484 -1344
rect 2478 -1356 2484 -1350
rect 2478 -1362 2484 -1356
rect 2478 -1368 2484 -1362
rect 2478 -1374 2484 -1368
rect 2478 -1380 2484 -1374
rect 2478 -1386 2484 -1380
rect 2478 -1392 2484 -1386
rect 2478 -1398 2484 -1392
rect 2478 -1404 2484 -1398
rect 2478 -1410 2484 -1404
rect 2478 -1416 2484 -1410
rect 2478 -1422 2484 -1416
rect 2478 -1428 2484 -1422
rect 2478 -1434 2484 -1428
rect 2478 -1440 2484 -1434
rect 2478 -1446 2484 -1440
rect 2478 -1452 2484 -1446
rect 2478 -1458 2484 -1452
rect 2478 -1464 2484 -1458
rect 2478 -1470 2484 -1464
rect 2478 -1476 2484 -1470
rect 2478 -1482 2484 -1476
rect 2478 -1488 2484 -1482
rect 2478 -1494 2484 -1488
rect 2478 -1500 2484 -1494
rect 2478 -1506 2484 -1500
rect 2478 -1512 2484 -1506
rect 2478 -1518 2484 -1512
rect 2478 -1524 2484 -1518
rect 2478 -1530 2484 -1524
rect 2478 -1536 2484 -1530
rect 2478 -1542 2484 -1536
rect 2478 -1548 2484 -1542
rect 2478 -1554 2484 -1548
rect 2478 -1560 2484 -1554
rect 2478 -1566 2484 -1560
rect 2478 -1572 2484 -1566
rect 2478 -1578 2484 -1572
rect 2478 -1584 2484 -1578
rect 2478 -1590 2484 -1584
rect 2478 -1596 2484 -1590
rect 2478 -1602 2484 -1596
rect 2478 -1608 2484 -1602
rect 2478 -1614 2484 -1608
rect 2478 -1620 2484 -1614
rect 2478 -1626 2484 -1620
rect 2478 -1632 2484 -1626
rect 2478 -1638 2484 -1632
rect 2478 -1644 2484 -1638
rect 2478 -1650 2484 -1644
rect 2478 -1656 2484 -1650
rect 2478 -1662 2484 -1656
rect 2478 -1668 2484 -1662
rect 2478 -1674 2484 -1668
rect 2478 -1680 2484 -1674
rect 2478 -1686 2484 -1680
rect 2478 -1692 2484 -1686
rect 2478 -1698 2484 -1692
rect 2478 -1704 2484 -1698
rect 2478 -1710 2484 -1704
rect 2478 -1716 2484 -1710
rect 2478 -1722 2484 -1716
rect 2478 -1728 2484 -1722
rect 2478 -1734 2484 -1728
rect 2478 -1740 2484 -1734
rect 2478 -1746 2484 -1740
rect 2478 -1752 2484 -1746
rect 2478 -1758 2484 -1752
rect 2478 -1764 2484 -1758
rect 2478 -1770 2484 -1764
rect 2478 -1776 2484 -1770
rect 2478 -1782 2484 -1776
rect 2478 -1788 2484 -1782
rect 2478 -1794 2484 -1788
rect 2478 -1800 2484 -1794
rect 2478 -1806 2484 -1800
rect 2478 -1812 2484 -1806
rect 2478 -1818 2484 -1812
rect 2478 -1824 2484 -1818
rect 2478 -1830 2484 -1824
rect 2478 -1836 2484 -1830
rect 2478 -1842 2484 -1836
rect 2478 -1848 2484 -1842
rect 2478 -1854 2484 -1848
rect 2478 -1860 2484 -1854
rect 2478 -1866 2484 -1860
rect 2478 -1872 2484 -1866
rect 2478 -1878 2484 -1872
rect 2478 -1884 2484 -1878
rect 2478 -1890 2484 -1884
rect 2478 -1896 2484 -1890
rect 2478 -1902 2484 -1896
rect 2478 -1908 2484 -1902
rect 2478 -1914 2484 -1908
rect 2478 -1920 2484 -1914
rect 2478 -1926 2484 -1920
rect 2478 -1932 2484 -1926
rect 2478 -1938 2484 -1932
rect 2478 -1944 2484 -1938
rect 2478 -1950 2484 -1944
rect 2478 -1956 2484 -1950
rect 2478 -1962 2484 -1956
rect 2478 -1968 2484 -1962
rect 2478 -1974 2484 -1968
rect 2478 -1980 2484 -1974
rect 2478 -1986 2484 -1980
rect 2478 -1992 2484 -1986
rect 2478 -1998 2484 -1992
rect 2478 -2004 2484 -1998
rect 2478 -2454 2484 -2448
rect 2478 -2460 2484 -2454
rect 2478 -2466 2484 -2460
rect 2478 -2472 2484 -2466
rect 2478 -2478 2484 -2472
rect 2478 -2484 2484 -2478
rect 2478 -2490 2484 -2484
rect 2478 -2496 2484 -2490
rect 2478 -2502 2484 -2496
rect 2478 -2508 2484 -2502
rect 2478 -2514 2484 -2508
rect 2478 -2520 2484 -2514
rect 2478 -2526 2484 -2520
rect 2478 -2532 2484 -2526
rect 2478 -2538 2484 -2532
rect 2478 -2544 2484 -2538
rect 2478 -2550 2484 -2544
rect 2478 -2556 2484 -2550
rect 2478 -2562 2484 -2556
rect 2478 -2568 2484 -2562
rect 2478 -2574 2484 -2568
rect 2478 -2580 2484 -2574
rect 2478 -2586 2484 -2580
rect 2478 -2592 2484 -2586
rect 2478 -2598 2484 -2592
rect 2478 -2604 2484 -2598
rect 2478 -2610 2484 -2604
rect 2478 -2616 2484 -2610
rect 2478 -2622 2484 -2616
rect 2478 -2628 2484 -2622
rect 2478 -2634 2484 -2628
rect 2478 -2640 2484 -2634
rect 2478 -2646 2484 -2640
rect 2478 -2652 2484 -2646
rect 2478 -2658 2484 -2652
rect 2478 -2664 2484 -2658
rect 2478 -2670 2484 -2664
rect 2478 -2676 2484 -2670
rect 2478 -2682 2484 -2676
rect 2478 -2688 2484 -2682
rect 2478 -2694 2484 -2688
rect 2478 -2700 2484 -2694
rect 2478 -2706 2484 -2700
rect 2478 -2712 2484 -2706
rect 2478 -2718 2484 -2712
rect 2478 -2724 2484 -2718
rect 2478 -2730 2484 -2724
rect 2478 -2736 2484 -2730
rect 2478 -2742 2484 -2736
rect 2478 -2748 2484 -2742
rect 2478 -2754 2484 -2748
rect 2478 -2760 2484 -2754
rect 2478 -2766 2484 -2760
rect 2478 -2772 2484 -2766
rect 2478 -2778 2484 -2772
rect 2478 -2784 2484 -2778
rect 2478 -2790 2484 -2784
rect 2478 -2796 2484 -2790
rect 2478 -2802 2484 -2796
rect 2478 -2808 2484 -2802
rect 2478 -2814 2484 -2808
rect 2478 -2820 2484 -2814
rect 2478 -2826 2484 -2820
rect 2478 -2832 2484 -2826
rect 2478 -2838 2484 -2832
rect 2484 -1320 2490 -1314
rect 2484 -1326 2490 -1320
rect 2484 -1332 2490 -1326
rect 2484 -1338 2490 -1332
rect 2484 -1344 2490 -1338
rect 2484 -1350 2490 -1344
rect 2484 -1356 2490 -1350
rect 2484 -1362 2490 -1356
rect 2484 -1368 2490 -1362
rect 2484 -1374 2490 -1368
rect 2484 -1380 2490 -1374
rect 2484 -1386 2490 -1380
rect 2484 -1392 2490 -1386
rect 2484 -1398 2490 -1392
rect 2484 -1404 2490 -1398
rect 2484 -1410 2490 -1404
rect 2484 -1416 2490 -1410
rect 2484 -1422 2490 -1416
rect 2484 -1428 2490 -1422
rect 2484 -1434 2490 -1428
rect 2484 -1440 2490 -1434
rect 2484 -1446 2490 -1440
rect 2484 -1452 2490 -1446
rect 2484 -1458 2490 -1452
rect 2484 -1464 2490 -1458
rect 2484 -1470 2490 -1464
rect 2484 -1476 2490 -1470
rect 2484 -1482 2490 -1476
rect 2484 -1488 2490 -1482
rect 2484 -1494 2490 -1488
rect 2484 -1500 2490 -1494
rect 2484 -1506 2490 -1500
rect 2484 -1512 2490 -1506
rect 2484 -1518 2490 -1512
rect 2484 -1524 2490 -1518
rect 2484 -1530 2490 -1524
rect 2484 -1536 2490 -1530
rect 2484 -1542 2490 -1536
rect 2484 -1548 2490 -1542
rect 2484 -1554 2490 -1548
rect 2484 -1560 2490 -1554
rect 2484 -1566 2490 -1560
rect 2484 -1572 2490 -1566
rect 2484 -1578 2490 -1572
rect 2484 -1584 2490 -1578
rect 2484 -1590 2490 -1584
rect 2484 -1596 2490 -1590
rect 2484 -1602 2490 -1596
rect 2484 -1608 2490 -1602
rect 2484 -1614 2490 -1608
rect 2484 -1620 2490 -1614
rect 2484 -1626 2490 -1620
rect 2484 -1632 2490 -1626
rect 2484 -1638 2490 -1632
rect 2484 -1644 2490 -1638
rect 2484 -1650 2490 -1644
rect 2484 -1656 2490 -1650
rect 2484 -1662 2490 -1656
rect 2484 -1668 2490 -1662
rect 2484 -1674 2490 -1668
rect 2484 -1680 2490 -1674
rect 2484 -1686 2490 -1680
rect 2484 -1692 2490 -1686
rect 2484 -1698 2490 -1692
rect 2484 -1704 2490 -1698
rect 2484 -1710 2490 -1704
rect 2484 -1716 2490 -1710
rect 2484 -1722 2490 -1716
rect 2484 -1728 2490 -1722
rect 2484 -1734 2490 -1728
rect 2484 -1740 2490 -1734
rect 2484 -1746 2490 -1740
rect 2484 -1752 2490 -1746
rect 2484 -1758 2490 -1752
rect 2484 -1764 2490 -1758
rect 2484 -1770 2490 -1764
rect 2484 -1776 2490 -1770
rect 2484 -1782 2490 -1776
rect 2484 -1788 2490 -1782
rect 2484 -1794 2490 -1788
rect 2484 -1800 2490 -1794
rect 2484 -1806 2490 -1800
rect 2484 -1812 2490 -1806
rect 2484 -1818 2490 -1812
rect 2484 -1824 2490 -1818
rect 2484 -1830 2490 -1824
rect 2484 -1836 2490 -1830
rect 2484 -1842 2490 -1836
rect 2484 -1848 2490 -1842
rect 2484 -1854 2490 -1848
rect 2484 -1860 2490 -1854
rect 2484 -1866 2490 -1860
rect 2484 -1872 2490 -1866
rect 2484 -1878 2490 -1872
rect 2484 -1884 2490 -1878
rect 2484 -1890 2490 -1884
rect 2484 -1896 2490 -1890
rect 2484 -1902 2490 -1896
rect 2484 -1908 2490 -1902
rect 2484 -1914 2490 -1908
rect 2484 -1920 2490 -1914
rect 2484 -1926 2490 -1920
rect 2484 -1932 2490 -1926
rect 2484 -1938 2490 -1932
rect 2484 -1944 2490 -1938
rect 2484 -1950 2490 -1944
rect 2484 -1956 2490 -1950
rect 2484 -1962 2490 -1956
rect 2484 -1968 2490 -1962
rect 2484 -1974 2490 -1968
rect 2484 -1980 2490 -1974
rect 2484 -1986 2490 -1980
rect 2484 -1992 2490 -1986
rect 2484 -2454 2490 -2448
rect 2484 -2460 2490 -2454
rect 2484 -2466 2490 -2460
rect 2484 -2472 2490 -2466
rect 2484 -2478 2490 -2472
rect 2484 -2484 2490 -2478
rect 2484 -2490 2490 -2484
rect 2484 -2496 2490 -2490
rect 2484 -2502 2490 -2496
rect 2484 -2508 2490 -2502
rect 2484 -2514 2490 -2508
rect 2484 -2520 2490 -2514
rect 2484 -2526 2490 -2520
rect 2484 -2532 2490 -2526
rect 2484 -2538 2490 -2532
rect 2484 -2544 2490 -2538
rect 2484 -2550 2490 -2544
rect 2484 -2556 2490 -2550
rect 2484 -2562 2490 -2556
rect 2484 -2568 2490 -2562
rect 2484 -2574 2490 -2568
rect 2484 -2580 2490 -2574
rect 2484 -2586 2490 -2580
rect 2484 -2592 2490 -2586
rect 2484 -2598 2490 -2592
rect 2484 -2604 2490 -2598
rect 2484 -2610 2490 -2604
rect 2484 -2616 2490 -2610
rect 2484 -2622 2490 -2616
rect 2484 -2628 2490 -2622
rect 2484 -2634 2490 -2628
rect 2484 -2640 2490 -2634
rect 2484 -2646 2490 -2640
rect 2484 -2652 2490 -2646
rect 2484 -2658 2490 -2652
rect 2484 -2664 2490 -2658
rect 2484 -2670 2490 -2664
rect 2484 -2676 2490 -2670
rect 2484 -2682 2490 -2676
rect 2484 -2688 2490 -2682
rect 2484 -2694 2490 -2688
rect 2484 -2700 2490 -2694
rect 2484 -2706 2490 -2700
rect 2484 -2712 2490 -2706
rect 2484 -2718 2490 -2712
rect 2484 -2724 2490 -2718
rect 2484 -2730 2490 -2724
rect 2484 -2736 2490 -2730
rect 2484 -2742 2490 -2736
rect 2484 -2748 2490 -2742
rect 2484 -2754 2490 -2748
rect 2484 -2760 2490 -2754
rect 2484 -2766 2490 -2760
rect 2484 -2772 2490 -2766
rect 2484 -2778 2490 -2772
rect 2484 -2784 2490 -2778
rect 2484 -2790 2490 -2784
rect 2484 -2796 2490 -2790
rect 2484 -2802 2490 -2796
rect 2484 -2808 2490 -2802
rect 2484 -2814 2490 -2808
rect 2484 -2820 2490 -2814
rect 2484 -2826 2490 -2820
rect 2484 -2832 2490 -2826
rect 2484 -2838 2490 -2832
rect 2490 -1314 2496 -1308
rect 2490 -1320 2496 -1314
rect 2490 -1326 2496 -1320
rect 2490 -1332 2496 -1326
rect 2490 -1338 2496 -1332
rect 2490 -1344 2496 -1338
rect 2490 -1350 2496 -1344
rect 2490 -1356 2496 -1350
rect 2490 -1362 2496 -1356
rect 2490 -1368 2496 -1362
rect 2490 -1374 2496 -1368
rect 2490 -1380 2496 -1374
rect 2490 -1386 2496 -1380
rect 2490 -1392 2496 -1386
rect 2490 -1398 2496 -1392
rect 2490 -1404 2496 -1398
rect 2490 -1410 2496 -1404
rect 2490 -1416 2496 -1410
rect 2490 -1422 2496 -1416
rect 2490 -1428 2496 -1422
rect 2490 -1434 2496 -1428
rect 2490 -1440 2496 -1434
rect 2490 -1446 2496 -1440
rect 2490 -1452 2496 -1446
rect 2490 -1458 2496 -1452
rect 2490 -1464 2496 -1458
rect 2490 -1470 2496 -1464
rect 2490 -1476 2496 -1470
rect 2490 -1482 2496 -1476
rect 2490 -1488 2496 -1482
rect 2490 -1494 2496 -1488
rect 2490 -1500 2496 -1494
rect 2490 -1506 2496 -1500
rect 2490 -1512 2496 -1506
rect 2490 -1518 2496 -1512
rect 2490 -1524 2496 -1518
rect 2490 -1530 2496 -1524
rect 2490 -1536 2496 -1530
rect 2490 -1542 2496 -1536
rect 2490 -1548 2496 -1542
rect 2490 -1554 2496 -1548
rect 2490 -1560 2496 -1554
rect 2490 -1566 2496 -1560
rect 2490 -1572 2496 -1566
rect 2490 -1578 2496 -1572
rect 2490 -1584 2496 -1578
rect 2490 -1590 2496 -1584
rect 2490 -1596 2496 -1590
rect 2490 -1602 2496 -1596
rect 2490 -1608 2496 -1602
rect 2490 -1614 2496 -1608
rect 2490 -1620 2496 -1614
rect 2490 -1626 2496 -1620
rect 2490 -1632 2496 -1626
rect 2490 -1638 2496 -1632
rect 2490 -1644 2496 -1638
rect 2490 -1650 2496 -1644
rect 2490 -1656 2496 -1650
rect 2490 -1662 2496 -1656
rect 2490 -1668 2496 -1662
rect 2490 -1674 2496 -1668
rect 2490 -1680 2496 -1674
rect 2490 -1686 2496 -1680
rect 2490 -1692 2496 -1686
rect 2490 -1698 2496 -1692
rect 2490 -1704 2496 -1698
rect 2490 -1710 2496 -1704
rect 2490 -1716 2496 -1710
rect 2490 -1722 2496 -1716
rect 2490 -1728 2496 -1722
rect 2490 -1734 2496 -1728
rect 2490 -1740 2496 -1734
rect 2490 -1746 2496 -1740
rect 2490 -1752 2496 -1746
rect 2490 -1758 2496 -1752
rect 2490 -1764 2496 -1758
rect 2490 -1770 2496 -1764
rect 2490 -1776 2496 -1770
rect 2490 -1782 2496 -1776
rect 2490 -1788 2496 -1782
rect 2490 -1794 2496 -1788
rect 2490 -1800 2496 -1794
rect 2490 -1806 2496 -1800
rect 2490 -1812 2496 -1806
rect 2490 -1818 2496 -1812
rect 2490 -1824 2496 -1818
rect 2490 -1830 2496 -1824
rect 2490 -1836 2496 -1830
rect 2490 -1842 2496 -1836
rect 2490 -1848 2496 -1842
rect 2490 -1854 2496 -1848
rect 2490 -1860 2496 -1854
rect 2490 -1866 2496 -1860
rect 2490 -1872 2496 -1866
rect 2490 -1878 2496 -1872
rect 2490 -1884 2496 -1878
rect 2490 -1890 2496 -1884
rect 2490 -1896 2496 -1890
rect 2490 -1902 2496 -1896
rect 2490 -1908 2496 -1902
rect 2490 -1914 2496 -1908
rect 2490 -1920 2496 -1914
rect 2490 -1926 2496 -1920
rect 2490 -1932 2496 -1926
rect 2490 -1938 2496 -1932
rect 2490 -1944 2496 -1938
rect 2490 -1950 2496 -1944
rect 2490 -1956 2496 -1950
rect 2490 -1962 2496 -1956
rect 2490 -1968 2496 -1962
rect 2490 -1974 2496 -1968
rect 2490 -1980 2496 -1974
rect 2490 -1986 2496 -1980
rect 2490 -2454 2496 -2448
rect 2490 -2460 2496 -2454
rect 2490 -2466 2496 -2460
rect 2490 -2472 2496 -2466
rect 2490 -2478 2496 -2472
rect 2490 -2484 2496 -2478
rect 2490 -2490 2496 -2484
rect 2490 -2496 2496 -2490
rect 2490 -2502 2496 -2496
rect 2490 -2508 2496 -2502
rect 2490 -2514 2496 -2508
rect 2490 -2520 2496 -2514
rect 2490 -2526 2496 -2520
rect 2490 -2532 2496 -2526
rect 2490 -2538 2496 -2532
rect 2490 -2544 2496 -2538
rect 2490 -2550 2496 -2544
rect 2490 -2556 2496 -2550
rect 2490 -2562 2496 -2556
rect 2490 -2568 2496 -2562
rect 2490 -2574 2496 -2568
rect 2490 -2580 2496 -2574
rect 2490 -2586 2496 -2580
rect 2490 -2592 2496 -2586
rect 2490 -2598 2496 -2592
rect 2490 -2604 2496 -2598
rect 2490 -2610 2496 -2604
rect 2490 -2616 2496 -2610
rect 2490 -2622 2496 -2616
rect 2490 -2628 2496 -2622
rect 2490 -2634 2496 -2628
rect 2490 -2640 2496 -2634
rect 2490 -2646 2496 -2640
rect 2490 -2652 2496 -2646
rect 2490 -2658 2496 -2652
rect 2490 -2664 2496 -2658
rect 2490 -2670 2496 -2664
rect 2490 -2676 2496 -2670
rect 2490 -2682 2496 -2676
rect 2490 -2688 2496 -2682
rect 2490 -2694 2496 -2688
rect 2490 -2700 2496 -2694
rect 2490 -2706 2496 -2700
rect 2490 -2712 2496 -2706
rect 2490 -2718 2496 -2712
rect 2490 -2724 2496 -2718
rect 2490 -2730 2496 -2724
rect 2490 -2736 2496 -2730
rect 2490 -2742 2496 -2736
rect 2490 -2748 2496 -2742
rect 2490 -2754 2496 -2748
rect 2490 -2760 2496 -2754
rect 2490 -2766 2496 -2760
rect 2490 -2772 2496 -2766
rect 2490 -2778 2496 -2772
rect 2490 -2784 2496 -2778
rect 2490 -2790 2496 -2784
rect 2490 -2796 2496 -2790
rect 2490 -2802 2496 -2796
rect 2490 -2808 2496 -2802
rect 2490 -2814 2496 -2808
rect 2490 -2820 2496 -2814
rect 2490 -2826 2496 -2820
rect 2490 -2832 2496 -2826
rect 2496 -1314 2502 -1308
rect 2496 -1320 2502 -1314
rect 2496 -1326 2502 -1320
rect 2496 -1332 2502 -1326
rect 2496 -1338 2502 -1332
rect 2496 -1344 2502 -1338
rect 2496 -1350 2502 -1344
rect 2496 -1356 2502 -1350
rect 2496 -1362 2502 -1356
rect 2496 -1368 2502 -1362
rect 2496 -1374 2502 -1368
rect 2496 -1380 2502 -1374
rect 2496 -1386 2502 -1380
rect 2496 -1392 2502 -1386
rect 2496 -1398 2502 -1392
rect 2496 -1404 2502 -1398
rect 2496 -1410 2502 -1404
rect 2496 -1416 2502 -1410
rect 2496 -1422 2502 -1416
rect 2496 -1428 2502 -1422
rect 2496 -1434 2502 -1428
rect 2496 -1440 2502 -1434
rect 2496 -1446 2502 -1440
rect 2496 -1452 2502 -1446
rect 2496 -1458 2502 -1452
rect 2496 -1464 2502 -1458
rect 2496 -1470 2502 -1464
rect 2496 -1476 2502 -1470
rect 2496 -1482 2502 -1476
rect 2496 -1488 2502 -1482
rect 2496 -1494 2502 -1488
rect 2496 -1500 2502 -1494
rect 2496 -1506 2502 -1500
rect 2496 -1512 2502 -1506
rect 2496 -1518 2502 -1512
rect 2496 -1524 2502 -1518
rect 2496 -1530 2502 -1524
rect 2496 -1536 2502 -1530
rect 2496 -1542 2502 -1536
rect 2496 -1548 2502 -1542
rect 2496 -1554 2502 -1548
rect 2496 -1560 2502 -1554
rect 2496 -1566 2502 -1560
rect 2496 -1572 2502 -1566
rect 2496 -1578 2502 -1572
rect 2496 -1584 2502 -1578
rect 2496 -1590 2502 -1584
rect 2496 -1596 2502 -1590
rect 2496 -1602 2502 -1596
rect 2496 -1608 2502 -1602
rect 2496 -1614 2502 -1608
rect 2496 -1620 2502 -1614
rect 2496 -1626 2502 -1620
rect 2496 -1632 2502 -1626
rect 2496 -1638 2502 -1632
rect 2496 -1644 2502 -1638
rect 2496 -1650 2502 -1644
rect 2496 -1656 2502 -1650
rect 2496 -1662 2502 -1656
rect 2496 -1668 2502 -1662
rect 2496 -1674 2502 -1668
rect 2496 -1680 2502 -1674
rect 2496 -1686 2502 -1680
rect 2496 -1692 2502 -1686
rect 2496 -1698 2502 -1692
rect 2496 -1704 2502 -1698
rect 2496 -1710 2502 -1704
rect 2496 -1716 2502 -1710
rect 2496 -1722 2502 -1716
rect 2496 -1728 2502 -1722
rect 2496 -1734 2502 -1728
rect 2496 -1740 2502 -1734
rect 2496 -1746 2502 -1740
rect 2496 -1752 2502 -1746
rect 2496 -1758 2502 -1752
rect 2496 -1764 2502 -1758
rect 2496 -1770 2502 -1764
rect 2496 -1776 2502 -1770
rect 2496 -1782 2502 -1776
rect 2496 -1788 2502 -1782
rect 2496 -1794 2502 -1788
rect 2496 -1800 2502 -1794
rect 2496 -1806 2502 -1800
rect 2496 -1812 2502 -1806
rect 2496 -1818 2502 -1812
rect 2496 -1824 2502 -1818
rect 2496 -1830 2502 -1824
rect 2496 -1836 2502 -1830
rect 2496 -1842 2502 -1836
rect 2496 -1848 2502 -1842
rect 2496 -1854 2502 -1848
rect 2496 -1860 2502 -1854
rect 2496 -1866 2502 -1860
rect 2496 -1872 2502 -1866
rect 2496 -1878 2502 -1872
rect 2496 -1884 2502 -1878
rect 2496 -1890 2502 -1884
rect 2496 -1896 2502 -1890
rect 2496 -1902 2502 -1896
rect 2496 -1908 2502 -1902
rect 2496 -1914 2502 -1908
rect 2496 -1920 2502 -1914
rect 2496 -1926 2502 -1920
rect 2496 -1932 2502 -1926
rect 2496 -1938 2502 -1932
rect 2496 -1944 2502 -1938
rect 2496 -1950 2502 -1944
rect 2496 -1956 2502 -1950
rect 2496 -1962 2502 -1956
rect 2496 -1968 2502 -1962
rect 2496 -1974 2502 -1968
rect 2496 -1980 2502 -1974
rect 2496 -2454 2502 -2448
rect 2496 -2460 2502 -2454
rect 2496 -2466 2502 -2460
rect 2496 -2472 2502 -2466
rect 2496 -2478 2502 -2472
rect 2496 -2484 2502 -2478
rect 2496 -2490 2502 -2484
rect 2496 -2496 2502 -2490
rect 2496 -2502 2502 -2496
rect 2496 -2508 2502 -2502
rect 2496 -2514 2502 -2508
rect 2496 -2520 2502 -2514
rect 2496 -2526 2502 -2520
rect 2496 -2532 2502 -2526
rect 2496 -2538 2502 -2532
rect 2496 -2544 2502 -2538
rect 2496 -2550 2502 -2544
rect 2496 -2556 2502 -2550
rect 2496 -2562 2502 -2556
rect 2496 -2568 2502 -2562
rect 2496 -2574 2502 -2568
rect 2496 -2580 2502 -2574
rect 2496 -2586 2502 -2580
rect 2496 -2592 2502 -2586
rect 2496 -2598 2502 -2592
rect 2496 -2604 2502 -2598
rect 2496 -2610 2502 -2604
rect 2496 -2616 2502 -2610
rect 2496 -2622 2502 -2616
rect 2496 -2628 2502 -2622
rect 2496 -2634 2502 -2628
rect 2496 -2640 2502 -2634
rect 2496 -2646 2502 -2640
rect 2496 -2652 2502 -2646
rect 2496 -2658 2502 -2652
rect 2496 -2664 2502 -2658
rect 2496 -2670 2502 -2664
rect 2496 -2676 2502 -2670
rect 2496 -2682 2502 -2676
rect 2496 -2688 2502 -2682
rect 2496 -2694 2502 -2688
rect 2496 -2700 2502 -2694
rect 2496 -2706 2502 -2700
rect 2496 -2712 2502 -2706
rect 2496 -2718 2502 -2712
rect 2496 -2724 2502 -2718
rect 2496 -2730 2502 -2724
rect 2496 -2736 2502 -2730
rect 2496 -2742 2502 -2736
rect 2496 -2748 2502 -2742
rect 2496 -2754 2502 -2748
rect 2496 -2760 2502 -2754
rect 2496 -2766 2502 -2760
rect 2496 -2772 2502 -2766
rect 2496 -2778 2502 -2772
rect 2496 -2784 2502 -2778
rect 2496 -2790 2502 -2784
rect 2496 -2796 2502 -2790
rect 2496 -2802 2502 -2796
rect 2496 -2808 2502 -2802
rect 2496 -2814 2502 -2808
rect 2496 -2820 2502 -2814
rect 2496 -2826 2502 -2820
rect 2502 -1308 2508 -1302
rect 2502 -1314 2508 -1308
rect 2502 -1320 2508 -1314
rect 2502 -1326 2508 -1320
rect 2502 -1332 2508 -1326
rect 2502 -1338 2508 -1332
rect 2502 -1344 2508 -1338
rect 2502 -1350 2508 -1344
rect 2502 -1356 2508 -1350
rect 2502 -1362 2508 -1356
rect 2502 -1368 2508 -1362
rect 2502 -1374 2508 -1368
rect 2502 -1380 2508 -1374
rect 2502 -1386 2508 -1380
rect 2502 -1392 2508 -1386
rect 2502 -1398 2508 -1392
rect 2502 -1404 2508 -1398
rect 2502 -1410 2508 -1404
rect 2502 -1416 2508 -1410
rect 2502 -1422 2508 -1416
rect 2502 -1428 2508 -1422
rect 2502 -1434 2508 -1428
rect 2502 -1440 2508 -1434
rect 2502 -1446 2508 -1440
rect 2502 -1452 2508 -1446
rect 2502 -1458 2508 -1452
rect 2502 -1464 2508 -1458
rect 2502 -1470 2508 -1464
rect 2502 -1476 2508 -1470
rect 2502 -1482 2508 -1476
rect 2502 -1488 2508 -1482
rect 2502 -1494 2508 -1488
rect 2502 -1500 2508 -1494
rect 2502 -1506 2508 -1500
rect 2502 -1512 2508 -1506
rect 2502 -1518 2508 -1512
rect 2502 -1524 2508 -1518
rect 2502 -1530 2508 -1524
rect 2502 -1536 2508 -1530
rect 2502 -1542 2508 -1536
rect 2502 -1548 2508 -1542
rect 2502 -1554 2508 -1548
rect 2502 -1560 2508 -1554
rect 2502 -1566 2508 -1560
rect 2502 -1572 2508 -1566
rect 2502 -1578 2508 -1572
rect 2502 -1584 2508 -1578
rect 2502 -1590 2508 -1584
rect 2502 -1596 2508 -1590
rect 2502 -1602 2508 -1596
rect 2502 -1608 2508 -1602
rect 2502 -1614 2508 -1608
rect 2502 -1620 2508 -1614
rect 2502 -1626 2508 -1620
rect 2502 -1632 2508 -1626
rect 2502 -1638 2508 -1632
rect 2502 -1644 2508 -1638
rect 2502 -1650 2508 -1644
rect 2502 -1656 2508 -1650
rect 2502 -1662 2508 -1656
rect 2502 -1668 2508 -1662
rect 2502 -1674 2508 -1668
rect 2502 -1680 2508 -1674
rect 2502 -1686 2508 -1680
rect 2502 -1692 2508 -1686
rect 2502 -1698 2508 -1692
rect 2502 -1704 2508 -1698
rect 2502 -1710 2508 -1704
rect 2502 -1716 2508 -1710
rect 2502 -1722 2508 -1716
rect 2502 -1728 2508 -1722
rect 2502 -1734 2508 -1728
rect 2502 -1740 2508 -1734
rect 2502 -1746 2508 -1740
rect 2502 -1752 2508 -1746
rect 2502 -1758 2508 -1752
rect 2502 -1764 2508 -1758
rect 2502 -1770 2508 -1764
rect 2502 -1776 2508 -1770
rect 2502 -1782 2508 -1776
rect 2502 -1788 2508 -1782
rect 2502 -1794 2508 -1788
rect 2502 -1800 2508 -1794
rect 2502 -1806 2508 -1800
rect 2502 -1812 2508 -1806
rect 2502 -1818 2508 -1812
rect 2502 -1824 2508 -1818
rect 2502 -1830 2508 -1824
rect 2502 -1836 2508 -1830
rect 2502 -1842 2508 -1836
rect 2502 -1848 2508 -1842
rect 2502 -1854 2508 -1848
rect 2502 -1860 2508 -1854
rect 2502 -1866 2508 -1860
rect 2502 -1872 2508 -1866
rect 2502 -1878 2508 -1872
rect 2502 -1884 2508 -1878
rect 2502 -1890 2508 -1884
rect 2502 -1896 2508 -1890
rect 2502 -1902 2508 -1896
rect 2502 -1908 2508 -1902
rect 2502 -1914 2508 -1908
rect 2502 -1920 2508 -1914
rect 2502 -1926 2508 -1920
rect 2502 -1932 2508 -1926
rect 2502 -1938 2508 -1932
rect 2502 -1944 2508 -1938
rect 2502 -1950 2508 -1944
rect 2502 -1956 2508 -1950
rect 2502 -1962 2508 -1956
rect 2502 -1968 2508 -1962
rect 2502 -1974 2508 -1968
rect 2502 -2448 2508 -2442
rect 2502 -2454 2508 -2448
rect 2502 -2460 2508 -2454
rect 2502 -2466 2508 -2460
rect 2502 -2472 2508 -2466
rect 2502 -2478 2508 -2472
rect 2502 -2484 2508 -2478
rect 2502 -2490 2508 -2484
rect 2502 -2496 2508 -2490
rect 2502 -2502 2508 -2496
rect 2502 -2508 2508 -2502
rect 2502 -2514 2508 -2508
rect 2502 -2520 2508 -2514
rect 2502 -2526 2508 -2520
rect 2502 -2532 2508 -2526
rect 2502 -2538 2508 -2532
rect 2502 -2544 2508 -2538
rect 2502 -2550 2508 -2544
rect 2502 -2556 2508 -2550
rect 2502 -2562 2508 -2556
rect 2502 -2568 2508 -2562
rect 2502 -2574 2508 -2568
rect 2502 -2580 2508 -2574
rect 2502 -2586 2508 -2580
rect 2502 -2592 2508 -2586
rect 2502 -2598 2508 -2592
rect 2502 -2604 2508 -2598
rect 2502 -2610 2508 -2604
rect 2502 -2616 2508 -2610
rect 2502 -2622 2508 -2616
rect 2502 -2628 2508 -2622
rect 2502 -2634 2508 -2628
rect 2502 -2640 2508 -2634
rect 2502 -2646 2508 -2640
rect 2502 -2652 2508 -2646
rect 2502 -2658 2508 -2652
rect 2502 -2664 2508 -2658
rect 2502 -2670 2508 -2664
rect 2502 -2676 2508 -2670
rect 2502 -2682 2508 -2676
rect 2502 -2688 2508 -2682
rect 2502 -2694 2508 -2688
rect 2502 -2700 2508 -2694
rect 2502 -2706 2508 -2700
rect 2502 -2712 2508 -2706
rect 2502 -2718 2508 -2712
rect 2502 -2724 2508 -2718
rect 2502 -2730 2508 -2724
rect 2502 -2736 2508 -2730
rect 2502 -2742 2508 -2736
rect 2502 -2748 2508 -2742
rect 2502 -2754 2508 -2748
rect 2502 -2760 2508 -2754
rect 2502 -2766 2508 -2760
rect 2502 -2772 2508 -2766
rect 2502 -2778 2508 -2772
rect 2502 -2784 2508 -2778
rect 2502 -2790 2508 -2784
rect 2502 -2796 2508 -2790
rect 2502 -2802 2508 -2796
rect 2502 -2808 2508 -2802
rect 2502 -2814 2508 -2808
rect 2502 -2820 2508 -2814
rect 2502 -2826 2508 -2820
rect 2508 -1302 2514 -1296
rect 2508 -1308 2514 -1302
rect 2508 -1314 2514 -1308
rect 2508 -1320 2514 -1314
rect 2508 -1326 2514 -1320
rect 2508 -1332 2514 -1326
rect 2508 -1338 2514 -1332
rect 2508 -1344 2514 -1338
rect 2508 -1350 2514 -1344
rect 2508 -1356 2514 -1350
rect 2508 -1362 2514 -1356
rect 2508 -1368 2514 -1362
rect 2508 -1374 2514 -1368
rect 2508 -1380 2514 -1374
rect 2508 -1386 2514 -1380
rect 2508 -1392 2514 -1386
rect 2508 -1398 2514 -1392
rect 2508 -1404 2514 -1398
rect 2508 -1410 2514 -1404
rect 2508 -1416 2514 -1410
rect 2508 -1422 2514 -1416
rect 2508 -1428 2514 -1422
rect 2508 -1434 2514 -1428
rect 2508 -1440 2514 -1434
rect 2508 -1446 2514 -1440
rect 2508 -1452 2514 -1446
rect 2508 -1458 2514 -1452
rect 2508 -1464 2514 -1458
rect 2508 -1470 2514 -1464
rect 2508 -1476 2514 -1470
rect 2508 -1482 2514 -1476
rect 2508 -1488 2514 -1482
rect 2508 -1494 2514 -1488
rect 2508 -1500 2514 -1494
rect 2508 -1506 2514 -1500
rect 2508 -1512 2514 -1506
rect 2508 -1518 2514 -1512
rect 2508 -1524 2514 -1518
rect 2508 -1530 2514 -1524
rect 2508 -1536 2514 -1530
rect 2508 -1542 2514 -1536
rect 2508 -1548 2514 -1542
rect 2508 -1554 2514 -1548
rect 2508 -1560 2514 -1554
rect 2508 -1566 2514 -1560
rect 2508 -1572 2514 -1566
rect 2508 -1578 2514 -1572
rect 2508 -1584 2514 -1578
rect 2508 -1590 2514 -1584
rect 2508 -1596 2514 -1590
rect 2508 -1602 2514 -1596
rect 2508 -1608 2514 -1602
rect 2508 -1614 2514 -1608
rect 2508 -1620 2514 -1614
rect 2508 -1626 2514 -1620
rect 2508 -1632 2514 -1626
rect 2508 -1638 2514 -1632
rect 2508 -1644 2514 -1638
rect 2508 -1650 2514 -1644
rect 2508 -1656 2514 -1650
rect 2508 -1662 2514 -1656
rect 2508 -1668 2514 -1662
rect 2508 -1674 2514 -1668
rect 2508 -1680 2514 -1674
rect 2508 -1686 2514 -1680
rect 2508 -1692 2514 -1686
rect 2508 -1698 2514 -1692
rect 2508 -1704 2514 -1698
rect 2508 -1710 2514 -1704
rect 2508 -1716 2514 -1710
rect 2508 -1722 2514 -1716
rect 2508 -1728 2514 -1722
rect 2508 -1734 2514 -1728
rect 2508 -1740 2514 -1734
rect 2508 -1746 2514 -1740
rect 2508 -1752 2514 -1746
rect 2508 -1758 2514 -1752
rect 2508 -1764 2514 -1758
rect 2508 -1770 2514 -1764
rect 2508 -1776 2514 -1770
rect 2508 -1782 2514 -1776
rect 2508 -1788 2514 -1782
rect 2508 -1794 2514 -1788
rect 2508 -1800 2514 -1794
rect 2508 -1806 2514 -1800
rect 2508 -1812 2514 -1806
rect 2508 -1818 2514 -1812
rect 2508 -1824 2514 -1818
rect 2508 -1830 2514 -1824
rect 2508 -1836 2514 -1830
rect 2508 -1842 2514 -1836
rect 2508 -1848 2514 -1842
rect 2508 -1854 2514 -1848
rect 2508 -1860 2514 -1854
rect 2508 -1866 2514 -1860
rect 2508 -1872 2514 -1866
rect 2508 -1878 2514 -1872
rect 2508 -1884 2514 -1878
rect 2508 -1890 2514 -1884
rect 2508 -1896 2514 -1890
rect 2508 -1902 2514 -1896
rect 2508 -1908 2514 -1902
rect 2508 -1914 2514 -1908
rect 2508 -1920 2514 -1914
rect 2508 -1926 2514 -1920
rect 2508 -1932 2514 -1926
rect 2508 -1938 2514 -1932
rect 2508 -1944 2514 -1938
rect 2508 -1950 2514 -1944
rect 2508 -1956 2514 -1950
rect 2508 -1962 2514 -1956
rect 2508 -2448 2514 -2442
rect 2508 -2454 2514 -2448
rect 2508 -2460 2514 -2454
rect 2508 -2466 2514 -2460
rect 2508 -2472 2514 -2466
rect 2508 -2478 2514 -2472
rect 2508 -2484 2514 -2478
rect 2508 -2490 2514 -2484
rect 2508 -2496 2514 -2490
rect 2508 -2502 2514 -2496
rect 2508 -2508 2514 -2502
rect 2508 -2514 2514 -2508
rect 2508 -2520 2514 -2514
rect 2508 -2526 2514 -2520
rect 2508 -2532 2514 -2526
rect 2508 -2538 2514 -2532
rect 2508 -2544 2514 -2538
rect 2508 -2550 2514 -2544
rect 2508 -2556 2514 -2550
rect 2508 -2562 2514 -2556
rect 2508 -2568 2514 -2562
rect 2508 -2574 2514 -2568
rect 2508 -2580 2514 -2574
rect 2508 -2586 2514 -2580
rect 2508 -2592 2514 -2586
rect 2508 -2598 2514 -2592
rect 2508 -2604 2514 -2598
rect 2508 -2610 2514 -2604
rect 2508 -2616 2514 -2610
rect 2508 -2622 2514 -2616
rect 2508 -2628 2514 -2622
rect 2508 -2634 2514 -2628
rect 2508 -2640 2514 -2634
rect 2508 -2646 2514 -2640
rect 2508 -2652 2514 -2646
rect 2508 -2658 2514 -2652
rect 2508 -2664 2514 -2658
rect 2508 -2670 2514 -2664
rect 2508 -2676 2514 -2670
rect 2508 -2682 2514 -2676
rect 2508 -2688 2514 -2682
rect 2508 -2694 2514 -2688
rect 2508 -2700 2514 -2694
rect 2508 -2706 2514 -2700
rect 2508 -2712 2514 -2706
rect 2508 -2718 2514 -2712
rect 2508 -2724 2514 -2718
rect 2508 -2730 2514 -2724
rect 2508 -2736 2514 -2730
rect 2508 -2742 2514 -2736
rect 2508 -2748 2514 -2742
rect 2508 -2754 2514 -2748
rect 2508 -2760 2514 -2754
rect 2508 -2766 2514 -2760
rect 2508 -2772 2514 -2766
rect 2508 -2778 2514 -2772
rect 2508 -2784 2514 -2778
rect 2508 -2790 2514 -2784
rect 2508 -2796 2514 -2790
rect 2508 -2802 2514 -2796
rect 2508 -2808 2514 -2802
rect 2508 -2814 2514 -2808
rect 2508 -2820 2514 -2814
rect 2514 -1296 2520 -1290
rect 2514 -1302 2520 -1296
rect 2514 -1308 2520 -1302
rect 2514 -1314 2520 -1308
rect 2514 -1320 2520 -1314
rect 2514 -1326 2520 -1320
rect 2514 -1332 2520 -1326
rect 2514 -1338 2520 -1332
rect 2514 -1344 2520 -1338
rect 2514 -1350 2520 -1344
rect 2514 -1356 2520 -1350
rect 2514 -1362 2520 -1356
rect 2514 -1368 2520 -1362
rect 2514 -1374 2520 -1368
rect 2514 -1380 2520 -1374
rect 2514 -1386 2520 -1380
rect 2514 -1392 2520 -1386
rect 2514 -1398 2520 -1392
rect 2514 -1404 2520 -1398
rect 2514 -1410 2520 -1404
rect 2514 -1416 2520 -1410
rect 2514 -1422 2520 -1416
rect 2514 -1428 2520 -1422
rect 2514 -1434 2520 -1428
rect 2514 -1440 2520 -1434
rect 2514 -1446 2520 -1440
rect 2514 -1452 2520 -1446
rect 2514 -1458 2520 -1452
rect 2514 -1464 2520 -1458
rect 2514 -1470 2520 -1464
rect 2514 -1476 2520 -1470
rect 2514 -1482 2520 -1476
rect 2514 -1488 2520 -1482
rect 2514 -1494 2520 -1488
rect 2514 -1500 2520 -1494
rect 2514 -1506 2520 -1500
rect 2514 -1512 2520 -1506
rect 2514 -1518 2520 -1512
rect 2514 -1524 2520 -1518
rect 2514 -1530 2520 -1524
rect 2514 -1536 2520 -1530
rect 2514 -1542 2520 -1536
rect 2514 -1548 2520 -1542
rect 2514 -1554 2520 -1548
rect 2514 -1560 2520 -1554
rect 2514 -1566 2520 -1560
rect 2514 -1572 2520 -1566
rect 2514 -1578 2520 -1572
rect 2514 -1584 2520 -1578
rect 2514 -1590 2520 -1584
rect 2514 -1596 2520 -1590
rect 2514 -1602 2520 -1596
rect 2514 -1608 2520 -1602
rect 2514 -1614 2520 -1608
rect 2514 -1620 2520 -1614
rect 2514 -1626 2520 -1620
rect 2514 -1632 2520 -1626
rect 2514 -1638 2520 -1632
rect 2514 -1644 2520 -1638
rect 2514 -1650 2520 -1644
rect 2514 -1656 2520 -1650
rect 2514 -1662 2520 -1656
rect 2514 -1668 2520 -1662
rect 2514 -1674 2520 -1668
rect 2514 -1680 2520 -1674
rect 2514 -1686 2520 -1680
rect 2514 -1692 2520 -1686
rect 2514 -1698 2520 -1692
rect 2514 -1704 2520 -1698
rect 2514 -1710 2520 -1704
rect 2514 -1716 2520 -1710
rect 2514 -1722 2520 -1716
rect 2514 -1728 2520 -1722
rect 2514 -1734 2520 -1728
rect 2514 -1740 2520 -1734
rect 2514 -1746 2520 -1740
rect 2514 -1752 2520 -1746
rect 2514 -1758 2520 -1752
rect 2514 -1764 2520 -1758
rect 2514 -1770 2520 -1764
rect 2514 -1776 2520 -1770
rect 2514 -1782 2520 -1776
rect 2514 -1788 2520 -1782
rect 2514 -1794 2520 -1788
rect 2514 -1800 2520 -1794
rect 2514 -1806 2520 -1800
rect 2514 -1812 2520 -1806
rect 2514 -1818 2520 -1812
rect 2514 -1824 2520 -1818
rect 2514 -1830 2520 -1824
rect 2514 -1836 2520 -1830
rect 2514 -1842 2520 -1836
rect 2514 -1848 2520 -1842
rect 2514 -1854 2520 -1848
rect 2514 -1860 2520 -1854
rect 2514 -1866 2520 -1860
rect 2514 -1872 2520 -1866
rect 2514 -1878 2520 -1872
rect 2514 -1884 2520 -1878
rect 2514 -1890 2520 -1884
rect 2514 -1896 2520 -1890
rect 2514 -1902 2520 -1896
rect 2514 -1908 2520 -1902
rect 2514 -1914 2520 -1908
rect 2514 -1920 2520 -1914
rect 2514 -1926 2520 -1920
rect 2514 -1932 2520 -1926
rect 2514 -1938 2520 -1932
rect 2514 -1944 2520 -1938
rect 2514 -1950 2520 -1944
rect 2514 -1956 2520 -1950
rect 2514 -2448 2520 -2442
rect 2514 -2454 2520 -2448
rect 2514 -2460 2520 -2454
rect 2514 -2466 2520 -2460
rect 2514 -2472 2520 -2466
rect 2514 -2478 2520 -2472
rect 2514 -2484 2520 -2478
rect 2514 -2490 2520 -2484
rect 2514 -2496 2520 -2490
rect 2514 -2502 2520 -2496
rect 2514 -2508 2520 -2502
rect 2514 -2514 2520 -2508
rect 2514 -2520 2520 -2514
rect 2514 -2526 2520 -2520
rect 2514 -2532 2520 -2526
rect 2514 -2538 2520 -2532
rect 2514 -2544 2520 -2538
rect 2514 -2550 2520 -2544
rect 2514 -2556 2520 -2550
rect 2514 -2562 2520 -2556
rect 2514 -2568 2520 -2562
rect 2514 -2574 2520 -2568
rect 2514 -2580 2520 -2574
rect 2514 -2586 2520 -2580
rect 2514 -2592 2520 -2586
rect 2514 -2598 2520 -2592
rect 2514 -2604 2520 -2598
rect 2514 -2610 2520 -2604
rect 2514 -2616 2520 -2610
rect 2514 -2622 2520 -2616
rect 2514 -2628 2520 -2622
rect 2514 -2634 2520 -2628
rect 2514 -2640 2520 -2634
rect 2514 -2646 2520 -2640
rect 2514 -2652 2520 -2646
rect 2514 -2658 2520 -2652
rect 2514 -2664 2520 -2658
rect 2514 -2670 2520 -2664
rect 2514 -2676 2520 -2670
rect 2514 -2682 2520 -2676
rect 2514 -2688 2520 -2682
rect 2514 -2694 2520 -2688
rect 2514 -2700 2520 -2694
rect 2514 -2706 2520 -2700
rect 2514 -2712 2520 -2706
rect 2514 -2718 2520 -2712
rect 2514 -2724 2520 -2718
rect 2514 -2730 2520 -2724
rect 2514 -2736 2520 -2730
rect 2514 -2742 2520 -2736
rect 2514 -2748 2520 -2742
rect 2514 -2754 2520 -2748
rect 2514 -2760 2520 -2754
rect 2514 -2766 2520 -2760
rect 2514 -2772 2520 -2766
rect 2514 -2778 2520 -2772
rect 2514 -2784 2520 -2778
rect 2514 -2790 2520 -2784
rect 2514 -2796 2520 -2790
rect 2514 -2802 2520 -2796
rect 2514 -2808 2520 -2802
rect 2514 -2814 2520 -2808
rect 2514 -2820 2520 -2814
rect 2520 -1296 2526 -1290
rect 2520 -1302 2526 -1296
rect 2520 -1308 2526 -1302
rect 2520 -1314 2526 -1308
rect 2520 -1320 2526 -1314
rect 2520 -1326 2526 -1320
rect 2520 -1332 2526 -1326
rect 2520 -1338 2526 -1332
rect 2520 -1344 2526 -1338
rect 2520 -1350 2526 -1344
rect 2520 -1356 2526 -1350
rect 2520 -1362 2526 -1356
rect 2520 -1368 2526 -1362
rect 2520 -1374 2526 -1368
rect 2520 -1380 2526 -1374
rect 2520 -1386 2526 -1380
rect 2520 -1392 2526 -1386
rect 2520 -1398 2526 -1392
rect 2520 -1404 2526 -1398
rect 2520 -1410 2526 -1404
rect 2520 -1416 2526 -1410
rect 2520 -1422 2526 -1416
rect 2520 -1428 2526 -1422
rect 2520 -1434 2526 -1428
rect 2520 -1440 2526 -1434
rect 2520 -1446 2526 -1440
rect 2520 -1452 2526 -1446
rect 2520 -1458 2526 -1452
rect 2520 -1464 2526 -1458
rect 2520 -1470 2526 -1464
rect 2520 -1476 2526 -1470
rect 2520 -1482 2526 -1476
rect 2520 -1488 2526 -1482
rect 2520 -1494 2526 -1488
rect 2520 -1500 2526 -1494
rect 2520 -1506 2526 -1500
rect 2520 -1512 2526 -1506
rect 2520 -1518 2526 -1512
rect 2520 -1524 2526 -1518
rect 2520 -1530 2526 -1524
rect 2520 -1536 2526 -1530
rect 2520 -1542 2526 -1536
rect 2520 -1548 2526 -1542
rect 2520 -1554 2526 -1548
rect 2520 -1560 2526 -1554
rect 2520 -1566 2526 -1560
rect 2520 -1572 2526 -1566
rect 2520 -1578 2526 -1572
rect 2520 -1584 2526 -1578
rect 2520 -1590 2526 -1584
rect 2520 -1596 2526 -1590
rect 2520 -1602 2526 -1596
rect 2520 -1608 2526 -1602
rect 2520 -1614 2526 -1608
rect 2520 -1620 2526 -1614
rect 2520 -1626 2526 -1620
rect 2520 -1632 2526 -1626
rect 2520 -1638 2526 -1632
rect 2520 -1644 2526 -1638
rect 2520 -1650 2526 -1644
rect 2520 -1656 2526 -1650
rect 2520 -1662 2526 -1656
rect 2520 -1668 2526 -1662
rect 2520 -1674 2526 -1668
rect 2520 -1680 2526 -1674
rect 2520 -1686 2526 -1680
rect 2520 -1692 2526 -1686
rect 2520 -1698 2526 -1692
rect 2520 -1704 2526 -1698
rect 2520 -1710 2526 -1704
rect 2520 -1716 2526 -1710
rect 2520 -1722 2526 -1716
rect 2520 -1728 2526 -1722
rect 2520 -1734 2526 -1728
rect 2520 -1740 2526 -1734
rect 2520 -1746 2526 -1740
rect 2520 -1752 2526 -1746
rect 2520 -1758 2526 -1752
rect 2520 -1764 2526 -1758
rect 2520 -1770 2526 -1764
rect 2520 -1776 2526 -1770
rect 2520 -1782 2526 -1776
rect 2520 -1788 2526 -1782
rect 2520 -1794 2526 -1788
rect 2520 -1800 2526 -1794
rect 2520 -1806 2526 -1800
rect 2520 -1812 2526 -1806
rect 2520 -1818 2526 -1812
rect 2520 -1824 2526 -1818
rect 2520 -1830 2526 -1824
rect 2520 -1836 2526 -1830
rect 2520 -1842 2526 -1836
rect 2520 -1848 2526 -1842
rect 2520 -1854 2526 -1848
rect 2520 -1860 2526 -1854
rect 2520 -1866 2526 -1860
rect 2520 -1872 2526 -1866
rect 2520 -1878 2526 -1872
rect 2520 -1884 2526 -1878
rect 2520 -1890 2526 -1884
rect 2520 -1896 2526 -1890
rect 2520 -1902 2526 -1896
rect 2520 -1908 2526 -1902
rect 2520 -1914 2526 -1908
rect 2520 -1920 2526 -1914
rect 2520 -1926 2526 -1920
rect 2520 -1932 2526 -1926
rect 2520 -1938 2526 -1932
rect 2520 -1944 2526 -1938
rect 2520 -1950 2526 -1944
rect 2520 -2442 2526 -2436
rect 2520 -2448 2526 -2442
rect 2520 -2454 2526 -2448
rect 2520 -2460 2526 -2454
rect 2520 -2466 2526 -2460
rect 2520 -2472 2526 -2466
rect 2520 -2478 2526 -2472
rect 2520 -2484 2526 -2478
rect 2520 -2490 2526 -2484
rect 2520 -2496 2526 -2490
rect 2520 -2502 2526 -2496
rect 2520 -2508 2526 -2502
rect 2520 -2514 2526 -2508
rect 2520 -2520 2526 -2514
rect 2520 -2526 2526 -2520
rect 2520 -2532 2526 -2526
rect 2520 -2538 2526 -2532
rect 2520 -2544 2526 -2538
rect 2520 -2550 2526 -2544
rect 2520 -2556 2526 -2550
rect 2520 -2562 2526 -2556
rect 2520 -2568 2526 -2562
rect 2520 -2574 2526 -2568
rect 2520 -2580 2526 -2574
rect 2520 -2586 2526 -2580
rect 2520 -2592 2526 -2586
rect 2520 -2598 2526 -2592
rect 2520 -2604 2526 -2598
rect 2520 -2610 2526 -2604
rect 2520 -2616 2526 -2610
rect 2520 -2622 2526 -2616
rect 2520 -2628 2526 -2622
rect 2520 -2634 2526 -2628
rect 2520 -2640 2526 -2634
rect 2520 -2646 2526 -2640
rect 2520 -2652 2526 -2646
rect 2520 -2658 2526 -2652
rect 2520 -2664 2526 -2658
rect 2520 -2670 2526 -2664
rect 2520 -2676 2526 -2670
rect 2520 -2682 2526 -2676
rect 2520 -2688 2526 -2682
rect 2520 -2694 2526 -2688
rect 2520 -2700 2526 -2694
rect 2520 -2706 2526 -2700
rect 2520 -2712 2526 -2706
rect 2520 -2718 2526 -2712
rect 2520 -2724 2526 -2718
rect 2520 -2730 2526 -2724
rect 2520 -2736 2526 -2730
rect 2520 -2742 2526 -2736
rect 2520 -2748 2526 -2742
rect 2520 -2754 2526 -2748
rect 2520 -2760 2526 -2754
rect 2520 -2766 2526 -2760
rect 2520 -2772 2526 -2766
rect 2520 -2778 2526 -2772
rect 2520 -2784 2526 -2778
rect 2520 -2790 2526 -2784
rect 2520 -2796 2526 -2790
rect 2520 -2802 2526 -2796
rect 2520 -2808 2526 -2802
rect 2520 -2814 2526 -2808
rect 2526 -1290 2532 -1284
rect 2526 -1296 2532 -1290
rect 2526 -1302 2532 -1296
rect 2526 -1308 2532 -1302
rect 2526 -1314 2532 -1308
rect 2526 -1320 2532 -1314
rect 2526 -1326 2532 -1320
rect 2526 -1332 2532 -1326
rect 2526 -1338 2532 -1332
rect 2526 -1344 2532 -1338
rect 2526 -1350 2532 -1344
rect 2526 -1356 2532 -1350
rect 2526 -1362 2532 -1356
rect 2526 -1368 2532 -1362
rect 2526 -1374 2532 -1368
rect 2526 -1380 2532 -1374
rect 2526 -1386 2532 -1380
rect 2526 -1392 2532 -1386
rect 2526 -1398 2532 -1392
rect 2526 -1404 2532 -1398
rect 2526 -1410 2532 -1404
rect 2526 -1416 2532 -1410
rect 2526 -1422 2532 -1416
rect 2526 -1428 2532 -1422
rect 2526 -1434 2532 -1428
rect 2526 -1440 2532 -1434
rect 2526 -1446 2532 -1440
rect 2526 -1452 2532 -1446
rect 2526 -1458 2532 -1452
rect 2526 -1464 2532 -1458
rect 2526 -1470 2532 -1464
rect 2526 -1476 2532 -1470
rect 2526 -1482 2532 -1476
rect 2526 -1488 2532 -1482
rect 2526 -1494 2532 -1488
rect 2526 -1500 2532 -1494
rect 2526 -1506 2532 -1500
rect 2526 -1512 2532 -1506
rect 2526 -1518 2532 -1512
rect 2526 -1524 2532 -1518
rect 2526 -1530 2532 -1524
rect 2526 -1536 2532 -1530
rect 2526 -1542 2532 -1536
rect 2526 -1548 2532 -1542
rect 2526 -1554 2532 -1548
rect 2526 -1560 2532 -1554
rect 2526 -1566 2532 -1560
rect 2526 -1572 2532 -1566
rect 2526 -1578 2532 -1572
rect 2526 -1584 2532 -1578
rect 2526 -1590 2532 -1584
rect 2526 -1596 2532 -1590
rect 2526 -1602 2532 -1596
rect 2526 -1608 2532 -1602
rect 2526 -1614 2532 -1608
rect 2526 -1620 2532 -1614
rect 2526 -1626 2532 -1620
rect 2526 -1632 2532 -1626
rect 2526 -1638 2532 -1632
rect 2526 -1644 2532 -1638
rect 2526 -1650 2532 -1644
rect 2526 -1656 2532 -1650
rect 2526 -1662 2532 -1656
rect 2526 -1668 2532 -1662
rect 2526 -1674 2532 -1668
rect 2526 -1680 2532 -1674
rect 2526 -1686 2532 -1680
rect 2526 -1692 2532 -1686
rect 2526 -1698 2532 -1692
rect 2526 -1704 2532 -1698
rect 2526 -1710 2532 -1704
rect 2526 -1716 2532 -1710
rect 2526 -1722 2532 -1716
rect 2526 -1728 2532 -1722
rect 2526 -1734 2532 -1728
rect 2526 -1740 2532 -1734
rect 2526 -1746 2532 -1740
rect 2526 -1752 2532 -1746
rect 2526 -1758 2532 -1752
rect 2526 -1764 2532 -1758
rect 2526 -1770 2532 -1764
rect 2526 -1776 2532 -1770
rect 2526 -1782 2532 -1776
rect 2526 -1788 2532 -1782
rect 2526 -1794 2532 -1788
rect 2526 -1800 2532 -1794
rect 2526 -1806 2532 -1800
rect 2526 -1812 2532 -1806
rect 2526 -1818 2532 -1812
rect 2526 -1824 2532 -1818
rect 2526 -1830 2532 -1824
rect 2526 -1836 2532 -1830
rect 2526 -1842 2532 -1836
rect 2526 -1848 2532 -1842
rect 2526 -1854 2532 -1848
rect 2526 -1860 2532 -1854
rect 2526 -1866 2532 -1860
rect 2526 -1872 2532 -1866
rect 2526 -1878 2532 -1872
rect 2526 -1884 2532 -1878
rect 2526 -1890 2532 -1884
rect 2526 -1896 2532 -1890
rect 2526 -1902 2532 -1896
rect 2526 -1908 2532 -1902
rect 2526 -1914 2532 -1908
rect 2526 -1920 2532 -1914
rect 2526 -1926 2532 -1920
rect 2526 -1932 2532 -1926
rect 2526 -1938 2532 -1932
rect 2526 -1944 2532 -1938
rect 2526 -2442 2532 -2436
rect 2526 -2448 2532 -2442
rect 2526 -2454 2532 -2448
rect 2526 -2460 2532 -2454
rect 2526 -2466 2532 -2460
rect 2526 -2472 2532 -2466
rect 2526 -2478 2532 -2472
rect 2526 -2484 2532 -2478
rect 2526 -2490 2532 -2484
rect 2526 -2496 2532 -2490
rect 2526 -2502 2532 -2496
rect 2526 -2508 2532 -2502
rect 2526 -2514 2532 -2508
rect 2526 -2520 2532 -2514
rect 2526 -2526 2532 -2520
rect 2526 -2532 2532 -2526
rect 2526 -2538 2532 -2532
rect 2526 -2544 2532 -2538
rect 2526 -2550 2532 -2544
rect 2526 -2556 2532 -2550
rect 2526 -2562 2532 -2556
rect 2526 -2568 2532 -2562
rect 2526 -2574 2532 -2568
rect 2526 -2580 2532 -2574
rect 2526 -2586 2532 -2580
rect 2526 -2592 2532 -2586
rect 2526 -2598 2532 -2592
rect 2526 -2604 2532 -2598
rect 2526 -2610 2532 -2604
rect 2526 -2616 2532 -2610
rect 2526 -2622 2532 -2616
rect 2526 -2628 2532 -2622
rect 2526 -2634 2532 -2628
rect 2526 -2640 2532 -2634
rect 2526 -2646 2532 -2640
rect 2526 -2652 2532 -2646
rect 2526 -2658 2532 -2652
rect 2526 -2664 2532 -2658
rect 2526 -2670 2532 -2664
rect 2526 -2676 2532 -2670
rect 2526 -2682 2532 -2676
rect 2526 -2688 2532 -2682
rect 2526 -2694 2532 -2688
rect 2526 -2700 2532 -2694
rect 2526 -2706 2532 -2700
rect 2526 -2712 2532 -2706
rect 2526 -2718 2532 -2712
rect 2526 -2724 2532 -2718
rect 2526 -2730 2532 -2724
rect 2526 -2736 2532 -2730
rect 2526 -2742 2532 -2736
rect 2526 -2748 2532 -2742
rect 2526 -2754 2532 -2748
rect 2526 -2760 2532 -2754
rect 2526 -2766 2532 -2760
rect 2526 -2772 2532 -2766
rect 2526 -2778 2532 -2772
rect 2526 -2784 2532 -2778
rect 2526 -2790 2532 -2784
rect 2526 -2796 2532 -2790
rect 2526 -2802 2532 -2796
rect 2526 -2808 2532 -2802
rect 2532 -1284 2538 -1278
rect 2532 -1290 2538 -1284
rect 2532 -1296 2538 -1290
rect 2532 -1302 2538 -1296
rect 2532 -1308 2538 -1302
rect 2532 -1314 2538 -1308
rect 2532 -1320 2538 -1314
rect 2532 -1326 2538 -1320
rect 2532 -1332 2538 -1326
rect 2532 -1338 2538 -1332
rect 2532 -1344 2538 -1338
rect 2532 -1350 2538 -1344
rect 2532 -1356 2538 -1350
rect 2532 -1362 2538 -1356
rect 2532 -1368 2538 -1362
rect 2532 -1374 2538 -1368
rect 2532 -1380 2538 -1374
rect 2532 -1386 2538 -1380
rect 2532 -1392 2538 -1386
rect 2532 -1398 2538 -1392
rect 2532 -1404 2538 -1398
rect 2532 -1410 2538 -1404
rect 2532 -1416 2538 -1410
rect 2532 -1422 2538 -1416
rect 2532 -1428 2538 -1422
rect 2532 -1434 2538 -1428
rect 2532 -1440 2538 -1434
rect 2532 -1446 2538 -1440
rect 2532 -1452 2538 -1446
rect 2532 -1458 2538 -1452
rect 2532 -1464 2538 -1458
rect 2532 -1470 2538 -1464
rect 2532 -1476 2538 -1470
rect 2532 -1482 2538 -1476
rect 2532 -1488 2538 -1482
rect 2532 -1494 2538 -1488
rect 2532 -1500 2538 -1494
rect 2532 -1506 2538 -1500
rect 2532 -1512 2538 -1506
rect 2532 -1518 2538 -1512
rect 2532 -1524 2538 -1518
rect 2532 -1530 2538 -1524
rect 2532 -1536 2538 -1530
rect 2532 -1542 2538 -1536
rect 2532 -1548 2538 -1542
rect 2532 -1554 2538 -1548
rect 2532 -1560 2538 -1554
rect 2532 -1566 2538 -1560
rect 2532 -1572 2538 -1566
rect 2532 -1578 2538 -1572
rect 2532 -1584 2538 -1578
rect 2532 -1590 2538 -1584
rect 2532 -1596 2538 -1590
rect 2532 -1602 2538 -1596
rect 2532 -1608 2538 -1602
rect 2532 -1614 2538 -1608
rect 2532 -1620 2538 -1614
rect 2532 -1626 2538 -1620
rect 2532 -1632 2538 -1626
rect 2532 -1638 2538 -1632
rect 2532 -1644 2538 -1638
rect 2532 -1650 2538 -1644
rect 2532 -1656 2538 -1650
rect 2532 -1662 2538 -1656
rect 2532 -1668 2538 -1662
rect 2532 -1674 2538 -1668
rect 2532 -1680 2538 -1674
rect 2532 -1686 2538 -1680
rect 2532 -1692 2538 -1686
rect 2532 -1698 2538 -1692
rect 2532 -1704 2538 -1698
rect 2532 -1710 2538 -1704
rect 2532 -1716 2538 -1710
rect 2532 -1722 2538 -1716
rect 2532 -1728 2538 -1722
rect 2532 -1734 2538 -1728
rect 2532 -1740 2538 -1734
rect 2532 -1746 2538 -1740
rect 2532 -1752 2538 -1746
rect 2532 -1758 2538 -1752
rect 2532 -1764 2538 -1758
rect 2532 -1770 2538 -1764
rect 2532 -1776 2538 -1770
rect 2532 -1782 2538 -1776
rect 2532 -1788 2538 -1782
rect 2532 -1794 2538 -1788
rect 2532 -1800 2538 -1794
rect 2532 -1806 2538 -1800
rect 2532 -1812 2538 -1806
rect 2532 -1818 2538 -1812
rect 2532 -1824 2538 -1818
rect 2532 -1830 2538 -1824
rect 2532 -1836 2538 -1830
rect 2532 -1842 2538 -1836
rect 2532 -1848 2538 -1842
rect 2532 -1854 2538 -1848
rect 2532 -1860 2538 -1854
rect 2532 -1866 2538 -1860
rect 2532 -1872 2538 -1866
rect 2532 -1878 2538 -1872
rect 2532 -1884 2538 -1878
rect 2532 -1890 2538 -1884
rect 2532 -1896 2538 -1890
rect 2532 -1902 2538 -1896
rect 2532 -1908 2538 -1902
rect 2532 -1914 2538 -1908
rect 2532 -1920 2538 -1914
rect 2532 -1926 2538 -1920
rect 2532 -1932 2538 -1926
rect 2532 -2442 2538 -2436
rect 2532 -2448 2538 -2442
rect 2532 -2454 2538 -2448
rect 2532 -2460 2538 -2454
rect 2532 -2466 2538 -2460
rect 2532 -2472 2538 -2466
rect 2532 -2478 2538 -2472
rect 2532 -2484 2538 -2478
rect 2532 -2490 2538 -2484
rect 2532 -2496 2538 -2490
rect 2532 -2502 2538 -2496
rect 2532 -2508 2538 -2502
rect 2532 -2514 2538 -2508
rect 2532 -2520 2538 -2514
rect 2532 -2526 2538 -2520
rect 2532 -2532 2538 -2526
rect 2532 -2538 2538 -2532
rect 2532 -2544 2538 -2538
rect 2532 -2550 2538 -2544
rect 2532 -2556 2538 -2550
rect 2532 -2562 2538 -2556
rect 2532 -2568 2538 -2562
rect 2532 -2574 2538 -2568
rect 2532 -2580 2538 -2574
rect 2532 -2586 2538 -2580
rect 2532 -2592 2538 -2586
rect 2532 -2598 2538 -2592
rect 2532 -2604 2538 -2598
rect 2532 -2610 2538 -2604
rect 2532 -2616 2538 -2610
rect 2532 -2622 2538 -2616
rect 2532 -2628 2538 -2622
rect 2532 -2634 2538 -2628
rect 2532 -2640 2538 -2634
rect 2532 -2646 2538 -2640
rect 2532 -2652 2538 -2646
rect 2532 -2658 2538 -2652
rect 2532 -2664 2538 -2658
rect 2532 -2670 2538 -2664
rect 2532 -2676 2538 -2670
rect 2532 -2682 2538 -2676
rect 2532 -2688 2538 -2682
rect 2532 -2694 2538 -2688
rect 2532 -2700 2538 -2694
rect 2532 -2706 2538 -2700
rect 2532 -2712 2538 -2706
rect 2532 -2718 2538 -2712
rect 2532 -2724 2538 -2718
rect 2532 -2730 2538 -2724
rect 2532 -2736 2538 -2730
rect 2532 -2742 2538 -2736
rect 2532 -2748 2538 -2742
rect 2532 -2754 2538 -2748
rect 2532 -2760 2538 -2754
rect 2532 -2766 2538 -2760
rect 2532 -2772 2538 -2766
rect 2532 -2778 2538 -2772
rect 2532 -2784 2538 -2778
rect 2532 -2790 2538 -2784
rect 2532 -2796 2538 -2790
rect 2532 -2802 2538 -2796
rect 2532 -2808 2538 -2802
rect 2538 -1278 2544 -1272
rect 2538 -1284 2544 -1278
rect 2538 -1290 2544 -1284
rect 2538 -1296 2544 -1290
rect 2538 -1302 2544 -1296
rect 2538 -1308 2544 -1302
rect 2538 -1314 2544 -1308
rect 2538 -1320 2544 -1314
rect 2538 -1326 2544 -1320
rect 2538 -1332 2544 -1326
rect 2538 -1338 2544 -1332
rect 2538 -1344 2544 -1338
rect 2538 -1350 2544 -1344
rect 2538 -1356 2544 -1350
rect 2538 -1362 2544 -1356
rect 2538 -1368 2544 -1362
rect 2538 -1374 2544 -1368
rect 2538 -1380 2544 -1374
rect 2538 -1386 2544 -1380
rect 2538 -1392 2544 -1386
rect 2538 -1398 2544 -1392
rect 2538 -1404 2544 -1398
rect 2538 -1410 2544 -1404
rect 2538 -1416 2544 -1410
rect 2538 -1422 2544 -1416
rect 2538 -1428 2544 -1422
rect 2538 -1434 2544 -1428
rect 2538 -1440 2544 -1434
rect 2538 -1446 2544 -1440
rect 2538 -1452 2544 -1446
rect 2538 -1458 2544 -1452
rect 2538 -1464 2544 -1458
rect 2538 -1470 2544 -1464
rect 2538 -1476 2544 -1470
rect 2538 -1482 2544 -1476
rect 2538 -1488 2544 -1482
rect 2538 -1494 2544 -1488
rect 2538 -1500 2544 -1494
rect 2538 -1506 2544 -1500
rect 2538 -1512 2544 -1506
rect 2538 -1518 2544 -1512
rect 2538 -1524 2544 -1518
rect 2538 -1530 2544 -1524
rect 2538 -1536 2544 -1530
rect 2538 -1542 2544 -1536
rect 2538 -1548 2544 -1542
rect 2538 -1554 2544 -1548
rect 2538 -1560 2544 -1554
rect 2538 -1566 2544 -1560
rect 2538 -1572 2544 -1566
rect 2538 -1578 2544 -1572
rect 2538 -1584 2544 -1578
rect 2538 -1590 2544 -1584
rect 2538 -1596 2544 -1590
rect 2538 -1602 2544 -1596
rect 2538 -1608 2544 -1602
rect 2538 -1614 2544 -1608
rect 2538 -1620 2544 -1614
rect 2538 -1626 2544 -1620
rect 2538 -1632 2544 -1626
rect 2538 -1638 2544 -1632
rect 2538 -1644 2544 -1638
rect 2538 -1650 2544 -1644
rect 2538 -1656 2544 -1650
rect 2538 -1662 2544 -1656
rect 2538 -1668 2544 -1662
rect 2538 -1674 2544 -1668
rect 2538 -1680 2544 -1674
rect 2538 -1686 2544 -1680
rect 2538 -1692 2544 -1686
rect 2538 -1698 2544 -1692
rect 2538 -1704 2544 -1698
rect 2538 -1710 2544 -1704
rect 2538 -1716 2544 -1710
rect 2538 -1722 2544 -1716
rect 2538 -1728 2544 -1722
rect 2538 -1734 2544 -1728
rect 2538 -1740 2544 -1734
rect 2538 -1746 2544 -1740
rect 2538 -1752 2544 -1746
rect 2538 -1758 2544 -1752
rect 2538 -1764 2544 -1758
rect 2538 -1770 2544 -1764
rect 2538 -1776 2544 -1770
rect 2538 -1782 2544 -1776
rect 2538 -1788 2544 -1782
rect 2538 -1794 2544 -1788
rect 2538 -1800 2544 -1794
rect 2538 -1806 2544 -1800
rect 2538 -1812 2544 -1806
rect 2538 -1818 2544 -1812
rect 2538 -1824 2544 -1818
rect 2538 -1830 2544 -1824
rect 2538 -1836 2544 -1830
rect 2538 -1842 2544 -1836
rect 2538 -1848 2544 -1842
rect 2538 -1854 2544 -1848
rect 2538 -1860 2544 -1854
rect 2538 -1866 2544 -1860
rect 2538 -1872 2544 -1866
rect 2538 -1878 2544 -1872
rect 2538 -1884 2544 -1878
rect 2538 -1890 2544 -1884
rect 2538 -1896 2544 -1890
rect 2538 -1902 2544 -1896
rect 2538 -1908 2544 -1902
rect 2538 -1914 2544 -1908
rect 2538 -1920 2544 -1914
rect 2538 -1926 2544 -1920
rect 2538 -2442 2544 -2436
rect 2538 -2448 2544 -2442
rect 2538 -2454 2544 -2448
rect 2538 -2460 2544 -2454
rect 2538 -2466 2544 -2460
rect 2538 -2472 2544 -2466
rect 2538 -2478 2544 -2472
rect 2538 -2484 2544 -2478
rect 2538 -2490 2544 -2484
rect 2538 -2496 2544 -2490
rect 2538 -2502 2544 -2496
rect 2538 -2508 2544 -2502
rect 2538 -2514 2544 -2508
rect 2538 -2520 2544 -2514
rect 2538 -2526 2544 -2520
rect 2538 -2532 2544 -2526
rect 2538 -2538 2544 -2532
rect 2538 -2544 2544 -2538
rect 2538 -2550 2544 -2544
rect 2538 -2556 2544 -2550
rect 2538 -2562 2544 -2556
rect 2538 -2568 2544 -2562
rect 2538 -2574 2544 -2568
rect 2538 -2580 2544 -2574
rect 2538 -2586 2544 -2580
rect 2538 -2592 2544 -2586
rect 2538 -2598 2544 -2592
rect 2538 -2604 2544 -2598
rect 2538 -2610 2544 -2604
rect 2538 -2616 2544 -2610
rect 2538 -2622 2544 -2616
rect 2538 -2628 2544 -2622
rect 2538 -2634 2544 -2628
rect 2538 -2640 2544 -2634
rect 2538 -2646 2544 -2640
rect 2538 -2652 2544 -2646
rect 2538 -2658 2544 -2652
rect 2538 -2664 2544 -2658
rect 2538 -2670 2544 -2664
rect 2538 -2676 2544 -2670
rect 2538 -2682 2544 -2676
rect 2538 -2688 2544 -2682
rect 2538 -2694 2544 -2688
rect 2538 -2700 2544 -2694
rect 2538 -2706 2544 -2700
rect 2538 -2712 2544 -2706
rect 2538 -2718 2544 -2712
rect 2538 -2724 2544 -2718
rect 2538 -2730 2544 -2724
rect 2538 -2736 2544 -2730
rect 2538 -2742 2544 -2736
rect 2538 -2748 2544 -2742
rect 2538 -2754 2544 -2748
rect 2538 -2760 2544 -2754
rect 2538 -2766 2544 -2760
rect 2538 -2772 2544 -2766
rect 2538 -2778 2544 -2772
rect 2538 -2784 2544 -2778
rect 2538 -2790 2544 -2784
rect 2538 -2796 2544 -2790
rect 2538 -2802 2544 -2796
rect 2544 -1278 2550 -1272
rect 2544 -1284 2550 -1278
rect 2544 -1290 2550 -1284
rect 2544 -1296 2550 -1290
rect 2544 -1302 2550 -1296
rect 2544 -1308 2550 -1302
rect 2544 -1314 2550 -1308
rect 2544 -1320 2550 -1314
rect 2544 -1326 2550 -1320
rect 2544 -1332 2550 -1326
rect 2544 -1338 2550 -1332
rect 2544 -1344 2550 -1338
rect 2544 -1350 2550 -1344
rect 2544 -1356 2550 -1350
rect 2544 -1362 2550 -1356
rect 2544 -1368 2550 -1362
rect 2544 -1374 2550 -1368
rect 2544 -1380 2550 -1374
rect 2544 -1386 2550 -1380
rect 2544 -1392 2550 -1386
rect 2544 -1398 2550 -1392
rect 2544 -1404 2550 -1398
rect 2544 -1410 2550 -1404
rect 2544 -1416 2550 -1410
rect 2544 -1422 2550 -1416
rect 2544 -1428 2550 -1422
rect 2544 -1434 2550 -1428
rect 2544 -1440 2550 -1434
rect 2544 -1446 2550 -1440
rect 2544 -1452 2550 -1446
rect 2544 -1458 2550 -1452
rect 2544 -1464 2550 -1458
rect 2544 -1470 2550 -1464
rect 2544 -1476 2550 -1470
rect 2544 -1482 2550 -1476
rect 2544 -1488 2550 -1482
rect 2544 -1494 2550 -1488
rect 2544 -1500 2550 -1494
rect 2544 -1506 2550 -1500
rect 2544 -1512 2550 -1506
rect 2544 -1518 2550 -1512
rect 2544 -1524 2550 -1518
rect 2544 -1530 2550 -1524
rect 2544 -1536 2550 -1530
rect 2544 -1542 2550 -1536
rect 2544 -1548 2550 -1542
rect 2544 -1554 2550 -1548
rect 2544 -1560 2550 -1554
rect 2544 -1566 2550 -1560
rect 2544 -1572 2550 -1566
rect 2544 -1578 2550 -1572
rect 2544 -1584 2550 -1578
rect 2544 -1590 2550 -1584
rect 2544 -1596 2550 -1590
rect 2544 -1602 2550 -1596
rect 2544 -1608 2550 -1602
rect 2544 -1614 2550 -1608
rect 2544 -1620 2550 -1614
rect 2544 -1626 2550 -1620
rect 2544 -1632 2550 -1626
rect 2544 -1638 2550 -1632
rect 2544 -1644 2550 -1638
rect 2544 -1650 2550 -1644
rect 2544 -1656 2550 -1650
rect 2544 -1662 2550 -1656
rect 2544 -1668 2550 -1662
rect 2544 -1674 2550 -1668
rect 2544 -1680 2550 -1674
rect 2544 -1686 2550 -1680
rect 2544 -1692 2550 -1686
rect 2544 -1698 2550 -1692
rect 2544 -1704 2550 -1698
rect 2544 -1710 2550 -1704
rect 2544 -1716 2550 -1710
rect 2544 -1722 2550 -1716
rect 2544 -1728 2550 -1722
rect 2544 -1734 2550 -1728
rect 2544 -1740 2550 -1734
rect 2544 -1746 2550 -1740
rect 2544 -1752 2550 -1746
rect 2544 -1758 2550 -1752
rect 2544 -1764 2550 -1758
rect 2544 -1770 2550 -1764
rect 2544 -1776 2550 -1770
rect 2544 -1782 2550 -1776
rect 2544 -1788 2550 -1782
rect 2544 -1794 2550 -1788
rect 2544 -1800 2550 -1794
rect 2544 -1806 2550 -1800
rect 2544 -1812 2550 -1806
rect 2544 -1818 2550 -1812
rect 2544 -1824 2550 -1818
rect 2544 -1830 2550 -1824
rect 2544 -1836 2550 -1830
rect 2544 -1842 2550 -1836
rect 2544 -1848 2550 -1842
rect 2544 -1854 2550 -1848
rect 2544 -1860 2550 -1854
rect 2544 -1866 2550 -1860
rect 2544 -1872 2550 -1866
rect 2544 -1878 2550 -1872
rect 2544 -1884 2550 -1878
rect 2544 -1890 2550 -1884
rect 2544 -1896 2550 -1890
rect 2544 -1902 2550 -1896
rect 2544 -1908 2550 -1902
rect 2544 -1914 2550 -1908
rect 2544 -1920 2550 -1914
rect 2544 -2436 2550 -2430
rect 2544 -2442 2550 -2436
rect 2544 -2448 2550 -2442
rect 2544 -2454 2550 -2448
rect 2544 -2460 2550 -2454
rect 2544 -2466 2550 -2460
rect 2544 -2472 2550 -2466
rect 2544 -2478 2550 -2472
rect 2544 -2484 2550 -2478
rect 2544 -2490 2550 -2484
rect 2544 -2496 2550 -2490
rect 2544 -2502 2550 -2496
rect 2544 -2508 2550 -2502
rect 2544 -2514 2550 -2508
rect 2544 -2520 2550 -2514
rect 2544 -2526 2550 -2520
rect 2544 -2532 2550 -2526
rect 2544 -2538 2550 -2532
rect 2544 -2544 2550 -2538
rect 2544 -2550 2550 -2544
rect 2544 -2556 2550 -2550
rect 2544 -2562 2550 -2556
rect 2544 -2568 2550 -2562
rect 2544 -2574 2550 -2568
rect 2544 -2580 2550 -2574
rect 2544 -2586 2550 -2580
rect 2544 -2592 2550 -2586
rect 2544 -2598 2550 -2592
rect 2544 -2604 2550 -2598
rect 2544 -2610 2550 -2604
rect 2544 -2616 2550 -2610
rect 2544 -2622 2550 -2616
rect 2544 -2628 2550 -2622
rect 2544 -2634 2550 -2628
rect 2544 -2640 2550 -2634
rect 2544 -2646 2550 -2640
rect 2544 -2652 2550 -2646
rect 2544 -2658 2550 -2652
rect 2544 -2664 2550 -2658
rect 2544 -2670 2550 -2664
rect 2544 -2676 2550 -2670
rect 2544 -2682 2550 -2676
rect 2544 -2688 2550 -2682
rect 2544 -2694 2550 -2688
rect 2544 -2700 2550 -2694
rect 2544 -2706 2550 -2700
rect 2544 -2712 2550 -2706
rect 2544 -2718 2550 -2712
rect 2544 -2724 2550 -2718
rect 2544 -2730 2550 -2724
rect 2544 -2736 2550 -2730
rect 2544 -2742 2550 -2736
rect 2544 -2748 2550 -2742
rect 2544 -2754 2550 -2748
rect 2544 -2760 2550 -2754
rect 2544 -2766 2550 -2760
rect 2544 -2772 2550 -2766
rect 2544 -2778 2550 -2772
rect 2544 -2784 2550 -2778
rect 2544 -2790 2550 -2784
rect 2544 -2796 2550 -2790
rect 2544 -2802 2550 -2796
rect 2550 -1272 2556 -1266
rect 2550 -1278 2556 -1272
rect 2550 -1284 2556 -1278
rect 2550 -1290 2556 -1284
rect 2550 -1296 2556 -1290
rect 2550 -1302 2556 -1296
rect 2550 -1308 2556 -1302
rect 2550 -1314 2556 -1308
rect 2550 -1320 2556 -1314
rect 2550 -1326 2556 -1320
rect 2550 -1332 2556 -1326
rect 2550 -1338 2556 -1332
rect 2550 -1344 2556 -1338
rect 2550 -1350 2556 -1344
rect 2550 -1356 2556 -1350
rect 2550 -1362 2556 -1356
rect 2550 -1368 2556 -1362
rect 2550 -1374 2556 -1368
rect 2550 -1380 2556 -1374
rect 2550 -1386 2556 -1380
rect 2550 -1392 2556 -1386
rect 2550 -1398 2556 -1392
rect 2550 -1404 2556 -1398
rect 2550 -1410 2556 -1404
rect 2550 -1416 2556 -1410
rect 2550 -1422 2556 -1416
rect 2550 -1428 2556 -1422
rect 2550 -1434 2556 -1428
rect 2550 -1440 2556 -1434
rect 2550 -1446 2556 -1440
rect 2550 -1452 2556 -1446
rect 2550 -1458 2556 -1452
rect 2550 -1464 2556 -1458
rect 2550 -1470 2556 -1464
rect 2550 -1476 2556 -1470
rect 2550 -1482 2556 -1476
rect 2550 -1488 2556 -1482
rect 2550 -1494 2556 -1488
rect 2550 -1500 2556 -1494
rect 2550 -1506 2556 -1500
rect 2550 -1512 2556 -1506
rect 2550 -1518 2556 -1512
rect 2550 -1524 2556 -1518
rect 2550 -1530 2556 -1524
rect 2550 -1536 2556 -1530
rect 2550 -1542 2556 -1536
rect 2550 -1548 2556 -1542
rect 2550 -1554 2556 -1548
rect 2550 -1560 2556 -1554
rect 2550 -1566 2556 -1560
rect 2550 -1572 2556 -1566
rect 2550 -1578 2556 -1572
rect 2550 -1584 2556 -1578
rect 2550 -1590 2556 -1584
rect 2550 -1596 2556 -1590
rect 2550 -1602 2556 -1596
rect 2550 -1608 2556 -1602
rect 2550 -1614 2556 -1608
rect 2550 -1620 2556 -1614
rect 2550 -1626 2556 -1620
rect 2550 -1632 2556 -1626
rect 2550 -1638 2556 -1632
rect 2550 -1644 2556 -1638
rect 2550 -1650 2556 -1644
rect 2550 -1656 2556 -1650
rect 2550 -1662 2556 -1656
rect 2550 -1668 2556 -1662
rect 2550 -1674 2556 -1668
rect 2550 -1680 2556 -1674
rect 2550 -1686 2556 -1680
rect 2550 -1692 2556 -1686
rect 2550 -1698 2556 -1692
rect 2550 -1704 2556 -1698
rect 2550 -1710 2556 -1704
rect 2550 -1716 2556 -1710
rect 2550 -1722 2556 -1716
rect 2550 -1728 2556 -1722
rect 2550 -1734 2556 -1728
rect 2550 -1740 2556 -1734
rect 2550 -1746 2556 -1740
rect 2550 -1752 2556 -1746
rect 2550 -1758 2556 -1752
rect 2550 -1764 2556 -1758
rect 2550 -1770 2556 -1764
rect 2550 -1776 2556 -1770
rect 2550 -1782 2556 -1776
rect 2550 -1788 2556 -1782
rect 2550 -1794 2556 -1788
rect 2550 -1800 2556 -1794
rect 2550 -1806 2556 -1800
rect 2550 -1812 2556 -1806
rect 2550 -1818 2556 -1812
rect 2550 -1824 2556 -1818
rect 2550 -1830 2556 -1824
rect 2550 -1836 2556 -1830
rect 2550 -1842 2556 -1836
rect 2550 -1848 2556 -1842
rect 2550 -1854 2556 -1848
rect 2550 -1860 2556 -1854
rect 2550 -1866 2556 -1860
rect 2550 -1872 2556 -1866
rect 2550 -1878 2556 -1872
rect 2550 -1884 2556 -1878
rect 2550 -1890 2556 -1884
rect 2550 -1896 2556 -1890
rect 2550 -1902 2556 -1896
rect 2550 -1908 2556 -1902
rect 2550 -1914 2556 -1908
rect 2550 -2436 2556 -2430
rect 2550 -2442 2556 -2436
rect 2550 -2448 2556 -2442
rect 2550 -2454 2556 -2448
rect 2550 -2460 2556 -2454
rect 2550 -2466 2556 -2460
rect 2550 -2472 2556 -2466
rect 2550 -2478 2556 -2472
rect 2550 -2484 2556 -2478
rect 2550 -2490 2556 -2484
rect 2550 -2496 2556 -2490
rect 2550 -2502 2556 -2496
rect 2550 -2508 2556 -2502
rect 2550 -2514 2556 -2508
rect 2550 -2520 2556 -2514
rect 2550 -2526 2556 -2520
rect 2550 -2532 2556 -2526
rect 2550 -2538 2556 -2532
rect 2550 -2544 2556 -2538
rect 2550 -2550 2556 -2544
rect 2550 -2556 2556 -2550
rect 2550 -2562 2556 -2556
rect 2550 -2568 2556 -2562
rect 2550 -2574 2556 -2568
rect 2550 -2580 2556 -2574
rect 2550 -2586 2556 -2580
rect 2550 -2592 2556 -2586
rect 2550 -2598 2556 -2592
rect 2550 -2604 2556 -2598
rect 2550 -2610 2556 -2604
rect 2550 -2616 2556 -2610
rect 2550 -2622 2556 -2616
rect 2550 -2628 2556 -2622
rect 2550 -2634 2556 -2628
rect 2550 -2640 2556 -2634
rect 2550 -2646 2556 -2640
rect 2550 -2652 2556 -2646
rect 2550 -2658 2556 -2652
rect 2550 -2664 2556 -2658
rect 2550 -2670 2556 -2664
rect 2550 -2676 2556 -2670
rect 2550 -2682 2556 -2676
rect 2550 -2688 2556 -2682
rect 2550 -2694 2556 -2688
rect 2550 -2700 2556 -2694
rect 2550 -2706 2556 -2700
rect 2550 -2712 2556 -2706
rect 2550 -2718 2556 -2712
rect 2550 -2724 2556 -2718
rect 2550 -2730 2556 -2724
rect 2550 -2736 2556 -2730
rect 2550 -2742 2556 -2736
rect 2550 -2748 2556 -2742
rect 2550 -2754 2556 -2748
rect 2550 -2760 2556 -2754
rect 2550 -2766 2556 -2760
rect 2550 -2772 2556 -2766
rect 2550 -2778 2556 -2772
rect 2550 -2784 2556 -2778
rect 2550 -2790 2556 -2784
rect 2550 -2796 2556 -2790
rect 2556 -1266 2562 -1260
rect 2556 -1272 2562 -1266
rect 2556 -1278 2562 -1272
rect 2556 -1284 2562 -1278
rect 2556 -1290 2562 -1284
rect 2556 -1296 2562 -1290
rect 2556 -1302 2562 -1296
rect 2556 -1308 2562 -1302
rect 2556 -1314 2562 -1308
rect 2556 -1320 2562 -1314
rect 2556 -1326 2562 -1320
rect 2556 -1332 2562 -1326
rect 2556 -1338 2562 -1332
rect 2556 -1344 2562 -1338
rect 2556 -1350 2562 -1344
rect 2556 -1356 2562 -1350
rect 2556 -1362 2562 -1356
rect 2556 -1368 2562 -1362
rect 2556 -1374 2562 -1368
rect 2556 -1380 2562 -1374
rect 2556 -1386 2562 -1380
rect 2556 -1392 2562 -1386
rect 2556 -1398 2562 -1392
rect 2556 -1404 2562 -1398
rect 2556 -1410 2562 -1404
rect 2556 -1416 2562 -1410
rect 2556 -1422 2562 -1416
rect 2556 -1428 2562 -1422
rect 2556 -1434 2562 -1428
rect 2556 -1440 2562 -1434
rect 2556 -1446 2562 -1440
rect 2556 -1452 2562 -1446
rect 2556 -1458 2562 -1452
rect 2556 -1464 2562 -1458
rect 2556 -1470 2562 -1464
rect 2556 -1476 2562 -1470
rect 2556 -1482 2562 -1476
rect 2556 -1488 2562 -1482
rect 2556 -1494 2562 -1488
rect 2556 -1500 2562 -1494
rect 2556 -1506 2562 -1500
rect 2556 -1512 2562 -1506
rect 2556 -1518 2562 -1512
rect 2556 -1524 2562 -1518
rect 2556 -1530 2562 -1524
rect 2556 -1536 2562 -1530
rect 2556 -1542 2562 -1536
rect 2556 -1548 2562 -1542
rect 2556 -1554 2562 -1548
rect 2556 -1560 2562 -1554
rect 2556 -1566 2562 -1560
rect 2556 -1572 2562 -1566
rect 2556 -1578 2562 -1572
rect 2556 -1584 2562 -1578
rect 2556 -1590 2562 -1584
rect 2556 -1596 2562 -1590
rect 2556 -1602 2562 -1596
rect 2556 -1608 2562 -1602
rect 2556 -1614 2562 -1608
rect 2556 -1620 2562 -1614
rect 2556 -1626 2562 -1620
rect 2556 -1632 2562 -1626
rect 2556 -1638 2562 -1632
rect 2556 -1644 2562 -1638
rect 2556 -1650 2562 -1644
rect 2556 -1656 2562 -1650
rect 2556 -1662 2562 -1656
rect 2556 -1668 2562 -1662
rect 2556 -1674 2562 -1668
rect 2556 -1680 2562 -1674
rect 2556 -1686 2562 -1680
rect 2556 -1692 2562 -1686
rect 2556 -1698 2562 -1692
rect 2556 -1704 2562 -1698
rect 2556 -1710 2562 -1704
rect 2556 -1716 2562 -1710
rect 2556 -1722 2562 -1716
rect 2556 -1728 2562 -1722
rect 2556 -1734 2562 -1728
rect 2556 -1740 2562 -1734
rect 2556 -1746 2562 -1740
rect 2556 -1752 2562 -1746
rect 2556 -1758 2562 -1752
rect 2556 -1764 2562 -1758
rect 2556 -1770 2562 -1764
rect 2556 -1776 2562 -1770
rect 2556 -1782 2562 -1776
rect 2556 -1788 2562 -1782
rect 2556 -1794 2562 -1788
rect 2556 -1800 2562 -1794
rect 2556 -1806 2562 -1800
rect 2556 -1812 2562 -1806
rect 2556 -1818 2562 -1812
rect 2556 -1824 2562 -1818
rect 2556 -1830 2562 -1824
rect 2556 -1836 2562 -1830
rect 2556 -1842 2562 -1836
rect 2556 -1848 2562 -1842
rect 2556 -1854 2562 -1848
rect 2556 -1860 2562 -1854
rect 2556 -1866 2562 -1860
rect 2556 -1872 2562 -1866
rect 2556 -1878 2562 -1872
rect 2556 -1884 2562 -1878
rect 2556 -1890 2562 -1884
rect 2556 -1896 2562 -1890
rect 2556 -1902 2562 -1896
rect 2556 -1908 2562 -1902
rect 2556 -2436 2562 -2430
rect 2556 -2442 2562 -2436
rect 2556 -2448 2562 -2442
rect 2556 -2454 2562 -2448
rect 2556 -2460 2562 -2454
rect 2556 -2466 2562 -2460
rect 2556 -2472 2562 -2466
rect 2556 -2478 2562 -2472
rect 2556 -2484 2562 -2478
rect 2556 -2490 2562 -2484
rect 2556 -2496 2562 -2490
rect 2556 -2502 2562 -2496
rect 2556 -2508 2562 -2502
rect 2556 -2514 2562 -2508
rect 2556 -2520 2562 -2514
rect 2556 -2526 2562 -2520
rect 2556 -2532 2562 -2526
rect 2556 -2538 2562 -2532
rect 2556 -2544 2562 -2538
rect 2556 -2550 2562 -2544
rect 2556 -2556 2562 -2550
rect 2556 -2562 2562 -2556
rect 2556 -2568 2562 -2562
rect 2556 -2574 2562 -2568
rect 2556 -2580 2562 -2574
rect 2556 -2586 2562 -2580
rect 2556 -2592 2562 -2586
rect 2556 -2598 2562 -2592
rect 2556 -2604 2562 -2598
rect 2556 -2610 2562 -2604
rect 2556 -2616 2562 -2610
rect 2556 -2622 2562 -2616
rect 2556 -2628 2562 -2622
rect 2556 -2634 2562 -2628
rect 2556 -2640 2562 -2634
rect 2556 -2646 2562 -2640
rect 2556 -2652 2562 -2646
rect 2556 -2658 2562 -2652
rect 2556 -2664 2562 -2658
rect 2556 -2670 2562 -2664
rect 2556 -2676 2562 -2670
rect 2556 -2682 2562 -2676
rect 2556 -2688 2562 -2682
rect 2556 -2694 2562 -2688
rect 2556 -2700 2562 -2694
rect 2556 -2706 2562 -2700
rect 2556 -2712 2562 -2706
rect 2556 -2718 2562 -2712
rect 2556 -2724 2562 -2718
rect 2556 -2730 2562 -2724
rect 2556 -2736 2562 -2730
rect 2556 -2742 2562 -2736
rect 2556 -2748 2562 -2742
rect 2556 -2754 2562 -2748
rect 2556 -2760 2562 -2754
rect 2556 -2766 2562 -2760
rect 2556 -2772 2562 -2766
rect 2556 -2778 2562 -2772
rect 2556 -2784 2562 -2778
rect 2556 -2790 2562 -2784
rect 2562 -1260 2568 -1254
rect 2562 -1266 2568 -1260
rect 2562 -1272 2568 -1266
rect 2562 -1278 2568 -1272
rect 2562 -1284 2568 -1278
rect 2562 -1290 2568 -1284
rect 2562 -1296 2568 -1290
rect 2562 -1302 2568 -1296
rect 2562 -1308 2568 -1302
rect 2562 -1314 2568 -1308
rect 2562 -1320 2568 -1314
rect 2562 -1326 2568 -1320
rect 2562 -1332 2568 -1326
rect 2562 -1338 2568 -1332
rect 2562 -1344 2568 -1338
rect 2562 -1350 2568 -1344
rect 2562 -1356 2568 -1350
rect 2562 -1362 2568 -1356
rect 2562 -1368 2568 -1362
rect 2562 -1374 2568 -1368
rect 2562 -1380 2568 -1374
rect 2562 -1386 2568 -1380
rect 2562 -1392 2568 -1386
rect 2562 -1398 2568 -1392
rect 2562 -1404 2568 -1398
rect 2562 -1410 2568 -1404
rect 2562 -1416 2568 -1410
rect 2562 -1422 2568 -1416
rect 2562 -1428 2568 -1422
rect 2562 -1434 2568 -1428
rect 2562 -1440 2568 -1434
rect 2562 -1446 2568 -1440
rect 2562 -1452 2568 -1446
rect 2562 -1458 2568 -1452
rect 2562 -1464 2568 -1458
rect 2562 -1470 2568 -1464
rect 2562 -1476 2568 -1470
rect 2562 -1482 2568 -1476
rect 2562 -1488 2568 -1482
rect 2562 -1494 2568 -1488
rect 2562 -1500 2568 -1494
rect 2562 -1506 2568 -1500
rect 2562 -1512 2568 -1506
rect 2562 -1518 2568 -1512
rect 2562 -1524 2568 -1518
rect 2562 -1530 2568 -1524
rect 2562 -1536 2568 -1530
rect 2562 -1542 2568 -1536
rect 2562 -1548 2568 -1542
rect 2562 -1554 2568 -1548
rect 2562 -1560 2568 -1554
rect 2562 -1566 2568 -1560
rect 2562 -1572 2568 -1566
rect 2562 -1578 2568 -1572
rect 2562 -1584 2568 -1578
rect 2562 -1590 2568 -1584
rect 2562 -1596 2568 -1590
rect 2562 -1602 2568 -1596
rect 2562 -1608 2568 -1602
rect 2562 -1614 2568 -1608
rect 2562 -1620 2568 -1614
rect 2562 -1626 2568 -1620
rect 2562 -1632 2568 -1626
rect 2562 -1638 2568 -1632
rect 2562 -1644 2568 -1638
rect 2562 -1650 2568 -1644
rect 2562 -1656 2568 -1650
rect 2562 -1662 2568 -1656
rect 2562 -1668 2568 -1662
rect 2562 -1674 2568 -1668
rect 2562 -1680 2568 -1674
rect 2562 -1686 2568 -1680
rect 2562 -1692 2568 -1686
rect 2562 -1698 2568 -1692
rect 2562 -1704 2568 -1698
rect 2562 -1710 2568 -1704
rect 2562 -1716 2568 -1710
rect 2562 -1722 2568 -1716
rect 2562 -1728 2568 -1722
rect 2562 -1734 2568 -1728
rect 2562 -1740 2568 -1734
rect 2562 -1746 2568 -1740
rect 2562 -1752 2568 -1746
rect 2562 -1758 2568 -1752
rect 2562 -1764 2568 -1758
rect 2562 -1770 2568 -1764
rect 2562 -1776 2568 -1770
rect 2562 -1782 2568 -1776
rect 2562 -1788 2568 -1782
rect 2562 -1794 2568 -1788
rect 2562 -1800 2568 -1794
rect 2562 -1806 2568 -1800
rect 2562 -1812 2568 -1806
rect 2562 -1818 2568 -1812
rect 2562 -1824 2568 -1818
rect 2562 -1830 2568 -1824
rect 2562 -1836 2568 -1830
rect 2562 -1842 2568 -1836
rect 2562 -1848 2568 -1842
rect 2562 -1854 2568 -1848
rect 2562 -1860 2568 -1854
rect 2562 -1866 2568 -1860
rect 2562 -1872 2568 -1866
rect 2562 -1878 2568 -1872
rect 2562 -1884 2568 -1878
rect 2562 -1890 2568 -1884
rect 2562 -1896 2568 -1890
rect 2562 -2436 2568 -2430
rect 2562 -2442 2568 -2436
rect 2562 -2448 2568 -2442
rect 2562 -2454 2568 -2448
rect 2562 -2460 2568 -2454
rect 2562 -2466 2568 -2460
rect 2562 -2472 2568 -2466
rect 2562 -2478 2568 -2472
rect 2562 -2484 2568 -2478
rect 2562 -2490 2568 -2484
rect 2562 -2496 2568 -2490
rect 2562 -2502 2568 -2496
rect 2562 -2508 2568 -2502
rect 2562 -2514 2568 -2508
rect 2562 -2520 2568 -2514
rect 2562 -2526 2568 -2520
rect 2562 -2532 2568 -2526
rect 2562 -2538 2568 -2532
rect 2562 -2544 2568 -2538
rect 2562 -2550 2568 -2544
rect 2562 -2556 2568 -2550
rect 2562 -2562 2568 -2556
rect 2562 -2568 2568 -2562
rect 2562 -2574 2568 -2568
rect 2562 -2580 2568 -2574
rect 2562 -2586 2568 -2580
rect 2562 -2592 2568 -2586
rect 2562 -2598 2568 -2592
rect 2562 -2604 2568 -2598
rect 2562 -2610 2568 -2604
rect 2562 -2616 2568 -2610
rect 2562 -2622 2568 -2616
rect 2562 -2628 2568 -2622
rect 2562 -2634 2568 -2628
rect 2562 -2640 2568 -2634
rect 2562 -2646 2568 -2640
rect 2562 -2652 2568 -2646
rect 2562 -2658 2568 -2652
rect 2562 -2664 2568 -2658
rect 2562 -2670 2568 -2664
rect 2562 -2676 2568 -2670
rect 2562 -2682 2568 -2676
rect 2562 -2688 2568 -2682
rect 2562 -2694 2568 -2688
rect 2562 -2700 2568 -2694
rect 2562 -2706 2568 -2700
rect 2562 -2712 2568 -2706
rect 2562 -2718 2568 -2712
rect 2562 -2724 2568 -2718
rect 2562 -2730 2568 -2724
rect 2562 -2736 2568 -2730
rect 2562 -2742 2568 -2736
rect 2562 -2748 2568 -2742
rect 2562 -2754 2568 -2748
rect 2562 -2760 2568 -2754
rect 2562 -2766 2568 -2760
rect 2562 -2772 2568 -2766
rect 2562 -2778 2568 -2772
rect 2562 -2784 2568 -2778
rect 2562 -2790 2568 -2784
rect 2568 -1260 2574 -1254
rect 2568 -1266 2574 -1260
rect 2568 -1272 2574 -1266
rect 2568 -1278 2574 -1272
rect 2568 -1284 2574 -1278
rect 2568 -1290 2574 -1284
rect 2568 -1296 2574 -1290
rect 2568 -1302 2574 -1296
rect 2568 -1308 2574 -1302
rect 2568 -1314 2574 -1308
rect 2568 -1320 2574 -1314
rect 2568 -1326 2574 -1320
rect 2568 -1332 2574 -1326
rect 2568 -1338 2574 -1332
rect 2568 -1344 2574 -1338
rect 2568 -1350 2574 -1344
rect 2568 -1356 2574 -1350
rect 2568 -1362 2574 -1356
rect 2568 -1368 2574 -1362
rect 2568 -1374 2574 -1368
rect 2568 -1380 2574 -1374
rect 2568 -1386 2574 -1380
rect 2568 -1392 2574 -1386
rect 2568 -1398 2574 -1392
rect 2568 -1404 2574 -1398
rect 2568 -1410 2574 -1404
rect 2568 -1416 2574 -1410
rect 2568 -1422 2574 -1416
rect 2568 -1428 2574 -1422
rect 2568 -1434 2574 -1428
rect 2568 -1440 2574 -1434
rect 2568 -1446 2574 -1440
rect 2568 -1452 2574 -1446
rect 2568 -1458 2574 -1452
rect 2568 -1464 2574 -1458
rect 2568 -1470 2574 -1464
rect 2568 -1476 2574 -1470
rect 2568 -1482 2574 -1476
rect 2568 -1488 2574 -1482
rect 2568 -1494 2574 -1488
rect 2568 -1500 2574 -1494
rect 2568 -1506 2574 -1500
rect 2568 -1512 2574 -1506
rect 2568 -1518 2574 -1512
rect 2568 -1524 2574 -1518
rect 2568 -1530 2574 -1524
rect 2568 -1536 2574 -1530
rect 2568 -1542 2574 -1536
rect 2568 -1548 2574 -1542
rect 2568 -1554 2574 -1548
rect 2568 -1560 2574 -1554
rect 2568 -1566 2574 -1560
rect 2568 -1572 2574 -1566
rect 2568 -1578 2574 -1572
rect 2568 -1584 2574 -1578
rect 2568 -1590 2574 -1584
rect 2568 -1596 2574 -1590
rect 2568 -1602 2574 -1596
rect 2568 -1608 2574 -1602
rect 2568 -1614 2574 -1608
rect 2568 -1620 2574 -1614
rect 2568 -1626 2574 -1620
rect 2568 -1632 2574 -1626
rect 2568 -1638 2574 -1632
rect 2568 -1644 2574 -1638
rect 2568 -1650 2574 -1644
rect 2568 -1656 2574 -1650
rect 2568 -1662 2574 -1656
rect 2568 -1668 2574 -1662
rect 2568 -1674 2574 -1668
rect 2568 -1680 2574 -1674
rect 2568 -1686 2574 -1680
rect 2568 -1692 2574 -1686
rect 2568 -1698 2574 -1692
rect 2568 -1704 2574 -1698
rect 2568 -1710 2574 -1704
rect 2568 -1716 2574 -1710
rect 2568 -1722 2574 -1716
rect 2568 -1728 2574 -1722
rect 2568 -1734 2574 -1728
rect 2568 -1740 2574 -1734
rect 2568 -1746 2574 -1740
rect 2568 -1752 2574 -1746
rect 2568 -1758 2574 -1752
rect 2568 -1764 2574 -1758
rect 2568 -1770 2574 -1764
rect 2568 -1776 2574 -1770
rect 2568 -1782 2574 -1776
rect 2568 -1788 2574 -1782
rect 2568 -1794 2574 -1788
rect 2568 -1800 2574 -1794
rect 2568 -1806 2574 -1800
rect 2568 -1812 2574 -1806
rect 2568 -1818 2574 -1812
rect 2568 -1824 2574 -1818
rect 2568 -1830 2574 -1824
rect 2568 -1836 2574 -1830
rect 2568 -1842 2574 -1836
rect 2568 -1848 2574 -1842
rect 2568 -1854 2574 -1848
rect 2568 -1860 2574 -1854
rect 2568 -1866 2574 -1860
rect 2568 -1872 2574 -1866
rect 2568 -1878 2574 -1872
rect 2568 -1884 2574 -1878
rect 2568 -1890 2574 -1884
rect 2568 -2430 2574 -2424
rect 2568 -2436 2574 -2430
rect 2568 -2442 2574 -2436
rect 2568 -2448 2574 -2442
rect 2568 -2454 2574 -2448
rect 2568 -2460 2574 -2454
rect 2568 -2466 2574 -2460
rect 2568 -2472 2574 -2466
rect 2568 -2478 2574 -2472
rect 2568 -2484 2574 -2478
rect 2568 -2490 2574 -2484
rect 2568 -2496 2574 -2490
rect 2568 -2502 2574 -2496
rect 2568 -2508 2574 -2502
rect 2568 -2514 2574 -2508
rect 2568 -2520 2574 -2514
rect 2568 -2526 2574 -2520
rect 2568 -2532 2574 -2526
rect 2568 -2538 2574 -2532
rect 2568 -2544 2574 -2538
rect 2568 -2550 2574 -2544
rect 2568 -2556 2574 -2550
rect 2568 -2562 2574 -2556
rect 2568 -2568 2574 -2562
rect 2568 -2574 2574 -2568
rect 2568 -2580 2574 -2574
rect 2568 -2586 2574 -2580
rect 2568 -2592 2574 -2586
rect 2568 -2598 2574 -2592
rect 2568 -2604 2574 -2598
rect 2568 -2610 2574 -2604
rect 2568 -2616 2574 -2610
rect 2568 -2622 2574 -2616
rect 2568 -2628 2574 -2622
rect 2568 -2634 2574 -2628
rect 2568 -2640 2574 -2634
rect 2568 -2646 2574 -2640
rect 2568 -2652 2574 -2646
rect 2568 -2658 2574 -2652
rect 2568 -2664 2574 -2658
rect 2568 -2670 2574 -2664
rect 2568 -2676 2574 -2670
rect 2568 -2682 2574 -2676
rect 2568 -2688 2574 -2682
rect 2568 -2694 2574 -2688
rect 2568 -2700 2574 -2694
rect 2568 -2706 2574 -2700
rect 2568 -2712 2574 -2706
rect 2568 -2718 2574 -2712
rect 2568 -2724 2574 -2718
rect 2568 -2730 2574 -2724
rect 2568 -2736 2574 -2730
rect 2568 -2742 2574 -2736
rect 2568 -2748 2574 -2742
rect 2568 -2754 2574 -2748
rect 2568 -2760 2574 -2754
rect 2568 -2766 2574 -2760
rect 2568 -2772 2574 -2766
rect 2568 -2778 2574 -2772
rect 2568 -2784 2574 -2778
rect 2574 -1254 2580 -1248
rect 2574 -1260 2580 -1254
rect 2574 -1266 2580 -1260
rect 2574 -1272 2580 -1266
rect 2574 -1278 2580 -1272
rect 2574 -1284 2580 -1278
rect 2574 -1290 2580 -1284
rect 2574 -1296 2580 -1290
rect 2574 -1302 2580 -1296
rect 2574 -1308 2580 -1302
rect 2574 -1314 2580 -1308
rect 2574 -1320 2580 -1314
rect 2574 -1326 2580 -1320
rect 2574 -1332 2580 -1326
rect 2574 -1338 2580 -1332
rect 2574 -1344 2580 -1338
rect 2574 -1350 2580 -1344
rect 2574 -1356 2580 -1350
rect 2574 -1362 2580 -1356
rect 2574 -1368 2580 -1362
rect 2574 -1374 2580 -1368
rect 2574 -1380 2580 -1374
rect 2574 -1386 2580 -1380
rect 2574 -1392 2580 -1386
rect 2574 -1398 2580 -1392
rect 2574 -1404 2580 -1398
rect 2574 -1410 2580 -1404
rect 2574 -1416 2580 -1410
rect 2574 -1422 2580 -1416
rect 2574 -1428 2580 -1422
rect 2574 -1434 2580 -1428
rect 2574 -1440 2580 -1434
rect 2574 -1446 2580 -1440
rect 2574 -1452 2580 -1446
rect 2574 -1458 2580 -1452
rect 2574 -1464 2580 -1458
rect 2574 -1470 2580 -1464
rect 2574 -1476 2580 -1470
rect 2574 -1482 2580 -1476
rect 2574 -1488 2580 -1482
rect 2574 -1494 2580 -1488
rect 2574 -1500 2580 -1494
rect 2574 -1506 2580 -1500
rect 2574 -1512 2580 -1506
rect 2574 -1518 2580 -1512
rect 2574 -1524 2580 -1518
rect 2574 -1530 2580 -1524
rect 2574 -1536 2580 -1530
rect 2574 -1542 2580 -1536
rect 2574 -1548 2580 -1542
rect 2574 -1554 2580 -1548
rect 2574 -1560 2580 -1554
rect 2574 -1566 2580 -1560
rect 2574 -1572 2580 -1566
rect 2574 -1578 2580 -1572
rect 2574 -1584 2580 -1578
rect 2574 -1590 2580 -1584
rect 2574 -1596 2580 -1590
rect 2574 -1602 2580 -1596
rect 2574 -1608 2580 -1602
rect 2574 -1614 2580 -1608
rect 2574 -1620 2580 -1614
rect 2574 -1626 2580 -1620
rect 2574 -1632 2580 -1626
rect 2574 -1638 2580 -1632
rect 2574 -1644 2580 -1638
rect 2574 -1650 2580 -1644
rect 2574 -1656 2580 -1650
rect 2574 -1662 2580 -1656
rect 2574 -1668 2580 -1662
rect 2574 -1674 2580 -1668
rect 2574 -1680 2580 -1674
rect 2574 -1686 2580 -1680
rect 2574 -1692 2580 -1686
rect 2574 -1698 2580 -1692
rect 2574 -1704 2580 -1698
rect 2574 -1710 2580 -1704
rect 2574 -1716 2580 -1710
rect 2574 -1722 2580 -1716
rect 2574 -1728 2580 -1722
rect 2574 -1734 2580 -1728
rect 2574 -1740 2580 -1734
rect 2574 -1746 2580 -1740
rect 2574 -1752 2580 -1746
rect 2574 -1758 2580 -1752
rect 2574 -1764 2580 -1758
rect 2574 -1770 2580 -1764
rect 2574 -1776 2580 -1770
rect 2574 -1782 2580 -1776
rect 2574 -1788 2580 -1782
rect 2574 -1794 2580 -1788
rect 2574 -1800 2580 -1794
rect 2574 -1806 2580 -1800
rect 2574 -1812 2580 -1806
rect 2574 -1818 2580 -1812
rect 2574 -1824 2580 -1818
rect 2574 -1830 2580 -1824
rect 2574 -1836 2580 -1830
rect 2574 -1842 2580 -1836
rect 2574 -1848 2580 -1842
rect 2574 -1854 2580 -1848
rect 2574 -1860 2580 -1854
rect 2574 -1866 2580 -1860
rect 2574 -1872 2580 -1866
rect 2574 -1878 2580 -1872
rect 2574 -1884 2580 -1878
rect 2574 -2430 2580 -2424
rect 2574 -2436 2580 -2430
rect 2574 -2442 2580 -2436
rect 2574 -2448 2580 -2442
rect 2574 -2454 2580 -2448
rect 2574 -2460 2580 -2454
rect 2574 -2466 2580 -2460
rect 2574 -2472 2580 -2466
rect 2574 -2478 2580 -2472
rect 2574 -2484 2580 -2478
rect 2574 -2490 2580 -2484
rect 2574 -2496 2580 -2490
rect 2574 -2502 2580 -2496
rect 2574 -2508 2580 -2502
rect 2574 -2514 2580 -2508
rect 2574 -2520 2580 -2514
rect 2574 -2526 2580 -2520
rect 2574 -2532 2580 -2526
rect 2574 -2538 2580 -2532
rect 2574 -2544 2580 -2538
rect 2574 -2550 2580 -2544
rect 2574 -2556 2580 -2550
rect 2574 -2562 2580 -2556
rect 2574 -2568 2580 -2562
rect 2574 -2574 2580 -2568
rect 2574 -2580 2580 -2574
rect 2574 -2586 2580 -2580
rect 2574 -2592 2580 -2586
rect 2574 -2598 2580 -2592
rect 2574 -2604 2580 -2598
rect 2574 -2610 2580 -2604
rect 2574 -2616 2580 -2610
rect 2574 -2622 2580 -2616
rect 2574 -2628 2580 -2622
rect 2574 -2634 2580 -2628
rect 2574 -2640 2580 -2634
rect 2574 -2646 2580 -2640
rect 2574 -2652 2580 -2646
rect 2574 -2658 2580 -2652
rect 2574 -2664 2580 -2658
rect 2574 -2670 2580 -2664
rect 2574 -2676 2580 -2670
rect 2574 -2682 2580 -2676
rect 2574 -2688 2580 -2682
rect 2574 -2694 2580 -2688
rect 2574 -2700 2580 -2694
rect 2574 -2706 2580 -2700
rect 2574 -2712 2580 -2706
rect 2574 -2718 2580 -2712
rect 2574 -2724 2580 -2718
rect 2574 -2730 2580 -2724
rect 2574 -2736 2580 -2730
rect 2574 -2742 2580 -2736
rect 2574 -2748 2580 -2742
rect 2574 -2754 2580 -2748
rect 2574 -2760 2580 -2754
rect 2574 -2766 2580 -2760
rect 2574 -2772 2580 -2766
rect 2574 -2778 2580 -2772
rect 2580 -1248 2586 -1242
rect 2580 -1254 2586 -1248
rect 2580 -1260 2586 -1254
rect 2580 -1266 2586 -1260
rect 2580 -1272 2586 -1266
rect 2580 -1278 2586 -1272
rect 2580 -1284 2586 -1278
rect 2580 -1290 2586 -1284
rect 2580 -1296 2586 -1290
rect 2580 -1302 2586 -1296
rect 2580 -1308 2586 -1302
rect 2580 -1314 2586 -1308
rect 2580 -1320 2586 -1314
rect 2580 -1326 2586 -1320
rect 2580 -1332 2586 -1326
rect 2580 -1338 2586 -1332
rect 2580 -1344 2586 -1338
rect 2580 -1350 2586 -1344
rect 2580 -1356 2586 -1350
rect 2580 -1362 2586 -1356
rect 2580 -1368 2586 -1362
rect 2580 -1374 2586 -1368
rect 2580 -1380 2586 -1374
rect 2580 -1386 2586 -1380
rect 2580 -1392 2586 -1386
rect 2580 -1398 2586 -1392
rect 2580 -1404 2586 -1398
rect 2580 -1410 2586 -1404
rect 2580 -1416 2586 -1410
rect 2580 -1422 2586 -1416
rect 2580 -1428 2586 -1422
rect 2580 -1434 2586 -1428
rect 2580 -1440 2586 -1434
rect 2580 -1446 2586 -1440
rect 2580 -1452 2586 -1446
rect 2580 -1458 2586 -1452
rect 2580 -1464 2586 -1458
rect 2580 -1470 2586 -1464
rect 2580 -1476 2586 -1470
rect 2580 -1482 2586 -1476
rect 2580 -1488 2586 -1482
rect 2580 -1494 2586 -1488
rect 2580 -1500 2586 -1494
rect 2580 -1506 2586 -1500
rect 2580 -1512 2586 -1506
rect 2580 -1518 2586 -1512
rect 2580 -1524 2586 -1518
rect 2580 -1530 2586 -1524
rect 2580 -1536 2586 -1530
rect 2580 -1542 2586 -1536
rect 2580 -1548 2586 -1542
rect 2580 -1554 2586 -1548
rect 2580 -1560 2586 -1554
rect 2580 -1566 2586 -1560
rect 2580 -1572 2586 -1566
rect 2580 -1578 2586 -1572
rect 2580 -1584 2586 -1578
rect 2580 -1590 2586 -1584
rect 2580 -1596 2586 -1590
rect 2580 -1602 2586 -1596
rect 2580 -1608 2586 -1602
rect 2580 -1614 2586 -1608
rect 2580 -1620 2586 -1614
rect 2580 -1626 2586 -1620
rect 2580 -1632 2586 -1626
rect 2580 -1638 2586 -1632
rect 2580 -1644 2586 -1638
rect 2580 -1650 2586 -1644
rect 2580 -1656 2586 -1650
rect 2580 -1662 2586 -1656
rect 2580 -1668 2586 -1662
rect 2580 -1674 2586 -1668
rect 2580 -1680 2586 -1674
rect 2580 -1686 2586 -1680
rect 2580 -1692 2586 -1686
rect 2580 -1698 2586 -1692
rect 2580 -1704 2586 -1698
rect 2580 -1710 2586 -1704
rect 2580 -1716 2586 -1710
rect 2580 -1722 2586 -1716
rect 2580 -1728 2586 -1722
rect 2580 -1734 2586 -1728
rect 2580 -1740 2586 -1734
rect 2580 -1746 2586 -1740
rect 2580 -1752 2586 -1746
rect 2580 -1758 2586 -1752
rect 2580 -1764 2586 -1758
rect 2580 -1770 2586 -1764
rect 2580 -1776 2586 -1770
rect 2580 -1782 2586 -1776
rect 2580 -1788 2586 -1782
rect 2580 -1794 2586 -1788
rect 2580 -1800 2586 -1794
rect 2580 -1806 2586 -1800
rect 2580 -1812 2586 -1806
rect 2580 -1818 2586 -1812
rect 2580 -1824 2586 -1818
rect 2580 -1830 2586 -1824
rect 2580 -1836 2586 -1830
rect 2580 -1842 2586 -1836
rect 2580 -1848 2586 -1842
rect 2580 -1854 2586 -1848
rect 2580 -1860 2586 -1854
rect 2580 -1866 2586 -1860
rect 2580 -1872 2586 -1866
rect 2580 -1878 2586 -1872
rect 2580 -2430 2586 -2424
rect 2580 -2436 2586 -2430
rect 2580 -2442 2586 -2436
rect 2580 -2448 2586 -2442
rect 2580 -2454 2586 -2448
rect 2580 -2460 2586 -2454
rect 2580 -2466 2586 -2460
rect 2580 -2472 2586 -2466
rect 2580 -2478 2586 -2472
rect 2580 -2484 2586 -2478
rect 2580 -2490 2586 -2484
rect 2580 -2496 2586 -2490
rect 2580 -2502 2586 -2496
rect 2580 -2508 2586 -2502
rect 2580 -2514 2586 -2508
rect 2580 -2520 2586 -2514
rect 2580 -2526 2586 -2520
rect 2580 -2532 2586 -2526
rect 2580 -2538 2586 -2532
rect 2580 -2544 2586 -2538
rect 2580 -2550 2586 -2544
rect 2580 -2556 2586 -2550
rect 2580 -2562 2586 -2556
rect 2580 -2568 2586 -2562
rect 2580 -2574 2586 -2568
rect 2580 -2580 2586 -2574
rect 2580 -2586 2586 -2580
rect 2580 -2592 2586 -2586
rect 2580 -2598 2586 -2592
rect 2580 -2604 2586 -2598
rect 2580 -2610 2586 -2604
rect 2580 -2616 2586 -2610
rect 2580 -2622 2586 -2616
rect 2580 -2628 2586 -2622
rect 2580 -2634 2586 -2628
rect 2580 -2640 2586 -2634
rect 2580 -2646 2586 -2640
rect 2580 -2652 2586 -2646
rect 2580 -2658 2586 -2652
rect 2580 -2664 2586 -2658
rect 2580 -2670 2586 -2664
rect 2580 -2676 2586 -2670
rect 2580 -2682 2586 -2676
rect 2580 -2688 2586 -2682
rect 2580 -2694 2586 -2688
rect 2580 -2700 2586 -2694
rect 2580 -2706 2586 -2700
rect 2580 -2712 2586 -2706
rect 2580 -2718 2586 -2712
rect 2580 -2724 2586 -2718
rect 2580 -2730 2586 -2724
rect 2580 -2736 2586 -2730
rect 2580 -2742 2586 -2736
rect 2580 -2748 2586 -2742
rect 2580 -2754 2586 -2748
rect 2580 -2760 2586 -2754
rect 2580 -2766 2586 -2760
rect 2580 -2772 2586 -2766
rect 2580 -2778 2586 -2772
rect 2586 -1242 2592 -1236
rect 2586 -1248 2592 -1242
rect 2586 -1254 2592 -1248
rect 2586 -1260 2592 -1254
rect 2586 -1266 2592 -1260
rect 2586 -1272 2592 -1266
rect 2586 -1278 2592 -1272
rect 2586 -1284 2592 -1278
rect 2586 -1290 2592 -1284
rect 2586 -1296 2592 -1290
rect 2586 -1302 2592 -1296
rect 2586 -1308 2592 -1302
rect 2586 -1314 2592 -1308
rect 2586 -1320 2592 -1314
rect 2586 -1326 2592 -1320
rect 2586 -1332 2592 -1326
rect 2586 -1338 2592 -1332
rect 2586 -1344 2592 -1338
rect 2586 -1350 2592 -1344
rect 2586 -1356 2592 -1350
rect 2586 -1362 2592 -1356
rect 2586 -1368 2592 -1362
rect 2586 -1374 2592 -1368
rect 2586 -1380 2592 -1374
rect 2586 -1386 2592 -1380
rect 2586 -1392 2592 -1386
rect 2586 -1398 2592 -1392
rect 2586 -1404 2592 -1398
rect 2586 -1410 2592 -1404
rect 2586 -1416 2592 -1410
rect 2586 -1422 2592 -1416
rect 2586 -1428 2592 -1422
rect 2586 -1434 2592 -1428
rect 2586 -1440 2592 -1434
rect 2586 -1446 2592 -1440
rect 2586 -1452 2592 -1446
rect 2586 -1458 2592 -1452
rect 2586 -1464 2592 -1458
rect 2586 -1470 2592 -1464
rect 2586 -1476 2592 -1470
rect 2586 -1482 2592 -1476
rect 2586 -1488 2592 -1482
rect 2586 -1494 2592 -1488
rect 2586 -1500 2592 -1494
rect 2586 -1506 2592 -1500
rect 2586 -1512 2592 -1506
rect 2586 -1518 2592 -1512
rect 2586 -1524 2592 -1518
rect 2586 -1530 2592 -1524
rect 2586 -1536 2592 -1530
rect 2586 -1542 2592 -1536
rect 2586 -1548 2592 -1542
rect 2586 -1554 2592 -1548
rect 2586 -1560 2592 -1554
rect 2586 -1566 2592 -1560
rect 2586 -1572 2592 -1566
rect 2586 -1578 2592 -1572
rect 2586 -1584 2592 -1578
rect 2586 -1590 2592 -1584
rect 2586 -1596 2592 -1590
rect 2586 -1602 2592 -1596
rect 2586 -1608 2592 -1602
rect 2586 -1614 2592 -1608
rect 2586 -1620 2592 -1614
rect 2586 -1626 2592 -1620
rect 2586 -1632 2592 -1626
rect 2586 -1638 2592 -1632
rect 2586 -1644 2592 -1638
rect 2586 -1650 2592 -1644
rect 2586 -1656 2592 -1650
rect 2586 -1662 2592 -1656
rect 2586 -1668 2592 -1662
rect 2586 -1674 2592 -1668
rect 2586 -1680 2592 -1674
rect 2586 -1686 2592 -1680
rect 2586 -1692 2592 -1686
rect 2586 -1698 2592 -1692
rect 2586 -1704 2592 -1698
rect 2586 -1710 2592 -1704
rect 2586 -1716 2592 -1710
rect 2586 -1722 2592 -1716
rect 2586 -1728 2592 -1722
rect 2586 -1734 2592 -1728
rect 2586 -1740 2592 -1734
rect 2586 -1746 2592 -1740
rect 2586 -1752 2592 -1746
rect 2586 -1758 2592 -1752
rect 2586 -1764 2592 -1758
rect 2586 -1770 2592 -1764
rect 2586 -1776 2592 -1770
rect 2586 -1782 2592 -1776
rect 2586 -1788 2592 -1782
rect 2586 -1794 2592 -1788
rect 2586 -1800 2592 -1794
rect 2586 -1806 2592 -1800
rect 2586 -1812 2592 -1806
rect 2586 -1818 2592 -1812
rect 2586 -1824 2592 -1818
rect 2586 -1830 2592 -1824
rect 2586 -1836 2592 -1830
rect 2586 -1842 2592 -1836
rect 2586 -1848 2592 -1842
rect 2586 -1854 2592 -1848
rect 2586 -1860 2592 -1854
rect 2586 -1866 2592 -1860
rect 2586 -2430 2592 -2424
rect 2586 -2436 2592 -2430
rect 2586 -2442 2592 -2436
rect 2586 -2448 2592 -2442
rect 2586 -2454 2592 -2448
rect 2586 -2460 2592 -2454
rect 2586 -2466 2592 -2460
rect 2586 -2472 2592 -2466
rect 2586 -2478 2592 -2472
rect 2586 -2484 2592 -2478
rect 2586 -2490 2592 -2484
rect 2586 -2496 2592 -2490
rect 2586 -2502 2592 -2496
rect 2586 -2508 2592 -2502
rect 2586 -2514 2592 -2508
rect 2586 -2520 2592 -2514
rect 2586 -2526 2592 -2520
rect 2586 -2532 2592 -2526
rect 2586 -2538 2592 -2532
rect 2586 -2544 2592 -2538
rect 2586 -2550 2592 -2544
rect 2586 -2556 2592 -2550
rect 2586 -2562 2592 -2556
rect 2586 -2568 2592 -2562
rect 2586 -2574 2592 -2568
rect 2586 -2580 2592 -2574
rect 2586 -2586 2592 -2580
rect 2586 -2592 2592 -2586
rect 2586 -2598 2592 -2592
rect 2586 -2604 2592 -2598
rect 2586 -2610 2592 -2604
rect 2586 -2616 2592 -2610
rect 2586 -2622 2592 -2616
rect 2586 -2628 2592 -2622
rect 2586 -2634 2592 -2628
rect 2586 -2640 2592 -2634
rect 2586 -2646 2592 -2640
rect 2586 -2652 2592 -2646
rect 2586 -2658 2592 -2652
rect 2586 -2664 2592 -2658
rect 2586 -2670 2592 -2664
rect 2586 -2676 2592 -2670
rect 2586 -2682 2592 -2676
rect 2586 -2688 2592 -2682
rect 2586 -2694 2592 -2688
rect 2586 -2700 2592 -2694
rect 2586 -2706 2592 -2700
rect 2586 -2712 2592 -2706
rect 2586 -2718 2592 -2712
rect 2586 -2724 2592 -2718
rect 2586 -2730 2592 -2724
rect 2586 -2736 2592 -2730
rect 2586 -2742 2592 -2736
rect 2586 -2748 2592 -2742
rect 2586 -2754 2592 -2748
rect 2586 -2760 2592 -2754
rect 2586 -2766 2592 -2760
rect 2586 -2772 2592 -2766
rect 2592 -1242 2598 -1236
rect 2592 -1248 2598 -1242
rect 2592 -1254 2598 -1248
rect 2592 -1260 2598 -1254
rect 2592 -1266 2598 -1260
rect 2592 -1272 2598 -1266
rect 2592 -1278 2598 -1272
rect 2592 -1284 2598 -1278
rect 2592 -1290 2598 -1284
rect 2592 -1296 2598 -1290
rect 2592 -1302 2598 -1296
rect 2592 -1308 2598 -1302
rect 2592 -1314 2598 -1308
rect 2592 -1320 2598 -1314
rect 2592 -1326 2598 -1320
rect 2592 -1332 2598 -1326
rect 2592 -1338 2598 -1332
rect 2592 -1344 2598 -1338
rect 2592 -1350 2598 -1344
rect 2592 -1356 2598 -1350
rect 2592 -1362 2598 -1356
rect 2592 -1368 2598 -1362
rect 2592 -1374 2598 -1368
rect 2592 -1380 2598 -1374
rect 2592 -1386 2598 -1380
rect 2592 -1392 2598 -1386
rect 2592 -1398 2598 -1392
rect 2592 -1404 2598 -1398
rect 2592 -1410 2598 -1404
rect 2592 -1416 2598 -1410
rect 2592 -1422 2598 -1416
rect 2592 -1428 2598 -1422
rect 2592 -1434 2598 -1428
rect 2592 -1440 2598 -1434
rect 2592 -1446 2598 -1440
rect 2592 -1452 2598 -1446
rect 2592 -1458 2598 -1452
rect 2592 -1464 2598 -1458
rect 2592 -1470 2598 -1464
rect 2592 -1476 2598 -1470
rect 2592 -1482 2598 -1476
rect 2592 -1488 2598 -1482
rect 2592 -1494 2598 -1488
rect 2592 -1500 2598 -1494
rect 2592 -1506 2598 -1500
rect 2592 -1512 2598 -1506
rect 2592 -1518 2598 -1512
rect 2592 -1524 2598 -1518
rect 2592 -1530 2598 -1524
rect 2592 -1536 2598 -1530
rect 2592 -1542 2598 -1536
rect 2592 -1548 2598 -1542
rect 2592 -1554 2598 -1548
rect 2592 -1560 2598 -1554
rect 2592 -1566 2598 -1560
rect 2592 -1572 2598 -1566
rect 2592 -1578 2598 -1572
rect 2592 -1584 2598 -1578
rect 2592 -1590 2598 -1584
rect 2592 -1596 2598 -1590
rect 2592 -1602 2598 -1596
rect 2592 -1608 2598 -1602
rect 2592 -1614 2598 -1608
rect 2592 -1620 2598 -1614
rect 2592 -1626 2598 -1620
rect 2592 -1632 2598 -1626
rect 2592 -1638 2598 -1632
rect 2592 -1644 2598 -1638
rect 2592 -1650 2598 -1644
rect 2592 -1656 2598 -1650
rect 2592 -1662 2598 -1656
rect 2592 -1668 2598 -1662
rect 2592 -1674 2598 -1668
rect 2592 -1680 2598 -1674
rect 2592 -1686 2598 -1680
rect 2592 -1692 2598 -1686
rect 2592 -1698 2598 -1692
rect 2592 -1704 2598 -1698
rect 2592 -1710 2598 -1704
rect 2592 -1716 2598 -1710
rect 2592 -1722 2598 -1716
rect 2592 -1728 2598 -1722
rect 2592 -1734 2598 -1728
rect 2592 -1740 2598 -1734
rect 2592 -1746 2598 -1740
rect 2592 -1752 2598 -1746
rect 2592 -1758 2598 -1752
rect 2592 -1764 2598 -1758
rect 2592 -1770 2598 -1764
rect 2592 -1776 2598 -1770
rect 2592 -1782 2598 -1776
rect 2592 -1788 2598 -1782
rect 2592 -1794 2598 -1788
rect 2592 -1800 2598 -1794
rect 2592 -1806 2598 -1800
rect 2592 -1812 2598 -1806
rect 2592 -1818 2598 -1812
rect 2592 -1824 2598 -1818
rect 2592 -1830 2598 -1824
rect 2592 -1836 2598 -1830
rect 2592 -1842 2598 -1836
rect 2592 -1848 2598 -1842
rect 2592 -1854 2598 -1848
rect 2592 -1860 2598 -1854
rect 2592 -2424 2598 -2418
rect 2592 -2430 2598 -2424
rect 2592 -2436 2598 -2430
rect 2592 -2442 2598 -2436
rect 2592 -2448 2598 -2442
rect 2592 -2454 2598 -2448
rect 2592 -2460 2598 -2454
rect 2592 -2466 2598 -2460
rect 2592 -2472 2598 -2466
rect 2592 -2478 2598 -2472
rect 2592 -2484 2598 -2478
rect 2592 -2490 2598 -2484
rect 2592 -2496 2598 -2490
rect 2592 -2502 2598 -2496
rect 2592 -2508 2598 -2502
rect 2592 -2514 2598 -2508
rect 2592 -2520 2598 -2514
rect 2592 -2526 2598 -2520
rect 2592 -2532 2598 -2526
rect 2592 -2538 2598 -2532
rect 2592 -2544 2598 -2538
rect 2592 -2550 2598 -2544
rect 2592 -2556 2598 -2550
rect 2592 -2562 2598 -2556
rect 2592 -2568 2598 -2562
rect 2592 -2574 2598 -2568
rect 2592 -2580 2598 -2574
rect 2592 -2586 2598 -2580
rect 2592 -2592 2598 -2586
rect 2592 -2598 2598 -2592
rect 2592 -2604 2598 -2598
rect 2592 -2610 2598 -2604
rect 2592 -2616 2598 -2610
rect 2592 -2622 2598 -2616
rect 2592 -2628 2598 -2622
rect 2592 -2634 2598 -2628
rect 2592 -2640 2598 -2634
rect 2592 -2646 2598 -2640
rect 2592 -2652 2598 -2646
rect 2592 -2658 2598 -2652
rect 2592 -2664 2598 -2658
rect 2592 -2670 2598 -2664
rect 2592 -2676 2598 -2670
rect 2592 -2682 2598 -2676
rect 2592 -2688 2598 -2682
rect 2592 -2694 2598 -2688
rect 2592 -2700 2598 -2694
rect 2592 -2706 2598 -2700
rect 2592 -2712 2598 -2706
rect 2592 -2718 2598 -2712
rect 2592 -2724 2598 -2718
rect 2592 -2730 2598 -2724
rect 2592 -2736 2598 -2730
rect 2592 -2742 2598 -2736
rect 2592 -2748 2598 -2742
rect 2592 -2754 2598 -2748
rect 2592 -2760 2598 -2754
rect 2592 -2766 2598 -2760
rect 2598 -1236 2604 -1230
rect 2598 -1242 2604 -1236
rect 2598 -1248 2604 -1242
rect 2598 -1254 2604 -1248
rect 2598 -1260 2604 -1254
rect 2598 -1266 2604 -1260
rect 2598 -1272 2604 -1266
rect 2598 -1278 2604 -1272
rect 2598 -1284 2604 -1278
rect 2598 -1290 2604 -1284
rect 2598 -1296 2604 -1290
rect 2598 -1302 2604 -1296
rect 2598 -1308 2604 -1302
rect 2598 -1314 2604 -1308
rect 2598 -1320 2604 -1314
rect 2598 -1326 2604 -1320
rect 2598 -1332 2604 -1326
rect 2598 -1338 2604 -1332
rect 2598 -1344 2604 -1338
rect 2598 -1350 2604 -1344
rect 2598 -1356 2604 -1350
rect 2598 -1362 2604 -1356
rect 2598 -1368 2604 -1362
rect 2598 -1374 2604 -1368
rect 2598 -1380 2604 -1374
rect 2598 -1386 2604 -1380
rect 2598 -1392 2604 -1386
rect 2598 -1398 2604 -1392
rect 2598 -1404 2604 -1398
rect 2598 -1410 2604 -1404
rect 2598 -1416 2604 -1410
rect 2598 -1422 2604 -1416
rect 2598 -1428 2604 -1422
rect 2598 -1434 2604 -1428
rect 2598 -1440 2604 -1434
rect 2598 -1446 2604 -1440
rect 2598 -1452 2604 -1446
rect 2598 -1458 2604 -1452
rect 2598 -1464 2604 -1458
rect 2598 -1470 2604 -1464
rect 2598 -1476 2604 -1470
rect 2598 -1482 2604 -1476
rect 2598 -1488 2604 -1482
rect 2598 -1494 2604 -1488
rect 2598 -1500 2604 -1494
rect 2598 -1506 2604 -1500
rect 2598 -1512 2604 -1506
rect 2598 -1518 2604 -1512
rect 2598 -1524 2604 -1518
rect 2598 -1530 2604 -1524
rect 2598 -1536 2604 -1530
rect 2598 -1542 2604 -1536
rect 2598 -1548 2604 -1542
rect 2598 -1554 2604 -1548
rect 2598 -1560 2604 -1554
rect 2598 -1566 2604 -1560
rect 2598 -1572 2604 -1566
rect 2598 -1578 2604 -1572
rect 2598 -1584 2604 -1578
rect 2598 -1590 2604 -1584
rect 2598 -1596 2604 -1590
rect 2598 -1602 2604 -1596
rect 2598 -1608 2604 -1602
rect 2598 -1614 2604 -1608
rect 2598 -1620 2604 -1614
rect 2598 -1626 2604 -1620
rect 2598 -1632 2604 -1626
rect 2598 -1638 2604 -1632
rect 2598 -1644 2604 -1638
rect 2598 -1650 2604 -1644
rect 2598 -1656 2604 -1650
rect 2598 -1662 2604 -1656
rect 2598 -1668 2604 -1662
rect 2598 -1674 2604 -1668
rect 2598 -1680 2604 -1674
rect 2598 -1686 2604 -1680
rect 2598 -1692 2604 -1686
rect 2598 -1698 2604 -1692
rect 2598 -1704 2604 -1698
rect 2598 -1710 2604 -1704
rect 2598 -1716 2604 -1710
rect 2598 -1722 2604 -1716
rect 2598 -1728 2604 -1722
rect 2598 -1734 2604 -1728
rect 2598 -1740 2604 -1734
rect 2598 -1746 2604 -1740
rect 2598 -1752 2604 -1746
rect 2598 -1758 2604 -1752
rect 2598 -1764 2604 -1758
rect 2598 -1770 2604 -1764
rect 2598 -1776 2604 -1770
rect 2598 -1782 2604 -1776
rect 2598 -1788 2604 -1782
rect 2598 -1794 2604 -1788
rect 2598 -1800 2604 -1794
rect 2598 -1806 2604 -1800
rect 2598 -1812 2604 -1806
rect 2598 -1818 2604 -1812
rect 2598 -1824 2604 -1818
rect 2598 -1830 2604 -1824
rect 2598 -1836 2604 -1830
rect 2598 -1842 2604 -1836
rect 2598 -1848 2604 -1842
rect 2598 -1854 2604 -1848
rect 2598 -2424 2604 -2418
rect 2598 -2430 2604 -2424
rect 2598 -2436 2604 -2430
rect 2598 -2442 2604 -2436
rect 2598 -2448 2604 -2442
rect 2598 -2454 2604 -2448
rect 2598 -2460 2604 -2454
rect 2598 -2466 2604 -2460
rect 2598 -2472 2604 -2466
rect 2598 -2478 2604 -2472
rect 2598 -2484 2604 -2478
rect 2598 -2490 2604 -2484
rect 2598 -2496 2604 -2490
rect 2598 -2502 2604 -2496
rect 2598 -2508 2604 -2502
rect 2598 -2514 2604 -2508
rect 2598 -2520 2604 -2514
rect 2598 -2526 2604 -2520
rect 2598 -2532 2604 -2526
rect 2598 -2538 2604 -2532
rect 2598 -2544 2604 -2538
rect 2598 -2550 2604 -2544
rect 2598 -2556 2604 -2550
rect 2598 -2562 2604 -2556
rect 2598 -2568 2604 -2562
rect 2598 -2574 2604 -2568
rect 2598 -2580 2604 -2574
rect 2598 -2586 2604 -2580
rect 2598 -2592 2604 -2586
rect 2598 -2598 2604 -2592
rect 2598 -2604 2604 -2598
rect 2598 -2610 2604 -2604
rect 2598 -2616 2604 -2610
rect 2598 -2622 2604 -2616
rect 2598 -2628 2604 -2622
rect 2598 -2634 2604 -2628
rect 2598 -2640 2604 -2634
rect 2598 -2646 2604 -2640
rect 2598 -2652 2604 -2646
rect 2598 -2658 2604 -2652
rect 2598 -2664 2604 -2658
rect 2598 -2670 2604 -2664
rect 2598 -2676 2604 -2670
rect 2598 -2682 2604 -2676
rect 2598 -2688 2604 -2682
rect 2598 -2694 2604 -2688
rect 2598 -2700 2604 -2694
rect 2598 -2706 2604 -2700
rect 2598 -2712 2604 -2706
rect 2598 -2718 2604 -2712
rect 2598 -2724 2604 -2718
rect 2598 -2730 2604 -2724
rect 2598 -2736 2604 -2730
rect 2598 -2742 2604 -2736
rect 2598 -2748 2604 -2742
rect 2598 -2754 2604 -2748
rect 2598 -2760 2604 -2754
rect 2598 -2766 2604 -2760
rect 2604 -1230 2610 -1224
rect 2604 -1236 2610 -1230
rect 2604 -1242 2610 -1236
rect 2604 -1248 2610 -1242
rect 2604 -1254 2610 -1248
rect 2604 -1260 2610 -1254
rect 2604 -1266 2610 -1260
rect 2604 -1272 2610 -1266
rect 2604 -1278 2610 -1272
rect 2604 -1284 2610 -1278
rect 2604 -1290 2610 -1284
rect 2604 -1296 2610 -1290
rect 2604 -1302 2610 -1296
rect 2604 -1308 2610 -1302
rect 2604 -1314 2610 -1308
rect 2604 -1320 2610 -1314
rect 2604 -1326 2610 -1320
rect 2604 -1332 2610 -1326
rect 2604 -1338 2610 -1332
rect 2604 -1344 2610 -1338
rect 2604 -1350 2610 -1344
rect 2604 -1356 2610 -1350
rect 2604 -1362 2610 -1356
rect 2604 -1368 2610 -1362
rect 2604 -1374 2610 -1368
rect 2604 -1380 2610 -1374
rect 2604 -1386 2610 -1380
rect 2604 -1392 2610 -1386
rect 2604 -1398 2610 -1392
rect 2604 -1404 2610 -1398
rect 2604 -1410 2610 -1404
rect 2604 -1416 2610 -1410
rect 2604 -1422 2610 -1416
rect 2604 -1428 2610 -1422
rect 2604 -1434 2610 -1428
rect 2604 -1440 2610 -1434
rect 2604 -1446 2610 -1440
rect 2604 -1452 2610 -1446
rect 2604 -1458 2610 -1452
rect 2604 -1464 2610 -1458
rect 2604 -1470 2610 -1464
rect 2604 -1476 2610 -1470
rect 2604 -1482 2610 -1476
rect 2604 -1488 2610 -1482
rect 2604 -1494 2610 -1488
rect 2604 -1500 2610 -1494
rect 2604 -1506 2610 -1500
rect 2604 -1512 2610 -1506
rect 2604 -1518 2610 -1512
rect 2604 -1524 2610 -1518
rect 2604 -1530 2610 -1524
rect 2604 -1536 2610 -1530
rect 2604 -1542 2610 -1536
rect 2604 -1548 2610 -1542
rect 2604 -1554 2610 -1548
rect 2604 -1560 2610 -1554
rect 2604 -1566 2610 -1560
rect 2604 -1572 2610 -1566
rect 2604 -1578 2610 -1572
rect 2604 -1584 2610 -1578
rect 2604 -1590 2610 -1584
rect 2604 -1596 2610 -1590
rect 2604 -1602 2610 -1596
rect 2604 -1608 2610 -1602
rect 2604 -1614 2610 -1608
rect 2604 -1620 2610 -1614
rect 2604 -1626 2610 -1620
rect 2604 -1632 2610 -1626
rect 2604 -1638 2610 -1632
rect 2604 -1644 2610 -1638
rect 2604 -1650 2610 -1644
rect 2604 -1656 2610 -1650
rect 2604 -1662 2610 -1656
rect 2604 -1668 2610 -1662
rect 2604 -1674 2610 -1668
rect 2604 -1680 2610 -1674
rect 2604 -1686 2610 -1680
rect 2604 -1692 2610 -1686
rect 2604 -1698 2610 -1692
rect 2604 -1704 2610 -1698
rect 2604 -1710 2610 -1704
rect 2604 -1716 2610 -1710
rect 2604 -1722 2610 -1716
rect 2604 -1728 2610 -1722
rect 2604 -1734 2610 -1728
rect 2604 -1740 2610 -1734
rect 2604 -1746 2610 -1740
rect 2604 -1752 2610 -1746
rect 2604 -1758 2610 -1752
rect 2604 -1764 2610 -1758
rect 2604 -1770 2610 -1764
rect 2604 -1776 2610 -1770
rect 2604 -1782 2610 -1776
rect 2604 -1788 2610 -1782
rect 2604 -1794 2610 -1788
rect 2604 -1800 2610 -1794
rect 2604 -1806 2610 -1800
rect 2604 -1812 2610 -1806
rect 2604 -1818 2610 -1812
rect 2604 -1824 2610 -1818
rect 2604 -1830 2610 -1824
rect 2604 -1836 2610 -1830
rect 2604 -1842 2610 -1836
rect 2604 -1848 2610 -1842
rect 2604 -2424 2610 -2418
rect 2604 -2430 2610 -2424
rect 2604 -2436 2610 -2430
rect 2604 -2442 2610 -2436
rect 2604 -2448 2610 -2442
rect 2604 -2454 2610 -2448
rect 2604 -2460 2610 -2454
rect 2604 -2466 2610 -2460
rect 2604 -2472 2610 -2466
rect 2604 -2478 2610 -2472
rect 2604 -2484 2610 -2478
rect 2604 -2490 2610 -2484
rect 2604 -2496 2610 -2490
rect 2604 -2502 2610 -2496
rect 2604 -2508 2610 -2502
rect 2604 -2514 2610 -2508
rect 2604 -2520 2610 -2514
rect 2604 -2526 2610 -2520
rect 2604 -2532 2610 -2526
rect 2604 -2538 2610 -2532
rect 2604 -2544 2610 -2538
rect 2604 -2550 2610 -2544
rect 2604 -2556 2610 -2550
rect 2604 -2562 2610 -2556
rect 2604 -2568 2610 -2562
rect 2604 -2574 2610 -2568
rect 2604 -2580 2610 -2574
rect 2604 -2586 2610 -2580
rect 2604 -2592 2610 -2586
rect 2604 -2598 2610 -2592
rect 2604 -2604 2610 -2598
rect 2604 -2610 2610 -2604
rect 2604 -2616 2610 -2610
rect 2604 -2622 2610 -2616
rect 2604 -2628 2610 -2622
rect 2604 -2634 2610 -2628
rect 2604 -2640 2610 -2634
rect 2604 -2646 2610 -2640
rect 2604 -2652 2610 -2646
rect 2604 -2658 2610 -2652
rect 2604 -2664 2610 -2658
rect 2604 -2670 2610 -2664
rect 2604 -2676 2610 -2670
rect 2604 -2682 2610 -2676
rect 2604 -2688 2610 -2682
rect 2604 -2694 2610 -2688
rect 2604 -2700 2610 -2694
rect 2604 -2706 2610 -2700
rect 2604 -2712 2610 -2706
rect 2604 -2718 2610 -2712
rect 2604 -2724 2610 -2718
rect 2604 -2730 2610 -2724
rect 2604 -2736 2610 -2730
rect 2604 -2742 2610 -2736
rect 2604 -2748 2610 -2742
rect 2604 -2754 2610 -2748
rect 2604 -2760 2610 -2754
rect 2610 -1224 2616 -1218
rect 2610 -1230 2616 -1224
rect 2610 -1236 2616 -1230
rect 2610 -1242 2616 -1236
rect 2610 -1248 2616 -1242
rect 2610 -1254 2616 -1248
rect 2610 -1260 2616 -1254
rect 2610 -1266 2616 -1260
rect 2610 -1272 2616 -1266
rect 2610 -1278 2616 -1272
rect 2610 -1284 2616 -1278
rect 2610 -1290 2616 -1284
rect 2610 -1296 2616 -1290
rect 2610 -1302 2616 -1296
rect 2610 -1308 2616 -1302
rect 2610 -1314 2616 -1308
rect 2610 -1320 2616 -1314
rect 2610 -1326 2616 -1320
rect 2610 -1332 2616 -1326
rect 2610 -1338 2616 -1332
rect 2610 -1344 2616 -1338
rect 2610 -1350 2616 -1344
rect 2610 -1356 2616 -1350
rect 2610 -1362 2616 -1356
rect 2610 -1368 2616 -1362
rect 2610 -1374 2616 -1368
rect 2610 -1380 2616 -1374
rect 2610 -1386 2616 -1380
rect 2610 -1392 2616 -1386
rect 2610 -1398 2616 -1392
rect 2610 -1404 2616 -1398
rect 2610 -1410 2616 -1404
rect 2610 -1416 2616 -1410
rect 2610 -1422 2616 -1416
rect 2610 -1428 2616 -1422
rect 2610 -1434 2616 -1428
rect 2610 -1440 2616 -1434
rect 2610 -1446 2616 -1440
rect 2610 -1452 2616 -1446
rect 2610 -1458 2616 -1452
rect 2610 -1464 2616 -1458
rect 2610 -1470 2616 -1464
rect 2610 -1476 2616 -1470
rect 2610 -1482 2616 -1476
rect 2610 -1488 2616 -1482
rect 2610 -1494 2616 -1488
rect 2610 -1500 2616 -1494
rect 2610 -1506 2616 -1500
rect 2610 -1512 2616 -1506
rect 2610 -1518 2616 -1512
rect 2610 -1524 2616 -1518
rect 2610 -1530 2616 -1524
rect 2610 -1536 2616 -1530
rect 2610 -1542 2616 -1536
rect 2610 -1548 2616 -1542
rect 2610 -1554 2616 -1548
rect 2610 -1560 2616 -1554
rect 2610 -1566 2616 -1560
rect 2610 -1572 2616 -1566
rect 2610 -1578 2616 -1572
rect 2610 -1584 2616 -1578
rect 2610 -1590 2616 -1584
rect 2610 -1596 2616 -1590
rect 2610 -1602 2616 -1596
rect 2610 -1608 2616 -1602
rect 2610 -1614 2616 -1608
rect 2610 -1620 2616 -1614
rect 2610 -1626 2616 -1620
rect 2610 -1632 2616 -1626
rect 2610 -1638 2616 -1632
rect 2610 -1644 2616 -1638
rect 2610 -1650 2616 -1644
rect 2610 -1656 2616 -1650
rect 2610 -1662 2616 -1656
rect 2610 -1668 2616 -1662
rect 2610 -1674 2616 -1668
rect 2610 -1680 2616 -1674
rect 2610 -1686 2616 -1680
rect 2610 -1692 2616 -1686
rect 2610 -1698 2616 -1692
rect 2610 -1704 2616 -1698
rect 2610 -1710 2616 -1704
rect 2610 -1716 2616 -1710
rect 2610 -1722 2616 -1716
rect 2610 -1728 2616 -1722
rect 2610 -1734 2616 -1728
rect 2610 -1740 2616 -1734
rect 2610 -1746 2616 -1740
rect 2610 -1752 2616 -1746
rect 2610 -1758 2616 -1752
rect 2610 -1764 2616 -1758
rect 2610 -1770 2616 -1764
rect 2610 -1776 2616 -1770
rect 2610 -1782 2616 -1776
rect 2610 -1788 2616 -1782
rect 2610 -1794 2616 -1788
rect 2610 -1800 2616 -1794
rect 2610 -1806 2616 -1800
rect 2610 -1812 2616 -1806
rect 2610 -1818 2616 -1812
rect 2610 -1824 2616 -1818
rect 2610 -1830 2616 -1824
rect 2610 -1836 2616 -1830
rect 2610 -2418 2616 -2412
rect 2610 -2424 2616 -2418
rect 2610 -2430 2616 -2424
rect 2610 -2436 2616 -2430
rect 2610 -2442 2616 -2436
rect 2610 -2448 2616 -2442
rect 2610 -2454 2616 -2448
rect 2610 -2460 2616 -2454
rect 2610 -2466 2616 -2460
rect 2610 -2472 2616 -2466
rect 2610 -2478 2616 -2472
rect 2610 -2484 2616 -2478
rect 2610 -2490 2616 -2484
rect 2610 -2496 2616 -2490
rect 2610 -2502 2616 -2496
rect 2610 -2508 2616 -2502
rect 2610 -2514 2616 -2508
rect 2610 -2520 2616 -2514
rect 2610 -2526 2616 -2520
rect 2610 -2532 2616 -2526
rect 2610 -2538 2616 -2532
rect 2610 -2544 2616 -2538
rect 2610 -2550 2616 -2544
rect 2610 -2556 2616 -2550
rect 2610 -2562 2616 -2556
rect 2610 -2568 2616 -2562
rect 2610 -2574 2616 -2568
rect 2610 -2580 2616 -2574
rect 2610 -2586 2616 -2580
rect 2610 -2592 2616 -2586
rect 2610 -2598 2616 -2592
rect 2610 -2604 2616 -2598
rect 2610 -2610 2616 -2604
rect 2610 -2616 2616 -2610
rect 2610 -2622 2616 -2616
rect 2610 -2628 2616 -2622
rect 2610 -2634 2616 -2628
rect 2610 -2640 2616 -2634
rect 2610 -2646 2616 -2640
rect 2610 -2652 2616 -2646
rect 2610 -2658 2616 -2652
rect 2610 -2664 2616 -2658
rect 2610 -2670 2616 -2664
rect 2610 -2676 2616 -2670
rect 2610 -2682 2616 -2676
rect 2610 -2688 2616 -2682
rect 2610 -2694 2616 -2688
rect 2610 -2700 2616 -2694
rect 2610 -2706 2616 -2700
rect 2610 -2712 2616 -2706
rect 2610 -2718 2616 -2712
rect 2610 -2724 2616 -2718
rect 2610 -2730 2616 -2724
rect 2610 -2736 2616 -2730
rect 2610 -2742 2616 -2736
rect 2610 -2748 2616 -2742
rect 2610 -2754 2616 -2748
rect 2616 -1224 2622 -1218
rect 2616 -1230 2622 -1224
rect 2616 -1236 2622 -1230
rect 2616 -1242 2622 -1236
rect 2616 -1248 2622 -1242
rect 2616 -1254 2622 -1248
rect 2616 -1260 2622 -1254
rect 2616 -1266 2622 -1260
rect 2616 -1272 2622 -1266
rect 2616 -1278 2622 -1272
rect 2616 -1284 2622 -1278
rect 2616 -1290 2622 -1284
rect 2616 -1296 2622 -1290
rect 2616 -1302 2622 -1296
rect 2616 -1308 2622 -1302
rect 2616 -1314 2622 -1308
rect 2616 -1320 2622 -1314
rect 2616 -1326 2622 -1320
rect 2616 -1332 2622 -1326
rect 2616 -1338 2622 -1332
rect 2616 -1344 2622 -1338
rect 2616 -1350 2622 -1344
rect 2616 -1356 2622 -1350
rect 2616 -1362 2622 -1356
rect 2616 -1368 2622 -1362
rect 2616 -1374 2622 -1368
rect 2616 -1380 2622 -1374
rect 2616 -1386 2622 -1380
rect 2616 -1392 2622 -1386
rect 2616 -1398 2622 -1392
rect 2616 -1404 2622 -1398
rect 2616 -1410 2622 -1404
rect 2616 -1416 2622 -1410
rect 2616 -1422 2622 -1416
rect 2616 -1428 2622 -1422
rect 2616 -1434 2622 -1428
rect 2616 -1440 2622 -1434
rect 2616 -1446 2622 -1440
rect 2616 -1452 2622 -1446
rect 2616 -1458 2622 -1452
rect 2616 -1464 2622 -1458
rect 2616 -1470 2622 -1464
rect 2616 -1476 2622 -1470
rect 2616 -1482 2622 -1476
rect 2616 -1488 2622 -1482
rect 2616 -1494 2622 -1488
rect 2616 -1500 2622 -1494
rect 2616 -1506 2622 -1500
rect 2616 -1512 2622 -1506
rect 2616 -1518 2622 -1512
rect 2616 -1524 2622 -1518
rect 2616 -1530 2622 -1524
rect 2616 -1536 2622 -1530
rect 2616 -1542 2622 -1536
rect 2616 -1548 2622 -1542
rect 2616 -1554 2622 -1548
rect 2616 -1560 2622 -1554
rect 2616 -1566 2622 -1560
rect 2616 -1572 2622 -1566
rect 2616 -1578 2622 -1572
rect 2616 -1584 2622 -1578
rect 2616 -1590 2622 -1584
rect 2616 -1596 2622 -1590
rect 2616 -1602 2622 -1596
rect 2616 -1608 2622 -1602
rect 2616 -1614 2622 -1608
rect 2616 -1620 2622 -1614
rect 2616 -1626 2622 -1620
rect 2616 -1632 2622 -1626
rect 2616 -1638 2622 -1632
rect 2616 -1644 2622 -1638
rect 2616 -1650 2622 -1644
rect 2616 -1656 2622 -1650
rect 2616 -1662 2622 -1656
rect 2616 -1668 2622 -1662
rect 2616 -1674 2622 -1668
rect 2616 -1680 2622 -1674
rect 2616 -1686 2622 -1680
rect 2616 -1692 2622 -1686
rect 2616 -1698 2622 -1692
rect 2616 -1704 2622 -1698
rect 2616 -1710 2622 -1704
rect 2616 -1716 2622 -1710
rect 2616 -1722 2622 -1716
rect 2616 -1728 2622 -1722
rect 2616 -1734 2622 -1728
rect 2616 -1740 2622 -1734
rect 2616 -1746 2622 -1740
rect 2616 -1752 2622 -1746
rect 2616 -1758 2622 -1752
rect 2616 -1764 2622 -1758
rect 2616 -1770 2622 -1764
rect 2616 -1776 2622 -1770
rect 2616 -1782 2622 -1776
rect 2616 -1788 2622 -1782
rect 2616 -1794 2622 -1788
rect 2616 -1800 2622 -1794
rect 2616 -1806 2622 -1800
rect 2616 -1812 2622 -1806
rect 2616 -1818 2622 -1812
rect 2616 -1824 2622 -1818
rect 2616 -1830 2622 -1824
rect 2616 -2418 2622 -2412
rect 2616 -2424 2622 -2418
rect 2616 -2430 2622 -2424
rect 2616 -2436 2622 -2430
rect 2616 -2442 2622 -2436
rect 2616 -2448 2622 -2442
rect 2616 -2454 2622 -2448
rect 2616 -2460 2622 -2454
rect 2616 -2466 2622 -2460
rect 2616 -2472 2622 -2466
rect 2616 -2478 2622 -2472
rect 2616 -2484 2622 -2478
rect 2616 -2490 2622 -2484
rect 2616 -2496 2622 -2490
rect 2616 -2502 2622 -2496
rect 2616 -2508 2622 -2502
rect 2616 -2514 2622 -2508
rect 2616 -2520 2622 -2514
rect 2616 -2526 2622 -2520
rect 2616 -2532 2622 -2526
rect 2616 -2538 2622 -2532
rect 2616 -2544 2622 -2538
rect 2616 -2550 2622 -2544
rect 2616 -2556 2622 -2550
rect 2616 -2562 2622 -2556
rect 2616 -2568 2622 -2562
rect 2616 -2574 2622 -2568
rect 2616 -2580 2622 -2574
rect 2616 -2586 2622 -2580
rect 2616 -2592 2622 -2586
rect 2616 -2598 2622 -2592
rect 2616 -2604 2622 -2598
rect 2616 -2610 2622 -2604
rect 2616 -2616 2622 -2610
rect 2616 -2622 2622 -2616
rect 2616 -2628 2622 -2622
rect 2616 -2634 2622 -2628
rect 2616 -2640 2622 -2634
rect 2616 -2646 2622 -2640
rect 2616 -2652 2622 -2646
rect 2616 -2658 2622 -2652
rect 2616 -2664 2622 -2658
rect 2616 -2670 2622 -2664
rect 2616 -2676 2622 -2670
rect 2616 -2682 2622 -2676
rect 2616 -2688 2622 -2682
rect 2616 -2694 2622 -2688
rect 2616 -2700 2622 -2694
rect 2616 -2706 2622 -2700
rect 2616 -2712 2622 -2706
rect 2616 -2718 2622 -2712
rect 2616 -2724 2622 -2718
rect 2616 -2730 2622 -2724
rect 2616 -2736 2622 -2730
rect 2616 -2742 2622 -2736
rect 2616 -2748 2622 -2742
rect 2616 -2754 2622 -2748
rect 2622 -1218 2628 -1212
rect 2622 -1224 2628 -1218
rect 2622 -1230 2628 -1224
rect 2622 -1236 2628 -1230
rect 2622 -1242 2628 -1236
rect 2622 -1248 2628 -1242
rect 2622 -1254 2628 -1248
rect 2622 -1260 2628 -1254
rect 2622 -1266 2628 -1260
rect 2622 -1272 2628 -1266
rect 2622 -1278 2628 -1272
rect 2622 -1284 2628 -1278
rect 2622 -1290 2628 -1284
rect 2622 -1296 2628 -1290
rect 2622 -1302 2628 -1296
rect 2622 -1308 2628 -1302
rect 2622 -1314 2628 -1308
rect 2622 -1320 2628 -1314
rect 2622 -1326 2628 -1320
rect 2622 -1332 2628 -1326
rect 2622 -1338 2628 -1332
rect 2622 -1344 2628 -1338
rect 2622 -1350 2628 -1344
rect 2622 -1356 2628 -1350
rect 2622 -1362 2628 -1356
rect 2622 -1368 2628 -1362
rect 2622 -1374 2628 -1368
rect 2622 -1380 2628 -1374
rect 2622 -1386 2628 -1380
rect 2622 -1392 2628 -1386
rect 2622 -1398 2628 -1392
rect 2622 -1404 2628 -1398
rect 2622 -1410 2628 -1404
rect 2622 -1416 2628 -1410
rect 2622 -1422 2628 -1416
rect 2622 -1428 2628 -1422
rect 2622 -1434 2628 -1428
rect 2622 -1440 2628 -1434
rect 2622 -1446 2628 -1440
rect 2622 -1452 2628 -1446
rect 2622 -1458 2628 -1452
rect 2622 -1464 2628 -1458
rect 2622 -1470 2628 -1464
rect 2622 -1476 2628 -1470
rect 2622 -1482 2628 -1476
rect 2622 -1488 2628 -1482
rect 2622 -1494 2628 -1488
rect 2622 -1500 2628 -1494
rect 2622 -1506 2628 -1500
rect 2622 -1512 2628 -1506
rect 2622 -1518 2628 -1512
rect 2622 -1524 2628 -1518
rect 2622 -1530 2628 -1524
rect 2622 -1536 2628 -1530
rect 2622 -1542 2628 -1536
rect 2622 -1548 2628 -1542
rect 2622 -1554 2628 -1548
rect 2622 -1560 2628 -1554
rect 2622 -1566 2628 -1560
rect 2622 -1572 2628 -1566
rect 2622 -1578 2628 -1572
rect 2622 -1584 2628 -1578
rect 2622 -1590 2628 -1584
rect 2622 -1596 2628 -1590
rect 2622 -1602 2628 -1596
rect 2622 -1608 2628 -1602
rect 2622 -1614 2628 -1608
rect 2622 -1620 2628 -1614
rect 2622 -1626 2628 -1620
rect 2622 -1632 2628 -1626
rect 2622 -1638 2628 -1632
rect 2622 -1644 2628 -1638
rect 2622 -1650 2628 -1644
rect 2622 -1656 2628 -1650
rect 2622 -1662 2628 -1656
rect 2622 -1668 2628 -1662
rect 2622 -1674 2628 -1668
rect 2622 -1680 2628 -1674
rect 2622 -1686 2628 -1680
rect 2622 -1692 2628 -1686
rect 2622 -1698 2628 -1692
rect 2622 -1704 2628 -1698
rect 2622 -1710 2628 -1704
rect 2622 -1716 2628 -1710
rect 2622 -1722 2628 -1716
rect 2622 -1728 2628 -1722
rect 2622 -1734 2628 -1728
rect 2622 -1740 2628 -1734
rect 2622 -1746 2628 -1740
rect 2622 -1752 2628 -1746
rect 2622 -1758 2628 -1752
rect 2622 -1764 2628 -1758
rect 2622 -1770 2628 -1764
rect 2622 -1776 2628 -1770
rect 2622 -1782 2628 -1776
rect 2622 -1788 2628 -1782
rect 2622 -1794 2628 -1788
rect 2622 -1800 2628 -1794
rect 2622 -1806 2628 -1800
rect 2622 -1812 2628 -1806
rect 2622 -1818 2628 -1812
rect 2622 -1824 2628 -1818
rect 2622 -2418 2628 -2412
rect 2622 -2424 2628 -2418
rect 2622 -2430 2628 -2424
rect 2622 -2436 2628 -2430
rect 2622 -2442 2628 -2436
rect 2622 -2448 2628 -2442
rect 2622 -2454 2628 -2448
rect 2622 -2460 2628 -2454
rect 2622 -2466 2628 -2460
rect 2622 -2472 2628 -2466
rect 2622 -2478 2628 -2472
rect 2622 -2484 2628 -2478
rect 2622 -2490 2628 -2484
rect 2622 -2496 2628 -2490
rect 2622 -2502 2628 -2496
rect 2622 -2508 2628 -2502
rect 2622 -2514 2628 -2508
rect 2622 -2520 2628 -2514
rect 2622 -2526 2628 -2520
rect 2622 -2532 2628 -2526
rect 2622 -2538 2628 -2532
rect 2622 -2544 2628 -2538
rect 2622 -2550 2628 -2544
rect 2622 -2556 2628 -2550
rect 2622 -2562 2628 -2556
rect 2622 -2568 2628 -2562
rect 2622 -2574 2628 -2568
rect 2622 -2580 2628 -2574
rect 2622 -2586 2628 -2580
rect 2622 -2592 2628 -2586
rect 2622 -2598 2628 -2592
rect 2622 -2604 2628 -2598
rect 2622 -2610 2628 -2604
rect 2622 -2616 2628 -2610
rect 2622 -2622 2628 -2616
rect 2622 -2628 2628 -2622
rect 2622 -2634 2628 -2628
rect 2622 -2640 2628 -2634
rect 2622 -2646 2628 -2640
rect 2622 -2652 2628 -2646
rect 2622 -2658 2628 -2652
rect 2622 -2664 2628 -2658
rect 2622 -2670 2628 -2664
rect 2622 -2676 2628 -2670
rect 2622 -2682 2628 -2676
rect 2622 -2688 2628 -2682
rect 2622 -2694 2628 -2688
rect 2622 -2700 2628 -2694
rect 2622 -2706 2628 -2700
rect 2622 -2712 2628 -2706
rect 2622 -2718 2628 -2712
rect 2622 -2724 2628 -2718
rect 2622 -2730 2628 -2724
rect 2622 -2736 2628 -2730
rect 2622 -2742 2628 -2736
rect 2622 -2748 2628 -2742
rect 2628 -1212 2634 -1206
rect 2628 -1218 2634 -1212
rect 2628 -1224 2634 -1218
rect 2628 -1230 2634 -1224
rect 2628 -1236 2634 -1230
rect 2628 -1242 2634 -1236
rect 2628 -1248 2634 -1242
rect 2628 -1254 2634 -1248
rect 2628 -1260 2634 -1254
rect 2628 -1266 2634 -1260
rect 2628 -1272 2634 -1266
rect 2628 -1278 2634 -1272
rect 2628 -1284 2634 -1278
rect 2628 -1290 2634 -1284
rect 2628 -1296 2634 -1290
rect 2628 -1302 2634 -1296
rect 2628 -1308 2634 -1302
rect 2628 -1314 2634 -1308
rect 2628 -1320 2634 -1314
rect 2628 -1326 2634 -1320
rect 2628 -1332 2634 -1326
rect 2628 -1338 2634 -1332
rect 2628 -1344 2634 -1338
rect 2628 -1350 2634 -1344
rect 2628 -1356 2634 -1350
rect 2628 -1362 2634 -1356
rect 2628 -1368 2634 -1362
rect 2628 -1374 2634 -1368
rect 2628 -1380 2634 -1374
rect 2628 -1386 2634 -1380
rect 2628 -1392 2634 -1386
rect 2628 -1398 2634 -1392
rect 2628 -1404 2634 -1398
rect 2628 -1410 2634 -1404
rect 2628 -1416 2634 -1410
rect 2628 -1422 2634 -1416
rect 2628 -1428 2634 -1422
rect 2628 -1434 2634 -1428
rect 2628 -1440 2634 -1434
rect 2628 -1446 2634 -1440
rect 2628 -1452 2634 -1446
rect 2628 -1458 2634 -1452
rect 2628 -1464 2634 -1458
rect 2628 -1470 2634 -1464
rect 2628 -1476 2634 -1470
rect 2628 -1482 2634 -1476
rect 2628 -1488 2634 -1482
rect 2628 -1494 2634 -1488
rect 2628 -1500 2634 -1494
rect 2628 -1506 2634 -1500
rect 2628 -1512 2634 -1506
rect 2628 -1518 2634 -1512
rect 2628 -1524 2634 -1518
rect 2628 -1530 2634 -1524
rect 2628 -1536 2634 -1530
rect 2628 -1542 2634 -1536
rect 2628 -1548 2634 -1542
rect 2628 -1554 2634 -1548
rect 2628 -1560 2634 -1554
rect 2628 -1566 2634 -1560
rect 2628 -1572 2634 -1566
rect 2628 -1578 2634 -1572
rect 2628 -1584 2634 -1578
rect 2628 -1590 2634 -1584
rect 2628 -1596 2634 -1590
rect 2628 -1602 2634 -1596
rect 2628 -1608 2634 -1602
rect 2628 -1614 2634 -1608
rect 2628 -1620 2634 -1614
rect 2628 -1626 2634 -1620
rect 2628 -1632 2634 -1626
rect 2628 -1638 2634 -1632
rect 2628 -1644 2634 -1638
rect 2628 -1650 2634 -1644
rect 2628 -1656 2634 -1650
rect 2628 -1662 2634 -1656
rect 2628 -1668 2634 -1662
rect 2628 -1674 2634 -1668
rect 2628 -1680 2634 -1674
rect 2628 -1686 2634 -1680
rect 2628 -1692 2634 -1686
rect 2628 -1698 2634 -1692
rect 2628 -1704 2634 -1698
rect 2628 -1710 2634 -1704
rect 2628 -1716 2634 -1710
rect 2628 -1722 2634 -1716
rect 2628 -1728 2634 -1722
rect 2628 -1734 2634 -1728
rect 2628 -1740 2634 -1734
rect 2628 -1746 2634 -1740
rect 2628 -1752 2634 -1746
rect 2628 -1758 2634 -1752
rect 2628 -1764 2634 -1758
rect 2628 -1770 2634 -1764
rect 2628 -1776 2634 -1770
rect 2628 -1782 2634 -1776
rect 2628 -1788 2634 -1782
rect 2628 -1794 2634 -1788
rect 2628 -1800 2634 -1794
rect 2628 -1806 2634 -1800
rect 2628 -1812 2634 -1806
rect 2628 -1818 2634 -1812
rect 2628 -2418 2634 -2412
rect 2628 -2424 2634 -2418
rect 2628 -2430 2634 -2424
rect 2628 -2436 2634 -2430
rect 2628 -2442 2634 -2436
rect 2628 -2448 2634 -2442
rect 2628 -2454 2634 -2448
rect 2628 -2460 2634 -2454
rect 2628 -2466 2634 -2460
rect 2628 -2472 2634 -2466
rect 2628 -2478 2634 -2472
rect 2628 -2484 2634 -2478
rect 2628 -2490 2634 -2484
rect 2628 -2496 2634 -2490
rect 2628 -2502 2634 -2496
rect 2628 -2508 2634 -2502
rect 2628 -2514 2634 -2508
rect 2628 -2520 2634 -2514
rect 2628 -2526 2634 -2520
rect 2628 -2532 2634 -2526
rect 2628 -2538 2634 -2532
rect 2628 -2544 2634 -2538
rect 2628 -2550 2634 -2544
rect 2628 -2556 2634 -2550
rect 2628 -2562 2634 -2556
rect 2628 -2568 2634 -2562
rect 2628 -2574 2634 -2568
rect 2628 -2580 2634 -2574
rect 2628 -2586 2634 -2580
rect 2628 -2592 2634 -2586
rect 2628 -2598 2634 -2592
rect 2628 -2604 2634 -2598
rect 2628 -2610 2634 -2604
rect 2628 -2616 2634 -2610
rect 2628 -2622 2634 -2616
rect 2628 -2628 2634 -2622
rect 2628 -2634 2634 -2628
rect 2628 -2640 2634 -2634
rect 2628 -2646 2634 -2640
rect 2628 -2652 2634 -2646
rect 2628 -2658 2634 -2652
rect 2628 -2664 2634 -2658
rect 2628 -2670 2634 -2664
rect 2628 -2676 2634 -2670
rect 2628 -2682 2634 -2676
rect 2628 -2688 2634 -2682
rect 2628 -2694 2634 -2688
rect 2628 -2700 2634 -2694
rect 2628 -2706 2634 -2700
rect 2628 -2712 2634 -2706
rect 2628 -2718 2634 -2712
rect 2628 -2724 2634 -2718
rect 2628 -2730 2634 -2724
rect 2628 -2736 2634 -2730
rect 2628 -2742 2634 -2736
rect 2628 -2748 2634 -2742
rect 2634 -1212 2640 -1206
rect 2634 -1218 2640 -1212
rect 2634 -1224 2640 -1218
rect 2634 -1230 2640 -1224
rect 2634 -1236 2640 -1230
rect 2634 -1242 2640 -1236
rect 2634 -1248 2640 -1242
rect 2634 -1254 2640 -1248
rect 2634 -1260 2640 -1254
rect 2634 -1266 2640 -1260
rect 2634 -1272 2640 -1266
rect 2634 -1278 2640 -1272
rect 2634 -1284 2640 -1278
rect 2634 -1290 2640 -1284
rect 2634 -1296 2640 -1290
rect 2634 -1302 2640 -1296
rect 2634 -1308 2640 -1302
rect 2634 -1314 2640 -1308
rect 2634 -1320 2640 -1314
rect 2634 -1326 2640 -1320
rect 2634 -1332 2640 -1326
rect 2634 -1338 2640 -1332
rect 2634 -1344 2640 -1338
rect 2634 -1350 2640 -1344
rect 2634 -1356 2640 -1350
rect 2634 -1362 2640 -1356
rect 2634 -1368 2640 -1362
rect 2634 -1374 2640 -1368
rect 2634 -1380 2640 -1374
rect 2634 -1386 2640 -1380
rect 2634 -1392 2640 -1386
rect 2634 -1398 2640 -1392
rect 2634 -1404 2640 -1398
rect 2634 -1410 2640 -1404
rect 2634 -1416 2640 -1410
rect 2634 -1422 2640 -1416
rect 2634 -1428 2640 -1422
rect 2634 -1434 2640 -1428
rect 2634 -1440 2640 -1434
rect 2634 -1446 2640 -1440
rect 2634 -1452 2640 -1446
rect 2634 -1458 2640 -1452
rect 2634 -1464 2640 -1458
rect 2634 -1470 2640 -1464
rect 2634 -1476 2640 -1470
rect 2634 -1482 2640 -1476
rect 2634 -1488 2640 -1482
rect 2634 -1494 2640 -1488
rect 2634 -1500 2640 -1494
rect 2634 -1506 2640 -1500
rect 2634 -1512 2640 -1506
rect 2634 -1518 2640 -1512
rect 2634 -1524 2640 -1518
rect 2634 -1530 2640 -1524
rect 2634 -1536 2640 -1530
rect 2634 -1542 2640 -1536
rect 2634 -1548 2640 -1542
rect 2634 -1554 2640 -1548
rect 2634 -1560 2640 -1554
rect 2634 -1566 2640 -1560
rect 2634 -1572 2640 -1566
rect 2634 -1578 2640 -1572
rect 2634 -1584 2640 -1578
rect 2634 -1590 2640 -1584
rect 2634 -1596 2640 -1590
rect 2634 -1602 2640 -1596
rect 2634 -1608 2640 -1602
rect 2634 -1614 2640 -1608
rect 2634 -1620 2640 -1614
rect 2634 -1626 2640 -1620
rect 2634 -1632 2640 -1626
rect 2634 -1638 2640 -1632
rect 2634 -1644 2640 -1638
rect 2634 -1650 2640 -1644
rect 2634 -1656 2640 -1650
rect 2634 -1662 2640 -1656
rect 2634 -1668 2640 -1662
rect 2634 -1674 2640 -1668
rect 2634 -1680 2640 -1674
rect 2634 -1686 2640 -1680
rect 2634 -1692 2640 -1686
rect 2634 -1698 2640 -1692
rect 2634 -1704 2640 -1698
rect 2634 -1710 2640 -1704
rect 2634 -1716 2640 -1710
rect 2634 -1722 2640 -1716
rect 2634 -1728 2640 -1722
rect 2634 -1734 2640 -1728
rect 2634 -1740 2640 -1734
rect 2634 -1746 2640 -1740
rect 2634 -1752 2640 -1746
rect 2634 -1758 2640 -1752
rect 2634 -1764 2640 -1758
rect 2634 -1770 2640 -1764
rect 2634 -1776 2640 -1770
rect 2634 -1782 2640 -1776
rect 2634 -1788 2640 -1782
rect 2634 -1794 2640 -1788
rect 2634 -1800 2640 -1794
rect 2634 -1806 2640 -1800
rect 2634 -2412 2640 -2406
rect 2634 -2418 2640 -2412
rect 2634 -2424 2640 -2418
rect 2634 -2430 2640 -2424
rect 2634 -2436 2640 -2430
rect 2634 -2442 2640 -2436
rect 2634 -2448 2640 -2442
rect 2634 -2454 2640 -2448
rect 2634 -2460 2640 -2454
rect 2634 -2466 2640 -2460
rect 2634 -2472 2640 -2466
rect 2634 -2478 2640 -2472
rect 2634 -2484 2640 -2478
rect 2634 -2490 2640 -2484
rect 2634 -2496 2640 -2490
rect 2634 -2502 2640 -2496
rect 2634 -2508 2640 -2502
rect 2634 -2514 2640 -2508
rect 2634 -2520 2640 -2514
rect 2634 -2526 2640 -2520
rect 2634 -2532 2640 -2526
rect 2634 -2538 2640 -2532
rect 2634 -2544 2640 -2538
rect 2634 -2550 2640 -2544
rect 2634 -2556 2640 -2550
rect 2634 -2562 2640 -2556
rect 2634 -2568 2640 -2562
rect 2634 -2574 2640 -2568
rect 2634 -2580 2640 -2574
rect 2634 -2586 2640 -2580
rect 2634 -2592 2640 -2586
rect 2634 -2598 2640 -2592
rect 2634 -2604 2640 -2598
rect 2634 -2610 2640 -2604
rect 2634 -2616 2640 -2610
rect 2634 -2622 2640 -2616
rect 2634 -2628 2640 -2622
rect 2634 -2634 2640 -2628
rect 2634 -2640 2640 -2634
rect 2634 -2646 2640 -2640
rect 2634 -2652 2640 -2646
rect 2634 -2658 2640 -2652
rect 2634 -2664 2640 -2658
rect 2634 -2670 2640 -2664
rect 2634 -2676 2640 -2670
rect 2634 -2682 2640 -2676
rect 2634 -2688 2640 -2682
rect 2634 -2694 2640 -2688
rect 2634 -2700 2640 -2694
rect 2634 -2706 2640 -2700
rect 2634 -2712 2640 -2706
rect 2634 -2718 2640 -2712
rect 2634 -2724 2640 -2718
rect 2634 -2730 2640 -2724
rect 2634 -2736 2640 -2730
rect 2634 -2742 2640 -2736
rect 2640 -1206 2646 -1200
rect 2640 -1212 2646 -1206
rect 2640 -1218 2646 -1212
rect 2640 -1224 2646 -1218
rect 2640 -1230 2646 -1224
rect 2640 -1236 2646 -1230
rect 2640 -1242 2646 -1236
rect 2640 -1248 2646 -1242
rect 2640 -1254 2646 -1248
rect 2640 -1260 2646 -1254
rect 2640 -1266 2646 -1260
rect 2640 -1272 2646 -1266
rect 2640 -1278 2646 -1272
rect 2640 -1284 2646 -1278
rect 2640 -1290 2646 -1284
rect 2640 -1296 2646 -1290
rect 2640 -1302 2646 -1296
rect 2640 -1308 2646 -1302
rect 2640 -1314 2646 -1308
rect 2640 -1320 2646 -1314
rect 2640 -1326 2646 -1320
rect 2640 -1332 2646 -1326
rect 2640 -1338 2646 -1332
rect 2640 -1344 2646 -1338
rect 2640 -1350 2646 -1344
rect 2640 -1356 2646 -1350
rect 2640 -1362 2646 -1356
rect 2640 -1368 2646 -1362
rect 2640 -1374 2646 -1368
rect 2640 -1380 2646 -1374
rect 2640 -1386 2646 -1380
rect 2640 -1392 2646 -1386
rect 2640 -1398 2646 -1392
rect 2640 -1404 2646 -1398
rect 2640 -1410 2646 -1404
rect 2640 -1416 2646 -1410
rect 2640 -1422 2646 -1416
rect 2640 -1428 2646 -1422
rect 2640 -1434 2646 -1428
rect 2640 -1440 2646 -1434
rect 2640 -1446 2646 -1440
rect 2640 -1452 2646 -1446
rect 2640 -1458 2646 -1452
rect 2640 -1464 2646 -1458
rect 2640 -1470 2646 -1464
rect 2640 -1476 2646 -1470
rect 2640 -1482 2646 -1476
rect 2640 -1488 2646 -1482
rect 2640 -1494 2646 -1488
rect 2640 -1500 2646 -1494
rect 2640 -1506 2646 -1500
rect 2640 -1512 2646 -1506
rect 2640 -1518 2646 -1512
rect 2640 -1524 2646 -1518
rect 2640 -1530 2646 -1524
rect 2640 -1536 2646 -1530
rect 2640 -1542 2646 -1536
rect 2640 -1548 2646 -1542
rect 2640 -1554 2646 -1548
rect 2640 -1560 2646 -1554
rect 2640 -1566 2646 -1560
rect 2640 -1572 2646 -1566
rect 2640 -1578 2646 -1572
rect 2640 -1584 2646 -1578
rect 2640 -1590 2646 -1584
rect 2640 -1596 2646 -1590
rect 2640 -1602 2646 -1596
rect 2640 -1608 2646 -1602
rect 2640 -1614 2646 -1608
rect 2640 -1620 2646 -1614
rect 2640 -1626 2646 -1620
rect 2640 -1632 2646 -1626
rect 2640 -1638 2646 -1632
rect 2640 -1644 2646 -1638
rect 2640 -1650 2646 -1644
rect 2640 -1656 2646 -1650
rect 2640 -1662 2646 -1656
rect 2640 -1668 2646 -1662
rect 2640 -1674 2646 -1668
rect 2640 -1680 2646 -1674
rect 2640 -1686 2646 -1680
rect 2640 -1692 2646 -1686
rect 2640 -1698 2646 -1692
rect 2640 -1704 2646 -1698
rect 2640 -1710 2646 -1704
rect 2640 -1716 2646 -1710
rect 2640 -1722 2646 -1716
rect 2640 -1728 2646 -1722
rect 2640 -1734 2646 -1728
rect 2640 -1740 2646 -1734
rect 2640 -1746 2646 -1740
rect 2640 -1752 2646 -1746
rect 2640 -1758 2646 -1752
rect 2640 -1764 2646 -1758
rect 2640 -1770 2646 -1764
rect 2640 -1776 2646 -1770
rect 2640 -1782 2646 -1776
rect 2640 -1788 2646 -1782
rect 2640 -1794 2646 -1788
rect 2640 -1800 2646 -1794
rect 2640 -2412 2646 -2406
rect 2640 -2418 2646 -2412
rect 2640 -2424 2646 -2418
rect 2640 -2430 2646 -2424
rect 2640 -2436 2646 -2430
rect 2640 -2442 2646 -2436
rect 2640 -2448 2646 -2442
rect 2640 -2454 2646 -2448
rect 2640 -2460 2646 -2454
rect 2640 -2466 2646 -2460
rect 2640 -2472 2646 -2466
rect 2640 -2478 2646 -2472
rect 2640 -2484 2646 -2478
rect 2640 -2490 2646 -2484
rect 2640 -2496 2646 -2490
rect 2640 -2502 2646 -2496
rect 2640 -2508 2646 -2502
rect 2640 -2514 2646 -2508
rect 2640 -2520 2646 -2514
rect 2640 -2526 2646 -2520
rect 2640 -2532 2646 -2526
rect 2640 -2538 2646 -2532
rect 2640 -2544 2646 -2538
rect 2640 -2550 2646 -2544
rect 2640 -2556 2646 -2550
rect 2640 -2562 2646 -2556
rect 2640 -2568 2646 -2562
rect 2640 -2574 2646 -2568
rect 2640 -2580 2646 -2574
rect 2640 -2586 2646 -2580
rect 2640 -2592 2646 -2586
rect 2640 -2598 2646 -2592
rect 2640 -2604 2646 -2598
rect 2640 -2610 2646 -2604
rect 2640 -2616 2646 -2610
rect 2640 -2622 2646 -2616
rect 2640 -2628 2646 -2622
rect 2640 -2634 2646 -2628
rect 2640 -2640 2646 -2634
rect 2640 -2646 2646 -2640
rect 2640 -2652 2646 -2646
rect 2640 -2658 2646 -2652
rect 2640 -2664 2646 -2658
rect 2640 -2670 2646 -2664
rect 2640 -2676 2646 -2670
rect 2640 -2682 2646 -2676
rect 2640 -2688 2646 -2682
rect 2640 -2694 2646 -2688
rect 2640 -2700 2646 -2694
rect 2640 -2706 2646 -2700
rect 2640 -2712 2646 -2706
rect 2640 -2718 2646 -2712
rect 2640 -2724 2646 -2718
rect 2640 -2730 2646 -2724
rect 2640 -2736 2646 -2730
rect 2646 -1200 2652 -1194
rect 2646 -1206 2652 -1200
rect 2646 -1212 2652 -1206
rect 2646 -1218 2652 -1212
rect 2646 -1224 2652 -1218
rect 2646 -1230 2652 -1224
rect 2646 -1236 2652 -1230
rect 2646 -1242 2652 -1236
rect 2646 -1248 2652 -1242
rect 2646 -1254 2652 -1248
rect 2646 -1260 2652 -1254
rect 2646 -1266 2652 -1260
rect 2646 -1272 2652 -1266
rect 2646 -1278 2652 -1272
rect 2646 -1284 2652 -1278
rect 2646 -1290 2652 -1284
rect 2646 -1296 2652 -1290
rect 2646 -1302 2652 -1296
rect 2646 -1308 2652 -1302
rect 2646 -1314 2652 -1308
rect 2646 -1320 2652 -1314
rect 2646 -1326 2652 -1320
rect 2646 -1332 2652 -1326
rect 2646 -1338 2652 -1332
rect 2646 -1344 2652 -1338
rect 2646 -1350 2652 -1344
rect 2646 -1356 2652 -1350
rect 2646 -1362 2652 -1356
rect 2646 -1368 2652 -1362
rect 2646 -1374 2652 -1368
rect 2646 -1380 2652 -1374
rect 2646 -1386 2652 -1380
rect 2646 -1392 2652 -1386
rect 2646 -1398 2652 -1392
rect 2646 -1404 2652 -1398
rect 2646 -1410 2652 -1404
rect 2646 -1416 2652 -1410
rect 2646 -1422 2652 -1416
rect 2646 -1428 2652 -1422
rect 2646 -1434 2652 -1428
rect 2646 -1440 2652 -1434
rect 2646 -1446 2652 -1440
rect 2646 -1452 2652 -1446
rect 2646 -1458 2652 -1452
rect 2646 -1464 2652 -1458
rect 2646 -1470 2652 -1464
rect 2646 -1476 2652 -1470
rect 2646 -1482 2652 -1476
rect 2646 -1488 2652 -1482
rect 2646 -1494 2652 -1488
rect 2646 -1500 2652 -1494
rect 2646 -1506 2652 -1500
rect 2646 -1512 2652 -1506
rect 2646 -1518 2652 -1512
rect 2646 -1524 2652 -1518
rect 2646 -1530 2652 -1524
rect 2646 -1536 2652 -1530
rect 2646 -1542 2652 -1536
rect 2646 -1548 2652 -1542
rect 2646 -1554 2652 -1548
rect 2646 -1560 2652 -1554
rect 2646 -1566 2652 -1560
rect 2646 -1572 2652 -1566
rect 2646 -1578 2652 -1572
rect 2646 -1584 2652 -1578
rect 2646 -1590 2652 -1584
rect 2646 -1596 2652 -1590
rect 2646 -1602 2652 -1596
rect 2646 -1608 2652 -1602
rect 2646 -1614 2652 -1608
rect 2646 -1620 2652 -1614
rect 2646 -1626 2652 -1620
rect 2646 -1632 2652 -1626
rect 2646 -1638 2652 -1632
rect 2646 -1644 2652 -1638
rect 2646 -1650 2652 -1644
rect 2646 -1656 2652 -1650
rect 2646 -1662 2652 -1656
rect 2646 -1668 2652 -1662
rect 2646 -1674 2652 -1668
rect 2646 -1680 2652 -1674
rect 2646 -1686 2652 -1680
rect 2646 -1692 2652 -1686
rect 2646 -1698 2652 -1692
rect 2646 -1704 2652 -1698
rect 2646 -1710 2652 -1704
rect 2646 -1716 2652 -1710
rect 2646 -1722 2652 -1716
rect 2646 -1728 2652 -1722
rect 2646 -1734 2652 -1728
rect 2646 -1740 2652 -1734
rect 2646 -1746 2652 -1740
rect 2646 -1752 2652 -1746
rect 2646 -1758 2652 -1752
rect 2646 -1764 2652 -1758
rect 2646 -1770 2652 -1764
rect 2646 -1776 2652 -1770
rect 2646 -1782 2652 -1776
rect 2646 -1788 2652 -1782
rect 2646 -1794 2652 -1788
rect 2646 -2412 2652 -2406
rect 2646 -2418 2652 -2412
rect 2646 -2424 2652 -2418
rect 2646 -2430 2652 -2424
rect 2646 -2436 2652 -2430
rect 2646 -2442 2652 -2436
rect 2646 -2448 2652 -2442
rect 2646 -2454 2652 -2448
rect 2646 -2460 2652 -2454
rect 2646 -2466 2652 -2460
rect 2646 -2472 2652 -2466
rect 2646 -2478 2652 -2472
rect 2646 -2484 2652 -2478
rect 2646 -2490 2652 -2484
rect 2646 -2496 2652 -2490
rect 2646 -2502 2652 -2496
rect 2646 -2508 2652 -2502
rect 2646 -2514 2652 -2508
rect 2646 -2520 2652 -2514
rect 2646 -2526 2652 -2520
rect 2646 -2532 2652 -2526
rect 2646 -2538 2652 -2532
rect 2646 -2544 2652 -2538
rect 2646 -2550 2652 -2544
rect 2646 -2556 2652 -2550
rect 2646 -2562 2652 -2556
rect 2646 -2568 2652 -2562
rect 2646 -2574 2652 -2568
rect 2646 -2580 2652 -2574
rect 2646 -2586 2652 -2580
rect 2646 -2592 2652 -2586
rect 2646 -2598 2652 -2592
rect 2646 -2604 2652 -2598
rect 2646 -2610 2652 -2604
rect 2646 -2616 2652 -2610
rect 2646 -2622 2652 -2616
rect 2646 -2628 2652 -2622
rect 2646 -2634 2652 -2628
rect 2646 -2640 2652 -2634
rect 2646 -2646 2652 -2640
rect 2646 -2652 2652 -2646
rect 2646 -2658 2652 -2652
rect 2646 -2664 2652 -2658
rect 2646 -2670 2652 -2664
rect 2646 -2676 2652 -2670
rect 2646 -2682 2652 -2676
rect 2646 -2688 2652 -2682
rect 2646 -2694 2652 -2688
rect 2646 -2700 2652 -2694
rect 2646 -2706 2652 -2700
rect 2646 -2712 2652 -2706
rect 2646 -2718 2652 -2712
rect 2646 -2724 2652 -2718
rect 2646 -2730 2652 -2724
rect 2646 -2736 2652 -2730
rect 2652 -1194 2658 -1188
rect 2652 -1200 2658 -1194
rect 2652 -1206 2658 -1200
rect 2652 -1212 2658 -1206
rect 2652 -1218 2658 -1212
rect 2652 -1224 2658 -1218
rect 2652 -1230 2658 -1224
rect 2652 -1236 2658 -1230
rect 2652 -1242 2658 -1236
rect 2652 -1248 2658 -1242
rect 2652 -1254 2658 -1248
rect 2652 -1260 2658 -1254
rect 2652 -1266 2658 -1260
rect 2652 -1272 2658 -1266
rect 2652 -1278 2658 -1272
rect 2652 -1284 2658 -1278
rect 2652 -1290 2658 -1284
rect 2652 -1296 2658 -1290
rect 2652 -1302 2658 -1296
rect 2652 -1308 2658 -1302
rect 2652 -1314 2658 -1308
rect 2652 -1320 2658 -1314
rect 2652 -1326 2658 -1320
rect 2652 -1332 2658 -1326
rect 2652 -1338 2658 -1332
rect 2652 -1344 2658 -1338
rect 2652 -1350 2658 -1344
rect 2652 -1356 2658 -1350
rect 2652 -1362 2658 -1356
rect 2652 -1368 2658 -1362
rect 2652 -1374 2658 -1368
rect 2652 -1380 2658 -1374
rect 2652 -1386 2658 -1380
rect 2652 -1392 2658 -1386
rect 2652 -1398 2658 -1392
rect 2652 -1404 2658 -1398
rect 2652 -1410 2658 -1404
rect 2652 -1416 2658 -1410
rect 2652 -1422 2658 -1416
rect 2652 -1428 2658 -1422
rect 2652 -1434 2658 -1428
rect 2652 -1440 2658 -1434
rect 2652 -1446 2658 -1440
rect 2652 -1452 2658 -1446
rect 2652 -1458 2658 -1452
rect 2652 -1464 2658 -1458
rect 2652 -1470 2658 -1464
rect 2652 -1476 2658 -1470
rect 2652 -1482 2658 -1476
rect 2652 -1488 2658 -1482
rect 2652 -1494 2658 -1488
rect 2652 -1500 2658 -1494
rect 2652 -1506 2658 -1500
rect 2652 -1512 2658 -1506
rect 2652 -1518 2658 -1512
rect 2652 -1524 2658 -1518
rect 2652 -1530 2658 -1524
rect 2652 -1536 2658 -1530
rect 2652 -1542 2658 -1536
rect 2652 -1548 2658 -1542
rect 2652 -1554 2658 -1548
rect 2652 -1560 2658 -1554
rect 2652 -1566 2658 -1560
rect 2652 -1572 2658 -1566
rect 2652 -1578 2658 -1572
rect 2652 -1584 2658 -1578
rect 2652 -1590 2658 -1584
rect 2652 -1596 2658 -1590
rect 2652 -1602 2658 -1596
rect 2652 -1608 2658 -1602
rect 2652 -1614 2658 -1608
rect 2652 -1620 2658 -1614
rect 2652 -1626 2658 -1620
rect 2652 -1632 2658 -1626
rect 2652 -1638 2658 -1632
rect 2652 -1644 2658 -1638
rect 2652 -1650 2658 -1644
rect 2652 -1656 2658 -1650
rect 2652 -1662 2658 -1656
rect 2652 -1668 2658 -1662
rect 2652 -1674 2658 -1668
rect 2652 -1680 2658 -1674
rect 2652 -1686 2658 -1680
rect 2652 -1692 2658 -1686
rect 2652 -1698 2658 -1692
rect 2652 -1704 2658 -1698
rect 2652 -1710 2658 -1704
rect 2652 -1716 2658 -1710
rect 2652 -1722 2658 -1716
rect 2652 -1728 2658 -1722
rect 2652 -1734 2658 -1728
rect 2652 -1740 2658 -1734
rect 2652 -1746 2658 -1740
rect 2652 -1752 2658 -1746
rect 2652 -1758 2658 -1752
rect 2652 -1764 2658 -1758
rect 2652 -1770 2658 -1764
rect 2652 -1776 2658 -1770
rect 2652 -1782 2658 -1776
rect 2652 -2412 2658 -2406
rect 2652 -2418 2658 -2412
rect 2652 -2424 2658 -2418
rect 2652 -2430 2658 -2424
rect 2652 -2436 2658 -2430
rect 2652 -2442 2658 -2436
rect 2652 -2448 2658 -2442
rect 2652 -2454 2658 -2448
rect 2652 -2460 2658 -2454
rect 2652 -2466 2658 -2460
rect 2652 -2472 2658 -2466
rect 2652 -2478 2658 -2472
rect 2652 -2484 2658 -2478
rect 2652 -2490 2658 -2484
rect 2652 -2496 2658 -2490
rect 2652 -2502 2658 -2496
rect 2652 -2508 2658 -2502
rect 2652 -2514 2658 -2508
rect 2652 -2520 2658 -2514
rect 2652 -2526 2658 -2520
rect 2652 -2532 2658 -2526
rect 2652 -2538 2658 -2532
rect 2652 -2544 2658 -2538
rect 2652 -2550 2658 -2544
rect 2652 -2556 2658 -2550
rect 2652 -2562 2658 -2556
rect 2652 -2568 2658 -2562
rect 2652 -2574 2658 -2568
rect 2652 -2580 2658 -2574
rect 2652 -2586 2658 -2580
rect 2652 -2592 2658 -2586
rect 2652 -2598 2658 -2592
rect 2652 -2604 2658 -2598
rect 2652 -2610 2658 -2604
rect 2652 -2616 2658 -2610
rect 2652 -2622 2658 -2616
rect 2652 -2628 2658 -2622
rect 2652 -2634 2658 -2628
rect 2652 -2640 2658 -2634
rect 2652 -2646 2658 -2640
rect 2652 -2652 2658 -2646
rect 2652 -2658 2658 -2652
rect 2652 -2664 2658 -2658
rect 2652 -2670 2658 -2664
rect 2652 -2676 2658 -2670
rect 2652 -2682 2658 -2676
rect 2652 -2688 2658 -2682
rect 2652 -2694 2658 -2688
rect 2652 -2700 2658 -2694
rect 2652 -2706 2658 -2700
rect 2652 -2712 2658 -2706
rect 2652 -2718 2658 -2712
rect 2652 -2724 2658 -2718
rect 2652 -2730 2658 -2724
rect 2658 -1194 2664 -1188
rect 2658 -1200 2664 -1194
rect 2658 -1206 2664 -1200
rect 2658 -1212 2664 -1206
rect 2658 -1218 2664 -1212
rect 2658 -1224 2664 -1218
rect 2658 -1230 2664 -1224
rect 2658 -1236 2664 -1230
rect 2658 -1242 2664 -1236
rect 2658 -1248 2664 -1242
rect 2658 -1254 2664 -1248
rect 2658 -1260 2664 -1254
rect 2658 -1266 2664 -1260
rect 2658 -1272 2664 -1266
rect 2658 -1278 2664 -1272
rect 2658 -1284 2664 -1278
rect 2658 -1290 2664 -1284
rect 2658 -1296 2664 -1290
rect 2658 -1302 2664 -1296
rect 2658 -1308 2664 -1302
rect 2658 -1314 2664 -1308
rect 2658 -1320 2664 -1314
rect 2658 -1326 2664 -1320
rect 2658 -1332 2664 -1326
rect 2658 -1338 2664 -1332
rect 2658 -1344 2664 -1338
rect 2658 -1350 2664 -1344
rect 2658 -1356 2664 -1350
rect 2658 -1362 2664 -1356
rect 2658 -1368 2664 -1362
rect 2658 -1374 2664 -1368
rect 2658 -1380 2664 -1374
rect 2658 -1386 2664 -1380
rect 2658 -1392 2664 -1386
rect 2658 -1398 2664 -1392
rect 2658 -1404 2664 -1398
rect 2658 -1410 2664 -1404
rect 2658 -1416 2664 -1410
rect 2658 -1422 2664 -1416
rect 2658 -1428 2664 -1422
rect 2658 -1434 2664 -1428
rect 2658 -1440 2664 -1434
rect 2658 -1446 2664 -1440
rect 2658 -1452 2664 -1446
rect 2658 -1458 2664 -1452
rect 2658 -1464 2664 -1458
rect 2658 -1470 2664 -1464
rect 2658 -1476 2664 -1470
rect 2658 -1482 2664 -1476
rect 2658 -1488 2664 -1482
rect 2658 -1494 2664 -1488
rect 2658 -1500 2664 -1494
rect 2658 -1506 2664 -1500
rect 2658 -1512 2664 -1506
rect 2658 -1518 2664 -1512
rect 2658 -1524 2664 -1518
rect 2658 -1530 2664 -1524
rect 2658 -1536 2664 -1530
rect 2658 -1542 2664 -1536
rect 2658 -1548 2664 -1542
rect 2658 -1554 2664 -1548
rect 2658 -1560 2664 -1554
rect 2658 -1566 2664 -1560
rect 2658 -1572 2664 -1566
rect 2658 -1578 2664 -1572
rect 2658 -1584 2664 -1578
rect 2658 -1590 2664 -1584
rect 2658 -1596 2664 -1590
rect 2658 -1602 2664 -1596
rect 2658 -1608 2664 -1602
rect 2658 -1614 2664 -1608
rect 2658 -1620 2664 -1614
rect 2658 -1626 2664 -1620
rect 2658 -1632 2664 -1626
rect 2658 -1638 2664 -1632
rect 2658 -1644 2664 -1638
rect 2658 -1650 2664 -1644
rect 2658 -1656 2664 -1650
rect 2658 -1662 2664 -1656
rect 2658 -1668 2664 -1662
rect 2658 -1674 2664 -1668
rect 2658 -1680 2664 -1674
rect 2658 -1686 2664 -1680
rect 2658 -1692 2664 -1686
rect 2658 -1698 2664 -1692
rect 2658 -1704 2664 -1698
rect 2658 -1710 2664 -1704
rect 2658 -1716 2664 -1710
rect 2658 -1722 2664 -1716
rect 2658 -1728 2664 -1722
rect 2658 -1734 2664 -1728
rect 2658 -1740 2664 -1734
rect 2658 -1746 2664 -1740
rect 2658 -1752 2664 -1746
rect 2658 -1758 2664 -1752
rect 2658 -1764 2664 -1758
rect 2658 -1770 2664 -1764
rect 2658 -1776 2664 -1770
rect 2658 -2406 2664 -2400
rect 2658 -2412 2664 -2406
rect 2658 -2418 2664 -2412
rect 2658 -2424 2664 -2418
rect 2658 -2430 2664 -2424
rect 2658 -2436 2664 -2430
rect 2658 -2442 2664 -2436
rect 2658 -2448 2664 -2442
rect 2658 -2454 2664 -2448
rect 2658 -2460 2664 -2454
rect 2658 -2466 2664 -2460
rect 2658 -2472 2664 -2466
rect 2658 -2478 2664 -2472
rect 2658 -2484 2664 -2478
rect 2658 -2490 2664 -2484
rect 2658 -2496 2664 -2490
rect 2658 -2502 2664 -2496
rect 2658 -2508 2664 -2502
rect 2658 -2514 2664 -2508
rect 2658 -2520 2664 -2514
rect 2658 -2526 2664 -2520
rect 2658 -2532 2664 -2526
rect 2658 -2538 2664 -2532
rect 2658 -2544 2664 -2538
rect 2658 -2550 2664 -2544
rect 2658 -2556 2664 -2550
rect 2658 -2562 2664 -2556
rect 2658 -2568 2664 -2562
rect 2658 -2574 2664 -2568
rect 2658 -2580 2664 -2574
rect 2658 -2586 2664 -2580
rect 2658 -2592 2664 -2586
rect 2658 -2598 2664 -2592
rect 2658 -2604 2664 -2598
rect 2658 -2610 2664 -2604
rect 2658 -2616 2664 -2610
rect 2658 -2622 2664 -2616
rect 2658 -2628 2664 -2622
rect 2658 -2634 2664 -2628
rect 2658 -2640 2664 -2634
rect 2658 -2646 2664 -2640
rect 2658 -2652 2664 -2646
rect 2658 -2658 2664 -2652
rect 2658 -2664 2664 -2658
rect 2658 -2670 2664 -2664
rect 2658 -2676 2664 -2670
rect 2658 -2682 2664 -2676
rect 2658 -2688 2664 -2682
rect 2658 -2694 2664 -2688
rect 2658 -2700 2664 -2694
rect 2658 -2706 2664 -2700
rect 2658 -2712 2664 -2706
rect 2658 -2718 2664 -2712
rect 2658 -2724 2664 -2718
rect 2664 -1188 2670 -1182
rect 2664 -1194 2670 -1188
rect 2664 -1200 2670 -1194
rect 2664 -1206 2670 -1200
rect 2664 -1212 2670 -1206
rect 2664 -1218 2670 -1212
rect 2664 -1224 2670 -1218
rect 2664 -1230 2670 -1224
rect 2664 -1236 2670 -1230
rect 2664 -1242 2670 -1236
rect 2664 -1248 2670 -1242
rect 2664 -1254 2670 -1248
rect 2664 -1260 2670 -1254
rect 2664 -1266 2670 -1260
rect 2664 -1272 2670 -1266
rect 2664 -1278 2670 -1272
rect 2664 -1284 2670 -1278
rect 2664 -1290 2670 -1284
rect 2664 -1296 2670 -1290
rect 2664 -1302 2670 -1296
rect 2664 -1308 2670 -1302
rect 2664 -1314 2670 -1308
rect 2664 -1320 2670 -1314
rect 2664 -1326 2670 -1320
rect 2664 -1332 2670 -1326
rect 2664 -1338 2670 -1332
rect 2664 -1344 2670 -1338
rect 2664 -1350 2670 -1344
rect 2664 -1356 2670 -1350
rect 2664 -1362 2670 -1356
rect 2664 -1368 2670 -1362
rect 2664 -1374 2670 -1368
rect 2664 -1380 2670 -1374
rect 2664 -1386 2670 -1380
rect 2664 -1392 2670 -1386
rect 2664 -1398 2670 -1392
rect 2664 -1404 2670 -1398
rect 2664 -1410 2670 -1404
rect 2664 -1416 2670 -1410
rect 2664 -1422 2670 -1416
rect 2664 -1428 2670 -1422
rect 2664 -1434 2670 -1428
rect 2664 -1440 2670 -1434
rect 2664 -1446 2670 -1440
rect 2664 -1452 2670 -1446
rect 2664 -1458 2670 -1452
rect 2664 -1464 2670 -1458
rect 2664 -1470 2670 -1464
rect 2664 -1476 2670 -1470
rect 2664 -1482 2670 -1476
rect 2664 -1488 2670 -1482
rect 2664 -1494 2670 -1488
rect 2664 -1500 2670 -1494
rect 2664 -1506 2670 -1500
rect 2664 -1512 2670 -1506
rect 2664 -1518 2670 -1512
rect 2664 -1524 2670 -1518
rect 2664 -1530 2670 -1524
rect 2664 -1536 2670 -1530
rect 2664 -1542 2670 -1536
rect 2664 -1548 2670 -1542
rect 2664 -1554 2670 -1548
rect 2664 -1560 2670 -1554
rect 2664 -1566 2670 -1560
rect 2664 -1572 2670 -1566
rect 2664 -1578 2670 -1572
rect 2664 -1584 2670 -1578
rect 2664 -1590 2670 -1584
rect 2664 -1596 2670 -1590
rect 2664 -1602 2670 -1596
rect 2664 -1608 2670 -1602
rect 2664 -1614 2670 -1608
rect 2664 -1620 2670 -1614
rect 2664 -1626 2670 -1620
rect 2664 -1632 2670 -1626
rect 2664 -1638 2670 -1632
rect 2664 -1644 2670 -1638
rect 2664 -1650 2670 -1644
rect 2664 -1656 2670 -1650
rect 2664 -1662 2670 -1656
rect 2664 -1668 2670 -1662
rect 2664 -1674 2670 -1668
rect 2664 -1680 2670 -1674
rect 2664 -1686 2670 -1680
rect 2664 -1692 2670 -1686
rect 2664 -1698 2670 -1692
rect 2664 -1704 2670 -1698
rect 2664 -1710 2670 -1704
rect 2664 -1716 2670 -1710
rect 2664 -1722 2670 -1716
rect 2664 -1728 2670 -1722
rect 2664 -1734 2670 -1728
rect 2664 -1740 2670 -1734
rect 2664 -1746 2670 -1740
rect 2664 -1752 2670 -1746
rect 2664 -1758 2670 -1752
rect 2664 -1764 2670 -1758
rect 2664 -1770 2670 -1764
rect 2664 -2406 2670 -2400
rect 2664 -2412 2670 -2406
rect 2664 -2418 2670 -2412
rect 2664 -2424 2670 -2418
rect 2664 -2430 2670 -2424
rect 2664 -2436 2670 -2430
rect 2664 -2442 2670 -2436
rect 2664 -2448 2670 -2442
rect 2664 -2454 2670 -2448
rect 2664 -2460 2670 -2454
rect 2664 -2466 2670 -2460
rect 2664 -2472 2670 -2466
rect 2664 -2478 2670 -2472
rect 2664 -2484 2670 -2478
rect 2664 -2490 2670 -2484
rect 2664 -2496 2670 -2490
rect 2664 -2502 2670 -2496
rect 2664 -2508 2670 -2502
rect 2664 -2514 2670 -2508
rect 2664 -2520 2670 -2514
rect 2664 -2526 2670 -2520
rect 2664 -2532 2670 -2526
rect 2664 -2538 2670 -2532
rect 2664 -2544 2670 -2538
rect 2664 -2550 2670 -2544
rect 2664 -2556 2670 -2550
rect 2664 -2562 2670 -2556
rect 2664 -2568 2670 -2562
rect 2664 -2574 2670 -2568
rect 2664 -2580 2670 -2574
rect 2664 -2586 2670 -2580
rect 2664 -2592 2670 -2586
rect 2664 -2598 2670 -2592
rect 2664 -2604 2670 -2598
rect 2664 -2610 2670 -2604
rect 2664 -2616 2670 -2610
rect 2664 -2622 2670 -2616
rect 2664 -2628 2670 -2622
rect 2664 -2634 2670 -2628
rect 2664 -2640 2670 -2634
rect 2664 -2646 2670 -2640
rect 2664 -2652 2670 -2646
rect 2664 -2658 2670 -2652
rect 2664 -2664 2670 -2658
rect 2664 -2670 2670 -2664
rect 2664 -2676 2670 -2670
rect 2664 -2682 2670 -2676
rect 2664 -2688 2670 -2682
rect 2664 -2694 2670 -2688
rect 2664 -2700 2670 -2694
rect 2664 -2706 2670 -2700
rect 2664 -2712 2670 -2706
rect 2664 -2718 2670 -2712
rect 2664 -2724 2670 -2718
rect 2670 -1182 2676 -1176
rect 2670 -1188 2676 -1182
rect 2670 -1194 2676 -1188
rect 2670 -1200 2676 -1194
rect 2670 -1206 2676 -1200
rect 2670 -1212 2676 -1206
rect 2670 -1218 2676 -1212
rect 2670 -1224 2676 -1218
rect 2670 -1230 2676 -1224
rect 2670 -1236 2676 -1230
rect 2670 -1242 2676 -1236
rect 2670 -1248 2676 -1242
rect 2670 -1254 2676 -1248
rect 2670 -1260 2676 -1254
rect 2670 -1266 2676 -1260
rect 2670 -1272 2676 -1266
rect 2670 -1278 2676 -1272
rect 2670 -1284 2676 -1278
rect 2670 -1290 2676 -1284
rect 2670 -1296 2676 -1290
rect 2670 -1302 2676 -1296
rect 2670 -1308 2676 -1302
rect 2670 -1314 2676 -1308
rect 2670 -1320 2676 -1314
rect 2670 -1326 2676 -1320
rect 2670 -1332 2676 -1326
rect 2670 -1338 2676 -1332
rect 2670 -1344 2676 -1338
rect 2670 -1350 2676 -1344
rect 2670 -1356 2676 -1350
rect 2670 -1362 2676 -1356
rect 2670 -1368 2676 -1362
rect 2670 -1374 2676 -1368
rect 2670 -1380 2676 -1374
rect 2670 -1386 2676 -1380
rect 2670 -1392 2676 -1386
rect 2670 -1398 2676 -1392
rect 2670 -1404 2676 -1398
rect 2670 -1410 2676 -1404
rect 2670 -1416 2676 -1410
rect 2670 -1422 2676 -1416
rect 2670 -1428 2676 -1422
rect 2670 -1434 2676 -1428
rect 2670 -1440 2676 -1434
rect 2670 -1446 2676 -1440
rect 2670 -1452 2676 -1446
rect 2670 -1458 2676 -1452
rect 2670 -1464 2676 -1458
rect 2670 -1470 2676 -1464
rect 2670 -1476 2676 -1470
rect 2670 -1482 2676 -1476
rect 2670 -1488 2676 -1482
rect 2670 -1494 2676 -1488
rect 2670 -1500 2676 -1494
rect 2670 -1506 2676 -1500
rect 2670 -1512 2676 -1506
rect 2670 -1518 2676 -1512
rect 2670 -1524 2676 -1518
rect 2670 -1530 2676 -1524
rect 2670 -1536 2676 -1530
rect 2670 -1542 2676 -1536
rect 2670 -1548 2676 -1542
rect 2670 -1554 2676 -1548
rect 2670 -1560 2676 -1554
rect 2670 -1566 2676 -1560
rect 2670 -1572 2676 -1566
rect 2670 -1578 2676 -1572
rect 2670 -1584 2676 -1578
rect 2670 -1590 2676 -1584
rect 2670 -1596 2676 -1590
rect 2670 -1602 2676 -1596
rect 2670 -1608 2676 -1602
rect 2670 -1614 2676 -1608
rect 2670 -1620 2676 -1614
rect 2670 -1626 2676 -1620
rect 2670 -1632 2676 -1626
rect 2670 -1638 2676 -1632
rect 2670 -1644 2676 -1638
rect 2670 -1650 2676 -1644
rect 2670 -1656 2676 -1650
rect 2670 -1662 2676 -1656
rect 2670 -1668 2676 -1662
rect 2670 -1674 2676 -1668
rect 2670 -1680 2676 -1674
rect 2670 -1686 2676 -1680
rect 2670 -1692 2676 -1686
rect 2670 -1698 2676 -1692
rect 2670 -1704 2676 -1698
rect 2670 -1710 2676 -1704
rect 2670 -1716 2676 -1710
rect 2670 -1722 2676 -1716
rect 2670 -1728 2676 -1722
rect 2670 -1734 2676 -1728
rect 2670 -1740 2676 -1734
rect 2670 -1746 2676 -1740
rect 2670 -1752 2676 -1746
rect 2670 -1758 2676 -1752
rect 2670 -1764 2676 -1758
rect 2670 -2406 2676 -2400
rect 2670 -2412 2676 -2406
rect 2670 -2418 2676 -2412
rect 2670 -2424 2676 -2418
rect 2670 -2430 2676 -2424
rect 2670 -2436 2676 -2430
rect 2670 -2442 2676 -2436
rect 2670 -2448 2676 -2442
rect 2670 -2454 2676 -2448
rect 2670 -2460 2676 -2454
rect 2670 -2466 2676 -2460
rect 2670 -2472 2676 -2466
rect 2670 -2478 2676 -2472
rect 2670 -2484 2676 -2478
rect 2670 -2490 2676 -2484
rect 2670 -2496 2676 -2490
rect 2670 -2502 2676 -2496
rect 2670 -2508 2676 -2502
rect 2670 -2514 2676 -2508
rect 2670 -2520 2676 -2514
rect 2670 -2526 2676 -2520
rect 2670 -2532 2676 -2526
rect 2670 -2538 2676 -2532
rect 2670 -2544 2676 -2538
rect 2670 -2550 2676 -2544
rect 2670 -2556 2676 -2550
rect 2670 -2562 2676 -2556
rect 2670 -2568 2676 -2562
rect 2670 -2574 2676 -2568
rect 2670 -2580 2676 -2574
rect 2670 -2586 2676 -2580
rect 2670 -2592 2676 -2586
rect 2670 -2598 2676 -2592
rect 2670 -2604 2676 -2598
rect 2670 -2610 2676 -2604
rect 2670 -2616 2676 -2610
rect 2670 -2622 2676 -2616
rect 2670 -2628 2676 -2622
rect 2670 -2634 2676 -2628
rect 2670 -2640 2676 -2634
rect 2670 -2646 2676 -2640
rect 2670 -2652 2676 -2646
rect 2670 -2658 2676 -2652
rect 2670 -2664 2676 -2658
rect 2670 -2670 2676 -2664
rect 2670 -2676 2676 -2670
rect 2670 -2682 2676 -2676
rect 2670 -2688 2676 -2682
rect 2670 -2694 2676 -2688
rect 2670 -2700 2676 -2694
rect 2670 -2706 2676 -2700
rect 2670 -2712 2676 -2706
rect 2670 -2718 2676 -2712
rect 2676 -1182 2682 -1176
rect 2676 -1188 2682 -1182
rect 2676 -1194 2682 -1188
rect 2676 -1200 2682 -1194
rect 2676 -1206 2682 -1200
rect 2676 -1212 2682 -1206
rect 2676 -1218 2682 -1212
rect 2676 -1224 2682 -1218
rect 2676 -1230 2682 -1224
rect 2676 -1236 2682 -1230
rect 2676 -1242 2682 -1236
rect 2676 -1248 2682 -1242
rect 2676 -1254 2682 -1248
rect 2676 -1260 2682 -1254
rect 2676 -1266 2682 -1260
rect 2676 -1272 2682 -1266
rect 2676 -1278 2682 -1272
rect 2676 -1284 2682 -1278
rect 2676 -1290 2682 -1284
rect 2676 -1296 2682 -1290
rect 2676 -1302 2682 -1296
rect 2676 -1308 2682 -1302
rect 2676 -1314 2682 -1308
rect 2676 -1320 2682 -1314
rect 2676 -1326 2682 -1320
rect 2676 -1332 2682 -1326
rect 2676 -1338 2682 -1332
rect 2676 -1344 2682 -1338
rect 2676 -1350 2682 -1344
rect 2676 -1356 2682 -1350
rect 2676 -1362 2682 -1356
rect 2676 -1368 2682 -1362
rect 2676 -1374 2682 -1368
rect 2676 -1380 2682 -1374
rect 2676 -1386 2682 -1380
rect 2676 -1392 2682 -1386
rect 2676 -1398 2682 -1392
rect 2676 -1404 2682 -1398
rect 2676 -1410 2682 -1404
rect 2676 -1416 2682 -1410
rect 2676 -1422 2682 -1416
rect 2676 -1428 2682 -1422
rect 2676 -1434 2682 -1428
rect 2676 -1440 2682 -1434
rect 2676 -1446 2682 -1440
rect 2676 -1452 2682 -1446
rect 2676 -1458 2682 -1452
rect 2676 -1464 2682 -1458
rect 2676 -1470 2682 -1464
rect 2676 -1476 2682 -1470
rect 2676 -1482 2682 -1476
rect 2676 -1488 2682 -1482
rect 2676 -1494 2682 -1488
rect 2676 -1500 2682 -1494
rect 2676 -1506 2682 -1500
rect 2676 -1512 2682 -1506
rect 2676 -1518 2682 -1512
rect 2676 -1524 2682 -1518
rect 2676 -1530 2682 -1524
rect 2676 -1536 2682 -1530
rect 2676 -1542 2682 -1536
rect 2676 -1548 2682 -1542
rect 2676 -1554 2682 -1548
rect 2676 -1560 2682 -1554
rect 2676 -1566 2682 -1560
rect 2676 -1572 2682 -1566
rect 2676 -1578 2682 -1572
rect 2676 -1584 2682 -1578
rect 2676 -1590 2682 -1584
rect 2676 -1596 2682 -1590
rect 2676 -1602 2682 -1596
rect 2676 -1608 2682 -1602
rect 2676 -1614 2682 -1608
rect 2676 -1620 2682 -1614
rect 2676 -1626 2682 -1620
rect 2676 -1632 2682 -1626
rect 2676 -1638 2682 -1632
rect 2676 -1644 2682 -1638
rect 2676 -1650 2682 -1644
rect 2676 -1656 2682 -1650
rect 2676 -1662 2682 -1656
rect 2676 -1668 2682 -1662
rect 2676 -1674 2682 -1668
rect 2676 -1680 2682 -1674
rect 2676 -1686 2682 -1680
rect 2676 -1692 2682 -1686
rect 2676 -1698 2682 -1692
rect 2676 -1704 2682 -1698
rect 2676 -1710 2682 -1704
rect 2676 -1716 2682 -1710
rect 2676 -1722 2682 -1716
rect 2676 -1728 2682 -1722
rect 2676 -1734 2682 -1728
rect 2676 -1740 2682 -1734
rect 2676 -1746 2682 -1740
rect 2676 -1752 2682 -1746
rect 2676 -2406 2682 -2400
rect 2676 -2412 2682 -2406
rect 2676 -2418 2682 -2412
rect 2676 -2424 2682 -2418
rect 2676 -2430 2682 -2424
rect 2676 -2436 2682 -2430
rect 2676 -2442 2682 -2436
rect 2676 -2448 2682 -2442
rect 2676 -2454 2682 -2448
rect 2676 -2460 2682 -2454
rect 2676 -2466 2682 -2460
rect 2676 -2472 2682 -2466
rect 2676 -2478 2682 -2472
rect 2676 -2484 2682 -2478
rect 2676 -2490 2682 -2484
rect 2676 -2496 2682 -2490
rect 2676 -2502 2682 -2496
rect 2676 -2508 2682 -2502
rect 2676 -2514 2682 -2508
rect 2676 -2520 2682 -2514
rect 2676 -2526 2682 -2520
rect 2676 -2532 2682 -2526
rect 2676 -2538 2682 -2532
rect 2676 -2544 2682 -2538
rect 2676 -2550 2682 -2544
rect 2676 -2556 2682 -2550
rect 2676 -2562 2682 -2556
rect 2676 -2568 2682 -2562
rect 2676 -2574 2682 -2568
rect 2676 -2580 2682 -2574
rect 2676 -2586 2682 -2580
rect 2676 -2592 2682 -2586
rect 2676 -2598 2682 -2592
rect 2676 -2604 2682 -2598
rect 2676 -2610 2682 -2604
rect 2676 -2616 2682 -2610
rect 2676 -2622 2682 -2616
rect 2676 -2628 2682 -2622
rect 2676 -2634 2682 -2628
rect 2676 -2640 2682 -2634
rect 2676 -2646 2682 -2640
rect 2676 -2652 2682 -2646
rect 2676 -2658 2682 -2652
rect 2676 -2664 2682 -2658
rect 2676 -2670 2682 -2664
rect 2676 -2676 2682 -2670
rect 2676 -2682 2682 -2676
rect 2676 -2688 2682 -2682
rect 2676 -2694 2682 -2688
rect 2676 -2700 2682 -2694
rect 2676 -2706 2682 -2700
rect 2676 -2712 2682 -2706
rect 2682 -1176 2688 -1170
rect 2682 -1182 2688 -1176
rect 2682 -1188 2688 -1182
rect 2682 -1194 2688 -1188
rect 2682 -1200 2688 -1194
rect 2682 -1206 2688 -1200
rect 2682 -1212 2688 -1206
rect 2682 -1218 2688 -1212
rect 2682 -1224 2688 -1218
rect 2682 -1230 2688 -1224
rect 2682 -1236 2688 -1230
rect 2682 -1242 2688 -1236
rect 2682 -1248 2688 -1242
rect 2682 -1254 2688 -1248
rect 2682 -1260 2688 -1254
rect 2682 -1266 2688 -1260
rect 2682 -1272 2688 -1266
rect 2682 -1278 2688 -1272
rect 2682 -1284 2688 -1278
rect 2682 -1290 2688 -1284
rect 2682 -1296 2688 -1290
rect 2682 -1302 2688 -1296
rect 2682 -1308 2688 -1302
rect 2682 -1314 2688 -1308
rect 2682 -1320 2688 -1314
rect 2682 -1326 2688 -1320
rect 2682 -1332 2688 -1326
rect 2682 -1338 2688 -1332
rect 2682 -1344 2688 -1338
rect 2682 -1350 2688 -1344
rect 2682 -1356 2688 -1350
rect 2682 -1362 2688 -1356
rect 2682 -1368 2688 -1362
rect 2682 -1374 2688 -1368
rect 2682 -1380 2688 -1374
rect 2682 -1386 2688 -1380
rect 2682 -1392 2688 -1386
rect 2682 -1398 2688 -1392
rect 2682 -1404 2688 -1398
rect 2682 -1410 2688 -1404
rect 2682 -1416 2688 -1410
rect 2682 -1422 2688 -1416
rect 2682 -1428 2688 -1422
rect 2682 -1434 2688 -1428
rect 2682 -1440 2688 -1434
rect 2682 -1446 2688 -1440
rect 2682 -1452 2688 -1446
rect 2682 -1458 2688 -1452
rect 2682 -1464 2688 -1458
rect 2682 -1470 2688 -1464
rect 2682 -1476 2688 -1470
rect 2682 -1482 2688 -1476
rect 2682 -1488 2688 -1482
rect 2682 -1494 2688 -1488
rect 2682 -1500 2688 -1494
rect 2682 -1506 2688 -1500
rect 2682 -1512 2688 -1506
rect 2682 -1518 2688 -1512
rect 2682 -1524 2688 -1518
rect 2682 -1530 2688 -1524
rect 2682 -1536 2688 -1530
rect 2682 -1542 2688 -1536
rect 2682 -1548 2688 -1542
rect 2682 -1554 2688 -1548
rect 2682 -1560 2688 -1554
rect 2682 -1566 2688 -1560
rect 2682 -1572 2688 -1566
rect 2682 -1578 2688 -1572
rect 2682 -1584 2688 -1578
rect 2682 -1590 2688 -1584
rect 2682 -1596 2688 -1590
rect 2682 -1602 2688 -1596
rect 2682 -1608 2688 -1602
rect 2682 -1614 2688 -1608
rect 2682 -1620 2688 -1614
rect 2682 -1626 2688 -1620
rect 2682 -1632 2688 -1626
rect 2682 -1638 2688 -1632
rect 2682 -1644 2688 -1638
rect 2682 -1650 2688 -1644
rect 2682 -1656 2688 -1650
rect 2682 -1662 2688 -1656
rect 2682 -1668 2688 -1662
rect 2682 -1674 2688 -1668
rect 2682 -1680 2688 -1674
rect 2682 -1686 2688 -1680
rect 2682 -1692 2688 -1686
rect 2682 -1698 2688 -1692
rect 2682 -1704 2688 -1698
rect 2682 -1710 2688 -1704
rect 2682 -1716 2688 -1710
rect 2682 -1722 2688 -1716
rect 2682 -1728 2688 -1722
rect 2682 -1734 2688 -1728
rect 2682 -1740 2688 -1734
rect 2682 -1746 2688 -1740
rect 2682 -2400 2688 -2394
rect 2682 -2406 2688 -2400
rect 2682 -2412 2688 -2406
rect 2682 -2418 2688 -2412
rect 2682 -2424 2688 -2418
rect 2682 -2430 2688 -2424
rect 2682 -2436 2688 -2430
rect 2682 -2442 2688 -2436
rect 2682 -2448 2688 -2442
rect 2682 -2454 2688 -2448
rect 2682 -2460 2688 -2454
rect 2682 -2466 2688 -2460
rect 2682 -2472 2688 -2466
rect 2682 -2478 2688 -2472
rect 2682 -2484 2688 -2478
rect 2682 -2490 2688 -2484
rect 2682 -2496 2688 -2490
rect 2682 -2502 2688 -2496
rect 2682 -2508 2688 -2502
rect 2682 -2514 2688 -2508
rect 2682 -2520 2688 -2514
rect 2682 -2526 2688 -2520
rect 2682 -2532 2688 -2526
rect 2682 -2538 2688 -2532
rect 2682 -2544 2688 -2538
rect 2682 -2550 2688 -2544
rect 2682 -2556 2688 -2550
rect 2682 -2562 2688 -2556
rect 2682 -2568 2688 -2562
rect 2682 -2574 2688 -2568
rect 2682 -2580 2688 -2574
rect 2682 -2586 2688 -2580
rect 2682 -2592 2688 -2586
rect 2682 -2598 2688 -2592
rect 2682 -2604 2688 -2598
rect 2682 -2610 2688 -2604
rect 2682 -2616 2688 -2610
rect 2682 -2622 2688 -2616
rect 2682 -2628 2688 -2622
rect 2682 -2634 2688 -2628
rect 2682 -2640 2688 -2634
rect 2682 -2646 2688 -2640
rect 2682 -2652 2688 -2646
rect 2682 -2658 2688 -2652
rect 2682 -2664 2688 -2658
rect 2682 -2670 2688 -2664
rect 2682 -2676 2688 -2670
rect 2682 -2682 2688 -2676
rect 2682 -2688 2688 -2682
rect 2682 -2694 2688 -2688
rect 2682 -2700 2688 -2694
rect 2682 -2706 2688 -2700
rect 2682 -2712 2688 -2706
rect 2688 -1170 2694 -1164
rect 2688 -1176 2694 -1170
rect 2688 -1182 2694 -1176
rect 2688 -1188 2694 -1182
rect 2688 -1194 2694 -1188
rect 2688 -1200 2694 -1194
rect 2688 -1206 2694 -1200
rect 2688 -1212 2694 -1206
rect 2688 -1218 2694 -1212
rect 2688 -1224 2694 -1218
rect 2688 -1230 2694 -1224
rect 2688 -1236 2694 -1230
rect 2688 -1242 2694 -1236
rect 2688 -1248 2694 -1242
rect 2688 -1254 2694 -1248
rect 2688 -1260 2694 -1254
rect 2688 -1266 2694 -1260
rect 2688 -1272 2694 -1266
rect 2688 -1278 2694 -1272
rect 2688 -1284 2694 -1278
rect 2688 -1290 2694 -1284
rect 2688 -1296 2694 -1290
rect 2688 -1302 2694 -1296
rect 2688 -1308 2694 -1302
rect 2688 -1314 2694 -1308
rect 2688 -1320 2694 -1314
rect 2688 -1326 2694 -1320
rect 2688 -1332 2694 -1326
rect 2688 -1338 2694 -1332
rect 2688 -1344 2694 -1338
rect 2688 -1350 2694 -1344
rect 2688 -1356 2694 -1350
rect 2688 -1362 2694 -1356
rect 2688 -1368 2694 -1362
rect 2688 -1374 2694 -1368
rect 2688 -1380 2694 -1374
rect 2688 -1386 2694 -1380
rect 2688 -1392 2694 -1386
rect 2688 -1398 2694 -1392
rect 2688 -1404 2694 -1398
rect 2688 -1410 2694 -1404
rect 2688 -1416 2694 -1410
rect 2688 -1422 2694 -1416
rect 2688 -1428 2694 -1422
rect 2688 -1434 2694 -1428
rect 2688 -1440 2694 -1434
rect 2688 -1446 2694 -1440
rect 2688 -1452 2694 -1446
rect 2688 -1458 2694 -1452
rect 2688 -1464 2694 -1458
rect 2688 -1470 2694 -1464
rect 2688 -1476 2694 -1470
rect 2688 -1482 2694 -1476
rect 2688 -1488 2694 -1482
rect 2688 -1494 2694 -1488
rect 2688 -1500 2694 -1494
rect 2688 -1506 2694 -1500
rect 2688 -1512 2694 -1506
rect 2688 -1518 2694 -1512
rect 2688 -1524 2694 -1518
rect 2688 -1530 2694 -1524
rect 2688 -1536 2694 -1530
rect 2688 -1542 2694 -1536
rect 2688 -1548 2694 -1542
rect 2688 -1554 2694 -1548
rect 2688 -1560 2694 -1554
rect 2688 -1566 2694 -1560
rect 2688 -1572 2694 -1566
rect 2688 -1578 2694 -1572
rect 2688 -1584 2694 -1578
rect 2688 -1590 2694 -1584
rect 2688 -1596 2694 -1590
rect 2688 -1602 2694 -1596
rect 2688 -1608 2694 -1602
rect 2688 -1614 2694 -1608
rect 2688 -1620 2694 -1614
rect 2688 -1626 2694 -1620
rect 2688 -1632 2694 -1626
rect 2688 -1638 2694 -1632
rect 2688 -1644 2694 -1638
rect 2688 -1650 2694 -1644
rect 2688 -1656 2694 -1650
rect 2688 -1662 2694 -1656
rect 2688 -1668 2694 -1662
rect 2688 -1674 2694 -1668
rect 2688 -1680 2694 -1674
rect 2688 -1686 2694 -1680
rect 2688 -1692 2694 -1686
rect 2688 -1698 2694 -1692
rect 2688 -1704 2694 -1698
rect 2688 -1710 2694 -1704
rect 2688 -1716 2694 -1710
rect 2688 -1722 2694 -1716
rect 2688 -1728 2694 -1722
rect 2688 -1734 2694 -1728
rect 2688 -1740 2694 -1734
rect 2688 -2400 2694 -2394
rect 2688 -2406 2694 -2400
rect 2688 -2412 2694 -2406
rect 2688 -2418 2694 -2412
rect 2688 -2424 2694 -2418
rect 2688 -2430 2694 -2424
rect 2688 -2436 2694 -2430
rect 2688 -2442 2694 -2436
rect 2688 -2448 2694 -2442
rect 2688 -2454 2694 -2448
rect 2688 -2460 2694 -2454
rect 2688 -2466 2694 -2460
rect 2688 -2472 2694 -2466
rect 2688 -2478 2694 -2472
rect 2688 -2484 2694 -2478
rect 2688 -2490 2694 -2484
rect 2688 -2496 2694 -2490
rect 2688 -2502 2694 -2496
rect 2688 -2508 2694 -2502
rect 2688 -2514 2694 -2508
rect 2688 -2520 2694 -2514
rect 2688 -2526 2694 -2520
rect 2688 -2532 2694 -2526
rect 2688 -2538 2694 -2532
rect 2688 -2544 2694 -2538
rect 2688 -2550 2694 -2544
rect 2688 -2556 2694 -2550
rect 2688 -2562 2694 -2556
rect 2688 -2568 2694 -2562
rect 2688 -2574 2694 -2568
rect 2688 -2580 2694 -2574
rect 2688 -2586 2694 -2580
rect 2688 -2592 2694 -2586
rect 2688 -2598 2694 -2592
rect 2688 -2604 2694 -2598
rect 2688 -2610 2694 -2604
rect 2688 -2616 2694 -2610
rect 2688 -2622 2694 -2616
rect 2688 -2628 2694 -2622
rect 2688 -2634 2694 -2628
rect 2688 -2640 2694 -2634
rect 2688 -2646 2694 -2640
rect 2688 -2652 2694 -2646
rect 2688 -2658 2694 -2652
rect 2688 -2664 2694 -2658
rect 2688 -2670 2694 -2664
rect 2688 -2676 2694 -2670
rect 2688 -2682 2694 -2676
rect 2688 -2688 2694 -2682
rect 2688 -2694 2694 -2688
rect 2688 -2700 2694 -2694
rect 2688 -2706 2694 -2700
rect 2694 -1170 2700 -1164
rect 2694 -1176 2700 -1170
rect 2694 -1182 2700 -1176
rect 2694 -1188 2700 -1182
rect 2694 -1194 2700 -1188
rect 2694 -1200 2700 -1194
rect 2694 -1206 2700 -1200
rect 2694 -1212 2700 -1206
rect 2694 -1218 2700 -1212
rect 2694 -1224 2700 -1218
rect 2694 -1230 2700 -1224
rect 2694 -1236 2700 -1230
rect 2694 -1242 2700 -1236
rect 2694 -1248 2700 -1242
rect 2694 -1254 2700 -1248
rect 2694 -1260 2700 -1254
rect 2694 -1266 2700 -1260
rect 2694 -1272 2700 -1266
rect 2694 -1278 2700 -1272
rect 2694 -1284 2700 -1278
rect 2694 -1290 2700 -1284
rect 2694 -1296 2700 -1290
rect 2694 -1302 2700 -1296
rect 2694 -1308 2700 -1302
rect 2694 -1314 2700 -1308
rect 2694 -1320 2700 -1314
rect 2694 -1326 2700 -1320
rect 2694 -1332 2700 -1326
rect 2694 -1338 2700 -1332
rect 2694 -1344 2700 -1338
rect 2694 -1350 2700 -1344
rect 2694 -1356 2700 -1350
rect 2694 -1362 2700 -1356
rect 2694 -1368 2700 -1362
rect 2694 -1374 2700 -1368
rect 2694 -1380 2700 -1374
rect 2694 -1386 2700 -1380
rect 2694 -1392 2700 -1386
rect 2694 -1398 2700 -1392
rect 2694 -1404 2700 -1398
rect 2694 -1410 2700 -1404
rect 2694 -1416 2700 -1410
rect 2694 -1422 2700 -1416
rect 2694 -1428 2700 -1422
rect 2694 -1434 2700 -1428
rect 2694 -1440 2700 -1434
rect 2694 -1446 2700 -1440
rect 2694 -1452 2700 -1446
rect 2694 -1458 2700 -1452
rect 2694 -1464 2700 -1458
rect 2694 -1470 2700 -1464
rect 2694 -1476 2700 -1470
rect 2694 -1482 2700 -1476
rect 2694 -1488 2700 -1482
rect 2694 -1494 2700 -1488
rect 2694 -1500 2700 -1494
rect 2694 -1506 2700 -1500
rect 2694 -1512 2700 -1506
rect 2694 -1518 2700 -1512
rect 2694 -1524 2700 -1518
rect 2694 -1530 2700 -1524
rect 2694 -1536 2700 -1530
rect 2694 -1542 2700 -1536
rect 2694 -1548 2700 -1542
rect 2694 -1554 2700 -1548
rect 2694 -1560 2700 -1554
rect 2694 -1566 2700 -1560
rect 2694 -1572 2700 -1566
rect 2694 -1578 2700 -1572
rect 2694 -1584 2700 -1578
rect 2694 -1590 2700 -1584
rect 2694 -1596 2700 -1590
rect 2694 -1602 2700 -1596
rect 2694 -1608 2700 -1602
rect 2694 -1614 2700 -1608
rect 2694 -1620 2700 -1614
rect 2694 -1626 2700 -1620
rect 2694 -1632 2700 -1626
rect 2694 -1638 2700 -1632
rect 2694 -1644 2700 -1638
rect 2694 -1650 2700 -1644
rect 2694 -1656 2700 -1650
rect 2694 -1662 2700 -1656
rect 2694 -1668 2700 -1662
rect 2694 -1674 2700 -1668
rect 2694 -1680 2700 -1674
rect 2694 -1686 2700 -1680
rect 2694 -1692 2700 -1686
rect 2694 -1698 2700 -1692
rect 2694 -1704 2700 -1698
rect 2694 -1710 2700 -1704
rect 2694 -1716 2700 -1710
rect 2694 -1722 2700 -1716
rect 2694 -1728 2700 -1722
rect 2694 -2400 2700 -2394
rect 2694 -2406 2700 -2400
rect 2694 -2412 2700 -2406
rect 2694 -2418 2700 -2412
rect 2694 -2424 2700 -2418
rect 2694 -2430 2700 -2424
rect 2694 -2436 2700 -2430
rect 2694 -2442 2700 -2436
rect 2694 -2448 2700 -2442
rect 2694 -2454 2700 -2448
rect 2694 -2460 2700 -2454
rect 2694 -2466 2700 -2460
rect 2694 -2472 2700 -2466
rect 2694 -2478 2700 -2472
rect 2694 -2484 2700 -2478
rect 2694 -2490 2700 -2484
rect 2694 -2496 2700 -2490
rect 2694 -2502 2700 -2496
rect 2694 -2508 2700 -2502
rect 2694 -2514 2700 -2508
rect 2694 -2520 2700 -2514
rect 2694 -2526 2700 -2520
rect 2694 -2532 2700 -2526
rect 2694 -2538 2700 -2532
rect 2694 -2544 2700 -2538
rect 2694 -2550 2700 -2544
rect 2694 -2556 2700 -2550
rect 2694 -2562 2700 -2556
rect 2694 -2568 2700 -2562
rect 2694 -2574 2700 -2568
rect 2694 -2580 2700 -2574
rect 2694 -2586 2700 -2580
rect 2694 -2592 2700 -2586
rect 2694 -2598 2700 -2592
rect 2694 -2604 2700 -2598
rect 2694 -2610 2700 -2604
rect 2694 -2616 2700 -2610
rect 2694 -2622 2700 -2616
rect 2694 -2628 2700 -2622
rect 2694 -2634 2700 -2628
rect 2694 -2640 2700 -2634
rect 2694 -2646 2700 -2640
rect 2694 -2652 2700 -2646
rect 2694 -2658 2700 -2652
rect 2694 -2664 2700 -2658
rect 2694 -2670 2700 -2664
rect 2694 -2676 2700 -2670
rect 2694 -2682 2700 -2676
rect 2694 -2688 2700 -2682
rect 2694 -2694 2700 -2688
rect 2694 -2700 2700 -2694
rect 2700 -1164 2706 -1158
rect 2700 -1170 2706 -1164
rect 2700 -1176 2706 -1170
rect 2700 -1182 2706 -1176
rect 2700 -1188 2706 -1182
rect 2700 -1194 2706 -1188
rect 2700 -1200 2706 -1194
rect 2700 -1206 2706 -1200
rect 2700 -1212 2706 -1206
rect 2700 -1218 2706 -1212
rect 2700 -1224 2706 -1218
rect 2700 -1230 2706 -1224
rect 2700 -1236 2706 -1230
rect 2700 -1242 2706 -1236
rect 2700 -1248 2706 -1242
rect 2700 -1254 2706 -1248
rect 2700 -1260 2706 -1254
rect 2700 -1266 2706 -1260
rect 2700 -1272 2706 -1266
rect 2700 -1278 2706 -1272
rect 2700 -1284 2706 -1278
rect 2700 -1290 2706 -1284
rect 2700 -1296 2706 -1290
rect 2700 -1302 2706 -1296
rect 2700 -1308 2706 -1302
rect 2700 -1314 2706 -1308
rect 2700 -1320 2706 -1314
rect 2700 -1326 2706 -1320
rect 2700 -1332 2706 -1326
rect 2700 -1338 2706 -1332
rect 2700 -1344 2706 -1338
rect 2700 -1350 2706 -1344
rect 2700 -1356 2706 -1350
rect 2700 -1362 2706 -1356
rect 2700 -1368 2706 -1362
rect 2700 -1374 2706 -1368
rect 2700 -1380 2706 -1374
rect 2700 -1386 2706 -1380
rect 2700 -1392 2706 -1386
rect 2700 -1398 2706 -1392
rect 2700 -1404 2706 -1398
rect 2700 -1410 2706 -1404
rect 2700 -1416 2706 -1410
rect 2700 -1422 2706 -1416
rect 2700 -1428 2706 -1422
rect 2700 -1434 2706 -1428
rect 2700 -1440 2706 -1434
rect 2700 -1446 2706 -1440
rect 2700 -1452 2706 -1446
rect 2700 -1458 2706 -1452
rect 2700 -1464 2706 -1458
rect 2700 -1470 2706 -1464
rect 2700 -1476 2706 -1470
rect 2700 -1482 2706 -1476
rect 2700 -1488 2706 -1482
rect 2700 -1494 2706 -1488
rect 2700 -1500 2706 -1494
rect 2700 -1506 2706 -1500
rect 2700 -1512 2706 -1506
rect 2700 -1518 2706 -1512
rect 2700 -1524 2706 -1518
rect 2700 -1530 2706 -1524
rect 2700 -1536 2706 -1530
rect 2700 -1542 2706 -1536
rect 2700 -1548 2706 -1542
rect 2700 -1554 2706 -1548
rect 2700 -1560 2706 -1554
rect 2700 -1566 2706 -1560
rect 2700 -1572 2706 -1566
rect 2700 -1578 2706 -1572
rect 2700 -1584 2706 -1578
rect 2700 -1590 2706 -1584
rect 2700 -1596 2706 -1590
rect 2700 -1602 2706 -1596
rect 2700 -1608 2706 -1602
rect 2700 -1614 2706 -1608
rect 2700 -1620 2706 -1614
rect 2700 -1626 2706 -1620
rect 2700 -1632 2706 -1626
rect 2700 -1638 2706 -1632
rect 2700 -1644 2706 -1638
rect 2700 -1650 2706 -1644
rect 2700 -1656 2706 -1650
rect 2700 -1662 2706 -1656
rect 2700 -1668 2706 -1662
rect 2700 -1674 2706 -1668
rect 2700 -1680 2706 -1674
rect 2700 -1686 2706 -1680
rect 2700 -1692 2706 -1686
rect 2700 -1698 2706 -1692
rect 2700 -1704 2706 -1698
rect 2700 -1710 2706 -1704
rect 2700 -1716 2706 -1710
rect 2700 -1722 2706 -1716
rect 2700 -2400 2706 -2394
rect 2700 -2406 2706 -2400
rect 2700 -2412 2706 -2406
rect 2700 -2418 2706 -2412
rect 2700 -2424 2706 -2418
rect 2700 -2430 2706 -2424
rect 2700 -2436 2706 -2430
rect 2700 -2442 2706 -2436
rect 2700 -2448 2706 -2442
rect 2700 -2454 2706 -2448
rect 2700 -2460 2706 -2454
rect 2700 -2466 2706 -2460
rect 2700 -2472 2706 -2466
rect 2700 -2478 2706 -2472
rect 2700 -2484 2706 -2478
rect 2700 -2490 2706 -2484
rect 2700 -2496 2706 -2490
rect 2700 -2502 2706 -2496
rect 2700 -2508 2706 -2502
rect 2700 -2514 2706 -2508
rect 2700 -2520 2706 -2514
rect 2700 -2526 2706 -2520
rect 2700 -2532 2706 -2526
rect 2700 -2538 2706 -2532
rect 2700 -2544 2706 -2538
rect 2700 -2550 2706 -2544
rect 2700 -2556 2706 -2550
rect 2700 -2562 2706 -2556
rect 2700 -2568 2706 -2562
rect 2700 -2574 2706 -2568
rect 2700 -2580 2706 -2574
rect 2700 -2586 2706 -2580
rect 2700 -2592 2706 -2586
rect 2700 -2598 2706 -2592
rect 2700 -2604 2706 -2598
rect 2700 -2610 2706 -2604
rect 2700 -2616 2706 -2610
rect 2700 -2622 2706 -2616
rect 2700 -2628 2706 -2622
rect 2700 -2634 2706 -2628
rect 2700 -2640 2706 -2634
rect 2700 -2646 2706 -2640
rect 2700 -2652 2706 -2646
rect 2700 -2658 2706 -2652
rect 2700 -2664 2706 -2658
rect 2700 -2670 2706 -2664
rect 2700 -2676 2706 -2670
rect 2700 -2682 2706 -2676
rect 2700 -2688 2706 -2682
rect 2700 -2694 2706 -2688
rect 2706 -1158 2712 -1152
rect 2706 -1164 2712 -1158
rect 2706 -1170 2712 -1164
rect 2706 -1176 2712 -1170
rect 2706 -1182 2712 -1176
rect 2706 -1188 2712 -1182
rect 2706 -1194 2712 -1188
rect 2706 -1200 2712 -1194
rect 2706 -1206 2712 -1200
rect 2706 -1212 2712 -1206
rect 2706 -1218 2712 -1212
rect 2706 -1224 2712 -1218
rect 2706 -1230 2712 -1224
rect 2706 -1236 2712 -1230
rect 2706 -1242 2712 -1236
rect 2706 -1248 2712 -1242
rect 2706 -1254 2712 -1248
rect 2706 -1260 2712 -1254
rect 2706 -1266 2712 -1260
rect 2706 -1272 2712 -1266
rect 2706 -1278 2712 -1272
rect 2706 -1284 2712 -1278
rect 2706 -1290 2712 -1284
rect 2706 -1296 2712 -1290
rect 2706 -1302 2712 -1296
rect 2706 -1308 2712 -1302
rect 2706 -1314 2712 -1308
rect 2706 -1320 2712 -1314
rect 2706 -1326 2712 -1320
rect 2706 -1332 2712 -1326
rect 2706 -1338 2712 -1332
rect 2706 -1344 2712 -1338
rect 2706 -1350 2712 -1344
rect 2706 -1356 2712 -1350
rect 2706 -1362 2712 -1356
rect 2706 -1368 2712 -1362
rect 2706 -1374 2712 -1368
rect 2706 -1380 2712 -1374
rect 2706 -1386 2712 -1380
rect 2706 -1392 2712 -1386
rect 2706 -1398 2712 -1392
rect 2706 -1404 2712 -1398
rect 2706 -1410 2712 -1404
rect 2706 -1416 2712 -1410
rect 2706 -1422 2712 -1416
rect 2706 -1428 2712 -1422
rect 2706 -1434 2712 -1428
rect 2706 -1440 2712 -1434
rect 2706 -1446 2712 -1440
rect 2706 -1452 2712 -1446
rect 2706 -1458 2712 -1452
rect 2706 -1464 2712 -1458
rect 2706 -1470 2712 -1464
rect 2706 -1476 2712 -1470
rect 2706 -1482 2712 -1476
rect 2706 -1488 2712 -1482
rect 2706 -1494 2712 -1488
rect 2706 -1500 2712 -1494
rect 2706 -1506 2712 -1500
rect 2706 -1512 2712 -1506
rect 2706 -1518 2712 -1512
rect 2706 -1524 2712 -1518
rect 2706 -1530 2712 -1524
rect 2706 -1536 2712 -1530
rect 2706 -1542 2712 -1536
rect 2706 -1548 2712 -1542
rect 2706 -1554 2712 -1548
rect 2706 -1560 2712 -1554
rect 2706 -1566 2712 -1560
rect 2706 -1572 2712 -1566
rect 2706 -1578 2712 -1572
rect 2706 -1584 2712 -1578
rect 2706 -1590 2712 -1584
rect 2706 -1596 2712 -1590
rect 2706 -1602 2712 -1596
rect 2706 -1608 2712 -1602
rect 2706 -1614 2712 -1608
rect 2706 -1620 2712 -1614
rect 2706 -1626 2712 -1620
rect 2706 -1632 2712 -1626
rect 2706 -1638 2712 -1632
rect 2706 -1644 2712 -1638
rect 2706 -1650 2712 -1644
rect 2706 -1656 2712 -1650
rect 2706 -1662 2712 -1656
rect 2706 -1668 2712 -1662
rect 2706 -1674 2712 -1668
rect 2706 -1680 2712 -1674
rect 2706 -1686 2712 -1680
rect 2706 -1692 2712 -1686
rect 2706 -1698 2712 -1692
rect 2706 -1704 2712 -1698
rect 2706 -1710 2712 -1704
rect 2706 -1716 2712 -1710
rect 2706 -2394 2712 -2388
rect 2706 -2400 2712 -2394
rect 2706 -2406 2712 -2400
rect 2706 -2412 2712 -2406
rect 2706 -2418 2712 -2412
rect 2706 -2424 2712 -2418
rect 2706 -2430 2712 -2424
rect 2706 -2436 2712 -2430
rect 2706 -2442 2712 -2436
rect 2706 -2448 2712 -2442
rect 2706 -2454 2712 -2448
rect 2706 -2460 2712 -2454
rect 2706 -2466 2712 -2460
rect 2706 -2472 2712 -2466
rect 2706 -2478 2712 -2472
rect 2706 -2484 2712 -2478
rect 2706 -2490 2712 -2484
rect 2706 -2496 2712 -2490
rect 2706 -2502 2712 -2496
rect 2706 -2508 2712 -2502
rect 2706 -2514 2712 -2508
rect 2706 -2520 2712 -2514
rect 2706 -2526 2712 -2520
rect 2706 -2532 2712 -2526
rect 2706 -2538 2712 -2532
rect 2706 -2544 2712 -2538
rect 2706 -2550 2712 -2544
rect 2706 -2556 2712 -2550
rect 2706 -2562 2712 -2556
rect 2706 -2568 2712 -2562
rect 2706 -2574 2712 -2568
rect 2706 -2580 2712 -2574
rect 2706 -2586 2712 -2580
rect 2706 -2592 2712 -2586
rect 2706 -2598 2712 -2592
rect 2706 -2604 2712 -2598
rect 2706 -2610 2712 -2604
rect 2706 -2616 2712 -2610
rect 2706 -2622 2712 -2616
rect 2706 -2628 2712 -2622
rect 2706 -2634 2712 -2628
rect 2706 -2640 2712 -2634
rect 2706 -2646 2712 -2640
rect 2706 -2652 2712 -2646
rect 2706 -2658 2712 -2652
rect 2706 -2664 2712 -2658
rect 2706 -2670 2712 -2664
rect 2706 -2676 2712 -2670
rect 2706 -2682 2712 -2676
rect 2706 -2688 2712 -2682
rect 2706 -2694 2712 -2688
rect 2712 -1152 2718 -1146
rect 2712 -1158 2718 -1152
rect 2712 -1164 2718 -1158
rect 2712 -1170 2718 -1164
rect 2712 -1176 2718 -1170
rect 2712 -1182 2718 -1176
rect 2712 -1188 2718 -1182
rect 2712 -1194 2718 -1188
rect 2712 -1200 2718 -1194
rect 2712 -1206 2718 -1200
rect 2712 -1212 2718 -1206
rect 2712 -1218 2718 -1212
rect 2712 -1224 2718 -1218
rect 2712 -1230 2718 -1224
rect 2712 -1236 2718 -1230
rect 2712 -1242 2718 -1236
rect 2712 -1248 2718 -1242
rect 2712 -1254 2718 -1248
rect 2712 -1260 2718 -1254
rect 2712 -1266 2718 -1260
rect 2712 -1272 2718 -1266
rect 2712 -1278 2718 -1272
rect 2712 -1284 2718 -1278
rect 2712 -1290 2718 -1284
rect 2712 -1296 2718 -1290
rect 2712 -1302 2718 -1296
rect 2712 -1308 2718 -1302
rect 2712 -1314 2718 -1308
rect 2712 -1320 2718 -1314
rect 2712 -1326 2718 -1320
rect 2712 -1332 2718 -1326
rect 2712 -1338 2718 -1332
rect 2712 -1344 2718 -1338
rect 2712 -1350 2718 -1344
rect 2712 -1356 2718 -1350
rect 2712 -1362 2718 -1356
rect 2712 -1368 2718 -1362
rect 2712 -1374 2718 -1368
rect 2712 -1380 2718 -1374
rect 2712 -1386 2718 -1380
rect 2712 -1392 2718 -1386
rect 2712 -1398 2718 -1392
rect 2712 -1404 2718 -1398
rect 2712 -1410 2718 -1404
rect 2712 -1416 2718 -1410
rect 2712 -1422 2718 -1416
rect 2712 -1428 2718 -1422
rect 2712 -1434 2718 -1428
rect 2712 -1440 2718 -1434
rect 2712 -1446 2718 -1440
rect 2712 -1452 2718 -1446
rect 2712 -1458 2718 -1452
rect 2712 -1464 2718 -1458
rect 2712 -1470 2718 -1464
rect 2712 -1476 2718 -1470
rect 2712 -1482 2718 -1476
rect 2712 -1488 2718 -1482
rect 2712 -1494 2718 -1488
rect 2712 -1500 2718 -1494
rect 2712 -1506 2718 -1500
rect 2712 -1512 2718 -1506
rect 2712 -1518 2718 -1512
rect 2712 -1524 2718 -1518
rect 2712 -1530 2718 -1524
rect 2712 -1536 2718 -1530
rect 2712 -1542 2718 -1536
rect 2712 -1548 2718 -1542
rect 2712 -1554 2718 -1548
rect 2712 -1560 2718 -1554
rect 2712 -1566 2718 -1560
rect 2712 -1572 2718 -1566
rect 2712 -1578 2718 -1572
rect 2712 -1584 2718 -1578
rect 2712 -1590 2718 -1584
rect 2712 -1596 2718 -1590
rect 2712 -1602 2718 -1596
rect 2712 -1608 2718 -1602
rect 2712 -1614 2718 -1608
rect 2712 -1620 2718 -1614
rect 2712 -1626 2718 -1620
rect 2712 -1632 2718 -1626
rect 2712 -1638 2718 -1632
rect 2712 -1644 2718 -1638
rect 2712 -1650 2718 -1644
rect 2712 -1656 2718 -1650
rect 2712 -1662 2718 -1656
rect 2712 -1668 2718 -1662
rect 2712 -1674 2718 -1668
rect 2712 -1680 2718 -1674
rect 2712 -1686 2718 -1680
rect 2712 -1692 2718 -1686
rect 2712 -1698 2718 -1692
rect 2712 -1704 2718 -1698
rect 2712 -1710 2718 -1704
rect 2712 -2394 2718 -2388
rect 2712 -2400 2718 -2394
rect 2712 -2406 2718 -2400
rect 2712 -2412 2718 -2406
rect 2712 -2418 2718 -2412
rect 2712 -2424 2718 -2418
rect 2712 -2430 2718 -2424
rect 2712 -2436 2718 -2430
rect 2712 -2442 2718 -2436
rect 2712 -2448 2718 -2442
rect 2712 -2454 2718 -2448
rect 2712 -2460 2718 -2454
rect 2712 -2466 2718 -2460
rect 2712 -2472 2718 -2466
rect 2712 -2478 2718 -2472
rect 2712 -2484 2718 -2478
rect 2712 -2490 2718 -2484
rect 2712 -2496 2718 -2490
rect 2712 -2502 2718 -2496
rect 2712 -2508 2718 -2502
rect 2712 -2514 2718 -2508
rect 2712 -2520 2718 -2514
rect 2712 -2526 2718 -2520
rect 2712 -2532 2718 -2526
rect 2712 -2538 2718 -2532
rect 2712 -2544 2718 -2538
rect 2712 -2550 2718 -2544
rect 2712 -2556 2718 -2550
rect 2712 -2562 2718 -2556
rect 2712 -2568 2718 -2562
rect 2712 -2574 2718 -2568
rect 2712 -2580 2718 -2574
rect 2712 -2586 2718 -2580
rect 2712 -2592 2718 -2586
rect 2712 -2598 2718 -2592
rect 2712 -2604 2718 -2598
rect 2712 -2610 2718 -2604
rect 2712 -2616 2718 -2610
rect 2712 -2622 2718 -2616
rect 2712 -2628 2718 -2622
rect 2712 -2634 2718 -2628
rect 2712 -2640 2718 -2634
rect 2712 -2646 2718 -2640
rect 2712 -2652 2718 -2646
rect 2712 -2658 2718 -2652
rect 2712 -2664 2718 -2658
rect 2712 -2670 2718 -2664
rect 2712 -2676 2718 -2670
rect 2712 -2682 2718 -2676
rect 2712 -2688 2718 -2682
rect 2718 -1152 2724 -1146
rect 2718 -1158 2724 -1152
rect 2718 -1164 2724 -1158
rect 2718 -1170 2724 -1164
rect 2718 -1176 2724 -1170
rect 2718 -1182 2724 -1176
rect 2718 -1188 2724 -1182
rect 2718 -1194 2724 -1188
rect 2718 -1200 2724 -1194
rect 2718 -1206 2724 -1200
rect 2718 -1212 2724 -1206
rect 2718 -1218 2724 -1212
rect 2718 -1224 2724 -1218
rect 2718 -1230 2724 -1224
rect 2718 -1236 2724 -1230
rect 2718 -1242 2724 -1236
rect 2718 -1248 2724 -1242
rect 2718 -1254 2724 -1248
rect 2718 -1260 2724 -1254
rect 2718 -1266 2724 -1260
rect 2718 -1272 2724 -1266
rect 2718 -1278 2724 -1272
rect 2718 -1284 2724 -1278
rect 2718 -1290 2724 -1284
rect 2718 -1296 2724 -1290
rect 2718 -1302 2724 -1296
rect 2718 -1308 2724 -1302
rect 2718 -1314 2724 -1308
rect 2718 -1320 2724 -1314
rect 2718 -1326 2724 -1320
rect 2718 -1332 2724 -1326
rect 2718 -1338 2724 -1332
rect 2718 -1344 2724 -1338
rect 2718 -1350 2724 -1344
rect 2718 -1356 2724 -1350
rect 2718 -1362 2724 -1356
rect 2718 -1368 2724 -1362
rect 2718 -1374 2724 -1368
rect 2718 -1380 2724 -1374
rect 2718 -1386 2724 -1380
rect 2718 -1392 2724 -1386
rect 2718 -1398 2724 -1392
rect 2718 -1404 2724 -1398
rect 2718 -1410 2724 -1404
rect 2718 -1416 2724 -1410
rect 2718 -1422 2724 -1416
rect 2718 -1428 2724 -1422
rect 2718 -1434 2724 -1428
rect 2718 -1440 2724 -1434
rect 2718 -1446 2724 -1440
rect 2718 -1452 2724 -1446
rect 2718 -1458 2724 -1452
rect 2718 -1464 2724 -1458
rect 2718 -1470 2724 -1464
rect 2718 -1476 2724 -1470
rect 2718 -1482 2724 -1476
rect 2718 -1488 2724 -1482
rect 2718 -1494 2724 -1488
rect 2718 -1500 2724 -1494
rect 2718 -1506 2724 -1500
rect 2718 -1512 2724 -1506
rect 2718 -1518 2724 -1512
rect 2718 -1524 2724 -1518
rect 2718 -1530 2724 -1524
rect 2718 -1536 2724 -1530
rect 2718 -1542 2724 -1536
rect 2718 -1548 2724 -1542
rect 2718 -1554 2724 -1548
rect 2718 -1560 2724 -1554
rect 2718 -1566 2724 -1560
rect 2718 -1572 2724 -1566
rect 2718 -1578 2724 -1572
rect 2718 -1584 2724 -1578
rect 2718 -1590 2724 -1584
rect 2718 -1596 2724 -1590
rect 2718 -1602 2724 -1596
rect 2718 -1608 2724 -1602
rect 2718 -1614 2724 -1608
rect 2718 -1620 2724 -1614
rect 2718 -1626 2724 -1620
rect 2718 -1632 2724 -1626
rect 2718 -1638 2724 -1632
rect 2718 -1644 2724 -1638
rect 2718 -1650 2724 -1644
rect 2718 -1656 2724 -1650
rect 2718 -1662 2724 -1656
rect 2718 -1668 2724 -1662
rect 2718 -1674 2724 -1668
rect 2718 -1680 2724 -1674
rect 2718 -1686 2724 -1680
rect 2718 -1692 2724 -1686
rect 2718 -1698 2724 -1692
rect 2718 -2394 2724 -2388
rect 2718 -2400 2724 -2394
rect 2718 -2406 2724 -2400
rect 2718 -2412 2724 -2406
rect 2718 -2418 2724 -2412
rect 2718 -2424 2724 -2418
rect 2718 -2430 2724 -2424
rect 2718 -2436 2724 -2430
rect 2718 -2442 2724 -2436
rect 2718 -2448 2724 -2442
rect 2718 -2454 2724 -2448
rect 2718 -2460 2724 -2454
rect 2718 -2466 2724 -2460
rect 2718 -2472 2724 -2466
rect 2718 -2478 2724 -2472
rect 2718 -2484 2724 -2478
rect 2718 -2490 2724 -2484
rect 2718 -2496 2724 -2490
rect 2718 -2502 2724 -2496
rect 2718 -2508 2724 -2502
rect 2718 -2514 2724 -2508
rect 2718 -2520 2724 -2514
rect 2718 -2526 2724 -2520
rect 2718 -2532 2724 -2526
rect 2718 -2538 2724 -2532
rect 2718 -2544 2724 -2538
rect 2718 -2550 2724 -2544
rect 2718 -2556 2724 -2550
rect 2718 -2562 2724 -2556
rect 2718 -2568 2724 -2562
rect 2718 -2574 2724 -2568
rect 2718 -2580 2724 -2574
rect 2718 -2586 2724 -2580
rect 2718 -2592 2724 -2586
rect 2718 -2598 2724 -2592
rect 2718 -2604 2724 -2598
rect 2718 -2610 2724 -2604
rect 2718 -2616 2724 -2610
rect 2718 -2622 2724 -2616
rect 2718 -2628 2724 -2622
rect 2718 -2634 2724 -2628
rect 2718 -2640 2724 -2634
rect 2718 -2646 2724 -2640
rect 2718 -2652 2724 -2646
rect 2718 -2658 2724 -2652
rect 2718 -2664 2724 -2658
rect 2718 -2670 2724 -2664
rect 2718 -2676 2724 -2670
rect 2718 -2682 2724 -2676
rect 2724 -1146 2730 -1140
rect 2724 -1152 2730 -1146
rect 2724 -1158 2730 -1152
rect 2724 -1164 2730 -1158
rect 2724 -1170 2730 -1164
rect 2724 -1176 2730 -1170
rect 2724 -1182 2730 -1176
rect 2724 -1188 2730 -1182
rect 2724 -1194 2730 -1188
rect 2724 -1200 2730 -1194
rect 2724 -1206 2730 -1200
rect 2724 -1212 2730 -1206
rect 2724 -1218 2730 -1212
rect 2724 -1224 2730 -1218
rect 2724 -1230 2730 -1224
rect 2724 -1236 2730 -1230
rect 2724 -1242 2730 -1236
rect 2724 -1248 2730 -1242
rect 2724 -1254 2730 -1248
rect 2724 -1260 2730 -1254
rect 2724 -1266 2730 -1260
rect 2724 -1272 2730 -1266
rect 2724 -1278 2730 -1272
rect 2724 -1284 2730 -1278
rect 2724 -1290 2730 -1284
rect 2724 -1296 2730 -1290
rect 2724 -1302 2730 -1296
rect 2724 -1308 2730 -1302
rect 2724 -1314 2730 -1308
rect 2724 -1320 2730 -1314
rect 2724 -1326 2730 -1320
rect 2724 -1332 2730 -1326
rect 2724 -1338 2730 -1332
rect 2724 -1344 2730 -1338
rect 2724 -1350 2730 -1344
rect 2724 -1356 2730 -1350
rect 2724 -1362 2730 -1356
rect 2724 -1368 2730 -1362
rect 2724 -1374 2730 -1368
rect 2724 -1380 2730 -1374
rect 2724 -1386 2730 -1380
rect 2724 -1392 2730 -1386
rect 2724 -1398 2730 -1392
rect 2724 -1404 2730 -1398
rect 2724 -1410 2730 -1404
rect 2724 -1416 2730 -1410
rect 2724 -1422 2730 -1416
rect 2724 -1428 2730 -1422
rect 2724 -1434 2730 -1428
rect 2724 -1440 2730 -1434
rect 2724 -1446 2730 -1440
rect 2724 -1452 2730 -1446
rect 2724 -1458 2730 -1452
rect 2724 -1464 2730 -1458
rect 2724 -1470 2730 -1464
rect 2724 -1476 2730 -1470
rect 2724 -1482 2730 -1476
rect 2724 -1488 2730 -1482
rect 2724 -1494 2730 -1488
rect 2724 -1500 2730 -1494
rect 2724 -1506 2730 -1500
rect 2724 -1512 2730 -1506
rect 2724 -1518 2730 -1512
rect 2724 -1524 2730 -1518
rect 2724 -1530 2730 -1524
rect 2724 -1536 2730 -1530
rect 2724 -1542 2730 -1536
rect 2724 -1548 2730 -1542
rect 2724 -1554 2730 -1548
rect 2724 -1560 2730 -1554
rect 2724 -1566 2730 -1560
rect 2724 -1572 2730 -1566
rect 2724 -1578 2730 -1572
rect 2724 -1584 2730 -1578
rect 2724 -1590 2730 -1584
rect 2724 -1596 2730 -1590
rect 2724 -1602 2730 -1596
rect 2724 -1608 2730 -1602
rect 2724 -1614 2730 -1608
rect 2724 -1620 2730 -1614
rect 2724 -1626 2730 -1620
rect 2724 -1632 2730 -1626
rect 2724 -1638 2730 -1632
rect 2724 -1644 2730 -1638
rect 2724 -1650 2730 -1644
rect 2724 -1656 2730 -1650
rect 2724 -1662 2730 -1656
rect 2724 -1668 2730 -1662
rect 2724 -1674 2730 -1668
rect 2724 -1680 2730 -1674
rect 2724 -1686 2730 -1680
rect 2724 -1692 2730 -1686
rect 2724 -2394 2730 -2388
rect 2724 -2400 2730 -2394
rect 2724 -2406 2730 -2400
rect 2724 -2412 2730 -2406
rect 2724 -2418 2730 -2412
rect 2724 -2424 2730 -2418
rect 2724 -2430 2730 -2424
rect 2724 -2436 2730 -2430
rect 2724 -2442 2730 -2436
rect 2724 -2448 2730 -2442
rect 2724 -2454 2730 -2448
rect 2724 -2460 2730 -2454
rect 2724 -2466 2730 -2460
rect 2724 -2472 2730 -2466
rect 2724 -2478 2730 -2472
rect 2724 -2484 2730 -2478
rect 2724 -2490 2730 -2484
rect 2724 -2496 2730 -2490
rect 2724 -2502 2730 -2496
rect 2724 -2508 2730 -2502
rect 2724 -2514 2730 -2508
rect 2724 -2520 2730 -2514
rect 2724 -2526 2730 -2520
rect 2724 -2532 2730 -2526
rect 2724 -2538 2730 -2532
rect 2724 -2544 2730 -2538
rect 2724 -2550 2730 -2544
rect 2724 -2556 2730 -2550
rect 2724 -2562 2730 -2556
rect 2724 -2568 2730 -2562
rect 2724 -2574 2730 -2568
rect 2724 -2580 2730 -2574
rect 2724 -2586 2730 -2580
rect 2724 -2592 2730 -2586
rect 2724 -2598 2730 -2592
rect 2724 -2604 2730 -2598
rect 2724 -2610 2730 -2604
rect 2724 -2616 2730 -2610
rect 2724 -2622 2730 -2616
rect 2724 -2628 2730 -2622
rect 2724 -2634 2730 -2628
rect 2724 -2640 2730 -2634
rect 2724 -2646 2730 -2640
rect 2724 -2652 2730 -2646
rect 2724 -2658 2730 -2652
rect 2724 -2664 2730 -2658
rect 2724 -2670 2730 -2664
rect 2724 -2676 2730 -2670
rect 2724 -2682 2730 -2676
rect 2730 -1140 2736 -1134
rect 2730 -1146 2736 -1140
rect 2730 -1152 2736 -1146
rect 2730 -1158 2736 -1152
rect 2730 -1164 2736 -1158
rect 2730 -1170 2736 -1164
rect 2730 -1176 2736 -1170
rect 2730 -1182 2736 -1176
rect 2730 -1188 2736 -1182
rect 2730 -1194 2736 -1188
rect 2730 -1200 2736 -1194
rect 2730 -1206 2736 -1200
rect 2730 -1212 2736 -1206
rect 2730 -1218 2736 -1212
rect 2730 -1224 2736 -1218
rect 2730 -1230 2736 -1224
rect 2730 -1236 2736 -1230
rect 2730 -1242 2736 -1236
rect 2730 -1248 2736 -1242
rect 2730 -1254 2736 -1248
rect 2730 -1260 2736 -1254
rect 2730 -1266 2736 -1260
rect 2730 -1272 2736 -1266
rect 2730 -1278 2736 -1272
rect 2730 -1284 2736 -1278
rect 2730 -1290 2736 -1284
rect 2730 -1296 2736 -1290
rect 2730 -1302 2736 -1296
rect 2730 -1308 2736 -1302
rect 2730 -1314 2736 -1308
rect 2730 -1320 2736 -1314
rect 2730 -1326 2736 -1320
rect 2730 -1332 2736 -1326
rect 2730 -1338 2736 -1332
rect 2730 -1344 2736 -1338
rect 2730 -1350 2736 -1344
rect 2730 -1356 2736 -1350
rect 2730 -1362 2736 -1356
rect 2730 -1368 2736 -1362
rect 2730 -1374 2736 -1368
rect 2730 -1380 2736 -1374
rect 2730 -1386 2736 -1380
rect 2730 -1392 2736 -1386
rect 2730 -1398 2736 -1392
rect 2730 -1404 2736 -1398
rect 2730 -1410 2736 -1404
rect 2730 -1416 2736 -1410
rect 2730 -1422 2736 -1416
rect 2730 -1428 2736 -1422
rect 2730 -1434 2736 -1428
rect 2730 -1440 2736 -1434
rect 2730 -1446 2736 -1440
rect 2730 -1452 2736 -1446
rect 2730 -1458 2736 -1452
rect 2730 -1464 2736 -1458
rect 2730 -1470 2736 -1464
rect 2730 -1476 2736 -1470
rect 2730 -1482 2736 -1476
rect 2730 -1488 2736 -1482
rect 2730 -1494 2736 -1488
rect 2730 -1500 2736 -1494
rect 2730 -1506 2736 -1500
rect 2730 -1512 2736 -1506
rect 2730 -1518 2736 -1512
rect 2730 -1524 2736 -1518
rect 2730 -1530 2736 -1524
rect 2730 -1536 2736 -1530
rect 2730 -1542 2736 -1536
rect 2730 -1548 2736 -1542
rect 2730 -1554 2736 -1548
rect 2730 -1560 2736 -1554
rect 2730 -1566 2736 -1560
rect 2730 -1572 2736 -1566
rect 2730 -1578 2736 -1572
rect 2730 -1584 2736 -1578
rect 2730 -1590 2736 -1584
rect 2730 -1596 2736 -1590
rect 2730 -1602 2736 -1596
rect 2730 -1608 2736 -1602
rect 2730 -1614 2736 -1608
rect 2730 -1620 2736 -1614
rect 2730 -1626 2736 -1620
rect 2730 -1632 2736 -1626
rect 2730 -1638 2736 -1632
rect 2730 -1644 2736 -1638
rect 2730 -1650 2736 -1644
rect 2730 -1656 2736 -1650
rect 2730 -1662 2736 -1656
rect 2730 -1668 2736 -1662
rect 2730 -1674 2736 -1668
rect 2730 -1680 2736 -1674
rect 2730 -2388 2736 -2382
rect 2730 -2394 2736 -2388
rect 2730 -2400 2736 -2394
rect 2730 -2406 2736 -2400
rect 2730 -2412 2736 -2406
rect 2730 -2418 2736 -2412
rect 2730 -2424 2736 -2418
rect 2730 -2430 2736 -2424
rect 2730 -2436 2736 -2430
rect 2730 -2442 2736 -2436
rect 2730 -2448 2736 -2442
rect 2730 -2454 2736 -2448
rect 2730 -2460 2736 -2454
rect 2730 -2466 2736 -2460
rect 2730 -2472 2736 -2466
rect 2730 -2478 2736 -2472
rect 2730 -2484 2736 -2478
rect 2730 -2490 2736 -2484
rect 2730 -2496 2736 -2490
rect 2730 -2502 2736 -2496
rect 2730 -2508 2736 -2502
rect 2730 -2514 2736 -2508
rect 2730 -2520 2736 -2514
rect 2730 -2526 2736 -2520
rect 2730 -2532 2736 -2526
rect 2730 -2538 2736 -2532
rect 2730 -2544 2736 -2538
rect 2730 -2550 2736 -2544
rect 2730 -2556 2736 -2550
rect 2730 -2562 2736 -2556
rect 2730 -2568 2736 -2562
rect 2730 -2574 2736 -2568
rect 2730 -2580 2736 -2574
rect 2730 -2586 2736 -2580
rect 2730 -2592 2736 -2586
rect 2730 -2598 2736 -2592
rect 2730 -2604 2736 -2598
rect 2730 -2610 2736 -2604
rect 2730 -2616 2736 -2610
rect 2730 -2622 2736 -2616
rect 2730 -2628 2736 -2622
rect 2730 -2634 2736 -2628
rect 2730 -2640 2736 -2634
rect 2730 -2646 2736 -2640
rect 2730 -2652 2736 -2646
rect 2730 -2658 2736 -2652
rect 2730 -2664 2736 -2658
rect 2730 -2670 2736 -2664
rect 2730 -2676 2736 -2670
rect 2736 -1140 2742 -1134
rect 2736 -1146 2742 -1140
rect 2736 -1152 2742 -1146
rect 2736 -1158 2742 -1152
rect 2736 -1164 2742 -1158
rect 2736 -1170 2742 -1164
rect 2736 -1176 2742 -1170
rect 2736 -1182 2742 -1176
rect 2736 -1188 2742 -1182
rect 2736 -1194 2742 -1188
rect 2736 -1200 2742 -1194
rect 2736 -1206 2742 -1200
rect 2736 -1212 2742 -1206
rect 2736 -1218 2742 -1212
rect 2736 -1224 2742 -1218
rect 2736 -1230 2742 -1224
rect 2736 -1236 2742 -1230
rect 2736 -1242 2742 -1236
rect 2736 -1248 2742 -1242
rect 2736 -1254 2742 -1248
rect 2736 -1260 2742 -1254
rect 2736 -1266 2742 -1260
rect 2736 -1272 2742 -1266
rect 2736 -1278 2742 -1272
rect 2736 -1284 2742 -1278
rect 2736 -1290 2742 -1284
rect 2736 -1296 2742 -1290
rect 2736 -1302 2742 -1296
rect 2736 -1308 2742 -1302
rect 2736 -1314 2742 -1308
rect 2736 -1320 2742 -1314
rect 2736 -1326 2742 -1320
rect 2736 -1332 2742 -1326
rect 2736 -1338 2742 -1332
rect 2736 -1344 2742 -1338
rect 2736 -1350 2742 -1344
rect 2736 -1356 2742 -1350
rect 2736 -1362 2742 -1356
rect 2736 -1368 2742 -1362
rect 2736 -1374 2742 -1368
rect 2736 -1380 2742 -1374
rect 2736 -1386 2742 -1380
rect 2736 -1392 2742 -1386
rect 2736 -1398 2742 -1392
rect 2736 -1404 2742 -1398
rect 2736 -1410 2742 -1404
rect 2736 -1416 2742 -1410
rect 2736 -1422 2742 -1416
rect 2736 -1428 2742 -1422
rect 2736 -1434 2742 -1428
rect 2736 -1440 2742 -1434
rect 2736 -1446 2742 -1440
rect 2736 -1452 2742 -1446
rect 2736 -1458 2742 -1452
rect 2736 -1464 2742 -1458
rect 2736 -1470 2742 -1464
rect 2736 -1476 2742 -1470
rect 2736 -1482 2742 -1476
rect 2736 -1488 2742 -1482
rect 2736 -1494 2742 -1488
rect 2736 -1500 2742 -1494
rect 2736 -1506 2742 -1500
rect 2736 -1512 2742 -1506
rect 2736 -1518 2742 -1512
rect 2736 -1524 2742 -1518
rect 2736 -1530 2742 -1524
rect 2736 -1536 2742 -1530
rect 2736 -1542 2742 -1536
rect 2736 -1548 2742 -1542
rect 2736 -1554 2742 -1548
rect 2736 -1560 2742 -1554
rect 2736 -1566 2742 -1560
rect 2736 -1572 2742 -1566
rect 2736 -1578 2742 -1572
rect 2736 -1584 2742 -1578
rect 2736 -1590 2742 -1584
rect 2736 -1596 2742 -1590
rect 2736 -1602 2742 -1596
rect 2736 -1608 2742 -1602
rect 2736 -1614 2742 -1608
rect 2736 -1620 2742 -1614
rect 2736 -1626 2742 -1620
rect 2736 -1632 2742 -1626
rect 2736 -1638 2742 -1632
rect 2736 -1644 2742 -1638
rect 2736 -1650 2742 -1644
rect 2736 -1656 2742 -1650
rect 2736 -1662 2742 -1656
rect 2736 -1668 2742 -1662
rect 2736 -1674 2742 -1668
rect 2736 -2388 2742 -2382
rect 2736 -2394 2742 -2388
rect 2736 -2400 2742 -2394
rect 2736 -2406 2742 -2400
rect 2736 -2412 2742 -2406
rect 2736 -2418 2742 -2412
rect 2736 -2424 2742 -2418
rect 2736 -2430 2742 -2424
rect 2736 -2436 2742 -2430
rect 2736 -2442 2742 -2436
rect 2736 -2448 2742 -2442
rect 2736 -2454 2742 -2448
rect 2736 -2460 2742 -2454
rect 2736 -2466 2742 -2460
rect 2736 -2472 2742 -2466
rect 2736 -2478 2742 -2472
rect 2736 -2484 2742 -2478
rect 2736 -2490 2742 -2484
rect 2736 -2496 2742 -2490
rect 2736 -2502 2742 -2496
rect 2736 -2508 2742 -2502
rect 2736 -2514 2742 -2508
rect 2736 -2520 2742 -2514
rect 2736 -2526 2742 -2520
rect 2736 -2532 2742 -2526
rect 2736 -2538 2742 -2532
rect 2736 -2544 2742 -2538
rect 2736 -2550 2742 -2544
rect 2736 -2556 2742 -2550
rect 2736 -2562 2742 -2556
rect 2736 -2568 2742 -2562
rect 2736 -2574 2742 -2568
rect 2736 -2580 2742 -2574
rect 2736 -2586 2742 -2580
rect 2736 -2592 2742 -2586
rect 2736 -2598 2742 -2592
rect 2736 -2604 2742 -2598
rect 2736 -2610 2742 -2604
rect 2736 -2616 2742 -2610
rect 2736 -2622 2742 -2616
rect 2736 -2628 2742 -2622
rect 2736 -2634 2742 -2628
rect 2736 -2640 2742 -2634
rect 2736 -2646 2742 -2640
rect 2736 -2652 2742 -2646
rect 2736 -2658 2742 -2652
rect 2736 -2664 2742 -2658
rect 2736 -2670 2742 -2664
rect 2742 -1134 2748 -1128
rect 2742 -1140 2748 -1134
rect 2742 -1146 2748 -1140
rect 2742 -1152 2748 -1146
rect 2742 -1158 2748 -1152
rect 2742 -1164 2748 -1158
rect 2742 -1170 2748 -1164
rect 2742 -1176 2748 -1170
rect 2742 -1182 2748 -1176
rect 2742 -1188 2748 -1182
rect 2742 -1194 2748 -1188
rect 2742 -1200 2748 -1194
rect 2742 -1206 2748 -1200
rect 2742 -1212 2748 -1206
rect 2742 -1218 2748 -1212
rect 2742 -1224 2748 -1218
rect 2742 -1230 2748 -1224
rect 2742 -1236 2748 -1230
rect 2742 -1242 2748 -1236
rect 2742 -1248 2748 -1242
rect 2742 -1254 2748 -1248
rect 2742 -1260 2748 -1254
rect 2742 -1266 2748 -1260
rect 2742 -1272 2748 -1266
rect 2742 -1278 2748 -1272
rect 2742 -1284 2748 -1278
rect 2742 -1290 2748 -1284
rect 2742 -1296 2748 -1290
rect 2742 -1302 2748 -1296
rect 2742 -1308 2748 -1302
rect 2742 -1314 2748 -1308
rect 2742 -1320 2748 -1314
rect 2742 -1326 2748 -1320
rect 2742 -1332 2748 -1326
rect 2742 -1338 2748 -1332
rect 2742 -1344 2748 -1338
rect 2742 -1350 2748 -1344
rect 2742 -1356 2748 -1350
rect 2742 -1362 2748 -1356
rect 2742 -1368 2748 -1362
rect 2742 -1374 2748 -1368
rect 2742 -1380 2748 -1374
rect 2742 -1386 2748 -1380
rect 2742 -1392 2748 -1386
rect 2742 -1398 2748 -1392
rect 2742 -1404 2748 -1398
rect 2742 -1410 2748 -1404
rect 2742 -1416 2748 -1410
rect 2742 -1422 2748 -1416
rect 2742 -1428 2748 -1422
rect 2742 -1434 2748 -1428
rect 2742 -1440 2748 -1434
rect 2742 -1446 2748 -1440
rect 2742 -1452 2748 -1446
rect 2742 -1458 2748 -1452
rect 2742 -1464 2748 -1458
rect 2742 -1470 2748 -1464
rect 2742 -1476 2748 -1470
rect 2742 -1482 2748 -1476
rect 2742 -1488 2748 -1482
rect 2742 -1494 2748 -1488
rect 2742 -1500 2748 -1494
rect 2742 -1506 2748 -1500
rect 2742 -1512 2748 -1506
rect 2742 -1518 2748 -1512
rect 2742 -1524 2748 -1518
rect 2742 -1530 2748 -1524
rect 2742 -1536 2748 -1530
rect 2742 -1542 2748 -1536
rect 2742 -1548 2748 -1542
rect 2742 -1554 2748 -1548
rect 2742 -1560 2748 -1554
rect 2742 -1566 2748 -1560
rect 2742 -1572 2748 -1566
rect 2742 -1578 2748 -1572
rect 2742 -1584 2748 -1578
rect 2742 -1590 2748 -1584
rect 2742 -1596 2748 -1590
rect 2742 -1602 2748 -1596
rect 2742 -1608 2748 -1602
rect 2742 -1614 2748 -1608
rect 2742 -1620 2748 -1614
rect 2742 -1626 2748 -1620
rect 2742 -1632 2748 -1626
rect 2742 -1638 2748 -1632
rect 2742 -1644 2748 -1638
rect 2742 -1650 2748 -1644
rect 2742 -1656 2748 -1650
rect 2742 -1662 2748 -1656
rect 2742 -1668 2748 -1662
rect 2742 -2388 2748 -2382
rect 2742 -2394 2748 -2388
rect 2742 -2400 2748 -2394
rect 2742 -2406 2748 -2400
rect 2742 -2412 2748 -2406
rect 2742 -2418 2748 -2412
rect 2742 -2424 2748 -2418
rect 2742 -2430 2748 -2424
rect 2742 -2436 2748 -2430
rect 2742 -2442 2748 -2436
rect 2742 -2448 2748 -2442
rect 2742 -2454 2748 -2448
rect 2742 -2460 2748 -2454
rect 2742 -2466 2748 -2460
rect 2742 -2472 2748 -2466
rect 2742 -2478 2748 -2472
rect 2742 -2484 2748 -2478
rect 2742 -2490 2748 -2484
rect 2742 -2496 2748 -2490
rect 2742 -2502 2748 -2496
rect 2742 -2508 2748 -2502
rect 2742 -2514 2748 -2508
rect 2742 -2520 2748 -2514
rect 2742 -2526 2748 -2520
rect 2742 -2532 2748 -2526
rect 2742 -2538 2748 -2532
rect 2742 -2544 2748 -2538
rect 2742 -2550 2748 -2544
rect 2742 -2556 2748 -2550
rect 2742 -2562 2748 -2556
rect 2742 -2568 2748 -2562
rect 2742 -2574 2748 -2568
rect 2742 -2580 2748 -2574
rect 2742 -2586 2748 -2580
rect 2742 -2592 2748 -2586
rect 2742 -2598 2748 -2592
rect 2742 -2604 2748 -2598
rect 2742 -2610 2748 -2604
rect 2742 -2616 2748 -2610
rect 2742 -2622 2748 -2616
rect 2742 -2628 2748 -2622
rect 2742 -2634 2748 -2628
rect 2742 -2640 2748 -2634
rect 2742 -2646 2748 -2640
rect 2742 -2652 2748 -2646
rect 2742 -2658 2748 -2652
rect 2742 -2664 2748 -2658
rect 2748 -1128 2754 -1122
rect 2748 -1134 2754 -1128
rect 2748 -1140 2754 -1134
rect 2748 -1146 2754 -1140
rect 2748 -1152 2754 -1146
rect 2748 -1158 2754 -1152
rect 2748 -1164 2754 -1158
rect 2748 -1170 2754 -1164
rect 2748 -1176 2754 -1170
rect 2748 -1182 2754 -1176
rect 2748 -1188 2754 -1182
rect 2748 -1194 2754 -1188
rect 2748 -1200 2754 -1194
rect 2748 -1206 2754 -1200
rect 2748 -1212 2754 -1206
rect 2748 -1218 2754 -1212
rect 2748 -1224 2754 -1218
rect 2748 -1230 2754 -1224
rect 2748 -1236 2754 -1230
rect 2748 -1242 2754 -1236
rect 2748 -1248 2754 -1242
rect 2748 -1254 2754 -1248
rect 2748 -1260 2754 -1254
rect 2748 -1266 2754 -1260
rect 2748 -1272 2754 -1266
rect 2748 -1278 2754 -1272
rect 2748 -1284 2754 -1278
rect 2748 -1290 2754 -1284
rect 2748 -1296 2754 -1290
rect 2748 -1302 2754 -1296
rect 2748 -1308 2754 -1302
rect 2748 -1314 2754 -1308
rect 2748 -1320 2754 -1314
rect 2748 -1326 2754 -1320
rect 2748 -1332 2754 -1326
rect 2748 -1338 2754 -1332
rect 2748 -1344 2754 -1338
rect 2748 -1350 2754 -1344
rect 2748 -1356 2754 -1350
rect 2748 -1362 2754 -1356
rect 2748 -1368 2754 -1362
rect 2748 -1374 2754 -1368
rect 2748 -1380 2754 -1374
rect 2748 -1386 2754 -1380
rect 2748 -1392 2754 -1386
rect 2748 -1398 2754 -1392
rect 2748 -1404 2754 -1398
rect 2748 -1410 2754 -1404
rect 2748 -1416 2754 -1410
rect 2748 -1422 2754 -1416
rect 2748 -1428 2754 -1422
rect 2748 -1434 2754 -1428
rect 2748 -1440 2754 -1434
rect 2748 -1446 2754 -1440
rect 2748 -1452 2754 -1446
rect 2748 -1458 2754 -1452
rect 2748 -1464 2754 -1458
rect 2748 -1470 2754 -1464
rect 2748 -1476 2754 -1470
rect 2748 -1482 2754 -1476
rect 2748 -1488 2754 -1482
rect 2748 -1494 2754 -1488
rect 2748 -1500 2754 -1494
rect 2748 -1506 2754 -1500
rect 2748 -1512 2754 -1506
rect 2748 -1518 2754 -1512
rect 2748 -1524 2754 -1518
rect 2748 -1530 2754 -1524
rect 2748 -1536 2754 -1530
rect 2748 -1542 2754 -1536
rect 2748 -1548 2754 -1542
rect 2748 -1554 2754 -1548
rect 2748 -1560 2754 -1554
rect 2748 -1566 2754 -1560
rect 2748 -1572 2754 -1566
rect 2748 -1578 2754 -1572
rect 2748 -1584 2754 -1578
rect 2748 -1590 2754 -1584
rect 2748 -1596 2754 -1590
rect 2748 -1602 2754 -1596
rect 2748 -1608 2754 -1602
rect 2748 -1614 2754 -1608
rect 2748 -1620 2754 -1614
rect 2748 -1626 2754 -1620
rect 2748 -1632 2754 -1626
rect 2748 -1638 2754 -1632
rect 2748 -1644 2754 -1638
rect 2748 -1650 2754 -1644
rect 2748 -1656 2754 -1650
rect 2748 -2388 2754 -2382
rect 2748 -2394 2754 -2388
rect 2748 -2400 2754 -2394
rect 2748 -2406 2754 -2400
rect 2748 -2412 2754 -2406
rect 2748 -2418 2754 -2412
rect 2748 -2424 2754 -2418
rect 2748 -2430 2754 -2424
rect 2748 -2436 2754 -2430
rect 2748 -2442 2754 -2436
rect 2748 -2448 2754 -2442
rect 2748 -2454 2754 -2448
rect 2748 -2460 2754 -2454
rect 2748 -2466 2754 -2460
rect 2748 -2472 2754 -2466
rect 2748 -2478 2754 -2472
rect 2748 -2484 2754 -2478
rect 2748 -2490 2754 -2484
rect 2748 -2496 2754 -2490
rect 2748 -2502 2754 -2496
rect 2748 -2508 2754 -2502
rect 2748 -2514 2754 -2508
rect 2748 -2520 2754 -2514
rect 2748 -2526 2754 -2520
rect 2748 -2532 2754 -2526
rect 2748 -2538 2754 -2532
rect 2748 -2544 2754 -2538
rect 2748 -2550 2754 -2544
rect 2748 -2556 2754 -2550
rect 2748 -2562 2754 -2556
rect 2748 -2568 2754 -2562
rect 2748 -2574 2754 -2568
rect 2748 -2580 2754 -2574
rect 2748 -2586 2754 -2580
rect 2748 -2592 2754 -2586
rect 2748 -2598 2754 -2592
rect 2748 -2604 2754 -2598
rect 2748 -2610 2754 -2604
rect 2748 -2616 2754 -2610
rect 2748 -2622 2754 -2616
rect 2748 -2628 2754 -2622
rect 2748 -2634 2754 -2628
rect 2748 -2640 2754 -2634
rect 2748 -2646 2754 -2640
rect 2748 -2652 2754 -2646
rect 2748 -2658 2754 -2652
rect 2748 -2664 2754 -2658
rect 2754 -1128 2760 -1122
rect 2754 -1134 2760 -1128
rect 2754 -1140 2760 -1134
rect 2754 -1146 2760 -1140
rect 2754 -1152 2760 -1146
rect 2754 -1158 2760 -1152
rect 2754 -1164 2760 -1158
rect 2754 -1170 2760 -1164
rect 2754 -1176 2760 -1170
rect 2754 -1182 2760 -1176
rect 2754 -1188 2760 -1182
rect 2754 -1194 2760 -1188
rect 2754 -1200 2760 -1194
rect 2754 -1206 2760 -1200
rect 2754 -1212 2760 -1206
rect 2754 -1218 2760 -1212
rect 2754 -1224 2760 -1218
rect 2754 -1230 2760 -1224
rect 2754 -1236 2760 -1230
rect 2754 -1242 2760 -1236
rect 2754 -1248 2760 -1242
rect 2754 -1254 2760 -1248
rect 2754 -1260 2760 -1254
rect 2754 -1266 2760 -1260
rect 2754 -1272 2760 -1266
rect 2754 -1278 2760 -1272
rect 2754 -1284 2760 -1278
rect 2754 -1290 2760 -1284
rect 2754 -1296 2760 -1290
rect 2754 -1302 2760 -1296
rect 2754 -1308 2760 -1302
rect 2754 -1314 2760 -1308
rect 2754 -1320 2760 -1314
rect 2754 -1326 2760 -1320
rect 2754 -1332 2760 -1326
rect 2754 -1338 2760 -1332
rect 2754 -1344 2760 -1338
rect 2754 -1350 2760 -1344
rect 2754 -1356 2760 -1350
rect 2754 -1362 2760 -1356
rect 2754 -1368 2760 -1362
rect 2754 -1374 2760 -1368
rect 2754 -1380 2760 -1374
rect 2754 -1386 2760 -1380
rect 2754 -1392 2760 -1386
rect 2754 -1398 2760 -1392
rect 2754 -1404 2760 -1398
rect 2754 -1410 2760 -1404
rect 2754 -1416 2760 -1410
rect 2754 -1422 2760 -1416
rect 2754 -1428 2760 -1422
rect 2754 -1434 2760 -1428
rect 2754 -1440 2760 -1434
rect 2754 -1446 2760 -1440
rect 2754 -1452 2760 -1446
rect 2754 -1458 2760 -1452
rect 2754 -1464 2760 -1458
rect 2754 -1470 2760 -1464
rect 2754 -1476 2760 -1470
rect 2754 -1482 2760 -1476
rect 2754 -1488 2760 -1482
rect 2754 -1494 2760 -1488
rect 2754 -1500 2760 -1494
rect 2754 -1506 2760 -1500
rect 2754 -1512 2760 -1506
rect 2754 -1518 2760 -1512
rect 2754 -1524 2760 -1518
rect 2754 -1530 2760 -1524
rect 2754 -1536 2760 -1530
rect 2754 -1542 2760 -1536
rect 2754 -1548 2760 -1542
rect 2754 -1554 2760 -1548
rect 2754 -1560 2760 -1554
rect 2754 -1566 2760 -1560
rect 2754 -1572 2760 -1566
rect 2754 -1578 2760 -1572
rect 2754 -1584 2760 -1578
rect 2754 -1590 2760 -1584
rect 2754 -1596 2760 -1590
rect 2754 -1602 2760 -1596
rect 2754 -1608 2760 -1602
rect 2754 -1614 2760 -1608
rect 2754 -1620 2760 -1614
rect 2754 -1626 2760 -1620
rect 2754 -1632 2760 -1626
rect 2754 -1638 2760 -1632
rect 2754 -1644 2760 -1638
rect 2754 -1650 2760 -1644
rect 2754 -2382 2760 -2376
rect 2754 -2388 2760 -2382
rect 2754 -2394 2760 -2388
rect 2754 -2400 2760 -2394
rect 2754 -2406 2760 -2400
rect 2754 -2412 2760 -2406
rect 2754 -2418 2760 -2412
rect 2754 -2424 2760 -2418
rect 2754 -2430 2760 -2424
rect 2754 -2436 2760 -2430
rect 2754 -2442 2760 -2436
rect 2754 -2448 2760 -2442
rect 2754 -2454 2760 -2448
rect 2754 -2460 2760 -2454
rect 2754 -2466 2760 -2460
rect 2754 -2472 2760 -2466
rect 2754 -2478 2760 -2472
rect 2754 -2484 2760 -2478
rect 2754 -2490 2760 -2484
rect 2754 -2496 2760 -2490
rect 2754 -2502 2760 -2496
rect 2754 -2508 2760 -2502
rect 2754 -2514 2760 -2508
rect 2754 -2520 2760 -2514
rect 2754 -2526 2760 -2520
rect 2754 -2532 2760 -2526
rect 2754 -2538 2760 -2532
rect 2754 -2544 2760 -2538
rect 2754 -2550 2760 -2544
rect 2754 -2556 2760 -2550
rect 2754 -2562 2760 -2556
rect 2754 -2568 2760 -2562
rect 2754 -2574 2760 -2568
rect 2754 -2580 2760 -2574
rect 2754 -2586 2760 -2580
rect 2754 -2592 2760 -2586
rect 2754 -2598 2760 -2592
rect 2754 -2604 2760 -2598
rect 2754 -2610 2760 -2604
rect 2754 -2616 2760 -2610
rect 2754 -2622 2760 -2616
rect 2754 -2628 2760 -2622
rect 2754 -2634 2760 -2628
rect 2754 -2640 2760 -2634
rect 2754 -2646 2760 -2640
rect 2754 -2652 2760 -2646
rect 2754 -2658 2760 -2652
rect 2760 -1122 2766 -1116
rect 2760 -1128 2766 -1122
rect 2760 -1134 2766 -1128
rect 2760 -1140 2766 -1134
rect 2760 -1146 2766 -1140
rect 2760 -1152 2766 -1146
rect 2760 -1158 2766 -1152
rect 2760 -1164 2766 -1158
rect 2760 -1170 2766 -1164
rect 2760 -1176 2766 -1170
rect 2760 -1182 2766 -1176
rect 2760 -1188 2766 -1182
rect 2760 -1194 2766 -1188
rect 2760 -1200 2766 -1194
rect 2760 -1206 2766 -1200
rect 2760 -1212 2766 -1206
rect 2760 -1218 2766 -1212
rect 2760 -1224 2766 -1218
rect 2760 -1230 2766 -1224
rect 2760 -1236 2766 -1230
rect 2760 -1242 2766 -1236
rect 2760 -1248 2766 -1242
rect 2760 -1254 2766 -1248
rect 2760 -1260 2766 -1254
rect 2760 -1266 2766 -1260
rect 2760 -1272 2766 -1266
rect 2760 -1278 2766 -1272
rect 2760 -1284 2766 -1278
rect 2760 -1290 2766 -1284
rect 2760 -1296 2766 -1290
rect 2760 -1302 2766 -1296
rect 2760 -1308 2766 -1302
rect 2760 -1314 2766 -1308
rect 2760 -1320 2766 -1314
rect 2760 -1326 2766 -1320
rect 2760 -1332 2766 -1326
rect 2760 -1338 2766 -1332
rect 2760 -1344 2766 -1338
rect 2760 -1350 2766 -1344
rect 2760 -1356 2766 -1350
rect 2760 -1362 2766 -1356
rect 2760 -1368 2766 -1362
rect 2760 -1374 2766 -1368
rect 2760 -1380 2766 -1374
rect 2760 -1386 2766 -1380
rect 2760 -1392 2766 -1386
rect 2760 -1398 2766 -1392
rect 2760 -1404 2766 -1398
rect 2760 -1410 2766 -1404
rect 2760 -1416 2766 -1410
rect 2760 -1422 2766 -1416
rect 2760 -1428 2766 -1422
rect 2760 -1434 2766 -1428
rect 2760 -1440 2766 -1434
rect 2760 -1446 2766 -1440
rect 2760 -1452 2766 -1446
rect 2760 -1458 2766 -1452
rect 2760 -1464 2766 -1458
rect 2760 -1470 2766 -1464
rect 2760 -1476 2766 -1470
rect 2760 -1482 2766 -1476
rect 2760 -1488 2766 -1482
rect 2760 -1494 2766 -1488
rect 2760 -1500 2766 -1494
rect 2760 -1506 2766 -1500
rect 2760 -1512 2766 -1506
rect 2760 -1518 2766 -1512
rect 2760 -1524 2766 -1518
rect 2760 -1530 2766 -1524
rect 2760 -1536 2766 -1530
rect 2760 -1542 2766 -1536
rect 2760 -1548 2766 -1542
rect 2760 -1554 2766 -1548
rect 2760 -1560 2766 -1554
rect 2760 -1566 2766 -1560
rect 2760 -1572 2766 -1566
rect 2760 -1578 2766 -1572
rect 2760 -1584 2766 -1578
rect 2760 -1590 2766 -1584
rect 2760 -1596 2766 -1590
rect 2760 -1602 2766 -1596
rect 2760 -1608 2766 -1602
rect 2760 -1614 2766 -1608
rect 2760 -1620 2766 -1614
rect 2760 -1626 2766 -1620
rect 2760 -1632 2766 -1626
rect 2760 -1638 2766 -1632
rect 2760 -2382 2766 -2376
rect 2760 -2388 2766 -2382
rect 2760 -2394 2766 -2388
rect 2760 -2400 2766 -2394
rect 2760 -2406 2766 -2400
rect 2760 -2412 2766 -2406
rect 2760 -2418 2766 -2412
rect 2760 -2424 2766 -2418
rect 2760 -2430 2766 -2424
rect 2760 -2436 2766 -2430
rect 2760 -2442 2766 -2436
rect 2760 -2448 2766 -2442
rect 2760 -2454 2766 -2448
rect 2760 -2460 2766 -2454
rect 2760 -2466 2766 -2460
rect 2760 -2472 2766 -2466
rect 2760 -2478 2766 -2472
rect 2760 -2484 2766 -2478
rect 2760 -2490 2766 -2484
rect 2760 -2496 2766 -2490
rect 2760 -2502 2766 -2496
rect 2760 -2508 2766 -2502
rect 2760 -2514 2766 -2508
rect 2760 -2520 2766 -2514
rect 2760 -2526 2766 -2520
rect 2760 -2532 2766 -2526
rect 2760 -2538 2766 -2532
rect 2760 -2544 2766 -2538
rect 2760 -2550 2766 -2544
rect 2760 -2556 2766 -2550
rect 2760 -2562 2766 -2556
rect 2760 -2568 2766 -2562
rect 2760 -2574 2766 -2568
rect 2760 -2580 2766 -2574
rect 2760 -2586 2766 -2580
rect 2760 -2592 2766 -2586
rect 2760 -2598 2766 -2592
rect 2760 -2604 2766 -2598
rect 2760 -2610 2766 -2604
rect 2760 -2616 2766 -2610
rect 2760 -2622 2766 -2616
rect 2760 -2628 2766 -2622
rect 2760 -2634 2766 -2628
rect 2760 -2640 2766 -2634
rect 2760 -2646 2766 -2640
rect 2760 -2652 2766 -2646
rect 2766 -1116 2772 -1110
rect 2766 -1122 2772 -1116
rect 2766 -1128 2772 -1122
rect 2766 -1134 2772 -1128
rect 2766 -1140 2772 -1134
rect 2766 -1146 2772 -1140
rect 2766 -1152 2772 -1146
rect 2766 -1158 2772 -1152
rect 2766 -1164 2772 -1158
rect 2766 -1170 2772 -1164
rect 2766 -1176 2772 -1170
rect 2766 -1182 2772 -1176
rect 2766 -1188 2772 -1182
rect 2766 -1194 2772 -1188
rect 2766 -1200 2772 -1194
rect 2766 -1206 2772 -1200
rect 2766 -1212 2772 -1206
rect 2766 -1218 2772 -1212
rect 2766 -1224 2772 -1218
rect 2766 -1230 2772 -1224
rect 2766 -1236 2772 -1230
rect 2766 -1242 2772 -1236
rect 2766 -1248 2772 -1242
rect 2766 -1254 2772 -1248
rect 2766 -1260 2772 -1254
rect 2766 -1266 2772 -1260
rect 2766 -1272 2772 -1266
rect 2766 -1278 2772 -1272
rect 2766 -1284 2772 -1278
rect 2766 -1290 2772 -1284
rect 2766 -1296 2772 -1290
rect 2766 -1302 2772 -1296
rect 2766 -1308 2772 -1302
rect 2766 -1314 2772 -1308
rect 2766 -1320 2772 -1314
rect 2766 -1326 2772 -1320
rect 2766 -1332 2772 -1326
rect 2766 -1338 2772 -1332
rect 2766 -1344 2772 -1338
rect 2766 -1350 2772 -1344
rect 2766 -1356 2772 -1350
rect 2766 -1362 2772 -1356
rect 2766 -1368 2772 -1362
rect 2766 -1374 2772 -1368
rect 2766 -1380 2772 -1374
rect 2766 -1386 2772 -1380
rect 2766 -1392 2772 -1386
rect 2766 -1398 2772 -1392
rect 2766 -1404 2772 -1398
rect 2766 -1410 2772 -1404
rect 2766 -1416 2772 -1410
rect 2766 -1422 2772 -1416
rect 2766 -1428 2772 -1422
rect 2766 -1434 2772 -1428
rect 2766 -1440 2772 -1434
rect 2766 -1446 2772 -1440
rect 2766 -1452 2772 -1446
rect 2766 -1458 2772 -1452
rect 2766 -1464 2772 -1458
rect 2766 -1470 2772 -1464
rect 2766 -1476 2772 -1470
rect 2766 -1482 2772 -1476
rect 2766 -1488 2772 -1482
rect 2766 -1494 2772 -1488
rect 2766 -1500 2772 -1494
rect 2766 -1506 2772 -1500
rect 2766 -1512 2772 -1506
rect 2766 -1518 2772 -1512
rect 2766 -1524 2772 -1518
rect 2766 -1530 2772 -1524
rect 2766 -1536 2772 -1530
rect 2766 -1542 2772 -1536
rect 2766 -1548 2772 -1542
rect 2766 -1554 2772 -1548
rect 2766 -1560 2772 -1554
rect 2766 -1566 2772 -1560
rect 2766 -1572 2772 -1566
rect 2766 -1578 2772 -1572
rect 2766 -1584 2772 -1578
rect 2766 -1590 2772 -1584
rect 2766 -1596 2772 -1590
rect 2766 -1602 2772 -1596
rect 2766 -1608 2772 -1602
rect 2766 -1614 2772 -1608
rect 2766 -1620 2772 -1614
rect 2766 -1626 2772 -1620
rect 2766 -1632 2772 -1626
rect 2766 -2382 2772 -2376
rect 2766 -2388 2772 -2382
rect 2766 -2394 2772 -2388
rect 2766 -2400 2772 -2394
rect 2766 -2406 2772 -2400
rect 2766 -2412 2772 -2406
rect 2766 -2418 2772 -2412
rect 2766 -2424 2772 -2418
rect 2766 -2430 2772 -2424
rect 2766 -2436 2772 -2430
rect 2766 -2442 2772 -2436
rect 2766 -2448 2772 -2442
rect 2766 -2454 2772 -2448
rect 2766 -2460 2772 -2454
rect 2766 -2466 2772 -2460
rect 2766 -2472 2772 -2466
rect 2766 -2478 2772 -2472
rect 2766 -2484 2772 -2478
rect 2766 -2490 2772 -2484
rect 2766 -2496 2772 -2490
rect 2766 -2502 2772 -2496
rect 2766 -2508 2772 -2502
rect 2766 -2514 2772 -2508
rect 2766 -2520 2772 -2514
rect 2766 -2526 2772 -2520
rect 2766 -2532 2772 -2526
rect 2766 -2538 2772 -2532
rect 2766 -2544 2772 -2538
rect 2766 -2550 2772 -2544
rect 2766 -2556 2772 -2550
rect 2766 -2562 2772 -2556
rect 2766 -2568 2772 -2562
rect 2766 -2574 2772 -2568
rect 2766 -2580 2772 -2574
rect 2766 -2586 2772 -2580
rect 2766 -2592 2772 -2586
rect 2766 -2598 2772 -2592
rect 2766 -2604 2772 -2598
rect 2766 -2610 2772 -2604
rect 2766 -2616 2772 -2610
rect 2766 -2622 2772 -2616
rect 2766 -2628 2772 -2622
rect 2766 -2634 2772 -2628
rect 2766 -2640 2772 -2634
rect 2766 -2646 2772 -2640
rect 2772 -1116 2778 -1110
rect 2772 -1122 2778 -1116
rect 2772 -1128 2778 -1122
rect 2772 -1134 2778 -1128
rect 2772 -1140 2778 -1134
rect 2772 -1146 2778 -1140
rect 2772 -1152 2778 -1146
rect 2772 -1158 2778 -1152
rect 2772 -1164 2778 -1158
rect 2772 -1170 2778 -1164
rect 2772 -1176 2778 -1170
rect 2772 -1182 2778 -1176
rect 2772 -1188 2778 -1182
rect 2772 -1194 2778 -1188
rect 2772 -1200 2778 -1194
rect 2772 -1206 2778 -1200
rect 2772 -1212 2778 -1206
rect 2772 -1218 2778 -1212
rect 2772 -1224 2778 -1218
rect 2772 -1230 2778 -1224
rect 2772 -1236 2778 -1230
rect 2772 -1242 2778 -1236
rect 2772 -1248 2778 -1242
rect 2772 -1254 2778 -1248
rect 2772 -1260 2778 -1254
rect 2772 -1266 2778 -1260
rect 2772 -1272 2778 -1266
rect 2772 -1278 2778 -1272
rect 2772 -1284 2778 -1278
rect 2772 -1290 2778 -1284
rect 2772 -1296 2778 -1290
rect 2772 -1302 2778 -1296
rect 2772 -1308 2778 -1302
rect 2772 -1314 2778 -1308
rect 2772 -1320 2778 -1314
rect 2772 -1326 2778 -1320
rect 2772 -1332 2778 -1326
rect 2772 -1338 2778 -1332
rect 2772 -1344 2778 -1338
rect 2772 -1350 2778 -1344
rect 2772 -1356 2778 -1350
rect 2772 -1362 2778 -1356
rect 2772 -1368 2778 -1362
rect 2772 -1374 2778 -1368
rect 2772 -1380 2778 -1374
rect 2772 -1386 2778 -1380
rect 2772 -1392 2778 -1386
rect 2772 -1398 2778 -1392
rect 2772 -1404 2778 -1398
rect 2772 -1410 2778 -1404
rect 2772 -1416 2778 -1410
rect 2772 -1422 2778 -1416
rect 2772 -1428 2778 -1422
rect 2772 -1434 2778 -1428
rect 2772 -1440 2778 -1434
rect 2772 -1446 2778 -1440
rect 2772 -1452 2778 -1446
rect 2772 -1458 2778 -1452
rect 2772 -1464 2778 -1458
rect 2772 -1470 2778 -1464
rect 2772 -1476 2778 -1470
rect 2772 -1482 2778 -1476
rect 2772 -1488 2778 -1482
rect 2772 -1494 2778 -1488
rect 2772 -1500 2778 -1494
rect 2772 -1506 2778 -1500
rect 2772 -1512 2778 -1506
rect 2772 -1518 2778 -1512
rect 2772 -1524 2778 -1518
rect 2772 -1530 2778 -1524
rect 2772 -1536 2778 -1530
rect 2772 -1542 2778 -1536
rect 2772 -1548 2778 -1542
rect 2772 -1554 2778 -1548
rect 2772 -1560 2778 -1554
rect 2772 -1566 2778 -1560
rect 2772 -1572 2778 -1566
rect 2772 -1578 2778 -1572
rect 2772 -1584 2778 -1578
rect 2772 -1590 2778 -1584
rect 2772 -1596 2778 -1590
rect 2772 -1602 2778 -1596
rect 2772 -1608 2778 -1602
rect 2772 -1614 2778 -1608
rect 2772 -1620 2778 -1614
rect 2772 -1626 2778 -1620
rect 2772 -2382 2778 -2376
rect 2772 -2388 2778 -2382
rect 2772 -2394 2778 -2388
rect 2772 -2400 2778 -2394
rect 2772 -2406 2778 -2400
rect 2772 -2412 2778 -2406
rect 2772 -2418 2778 -2412
rect 2772 -2424 2778 -2418
rect 2772 -2430 2778 -2424
rect 2772 -2436 2778 -2430
rect 2772 -2442 2778 -2436
rect 2772 -2448 2778 -2442
rect 2772 -2454 2778 -2448
rect 2772 -2460 2778 -2454
rect 2772 -2466 2778 -2460
rect 2772 -2472 2778 -2466
rect 2772 -2478 2778 -2472
rect 2772 -2484 2778 -2478
rect 2772 -2490 2778 -2484
rect 2772 -2496 2778 -2490
rect 2772 -2502 2778 -2496
rect 2772 -2508 2778 -2502
rect 2772 -2514 2778 -2508
rect 2772 -2520 2778 -2514
rect 2772 -2526 2778 -2520
rect 2772 -2532 2778 -2526
rect 2772 -2538 2778 -2532
rect 2772 -2544 2778 -2538
rect 2772 -2550 2778 -2544
rect 2772 -2556 2778 -2550
rect 2772 -2562 2778 -2556
rect 2772 -2568 2778 -2562
rect 2772 -2574 2778 -2568
rect 2772 -2580 2778 -2574
rect 2772 -2586 2778 -2580
rect 2772 -2592 2778 -2586
rect 2772 -2598 2778 -2592
rect 2772 -2604 2778 -2598
rect 2772 -2610 2778 -2604
rect 2772 -2616 2778 -2610
rect 2772 -2622 2778 -2616
rect 2772 -2628 2778 -2622
rect 2772 -2634 2778 -2628
rect 2772 -2640 2778 -2634
rect 2778 -1110 2784 -1104
rect 2778 -1116 2784 -1110
rect 2778 -1122 2784 -1116
rect 2778 -1128 2784 -1122
rect 2778 -1134 2784 -1128
rect 2778 -1140 2784 -1134
rect 2778 -1146 2784 -1140
rect 2778 -1152 2784 -1146
rect 2778 -1158 2784 -1152
rect 2778 -1164 2784 -1158
rect 2778 -1170 2784 -1164
rect 2778 -1176 2784 -1170
rect 2778 -1182 2784 -1176
rect 2778 -1188 2784 -1182
rect 2778 -1194 2784 -1188
rect 2778 -1200 2784 -1194
rect 2778 -1206 2784 -1200
rect 2778 -1212 2784 -1206
rect 2778 -1218 2784 -1212
rect 2778 -1224 2784 -1218
rect 2778 -1230 2784 -1224
rect 2778 -1236 2784 -1230
rect 2778 -1242 2784 -1236
rect 2778 -1248 2784 -1242
rect 2778 -1254 2784 -1248
rect 2778 -1260 2784 -1254
rect 2778 -1266 2784 -1260
rect 2778 -1272 2784 -1266
rect 2778 -1278 2784 -1272
rect 2778 -1284 2784 -1278
rect 2778 -1290 2784 -1284
rect 2778 -1296 2784 -1290
rect 2778 -1302 2784 -1296
rect 2778 -1308 2784 -1302
rect 2778 -1314 2784 -1308
rect 2778 -1320 2784 -1314
rect 2778 -1326 2784 -1320
rect 2778 -1332 2784 -1326
rect 2778 -1338 2784 -1332
rect 2778 -1344 2784 -1338
rect 2778 -1350 2784 -1344
rect 2778 -1356 2784 -1350
rect 2778 -1362 2784 -1356
rect 2778 -1368 2784 -1362
rect 2778 -1374 2784 -1368
rect 2778 -1380 2784 -1374
rect 2778 -1386 2784 -1380
rect 2778 -1392 2784 -1386
rect 2778 -1398 2784 -1392
rect 2778 -1404 2784 -1398
rect 2778 -1410 2784 -1404
rect 2778 -1416 2784 -1410
rect 2778 -1422 2784 -1416
rect 2778 -1428 2784 -1422
rect 2778 -1434 2784 -1428
rect 2778 -1440 2784 -1434
rect 2778 -1446 2784 -1440
rect 2778 -1452 2784 -1446
rect 2778 -1458 2784 -1452
rect 2778 -1464 2784 -1458
rect 2778 -1470 2784 -1464
rect 2778 -1476 2784 -1470
rect 2778 -1482 2784 -1476
rect 2778 -1488 2784 -1482
rect 2778 -1494 2784 -1488
rect 2778 -1500 2784 -1494
rect 2778 -1506 2784 -1500
rect 2778 -1512 2784 -1506
rect 2778 -1518 2784 -1512
rect 2778 -1524 2784 -1518
rect 2778 -1530 2784 -1524
rect 2778 -1536 2784 -1530
rect 2778 -1542 2784 -1536
rect 2778 -1548 2784 -1542
rect 2778 -1554 2784 -1548
rect 2778 -1560 2784 -1554
rect 2778 -1566 2784 -1560
rect 2778 -1572 2784 -1566
rect 2778 -1578 2784 -1572
rect 2778 -1584 2784 -1578
rect 2778 -1590 2784 -1584
rect 2778 -1596 2784 -1590
rect 2778 -1602 2784 -1596
rect 2778 -1608 2784 -1602
rect 2778 -1614 2784 -1608
rect 2778 -2376 2784 -2370
rect 2778 -2382 2784 -2376
rect 2778 -2388 2784 -2382
rect 2778 -2394 2784 -2388
rect 2778 -2400 2784 -2394
rect 2778 -2406 2784 -2400
rect 2778 -2412 2784 -2406
rect 2778 -2418 2784 -2412
rect 2778 -2424 2784 -2418
rect 2778 -2430 2784 -2424
rect 2778 -2436 2784 -2430
rect 2778 -2442 2784 -2436
rect 2778 -2448 2784 -2442
rect 2778 -2454 2784 -2448
rect 2778 -2460 2784 -2454
rect 2778 -2466 2784 -2460
rect 2778 -2472 2784 -2466
rect 2778 -2478 2784 -2472
rect 2778 -2484 2784 -2478
rect 2778 -2490 2784 -2484
rect 2778 -2496 2784 -2490
rect 2778 -2502 2784 -2496
rect 2778 -2508 2784 -2502
rect 2778 -2514 2784 -2508
rect 2778 -2520 2784 -2514
rect 2778 -2526 2784 -2520
rect 2778 -2532 2784 -2526
rect 2778 -2538 2784 -2532
rect 2778 -2544 2784 -2538
rect 2778 -2550 2784 -2544
rect 2778 -2556 2784 -2550
rect 2778 -2562 2784 -2556
rect 2778 -2568 2784 -2562
rect 2778 -2574 2784 -2568
rect 2778 -2580 2784 -2574
rect 2778 -2586 2784 -2580
rect 2778 -2592 2784 -2586
rect 2778 -2598 2784 -2592
rect 2778 -2604 2784 -2598
rect 2778 -2610 2784 -2604
rect 2778 -2616 2784 -2610
rect 2778 -2622 2784 -2616
rect 2778 -2628 2784 -2622
rect 2778 -2634 2784 -2628
rect 2778 -2640 2784 -2634
rect 2784 -1104 2790 -1098
rect 2784 -1110 2790 -1104
rect 2784 -1116 2790 -1110
rect 2784 -1122 2790 -1116
rect 2784 -1128 2790 -1122
rect 2784 -1134 2790 -1128
rect 2784 -1140 2790 -1134
rect 2784 -1146 2790 -1140
rect 2784 -1152 2790 -1146
rect 2784 -1158 2790 -1152
rect 2784 -1164 2790 -1158
rect 2784 -1170 2790 -1164
rect 2784 -1176 2790 -1170
rect 2784 -1182 2790 -1176
rect 2784 -1188 2790 -1182
rect 2784 -1194 2790 -1188
rect 2784 -1200 2790 -1194
rect 2784 -1206 2790 -1200
rect 2784 -1212 2790 -1206
rect 2784 -1218 2790 -1212
rect 2784 -1224 2790 -1218
rect 2784 -1230 2790 -1224
rect 2784 -1236 2790 -1230
rect 2784 -1242 2790 -1236
rect 2784 -1248 2790 -1242
rect 2784 -1254 2790 -1248
rect 2784 -1260 2790 -1254
rect 2784 -1266 2790 -1260
rect 2784 -1272 2790 -1266
rect 2784 -1278 2790 -1272
rect 2784 -1284 2790 -1278
rect 2784 -1290 2790 -1284
rect 2784 -1296 2790 -1290
rect 2784 -1302 2790 -1296
rect 2784 -1308 2790 -1302
rect 2784 -1314 2790 -1308
rect 2784 -1320 2790 -1314
rect 2784 -1326 2790 -1320
rect 2784 -1332 2790 -1326
rect 2784 -1338 2790 -1332
rect 2784 -1344 2790 -1338
rect 2784 -1350 2790 -1344
rect 2784 -1356 2790 -1350
rect 2784 -1362 2790 -1356
rect 2784 -1368 2790 -1362
rect 2784 -1374 2790 -1368
rect 2784 -1380 2790 -1374
rect 2784 -1386 2790 -1380
rect 2784 -1392 2790 -1386
rect 2784 -1398 2790 -1392
rect 2784 -1404 2790 -1398
rect 2784 -1410 2790 -1404
rect 2784 -1416 2790 -1410
rect 2784 -1422 2790 -1416
rect 2784 -1428 2790 -1422
rect 2784 -1434 2790 -1428
rect 2784 -1440 2790 -1434
rect 2784 -1446 2790 -1440
rect 2784 -1452 2790 -1446
rect 2784 -1458 2790 -1452
rect 2784 -1464 2790 -1458
rect 2784 -1470 2790 -1464
rect 2784 -1476 2790 -1470
rect 2784 -1482 2790 -1476
rect 2784 -1488 2790 -1482
rect 2784 -1494 2790 -1488
rect 2784 -1500 2790 -1494
rect 2784 -1506 2790 -1500
rect 2784 -1512 2790 -1506
rect 2784 -1518 2790 -1512
rect 2784 -1524 2790 -1518
rect 2784 -1530 2790 -1524
rect 2784 -1536 2790 -1530
rect 2784 -1542 2790 -1536
rect 2784 -1548 2790 -1542
rect 2784 -1554 2790 -1548
rect 2784 -1560 2790 -1554
rect 2784 -1566 2790 -1560
rect 2784 -1572 2790 -1566
rect 2784 -1578 2790 -1572
rect 2784 -1584 2790 -1578
rect 2784 -1590 2790 -1584
rect 2784 -1596 2790 -1590
rect 2784 -1602 2790 -1596
rect 2784 -1608 2790 -1602
rect 2784 -2376 2790 -2370
rect 2784 -2382 2790 -2376
rect 2784 -2388 2790 -2382
rect 2784 -2394 2790 -2388
rect 2784 -2400 2790 -2394
rect 2784 -2406 2790 -2400
rect 2784 -2412 2790 -2406
rect 2784 -2418 2790 -2412
rect 2784 -2424 2790 -2418
rect 2784 -2430 2790 -2424
rect 2784 -2436 2790 -2430
rect 2784 -2442 2790 -2436
rect 2784 -2448 2790 -2442
rect 2784 -2454 2790 -2448
rect 2784 -2460 2790 -2454
rect 2784 -2466 2790 -2460
rect 2784 -2472 2790 -2466
rect 2784 -2478 2790 -2472
rect 2784 -2484 2790 -2478
rect 2784 -2490 2790 -2484
rect 2784 -2496 2790 -2490
rect 2784 -2502 2790 -2496
rect 2784 -2508 2790 -2502
rect 2784 -2514 2790 -2508
rect 2784 -2520 2790 -2514
rect 2784 -2526 2790 -2520
rect 2784 -2532 2790 -2526
rect 2784 -2538 2790 -2532
rect 2784 -2544 2790 -2538
rect 2784 -2550 2790 -2544
rect 2784 -2556 2790 -2550
rect 2784 -2562 2790 -2556
rect 2784 -2568 2790 -2562
rect 2784 -2574 2790 -2568
rect 2784 -2580 2790 -2574
rect 2784 -2586 2790 -2580
rect 2784 -2592 2790 -2586
rect 2784 -2598 2790 -2592
rect 2784 -2604 2790 -2598
rect 2784 -2610 2790 -2604
rect 2784 -2616 2790 -2610
rect 2784 -2622 2790 -2616
rect 2784 -2628 2790 -2622
rect 2784 -2634 2790 -2628
rect 2790 -1104 2796 -1098
rect 2790 -1110 2796 -1104
rect 2790 -1116 2796 -1110
rect 2790 -1122 2796 -1116
rect 2790 -1128 2796 -1122
rect 2790 -1134 2796 -1128
rect 2790 -1140 2796 -1134
rect 2790 -1146 2796 -1140
rect 2790 -1152 2796 -1146
rect 2790 -1158 2796 -1152
rect 2790 -1164 2796 -1158
rect 2790 -1170 2796 -1164
rect 2790 -1176 2796 -1170
rect 2790 -1182 2796 -1176
rect 2790 -1188 2796 -1182
rect 2790 -1194 2796 -1188
rect 2790 -1200 2796 -1194
rect 2790 -1206 2796 -1200
rect 2790 -1212 2796 -1206
rect 2790 -1218 2796 -1212
rect 2790 -1224 2796 -1218
rect 2790 -1230 2796 -1224
rect 2790 -1236 2796 -1230
rect 2790 -1242 2796 -1236
rect 2790 -1248 2796 -1242
rect 2790 -1254 2796 -1248
rect 2790 -1260 2796 -1254
rect 2790 -1266 2796 -1260
rect 2790 -1272 2796 -1266
rect 2790 -1278 2796 -1272
rect 2790 -1284 2796 -1278
rect 2790 -1290 2796 -1284
rect 2790 -1296 2796 -1290
rect 2790 -1302 2796 -1296
rect 2790 -1308 2796 -1302
rect 2790 -1314 2796 -1308
rect 2790 -1320 2796 -1314
rect 2790 -1326 2796 -1320
rect 2790 -1332 2796 -1326
rect 2790 -1338 2796 -1332
rect 2790 -1344 2796 -1338
rect 2790 -1350 2796 -1344
rect 2790 -1356 2796 -1350
rect 2790 -1362 2796 -1356
rect 2790 -1368 2796 -1362
rect 2790 -1374 2796 -1368
rect 2790 -1380 2796 -1374
rect 2790 -1386 2796 -1380
rect 2790 -1392 2796 -1386
rect 2790 -1398 2796 -1392
rect 2790 -1404 2796 -1398
rect 2790 -1410 2796 -1404
rect 2790 -1416 2796 -1410
rect 2790 -1422 2796 -1416
rect 2790 -1428 2796 -1422
rect 2790 -1434 2796 -1428
rect 2790 -1440 2796 -1434
rect 2790 -1446 2796 -1440
rect 2790 -1452 2796 -1446
rect 2790 -1458 2796 -1452
rect 2790 -1464 2796 -1458
rect 2790 -1470 2796 -1464
rect 2790 -1476 2796 -1470
rect 2790 -1482 2796 -1476
rect 2790 -1488 2796 -1482
rect 2790 -1494 2796 -1488
rect 2790 -1500 2796 -1494
rect 2790 -1506 2796 -1500
rect 2790 -1512 2796 -1506
rect 2790 -1518 2796 -1512
rect 2790 -1524 2796 -1518
rect 2790 -1530 2796 -1524
rect 2790 -1536 2796 -1530
rect 2790 -1542 2796 -1536
rect 2790 -1548 2796 -1542
rect 2790 -1554 2796 -1548
rect 2790 -1560 2796 -1554
rect 2790 -1566 2796 -1560
rect 2790 -1572 2796 -1566
rect 2790 -1578 2796 -1572
rect 2790 -1584 2796 -1578
rect 2790 -1590 2796 -1584
rect 2790 -1596 2796 -1590
rect 2790 -2376 2796 -2370
rect 2790 -2382 2796 -2376
rect 2790 -2388 2796 -2382
rect 2790 -2394 2796 -2388
rect 2790 -2400 2796 -2394
rect 2790 -2406 2796 -2400
rect 2790 -2412 2796 -2406
rect 2790 -2418 2796 -2412
rect 2790 -2424 2796 -2418
rect 2790 -2430 2796 -2424
rect 2790 -2436 2796 -2430
rect 2790 -2442 2796 -2436
rect 2790 -2448 2796 -2442
rect 2790 -2454 2796 -2448
rect 2790 -2460 2796 -2454
rect 2790 -2466 2796 -2460
rect 2790 -2472 2796 -2466
rect 2790 -2478 2796 -2472
rect 2790 -2484 2796 -2478
rect 2790 -2490 2796 -2484
rect 2790 -2496 2796 -2490
rect 2790 -2502 2796 -2496
rect 2790 -2508 2796 -2502
rect 2790 -2514 2796 -2508
rect 2790 -2520 2796 -2514
rect 2790 -2526 2796 -2520
rect 2790 -2532 2796 -2526
rect 2790 -2538 2796 -2532
rect 2790 -2544 2796 -2538
rect 2790 -2550 2796 -2544
rect 2790 -2556 2796 -2550
rect 2790 -2562 2796 -2556
rect 2790 -2568 2796 -2562
rect 2790 -2574 2796 -2568
rect 2790 -2580 2796 -2574
rect 2790 -2586 2796 -2580
rect 2790 -2592 2796 -2586
rect 2790 -2598 2796 -2592
rect 2790 -2604 2796 -2598
rect 2790 -2610 2796 -2604
rect 2790 -2616 2796 -2610
rect 2790 -2622 2796 -2616
rect 2790 -2628 2796 -2622
rect 2796 -1098 2802 -1092
rect 2796 -1104 2802 -1098
rect 2796 -1110 2802 -1104
rect 2796 -1116 2802 -1110
rect 2796 -1122 2802 -1116
rect 2796 -1128 2802 -1122
rect 2796 -1134 2802 -1128
rect 2796 -1140 2802 -1134
rect 2796 -1146 2802 -1140
rect 2796 -1152 2802 -1146
rect 2796 -1158 2802 -1152
rect 2796 -1164 2802 -1158
rect 2796 -1170 2802 -1164
rect 2796 -1176 2802 -1170
rect 2796 -1182 2802 -1176
rect 2796 -1188 2802 -1182
rect 2796 -1194 2802 -1188
rect 2796 -1200 2802 -1194
rect 2796 -1206 2802 -1200
rect 2796 -1212 2802 -1206
rect 2796 -1218 2802 -1212
rect 2796 -1224 2802 -1218
rect 2796 -1230 2802 -1224
rect 2796 -1236 2802 -1230
rect 2796 -1242 2802 -1236
rect 2796 -1248 2802 -1242
rect 2796 -1254 2802 -1248
rect 2796 -1260 2802 -1254
rect 2796 -1266 2802 -1260
rect 2796 -1272 2802 -1266
rect 2796 -1278 2802 -1272
rect 2796 -1284 2802 -1278
rect 2796 -1290 2802 -1284
rect 2796 -1296 2802 -1290
rect 2796 -1302 2802 -1296
rect 2796 -1308 2802 -1302
rect 2796 -1314 2802 -1308
rect 2796 -1320 2802 -1314
rect 2796 -1326 2802 -1320
rect 2796 -1332 2802 -1326
rect 2796 -1338 2802 -1332
rect 2796 -1344 2802 -1338
rect 2796 -1350 2802 -1344
rect 2796 -1356 2802 -1350
rect 2796 -1362 2802 -1356
rect 2796 -1368 2802 -1362
rect 2796 -1374 2802 -1368
rect 2796 -1380 2802 -1374
rect 2796 -1386 2802 -1380
rect 2796 -1392 2802 -1386
rect 2796 -1398 2802 -1392
rect 2796 -1404 2802 -1398
rect 2796 -1410 2802 -1404
rect 2796 -1416 2802 -1410
rect 2796 -1422 2802 -1416
rect 2796 -1428 2802 -1422
rect 2796 -1434 2802 -1428
rect 2796 -1440 2802 -1434
rect 2796 -1446 2802 -1440
rect 2796 -1452 2802 -1446
rect 2796 -1458 2802 -1452
rect 2796 -1464 2802 -1458
rect 2796 -1470 2802 -1464
rect 2796 -1476 2802 -1470
rect 2796 -1482 2802 -1476
rect 2796 -1488 2802 -1482
rect 2796 -1494 2802 -1488
rect 2796 -1500 2802 -1494
rect 2796 -1506 2802 -1500
rect 2796 -1512 2802 -1506
rect 2796 -1518 2802 -1512
rect 2796 -1524 2802 -1518
rect 2796 -1530 2802 -1524
rect 2796 -1536 2802 -1530
rect 2796 -1542 2802 -1536
rect 2796 -1548 2802 -1542
rect 2796 -1554 2802 -1548
rect 2796 -1560 2802 -1554
rect 2796 -1566 2802 -1560
rect 2796 -1572 2802 -1566
rect 2796 -1578 2802 -1572
rect 2796 -1584 2802 -1578
rect 2796 -1590 2802 -1584
rect 2796 -2376 2802 -2370
rect 2796 -2382 2802 -2376
rect 2796 -2388 2802 -2382
rect 2796 -2394 2802 -2388
rect 2796 -2400 2802 -2394
rect 2796 -2406 2802 -2400
rect 2796 -2412 2802 -2406
rect 2796 -2418 2802 -2412
rect 2796 -2424 2802 -2418
rect 2796 -2430 2802 -2424
rect 2796 -2436 2802 -2430
rect 2796 -2442 2802 -2436
rect 2796 -2448 2802 -2442
rect 2796 -2454 2802 -2448
rect 2796 -2460 2802 -2454
rect 2796 -2466 2802 -2460
rect 2796 -2472 2802 -2466
rect 2796 -2478 2802 -2472
rect 2796 -2484 2802 -2478
rect 2796 -2490 2802 -2484
rect 2796 -2496 2802 -2490
rect 2796 -2502 2802 -2496
rect 2796 -2508 2802 -2502
rect 2796 -2514 2802 -2508
rect 2796 -2520 2802 -2514
rect 2796 -2526 2802 -2520
rect 2796 -2532 2802 -2526
rect 2796 -2538 2802 -2532
rect 2796 -2544 2802 -2538
rect 2796 -2550 2802 -2544
rect 2796 -2556 2802 -2550
rect 2796 -2562 2802 -2556
rect 2796 -2568 2802 -2562
rect 2796 -2574 2802 -2568
rect 2796 -2580 2802 -2574
rect 2796 -2586 2802 -2580
rect 2796 -2592 2802 -2586
rect 2796 -2598 2802 -2592
rect 2796 -2604 2802 -2598
rect 2796 -2610 2802 -2604
rect 2796 -2616 2802 -2610
rect 2796 -2622 2802 -2616
rect 2802 -1092 2808 -1086
rect 2802 -1098 2808 -1092
rect 2802 -1104 2808 -1098
rect 2802 -1110 2808 -1104
rect 2802 -1116 2808 -1110
rect 2802 -1122 2808 -1116
rect 2802 -1128 2808 -1122
rect 2802 -1134 2808 -1128
rect 2802 -1140 2808 -1134
rect 2802 -1146 2808 -1140
rect 2802 -1152 2808 -1146
rect 2802 -1158 2808 -1152
rect 2802 -1164 2808 -1158
rect 2802 -1170 2808 -1164
rect 2802 -1176 2808 -1170
rect 2802 -1182 2808 -1176
rect 2802 -1188 2808 -1182
rect 2802 -1194 2808 -1188
rect 2802 -1200 2808 -1194
rect 2802 -1206 2808 -1200
rect 2802 -1212 2808 -1206
rect 2802 -1218 2808 -1212
rect 2802 -1224 2808 -1218
rect 2802 -1230 2808 -1224
rect 2802 -1236 2808 -1230
rect 2802 -1242 2808 -1236
rect 2802 -1248 2808 -1242
rect 2802 -1254 2808 -1248
rect 2802 -1260 2808 -1254
rect 2802 -1266 2808 -1260
rect 2802 -1272 2808 -1266
rect 2802 -1278 2808 -1272
rect 2802 -1284 2808 -1278
rect 2802 -1290 2808 -1284
rect 2802 -1296 2808 -1290
rect 2802 -1302 2808 -1296
rect 2802 -1308 2808 -1302
rect 2802 -1314 2808 -1308
rect 2802 -1320 2808 -1314
rect 2802 -1326 2808 -1320
rect 2802 -1332 2808 -1326
rect 2802 -1338 2808 -1332
rect 2802 -1344 2808 -1338
rect 2802 -1350 2808 -1344
rect 2802 -1356 2808 -1350
rect 2802 -1362 2808 -1356
rect 2802 -1368 2808 -1362
rect 2802 -1374 2808 -1368
rect 2802 -1380 2808 -1374
rect 2802 -1386 2808 -1380
rect 2802 -1392 2808 -1386
rect 2802 -1398 2808 -1392
rect 2802 -1404 2808 -1398
rect 2802 -1410 2808 -1404
rect 2802 -1416 2808 -1410
rect 2802 -1422 2808 -1416
rect 2802 -1428 2808 -1422
rect 2802 -1434 2808 -1428
rect 2802 -1440 2808 -1434
rect 2802 -1446 2808 -1440
rect 2802 -1452 2808 -1446
rect 2802 -1458 2808 -1452
rect 2802 -1464 2808 -1458
rect 2802 -1470 2808 -1464
rect 2802 -1476 2808 -1470
rect 2802 -1482 2808 -1476
rect 2802 -1488 2808 -1482
rect 2802 -1494 2808 -1488
rect 2802 -1500 2808 -1494
rect 2802 -1506 2808 -1500
rect 2802 -1512 2808 -1506
rect 2802 -1518 2808 -1512
rect 2802 -1524 2808 -1518
rect 2802 -1530 2808 -1524
rect 2802 -1536 2808 -1530
rect 2802 -1542 2808 -1536
rect 2802 -1548 2808 -1542
rect 2802 -1554 2808 -1548
rect 2802 -1560 2808 -1554
rect 2802 -1566 2808 -1560
rect 2802 -1572 2808 -1566
rect 2802 -1578 2808 -1572
rect 2802 -2370 2808 -2364
rect 2802 -2376 2808 -2370
rect 2802 -2382 2808 -2376
rect 2802 -2388 2808 -2382
rect 2802 -2394 2808 -2388
rect 2802 -2400 2808 -2394
rect 2802 -2406 2808 -2400
rect 2802 -2412 2808 -2406
rect 2802 -2418 2808 -2412
rect 2802 -2424 2808 -2418
rect 2802 -2430 2808 -2424
rect 2802 -2436 2808 -2430
rect 2802 -2442 2808 -2436
rect 2802 -2448 2808 -2442
rect 2802 -2454 2808 -2448
rect 2802 -2460 2808 -2454
rect 2802 -2466 2808 -2460
rect 2802 -2472 2808 -2466
rect 2802 -2478 2808 -2472
rect 2802 -2484 2808 -2478
rect 2802 -2490 2808 -2484
rect 2802 -2496 2808 -2490
rect 2802 -2502 2808 -2496
rect 2802 -2508 2808 -2502
rect 2802 -2514 2808 -2508
rect 2802 -2520 2808 -2514
rect 2802 -2526 2808 -2520
rect 2802 -2532 2808 -2526
rect 2802 -2538 2808 -2532
rect 2802 -2544 2808 -2538
rect 2802 -2550 2808 -2544
rect 2802 -2556 2808 -2550
rect 2802 -2562 2808 -2556
rect 2802 -2568 2808 -2562
rect 2802 -2574 2808 -2568
rect 2802 -2580 2808 -2574
rect 2802 -2586 2808 -2580
rect 2802 -2592 2808 -2586
rect 2802 -2598 2808 -2592
rect 2802 -2604 2808 -2598
rect 2802 -2610 2808 -2604
rect 2802 -2616 2808 -2610
rect 2808 -1092 2814 -1086
rect 2808 -1098 2814 -1092
rect 2808 -1104 2814 -1098
rect 2808 -1110 2814 -1104
rect 2808 -1116 2814 -1110
rect 2808 -1122 2814 -1116
rect 2808 -1128 2814 -1122
rect 2808 -1134 2814 -1128
rect 2808 -1140 2814 -1134
rect 2808 -1146 2814 -1140
rect 2808 -1152 2814 -1146
rect 2808 -1158 2814 -1152
rect 2808 -1164 2814 -1158
rect 2808 -1170 2814 -1164
rect 2808 -1176 2814 -1170
rect 2808 -1182 2814 -1176
rect 2808 -1188 2814 -1182
rect 2808 -1194 2814 -1188
rect 2808 -1200 2814 -1194
rect 2808 -1206 2814 -1200
rect 2808 -1212 2814 -1206
rect 2808 -1218 2814 -1212
rect 2808 -1224 2814 -1218
rect 2808 -1230 2814 -1224
rect 2808 -1236 2814 -1230
rect 2808 -1242 2814 -1236
rect 2808 -1248 2814 -1242
rect 2808 -1254 2814 -1248
rect 2808 -1260 2814 -1254
rect 2808 -1266 2814 -1260
rect 2808 -1272 2814 -1266
rect 2808 -1278 2814 -1272
rect 2808 -1284 2814 -1278
rect 2808 -1290 2814 -1284
rect 2808 -1296 2814 -1290
rect 2808 -1302 2814 -1296
rect 2808 -1308 2814 -1302
rect 2808 -1314 2814 -1308
rect 2808 -1320 2814 -1314
rect 2808 -1326 2814 -1320
rect 2808 -1332 2814 -1326
rect 2808 -1338 2814 -1332
rect 2808 -1344 2814 -1338
rect 2808 -1350 2814 -1344
rect 2808 -1356 2814 -1350
rect 2808 -1362 2814 -1356
rect 2808 -1368 2814 -1362
rect 2808 -1374 2814 -1368
rect 2808 -1380 2814 -1374
rect 2808 -1386 2814 -1380
rect 2808 -1392 2814 -1386
rect 2808 -1398 2814 -1392
rect 2808 -1404 2814 -1398
rect 2808 -1410 2814 -1404
rect 2808 -1416 2814 -1410
rect 2808 -1422 2814 -1416
rect 2808 -1428 2814 -1422
rect 2808 -1434 2814 -1428
rect 2808 -1440 2814 -1434
rect 2808 -1446 2814 -1440
rect 2808 -1452 2814 -1446
rect 2808 -1458 2814 -1452
rect 2808 -1464 2814 -1458
rect 2808 -1470 2814 -1464
rect 2808 -1476 2814 -1470
rect 2808 -1482 2814 -1476
rect 2808 -1488 2814 -1482
rect 2808 -1494 2814 -1488
rect 2808 -1500 2814 -1494
rect 2808 -1506 2814 -1500
rect 2808 -1512 2814 -1506
rect 2808 -1518 2814 -1512
rect 2808 -1524 2814 -1518
rect 2808 -1530 2814 -1524
rect 2808 -1536 2814 -1530
rect 2808 -1542 2814 -1536
rect 2808 -1548 2814 -1542
rect 2808 -1554 2814 -1548
rect 2808 -1560 2814 -1554
rect 2808 -1566 2814 -1560
rect 2808 -2370 2814 -2364
rect 2808 -2376 2814 -2370
rect 2808 -2382 2814 -2376
rect 2808 -2388 2814 -2382
rect 2808 -2394 2814 -2388
rect 2808 -2400 2814 -2394
rect 2808 -2406 2814 -2400
rect 2808 -2412 2814 -2406
rect 2808 -2418 2814 -2412
rect 2808 -2424 2814 -2418
rect 2808 -2430 2814 -2424
rect 2808 -2436 2814 -2430
rect 2808 -2442 2814 -2436
rect 2808 -2448 2814 -2442
rect 2808 -2454 2814 -2448
rect 2808 -2460 2814 -2454
rect 2808 -2466 2814 -2460
rect 2808 -2472 2814 -2466
rect 2808 -2478 2814 -2472
rect 2808 -2484 2814 -2478
rect 2808 -2490 2814 -2484
rect 2808 -2496 2814 -2490
rect 2808 -2502 2814 -2496
rect 2808 -2508 2814 -2502
rect 2808 -2514 2814 -2508
rect 2808 -2520 2814 -2514
rect 2808 -2526 2814 -2520
rect 2808 -2532 2814 -2526
rect 2808 -2538 2814 -2532
rect 2808 -2544 2814 -2538
rect 2808 -2550 2814 -2544
rect 2808 -2556 2814 -2550
rect 2808 -2562 2814 -2556
rect 2808 -2568 2814 -2562
rect 2808 -2574 2814 -2568
rect 2808 -2580 2814 -2574
rect 2808 -2586 2814 -2580
rect 2808 -2592 2814 -2586
rect 2808 -2598 2814 -2592
rect 2808 -2604 2814 -2598
rect 2808 -2610 2814 -2604
rect 2814 -1086 2820 -1080
rect 2814 -1092 2820 -1086
rect 2814 -1098 2820 -1092
rect 2814 -1104 2820 -1098
rect 2814 -1110 2820 -1104
rect 2814 -1116 2820 -1110
rect 2814 -1122 2820 -1116
rect 2814 -1128 2820 -1122
rect 2814 -1134 2820 -1128
rect 2814 -1140 2820 -1134
rect 2814 -1146 2820 -1140
rect 2814 -1152 2820 -1146
rect 2814 -1158 2820 -1152
rect 2814 -1164 2820 -1158
rect 2814 -1170 2820 -1164
rect 2814 -1176 2820 -1170
rect 2814 -1182 2820 -1176
rect 2814 -1188 2820 -1182
rect 2814 -1194 2820 -1188
rect 2814 -1200 2820 -1194
rect 2814 -1206 2820 -1200
rect 2814 -1212 2820 -1206
rect 2814 -1218 2820 -1212
rect 2814 -1224 2820 -1218
rect 2814 -1230 2820 -1224
rect 2814 -1236 2820 -1230
rect 2814 -1242 2820 -1236
rect 2814 -1248 2820 -1242
rect 2814 -1254 2820 -1248
rect 2814 -1260 2820 -1254
rect 2814 -1266 2820 -1260
rect 2814 -1272 2820 -1266
rect 2814 -1278 2820 -1272
rect 2814 -1284 2820 -1278
rect 2814 -1290 2820 -1284
rect 2814 -1296 2820 -1290
rect 2814 -1302 2820 -1296
rect 2814 -1308 2820 -1302
rect 2814 -1314 2820 -1308
rect 2814 -1320 2820 -1314
rect 2814 -1326 2820 -1320
rect 2814 -1332 2820 -1326
rect 2814 -1338 2820 -1332
rect 2814 -1344 2820 -1338
rect 2814 -1350 2820 -1344
rect 2814 -1356 2820 -1350
rect 2814 -1362 2820 -1356
rect 2814 -1368 2820 -1362
rect 2814 -1374 2820 -1368
rect 2814 -1380 2820 -1374
rect 2814 -1386 2820 -1380
rect 2814 -1392 2820 -1386
rect 2814 -1398 2820 -1392
rect 2814 -1404 2820 -1398
rect 2814 -1410 2820 -1404
rect 2814 -1416 2820 -1410
rect 2814 -1422 2820 -1416
rect 2814 -1428 2820 -1422
rect 2814 -1434 2820 -1428
rect 2814 -1440 2820 -1434
rect 2814 -1446 2820 -1440
rect 2814 -1452 2820 -1446
rect 2814 -1458 2820 -1452
rect 2814 -1464 2820 -1458
rect 2814 -1470 2820 -1464
rect 2814 -1476 2820 -1470
rect 2814 -1482 2820 -1476
rect 2814 -1488 2820 -1482
rect 2814 -1494 2820 -1488
rect 2814 -1500 2820 -1494
rect 2814 -1506 2820 -1500
rect 2814 -1512 2820 -1506
rect 2814 -1518 2820 -1512
rect 2814 -1524 2820 -1518
rect 2814 -1530 2820 -1524
rect 2814 -1536 2820 -1530
rect 2814 -1542 2820 -1536
rect 2814 -1548 2820 -1542
rect 2814 -1554 2820 -1548
rect 2814 -1560 2820 -1554
rect 2814 -2370 2820 -2364
rect 2814 -2376 2820 -2370
rect 2814 -2382 2820 -2376
rect 2814 -2388 2820 -2382
rect 2814 -2394 2820 -2388
rect 2814 -2400 2820 -2394
rect 2814 -2406 2820 -2400
rect 2814 -2412 2820 -2406
rect 2814 -2418 2820 -2412
rect 2814 -2424 2820 -2418
rect 2814 -2430 2820 -2424
rect 2814 -2436 2820 -2430
rect 2814 -2442 2820 -2436
rect 2814 -2448 2820 -2442
rect 2814 -2454 2820 -2448
rect 2814 -2460 2820 -2454
rect 2814 -2466 2820 -2460
rect 2814 -2472 2820 -2466
rect 2814 -2478 2820 -2472
rect 2814 -2484 2820 -2478
rect 2814 -2490 2820 -2484
rect 2814 -2496 2820 -2490
rect 2814 -2502 2820 -2496
rect 2814 -2508 2820 -2502
rect 2814 -2514 2820 -2508
rect 2814 -2520 2820 -2514
rect 2814 -2526 2820 -2520
rect 2814 -2532 2820 -2526
rect 2814 -2538 2820 -2532
rect 2814 -2544 2820 -2538
rect 2814 -2550 2820 -2544
rect 2814 -2556 2820 -2550
rect 2814 -2562 2820 -2556
rect 2814 -2568 2820 -2562
rect 2814 -2574 2820 -2568
rect 2814 -2580 2820 -2574
rect 2814 -2586 2820 -2580
rect 2814 -2592 2820 -2586
rect 2814 -2598 2820 -2592
rect 2814 -2604 2820 -2598
rect 2814 -2610 2820 -2604
rect 2820 -1080 2826 -1074
rect 2820 -1086 2826 -1080
rect 2820 -1092 2826 -1086
rect 2820 -1098 2826 -1092
rect 2820 -1104 2826 -1098
rect 2820 -1110 2826 -1104
rect 2820 -1116 2826 -1110
rect 2820 -1122 2826 -1116
rect 2820 -1128 2826 -1122
rect 2820 -1134 2826 -1128
rect 2820 -1140 2826 -1134
rect 2820 -1146 2826 -1140
rect 2820 -1152 2826 -1146
rect 2820 -1158 2826 -1152
rect 2820 -1164 2826 -1158
rect 2820 -1170 2826 -1164
rect 2820 -1176 2826 -1170
rect 2820 -1182 2826 -1176
rect 2820 -1188 2826 -1182
rect 2820 -1194 2826 -1188
rect 2820 -1200 2826 -1194
rect 2820 -1206 2826 -1200
rect 2820 -1212 2826 -1206
rect 2820 -1218 2826 -1212
rect 2820 -1224 2826 -1218
rect 2820 -1230 2826 -1224
rect 2820 -1236 2826 -1230
rect 2820 -1242 2826 -1236
rect 2820 -1248 2826 -1242
rect 2820 -1254 2826 -1248
rect 2820 -1260 2826 -1254
rect 2820 -1266 2826 -1260
rect 2820 -1272 2826 -1266
rect 2820 -1278 2826 -1272
rect 2820 -1284 2826 -1278
rect 2820 -1290 2826 -1284
rect 2820 -1296 2826 -1290
rect 2820 -1302 2826 -1296
rect 2820 -1308 2826 -1302
rect 2820 -1314 2826 -1308
rect 2820 -1320 2826 -1314
rect 2820 -1326 2826 -1320
rect 2820 -1332 2826 -1326
rect 2820 -1338 2826 -1332
rect 2820 -1344 2826 -1338
rect 2820 -1350 2826 -1344
rect 2820 -1356 2826 -1350
rect 2820 -1362 2826 -1356
rect 2820 -1368 2826 -1362
rect 2820 -1374 2826 -1368
rect 2820 -1380 2826 -1374
rect 2820 -1386 2826 -1380
rect 2820 -1392 2826 -1386
rect 2820 -1398 2826 -1392
rect 2820 -1404 2826 -1398
rect 2820 -1410 2826 -1404
rect 2820 -1416 2826 -1410
rect 2820 -1422 2826 -1416
rect 2820 -1428 2826 -1422
rect 2820 -1434 2826 -1428
rect 2820 -1440 2826 -1434
rect 2820 -1446 2826 -1440
rect 2820 -1452 2826 -1446
rect 2820 -1458 2826 -1452
rect 2820 -1464 2826 -1458
rect 2820 -1470 2826 -1464
rect 2820 -1476 2826 -1470
rect 2820 -1482 2826 -1476
rect 2820 -1488 2826 -1482
rect 2820 -1494 2826 -1488
rect 2820 -1500 2826 -1494
rect 2820 -1506 2826 -1500
rect 2820 -1512 2826 -1506
rect 2820 -1518 2826 -1512
rect 2820 -1524 2826 -1518
rect 2820 -1530 2826 -1524
rect 2820 -1536 2826 -1530
rect 2820 -1542 2826 -1536
rect 2820 -1548 2826 -1542
rect 2820 -2370 2826 -2364
rect 2820 -2376 2826 -2370
rect 2820 -2382 2826 -2376
rect 2820 -2388 2826 -2382
rect 2820 -2394 2826 -2388
rect 2820 -2400 2826 -2394
rect 2820 -2406 2826 -2400
rect 2820 -2412 2826 -2406
rect 2820 -2418 2826 -2412
rect 2820 -2424 2826 -2418
rect 2820 -2430 2826 -2424
rect 2820 -2436 2826 -2430
rect 2820 -2442 2826 -2436
rect 2820 -2448 2826 -2442
rect 2820 -2454 2826 -2448
rect 2820 -2460 2826 -2454
rect 2820 -2466 2826 -2460
rect 2820 -2472 2826 -2466
rect 2820 -2478 2826 -2472
rect 2820 -2484 2826 -2478
rect 2820 -2490 2826 -2484
rect 2820 -2496 2826 -2490
rect 2820 -2502 2826 -2496
rect 2820 -2508 2826 -2502
rect 2820 -2514 2826 -2508
rect 2820 -2520 2826 -2514
rect 2820 -2526 2826 -2520
rect 2820 -2532 2826 -2526
rect 2820 -2538 2826 -2532
rect 2820 -2544 2826 -2538
rect 2820 -2550 2826 -2544
rect 2820 -2556 2826 -2550
rect 2820 -2562 2826 -2556
rect 2820 -2568 2826 -2562
rect 2820 -2574 2826 -2568
rect 2820 -2580 2826 -2574
rect 2820 -2586 2826 -2580
rect 2820 -2592 2826 -2586
rect 2820 -2598 2826 -2592
rect 2820 -2604 2826 -2598
rect 2826 -1080 2832 -1074
rect 2826 -1086 2832 -1080
rect 2826 -1092 2832 -1086
rect 2826 -1098 2832 -1092
rect 2826 -1104 2832 -1098
rect 2826 -1110 2832 -1104
rect 2826 -1116 2832 -1110
rect 2826 -1122 2832 -1116
rect 2826 -1128 2832 -1122
rect 2826 -1134 2832 -1128
rect 2826 -1140 2832 -1134
rect 2826 -1146 2832 -1140
rect 2826 -1152 2832 -1146
rect 2826 -1158 2832 -1152
rect 2826 -1164 2832 -1158
rect 2826 -1170 2832 -1164
rect 2826 -1176 2832 -1170
rect 2826 -1182 2832 -1176
rect 2826 -1188 2832 -1182
rect 2826 -1194 2832 -1188
rect 2826 -1200 2832 -1194
rect 2826 -1206 2832 -1200
rect 2826 -1212 2832 -1206
rect 2826 -1218 2832 -1212
rect 2826 -1224 2832 -1218
rect 2826 -1230 2832 -1224
rect 2826 -1236 2832 -1230
rect 2826 -1242 2832 -1236
rect 2826 -1248 2832 -1242
rect 2826 -1254 2832 -1248
rect 2826 -1260 2832 -1254
rect 2826 -1266 2832 -1260
rect 2826 -1272 2832 -1266
rect 2826 -1278 2832 -1272
rect 2826 -1284 2832 -1278
rect 2826 -1290 2832 -1284
rect 2826 -1296 2832 -1290
rect 2826 -1302 2832 -1296
rect 2826 -1308 2832 -1302
rect 2826 -1314 2832 -1308
rect 2826 -1320 2832 -1314
rect 2826 -1326 2832 -1320
rect 2826 -1332 2832 -1326
rect 2826 -1338 2832 -1332
rect 2826 -1344 2832 -1338
rect 2826 -1350 2832 -1344
rect 2826 -1356 2832 -1350
rect 2826 -1362 2832 -1356
rect 2826 -1368 2832 -1362
rect 2826 -1374 2832 -1368
rect 2826 -1380 2832 -1374
rect 2826 -1386 2832 -1380
rect 2826 -1392 2832 -1386
rect 2826 -1398 2832 -1392
rect 2826 -1404 2832 -1398
rect 2826 -1410 2832 -1404
rect 2826 -1416 2832 -1410
rect 2826 -1422 2832 -1416
rect 2826 -1428 2832 -1422
rect 2826 -1434 2832 -1428
rect 2826 -1440 2832 -1434
rect 2826 -1446 2832 -1440
rect 2826 -1452 2832 -1446
rect 2826 -1458 2832 -1452
rect 2826 -1464 2832 -1458
rect 2826 -1470 2832 -1464
rect 2826 -1476 2832 -1470
rect 2826 -1482 2832 -1476
rect 2826 -1488 2832 -1482
rect 2826 -1494 2832 -1488
rect 2826 -1500 2832 -1494
rect 2826 -1506 2832 -1500
rect 2826 -1512 2832 -1506
rect 2826 -1518 2832 -1512
rect 2826 -1524 2832 -1518
rect 2826 -1530 2832 -1524
rect 2826 -1536 2832 -1530
rect 2826 -2364 2832 -2358
rect 2826 -2370 2832 -2364
rect 2826 -2376 2832 -2370
rect 2826 -2382 2832 -2376
rect 2826 -2388 2832 -2382
rect 2826 -2394 2832 -2388
rect 2826 -2400 2832 -2394
rect 2826 -2406 2832 -2400
rect 2826 -2412 2832 -2406
rect 2826 -2418 2832 -2412
rect 2826 -2424 2832 -2418
rect 2826 -2430 2832 -2424
rect 2826 -2436 2832 -2430
rect 2826 -2442 2832 -2436
rect 2826 -2448 2832 -2442
rect 2826 -2454 2832 -2448
rect 2826 -2460 2832 -2454
rect 2826 -2466 2832 -2460
rect 2826 -2472 2832 -2466
rect 2826 -2478 2832 -2472
rect 2826 -2484 2832 -2478
rect 2826 -2490 2832 -2484
rect 2826 -2496 2832 -2490
rect 2826 -2502 2832 -2496
rect 2826 -2508 2832 -2502
rect 2826 -2514 2832 -2508
rect 2826 -2520 2832 -2514
rect 2826 -2526 2832 -2520
rect 2826 -2532 2832 -2526
rect 2826 -2538 2832 -2532
rect 2826 -2544 2832 -2538
rect 2826 -2550 2832 -2544
rect 2826 -2556 2832 -2550
rect 2826 -2562 2832 -2556
rect 2826 -2568 2832 -2562
rect 2826 -2574 2832 -2568
rect 2826 -2580 2832 -2574
rect 2826 -2586 2832 -2580
rect 2826 -2592 2832 -2586
rect 2826 -2598 2832 -2592
rect 2832 -1074 2838 -1068
rect 2832 -1080 2838 -1074
rect 2832 -1086 2838 -1080
rect 2832 -1092 2838 -1086
rect 2832 -1098 2838 -1092
rect 2832 -1104 2838 -1098
rect 2832 -1110 2838 -1104
rect 2832 -1116 2838 -1110
rect 2832 -1122 2838 -1116
rect 2832 -1128 2838 -1122
rect 2832 -1134 2838 -1128
rect 2832 -1140 2838 -1134
rect 2832 -1146 2838 -1140
rect 2832 -1152 2838 -1146
rect 2832 -1158 2838 -1152
rect 2832 -1164 2838 -1158
rect 2832 -1170 2838 -1164
rect 2832 -1176 2838 -1170
rect 2832 -1182 2838 -1176
rect 2832 -1188 2838 -1182
rect 2832 -1194 2838 -1188
rect 2832 -1200 2838 -1194
rect 2832 -1206 2838 -1200
rect 2832 -1212 2838 -1206
rect 2832 -1218 2838 -1212
rect 2832 -1224 2838 -1218
rect 2832 -1230 2838 -1224
rect 2832 -1236 2838 -1230
rect 2832 -1242 2838 -1236
rect 2832 -1248 2838 -1242
rect 2832 -1254 2838 -1248
rect 2832 -1260 2838 -1254
rect 2832 -1266 2838 -1260
rect 2832 -1272 2838 -1266
rect 2832 -1278 2838 -1272
rect 2832 -1284 2838 -1278
rect 2832 -1290 2838 -1284
rect 2832 -1296 2838 -1290
rect 2832 -1302 2838 -1296
rect 2832 -1308 2838 -1302
rect 2832 -1314 2838 -1308
rect 2832 -1320 2838 -1314
rect 2832 -1326 2838 -1320
rect 2832 -1332 2838 -1326
rect 2832 -1338 2838 -1332
rect 2832 -1344 2838 -1338
rect 2832 -1350 2838 -1344
rect 2832 -1356 2838 -1350
rect 2832 -1362 2838 -1356
rect 2832 -1368 2838 -1362
rect 2832 -1374 2838 -1368
rect 2832 -1380 2838 -1374
rect 2832 -1386 2838 -1380
rect 2832 -1392 2838 -1386
rect 2832 -1398 2838 -1392
rect 2832 -1404 2838 -1398
rect 2832 -1410 2838 -1404
rect 2832 -1416 2838 -1410
rect 2832 -1422 2838 -1416
rect 2832 -1428 2838 -1422
rect 2832 -1434 2838 -1428
rect 2832 -1440 2838 -1434
rect 2832 -1446 2838 -1440
rect 2832 -1452 2838 -1446
rect 2832 -1458 2838 -1452
rect 2832 -1464 2838 -1458
rect 2832 -1470 2838 -1464
rect 2832 -1476 2838 -1470
rect 2832 -1482 2838 -1476
rect 2832 -1488 2838 -1482
rect 2832 -1494 2838 -1488
rect 2832 -1500 2838 -1494
rect 2832 -1506 2838 -1500
rect 2832 -1512 2838 -1506
rect 2832 -1518 2838 -1512
rect 2832 -1524 2838 -1518
rect 2832 -1530 2838 -1524
rect 2832 -2364 2838 -2358
rect 2832 -2370 2838 -2364
rect 2832 -2376 2838 -2370
rect 2832 -2382 2838 -2376
rect 2832 -2388 2838 -2382
rect 2832 -2394 2838 -2388
rect 2832 -2400 2838 -2394
rect 2832 -2406 2838 -2400
rect 2832 -2412 2838 -2406
rect 2832 -2418 2838 -2412
rect 2832 -2424 2838 -2418
rect 2832 -2430 2838 -2424
rect 2832 -2436 2838 -2430
rect 2832 -2442 2838 -2436
rect 2832 -2448 2838 -2442
rect 2832 -2454 2838 -2448
rect 2832 -2460 2838 -2454
rect 2832 -2466 2838 -2460
rect 2832 -2472 2838 -2466
rect 2832 -2478 2838 -2472
rect 2832 -2484 2838 -2478
rect 2832 -2490 2838 -2484
rect 2832 -2496 2838 -2490
rect 2832 -2502 2838 -2496
rect 2832 -2508 2838 -2502
rect 2832 -2514 2838 -2508
rect 2832 -2520 2838 -2514
rect 2832 -2526 2838 -2520
rect 2832 -2532 2838 -2526
rect 2832 -2538 2838 -2532
rect 2832 -2544 2838 -2538
rect 2832 -2550 2838 -2544
rect 2832 -2556 2838 -2550
rect 2832 -2562 2838 -2556
rect 2832 -2568 2838 -2562
rect 2832 -2574 2838 -2568
rect 2832 -2580 2838 -2574
rect 2832 -2586 2838 -2580
rect 2832 -2592 2838 -2586
rect 2838 -1068 2844 -1062
rect 2838 -1074 2844 -1068
rect 2838 -1080 2844 -1074
rect 2838 -1086 2844 -1080
rect 2838 -1092 2844 -1086
rect 2838 -1098 2844 -1092
rect 2838 -1104 2844 -1098
rect 2838 -1110 2844 -1104
rect 2838 -1116 2844 -1110
rect 2838 -1122 2844 -1116
rect 2838 -1128 2844 -1122
rect 2838 -1134 2844 -1128
rect 2838 -1140 2844 -1134
rect 2838 -1146 2844 -1140
rect 2838 -1152 2844 -1146
rect 2838 -1158 2844 -1152
rect 2838 -1164 2844 -1158
rect 2838 -1170 2844 -1164
rect 2838 -1176 2844 -1170
rect 2838 -1182 2844 -1176
rect 2838 -1188 2844 -1182
rect 2838 -1194 2844 -1188
rect 2838 -1200 2844 -1194
rect 2838 -1206 2844 -1200
rect 2838 -1212 2844 -1206
rect 2838 -1218 2844 -1212
rect 2838 -1224 2844 -1218
rect 2838 -1230 2844 -1224
rect 2838 -1236 2844 -1230
rect 2838 -1242 2844 -1236
rect 2838 -1248 2844 -1242
rect 2838 -1254 2844 -1248
rect 2838 -1260 2844 -1254
rect 2838 -1266 2844 -1260
rect 2838 -1272 2844 -1266
rect 2838 -1278 2844 -1272
rect 2838 -1284 2844 -1278
rect 2838 -1290 2844 -1284
rect 2838 -1296 2844 -1290
rect 2838 -1302 2844 -1296
rect 2838 -1308 2844 -1302
rect 2838 -1314 2844 -1308
rect 2838 -1320 2844 -1314
rect 2838 -1326 2844 -1320
rect 2838 -1332 2844 -1326
rect 2838 -1338 2844 -1332
rect 2838 -1344 2844 -1338
rect 2838 -1350 2844 -1344
rect 2838 -1356 2844 -1350
rect 2838 -1362 2844 -1356
rect 2838 -1368 2844 -1362
rect 2838 -1374 2844 -1368
rect 2838 -1380 2844 -1374
rect 2838 -1386 2844 -1380
rect 2838 -1392 2844 -1386
rect 2838 -1398 2844 -1392
rect 2838 -1404 2844 -1398
rect 2838 -1410 2844 -1404
rect 2838 -1416 2844 -1410
rect 2838 -1422 2844 -1416
rect 2838 -1428 2844 -1422
rect 2838 -1434 2844 -1428
rect 2838 -1440 2844 -1434
rect 2838 -1446 2844 -1440
rect 2838 -1452 2844 -1446
rect 2838 -1458 2844 -1452
rect 2838 -1464 2844 -1458
rect 2838 -1470 2844 -1464
rect 2838 -1476 2844 -1470
rect 2838 -1482 2844 -1476
rect 2838 -1488 2844 -1482
rect 2838 -1494 2844 -1488
rect 2838 -1500 2844 -1494
rect 2838 -1506 2844 -1500
rect 2838 -1512 2844 -1506
rect 2838 -1518 2844 -1512
rect 2838 -2364 2844 -2358
rect 2838 -2370 2844 -2364
rect 2838 -2376 2844 -2370
rect 2838 -2382 2844 -2376
rect 2838 -2388 2844 -2382
rect 2838 -2394 2844 -2388
rect 2838 -2400 2844 -2394
rect 2838 -2406 2844 -2400
rect 2838 -2412 2844 -2406
rect 2838 -2418 2844 -2412
rect 2838 -2424 2844 -2418
rect 2838 -2430 2844 -2424
rect 2838 -2436 2844 -2430
rect 2838 -2442 2844 -2436
rect 2838 -2448 2844 -2442
rect 2838 -2454 2844 -2448
rect 2838 -2460 2844 -2454
rect 2838 -2466 2844 -2460
rect 2838 -2472 2844 -2466
rect 2838 -2478 2844 -2472
rect 2838 -2484 2844 -2478
rect 2838 -2490 2844 -2484
rect 2838 -2496 2844 -2490
rect 2838 -2502 2844 -2496
rect 2838 -2508 2844 -2502
rect 2838 -2514 2844 -2508
rect 2838 -2520 2844 -2514
rect 2838 -2526 2844 -2520
rect 2838 -2532 2844 -2526
rect 2838 -2538 2844 -2532
rect 2838 -2544 2844 -2538
rect 2838 -2550 2844 -2544
rect 2838 -2556 2844 -2550
rect 2838 -2562 2844 -2556
rect 2838 -2568 2844 -2562
rect 2838 -2574 2844 -2568
rect 2838 -2580 2844 -2574
rect 2838 -2586 2844 -2580
rect 2844 -1068 2850 -1062
rect 2844 -1074 2850 -1068
rect 2844 -1080 2850 -1074
rect 2844 -1086 2850 -1080
rect 2844 -1092 2850 -1086
rect 2844 -1098 2850 -1092
rect 2844 -1104 2850 -1098
rect 2844 -1110 2850 -1104
rect 2844 -1116 2850 -1110
rect 2844 -1122 2850 -1116
rect 2844 -1128 2850 -1122
rect 2844 -1134 2850 -1128
rect 2844 -1140 2850 -1134
rect 2844 -1146 2850 -1140
rect 2844 -1152 2850 -1146
rect 2844 -1158 2850 -1152
rect 2844 -1164 2850 -1158
rect 2844 -1170 2850 -1164
rect 2844 -1176 2850 -1170
rect 2844 -1182 2850 -1176
rect 2844 -1188 2850 -1182
rect 2844 -1194 2850 -1188
rect 2844 -1200 2850 -1194
rect 2844 -1206 2850 -1200
rect 2844 -1212 2850 -1206
rect 2844 -1218 2850 -1212
rect 2844 -1224 2850 -1218
rect 2844 -1230 2850 -1224
rect 2844 -1236 2850 -1230
rect 2844 -1242 2850 -1236
rect 2844 -1248 2850 -1242
rect 2844 -1254 2850 -1248
rect 2844 -1260 2850 -1254
rect 2844 -1266 2850 -1260
rect 2844 -1272 2850 -1266
rect 2844 -1278 2850 -1272
rect 2844 -1284 2850 -1278
rect 2844 -1290 2850 -1284
rect 2844 -1296 2850 -1290
rect 2844 -1302 2850 -1296
rect 2844 -1308 2850 -1302
rect 2844 -1314 2850 -1308
rect 2844 -1320 2850 -1314
rect 2844 -1326 2850 -1320
rect 2844 -1332 2850 -1326
rect 2844 -1338 2850 -1332
rect 2844 -1344 2850 -1338
rect 2844 -1350 2850 -1344
rect 2844 -1356 2850 -1350
rect 2844 -1362 2850 -1356
rect 2844 -1368 2850 -1362
rect 2844 -1374 2850 -1368
rect 2844 -1380 2850 -1374
rect 2844 -1386 2850 -1380
rect 2844 -1392 2850 -1386
rect 2844 -1398 2850 -1392
rect 2844 -1404 2850 -1398
rect 2844 -1410 2850 -1404
rect 2844 -1416 2850 -1410
rect 2844 -1422 2850 -1416
rect 2844 -1428 2850 -1422
rect 2844 -1434 2850 -1428
rect 2844 -1440 2850 -1434
rect 2844 -1446 2850 -1440
rect 2844 -1452 2850 -1446
rect 2844 -1458 2850 -1452
rect 2844 -1464 2850 -1458
rect 2844 -1470 2850 -1464
rect 2844 -1476 2850 -1470
rect 2844 -1482 2850 -1476
rect 2844 -1488 2850 -1482
rect 2844 -1494 2850 -1488
rect 2844 -1500 2850 -1494
rect 2844 -1506 2850 -1500
rect 2844 -2364 2850 -2358
rect 2844 -2370 2850 -2364
rect 2844 -2376 2850 -2370
rect 2844 -2382 2850 -2376
rect 2844 -2388 2850 -2382
rect 2844 -2394 2850 -2388
rect 2844 -2400 2850 -2394
rect 2844 -2406 2850 -2400
rect 2844 -2412 2850 -2406
rect 2844 -2418 2850 -2412
rect 2844 -2424 2850 -2418
rect 2844 -2430 2850 -2424
rect 2844 -2436 2850 -2430
rect 2844 -2442 2850 -2436
rect 2844 -2448 2850 -2442
rect 2844 -2454 2850 -2448
rect 2844 -2460 2850 -2454
rect 2844 -2466 2850 -2460
rect 2844 -2472 2850 -2466
rect 2844 -2478 2850 -2472
rect 2844 -2484 2850 -2478
rect 2844 -2490 2850 -2484
rect 2844 -2496 2850 -2490
rect 2844 -2502 2850 -2496
rect 2844 -2508 2850 -2502
rect 2844 -2514 2850 -2508
rect 2844 -2520 2850 -2514
rect 2844 -2526 2850 -2520
rect 2844 -2532 2850 -2526
rect 2844 -2538 2850 -2532
rect 2844 -2544 2850 -2538
rect 2844 -2550 2850 -2544
rect 2844 -2556 2850 -2550
rect 2844 -2562 2850 -2556
rect 2844 -2568 2850 -2562
rect 2844 -2574 2850 -2568
rect 2844 -2580 2850 -2574
rect 2850 -1062 2856 -1056
rect 2850 -1068 2856 -1062
rect 2850 -1074 2856 -1068
rect 2850 -1080 2856 -1074
rect 2850 -1086 2856 -1080
rect 2850 -1092 2856 -1086
rect 2850 -1098 2856 -1092
rect 2850 -1104 2856 -1098
rect 2850 -1110 2856 -1104
rect 2850 -1116 2856 -1110
rect 2850 -1122 2856 -1116
rect 2850 -1128 2856 -1122
rect 2850 -1134 2856 -1128
rect 2850 -1140 2856 -1134
rect 2850 -1146 2856 -1140
rect 2850 -1152 2856 -1146
rect 2850 -1158 2856 -1152
rect 2850 -1164 2856 -1158
rect 2850 -1170 2856 -1164
rect 2850 -1176 2856 -1170
rect 2850 -1182 2856 -1176
rect 2850 -1188 2856 -1182
rect 2850 -1194 2856 -1188
rect 2850 -1200 2856 -1194
rect 2850 -1206 2856 -1200
rect 2850 -1212 2856 -1206
rect 2850 -1218 2856 -1212
rect 2850 -1224 2856 -1218
rect 2850 -1230 2856 -1224
rect 2850 -1236 2856 -1230
rect 2850 -1242 2856 -1236
rect 2850 -1248 2856 -1242
rect 2850 -1254 2856 -1248
rect 2850 -1260 2856 -1254
rect 2850 -1266 2856 -1260
rect 2850 -1272 2856 -1266
rect 2850 -1278 2856 -1272
rect 2850 -1284 2856 -1278
rect 2850 -1290 2856 -1284
rect 2850 -1296 2856 -1290
rect 2850 -1302 2856 -1296
rect 2850 -1308 2856 -1302
rect 2850 -1314 2856 -1308
rect 2850 -1320 2856 -1314
rect 2850 -1326 2856 -1320
rect 2850 -1332 2856 -1326
rect 2850 -1338 2856 -1332
rect 2850 -1344 2856 -1338
rect 2850 -1350 2856 -1344
rect 2850 -1356 2856 -1350
rect 2850 -1362 2856 -1356
rect 2850 -1368 2856 -1362
rect 2850 -1374 2856 -1368
rect 2850 -1380 2856 -1374
rect 2850 -1386 2856 -1380
rect 2850 -1392 2856 -1386
rect 2850 -1398 2856 -1392
rect 2850 -1404 2856 -1398
rect 2850 -1410 2856 -1404
rect 2850 -1416 2856 -1410
rect 2850 -1422 2856 -1416
rect 2850 -1428 2856 -1422
rect 2850 -1434 2856 -1428
rect 2850 -1440 2856 -1434
rect 2850 -1446 2856 -1440
rect 2850 -1452 2856 -1446
rect 2850 -1458 2856 -1452
rect 2850 -1464 2856 -1458
rect 2850 -1470 2856 -1464
rect 2850 -1476 2856 -1470
rect 2850 -1482 2856 -1476
rect 2850 -1488 2856 -1482
rect 2850 -1494 2856 -1488
rect 2850 -1500 2856 -1494
rect 2850 -2358 2856 -2352
rect 2850 -2364 2856 -2358
rect 2850 -2370 2856 -2364
rect 2850 -2376 2856 -2370
rect 2850 -2382 2856 -2376
rect 2850 -2388 2856 -2382
rect 2850 -2394 2856 -2388
rect 2850 -2400 2856 -2394
rect 2850 -2406 2856 -2400
rect 2850 -2412 2856 -2406
rect 2850 -2418 2856 -2412
rect 2850 -2424 2856 -2418
rect 2850 -2430 2856 -2424
rect 2850 -2436 2856 -2430
rect 2850 -2442 2856 -2436
rect 2850 -2448 2856 -2442
rect 2850 -2454 2856 -2448
rect 2850 -2460 2856 -2454
rect 2850 -2466 2856 -2460
rect 2850 -2472 2856 -2466
rect 2850 -2478 2856 -2472
rect 2850 -2484 2856 -2478
rect 2850 -2490 2856 -2484
rect 2850 -2496 2856 -2490
rect 2850 -2502 2856 -2496
rect 2850 -2508 2856 -2502
rect 2850 -2514 2856 -2508
rect 2850 -2520 2856 -2514
rect 2850 -2526 2856 -2520
rect 2850 -2532 2856 -2526
rect 2850 -2538 2856 -2532
rect 2850 -2544 2856 -2538
rect 2850 -2550 2856 -2544
rect 2850 -2556 2856 -2550
rect 2850 -2562 2856 -2556
rect 2850 -2568 2856 -2562
rect 2850 -2574 2856 -2568
rect 2856 -1062 2862 -1056
rect 2856 -1068 2862 -1062
rect 2856 -1074 2862 -1068
rect 2856 -1080 2862 -1074
rect 2856 -1086 2862 -1080
rect 2856 -1092 2862 -1086
rect 2856 -1098 2862 -1092
rect 2856 -1104 2862 -1098
rect 2856 -1110 2862 -1104
rect 2856 -1116 2862 -1110
rect 2856 -1122 2862 -1116
rect 2856 -1128 2862 -1122
rect 2856 -1134 2862 -1128
rect 2856 -1140 2862 -1134
rect 2856 -1146 2862 -1140
rect 2856 -1152 2862 -1146
rect 2856 -1158 2862 -1152
rect 2856 -1164 2862 -1158
rect 2856 -1170 2862 -1164
rect 2856 -1176 2862 -1170
rect 2856 -1182 2862 -1176
rect 2856 -1188 2862 -1182
rect 2856 -1194 2862 -1188
rect 2856 -1200 2862 -1194
rect 2856 -1206 2862 -1200
rect 2856 -1212 2862 -1206
rect 2856 -1218 2862 -1212
rect 2856 -1224 2862 -1218
rect 2856 -1230 2862 -1224
rect 2856 -1236 2862 -1230
rect 2856 -1242 2862 -1236
rect 2856 -1248 2862 -1242
rect 2856 -1254 2862 -1248
rect 2856 -1260 2862 -1254
rect 2856 -1266 2862 -1260
rect 2856 -1272 2862 -1266
rect 2856 -1278 2862 -1272
rect 2856 -1284 2862 -1278
rect 2856 -1290 2862 -1284
rect 2856 -1296 2862 -1290
rect 2856 -1302 2862 -1296
rect 2856 -1308 2862 -1302
rect 2856 -1314 2862 -1308
rect 2856 -1320 2862 -1314
rect 2856 -1326 2862 -1320
rect 2856 -1332 2862 -1326
rect 2856 -1338 2862 -1332
rect 2856 -1344 2862 -1338
rect 2856 -1350 2862 -1344
rect 2856 -1356 2862 -1350
rect 2856 -1362 2862 -1356
rect 2856 -1368 2862 -1362
rect 2856 -1374 2862 -1368
rect 2856 -1380 2862 -1374
rect 2856 -1386 2862 -1380
rect 2856 -1392 2862 -1386
rect 2856 -1398 2862 -1392
rect 2856 -1404 2862 -1398
rect 2856 -1410 2862 -1404
rect 2856 -1416 2862 -1410
rect 2856 -1422 2862 -1416
rect 2856 -1428 2862 -1422
rect 2856 -1434 2862 -1428
rect 2856 -1440 2862 -1434
rect 2856 -1446 2862 -1440
rect 2856 -1452 2862 -1446
rect 2856 -1458 2862 -1452
rect 2856 -1464 2862 -1458
rect 2856 -1470 2862 -1464
rect 2856 -1476 2862 -1470
rect 2856 -1482 2862 -1476
rect 2856 -1488 2862 -1482
rect 2856 -2358 2862 -2352
rect 2856 -2364 2862 -2358
rect 2856 -2370 2862 -2364
rect 2856 -2376 2862 -2370
rect 2856 -2382 2862 -2376
rect 2856 -2388 2862 -2382
rect 2856 -2394 2862 -2388
rect 2856 -2400 2862 -2394
rect 2856 -2406 2862 -2400
rect 2856 -2412 2862 -2406
rect 2856 -2418 2862 -2412
rect 2856 -2424 2862 -2418
rect 2856 -2430 2862 -2424
rect 2856 -2436 2862 -2430
rect 2856 -2442 2862 -2436
rect 2856 -2448 2862 -2442
rect 2856 -2454 2862 -2448
rect 2856 -2460 2862 -2454
rect 2856 -2466 2862 -2460
rect 2856 -2472 2862 -2466
rect 2856 -2478 2862 -2472
rect 2856 -2484 2862 -2478
rect 2856 -2490 2862 -2484
rect 2856 -2496 2862 -2490
rect 2856 -2502 2862 -2496
rect 2856 -2508 2862 -2502
rect 2856 -2514 2862 -2508
rect 2856 -2520 2862 -2514
rect 2856 -2526 2862 -2520
rect 2856 -2532 2862 -2526
rect 2856 -2538 2862 -2532
rect 2856 -2544 2862 -2538
rect 2856 -2550 2862 -2544
rect 2856 -2556 2862 -2550
rect 2856 -2562 2862 -2556
rect 2856 -2568 2862 -2562
rect 2862 -1056 2868 -1050
rect 2862 -1062 2868 -1056
rect 2862 -1068 2868 -1062
rect 2862 -1074 2868 -1068
rect 2862 -1080 2868 -1074
rect 2862 -1086 2868 -1080
rect 2862 -1092 2868 -1086
rect 2862 -1098 2868 -1092
rect 2862 -1104 2868 -1098
rect 2862 -1110 2868 -1104
rect 2862 -1116 2868 -1110
rect 2862 -1122 2868 -1116
rect 2862 -1128 2868 -1122
rect 2862 -1134 2868 -1128
rect 2862 -1140 2868 -1134
rect 2862 -1146 2868 -1140
rect 2862 -1152 2868 -1146
rect 2862 -1158 2868 -1152
rect 2862 -1164 2868 -1158
rect 2862 -1170 2868 -1164
rect 2862 -1176 2868 -1170
rect 2862 -1182 2868 -1176
rect 2862 -1188 2868 -1182
rect 2862 -1194 2868 -1188
rect 2862 -1200 2868 -1194
rect 2862 -1206 2868 -1200
rect 2862 -1212 2868 -1206
rect 2862 -1218 2868 -1212
rect 2862 -1224 2868 -1218
rect 2862 -1230 2868 -1224
rect 2862 -1236 2868 -1230
rect 2862 -1242 2868 -1236
rect 2862 -1248 2868 -1242
rect 2862 -1254 2868 -1248
rect 2862 -1260 2868 -1254
rect 2862 -1266 2868 -1260
rect 2862 -1272 2868 -1266
rect 2862 -1278 2868 -1272
rect 2862 -1284 2868 -1278
rect 2862 -1290 2868 -1284
rect 2862 -1296 2868 -1290
rect 2862 -1302 2868 -1296
rect 2862 -1308 2868 -1302
rect 2862 -1314 2868 -1308
rect 2862 -1320 2868 -1314
rect 2862 -1326 2868 -1320
rect 2862 -1332 2868 -1326
rect 2862 -1338 2868 -1332
rect 2862 -1344 2868 -1338
rect 2862 -1350 2868 -1344
rect 2862 -1356 2868 -1350
rect 2862 -1362 2868 -1356
rect 2862 -1368 2868 -1362
rect 2862 -1374 2868 -1368
rect 2862 -1380 2868 -1374
rect 2862 -1386 2868 -1380
rect 2862 -1392 2868 -1386
rect 2862 -1398 2868 -1392
rect 2862 -1404 2868 -1398
rect 2862 -1410 2868 -1404
rect 2862 -1416 2868 -1410
rect 2862 -1422 2868 -1416
rect 2862 -1428 2868 -1422
rect 2862 -1434 2868 -1428
rect 2862 -1440 2868 -1434
rect 2862 -1446 2868 -1440
rect 2862 -1452 2868 -1446
rect 2862 -1458 2868 -1452
rect 2862 -1464 2868 -1458
rect 2862 -1470 2868 -1464
rect 2862 -2358 2868 -2352
rect 2862 -2364 2868 -2358
rect 2862 -2370 2868 -2364
rect 2862 -2376 2868 -2370
rect 2862 -2382 2868 -2376
rect 2862 -2388 2868 -2382
rect 2862 -2394 2868 -2388
rect 2862 -2400 2868 -2394
rect 2862 -2406 2868 -2400
rect 2862 -2412 2868 -2406
rect 2862 -2418 2868 -2412
rect 2862 -2424 2868 -2418
rect 2862 -2430 2868 -2424
rect 2862 -2436 2868 -2430
rect 2862 -2442 2868 -2436
rect 2862 -2448 2868 -2442
rect 2862 -2454 2868 -2448
rect 2862 -2460 2868 -2454
rect 2862 -2466 2868 -2460
rect 2862 -2472 2868 -2466
rect 2862 -2478 2868 -2472
rect 2862 -2484 2868 -2478
rect 2862 -2490 2868 -2484
rect 2862 -2496 2868 -2490
rect 2862 -2502 2868 -2496
rect 2862 -2508 2868 -2502
rect 2862 -2514 2868 -2508
rect 2862 -2520 2868 -2514
rect 2862 -2526 2868 -2520
rect 2862 -2532 2868 -2526
rect 2862 -2538 2868 -2532
rect 2862 -2544 2868 -2538
rect 2862 -2550 2868 -2544
rect 2862 -2556 2868 -2550
rect 2868 -1050 2874 -1044
rect 2868 -1056 2874 -1050
rect 2868 -1062 2874 -1056
rect 2868 -1068 2874 -1062
rect 2868 -1074 2874 -1068
rect 2868 -1080 2874 -1074
rect 2868 -1086 2874 -1080
rect 2868 -1092 2874 -1086
rect 2868 -1098 2874 -1092
rect 2868 -1104 2874 -1098
rect 2868 -1110 2874 -1104
rect 2868 -1116 2874 -1110
rect 2868 -1122 2874 -1116
rect 2868 -1128 2874 -1122
rect 2868 -1134 2874 -1128
rect 2868 -1140 2874 -1134
rect 2868 -1146 2874 -1140
rect 2868 -1152 2874 -1146
rect 2868 -1158 2874 -1152
rect 2868 -1164 2874 -1158
rect 2868 -1170 2874 -1164
rect 2868 -1176 2874 -1170
rect 2868 -1182 2874 -1176
rect 2868 -1188 2874 -1182
rect 2868 -1194 2874 -1188
rect 2868 -1200 2874 -1194
rect 2868 -1206 2874 -1200
rect 2868 -1212 2874 -1206
rect 2868 -1218 2874 -1212
rect 2868 -1224 2874 -1218
rect 2868 -1230 2874 -1224
rect 2868 -1236 2874 -1230
rect 2868 -1242 2874 -1236
rect 2868 -1248 2874 -1242
rect 2868 -1254 2874 -1248
rect 2868 -1260 2874 -1254
rect 2868 -1266 2874 -1260
rect 2868 -1272 2874 -1266
rect 2868 -1278 2874 -1272
rect 2868 -1284 2874 -1278
rect 2868 -1290 2874 -1284
rect 2868 -1296 2874 -1290
rect 2868 -1302 2874 -1296
rect 2868 -1308 2874 -1302
rect 2868 -1314 2874 -1308
rect 2868 -1320 2874 -1314
rect 2868 -1326 2874 -1320
rect 2868 -1332 2874 -1326
rect 2868 -1338 2874 -1332
rect 2868 -1344 2874 -1338
rect 2868 -1350 2874 -1344
rect 2868 -1356 2874 -1350
rect 2868 -1362 2874 -1356
rect 2868 -1368 2874 -1362
rect 2868 -1374 2874 -1368
rect 2868 -1380 2874 -1374
rect 2868 -1386 2874 -1380
rect 2868 -1392 2874 -1386
rect 2868 -1398 2874 -1392
rect 2868 -1404 2874 -1398
rect 2868 -1410 2874 -1404
rect 2868 -1416 2874 -1410
rect 2868 -1422 2874 -1416
rect 2868 -1428 2874 -1422
rect 2868 -1434 2874 -1428
rect 2868 -1440 2874 -1434
rect 2868 -1446 2874 -1440
rect 2868 -1452 2874 -1446
rect 2868 -1458 2874 -1452
rect 2868 -2358 2874 -2352
rect 2868 -2364 2874 -2358
rect 2868 -2370 2874 -2364
rect 2868 -2376 2874 -2370
rect 2868 -2382 2874 -2376
rect 2868 -2388 2874 -2382
rect 2868 -2394 2874 -2388
rect 2868 -2400 2874 -2394
rect 2868 -2406 2874 -2400
rect 2868 -2412 2874 -2406
rect 2868 -2418 2874 -2412
rect 2868 -2424 2874 -2418
rect 2868 -2430 2874 -2424
rect 2868 -2436 2874 -2430
rect 2868 -2442 2874 -2436
rect 2868 -2448 2874 -2442
rect 2868 -2454 2874 -2448
rect 2868 -2460 2874 -2454
rect 2868 -2466 2874 -2460
rect 2868 -2472 2874 -2466
rect 2868 -2478 2874 -2472
rect 2868 -2484 2874 -2478
rect 2868 -2490 2874 -2484
rect 2868 -2496 2874 -2490
rect 2868 -2502 2874 -2496
rect 2868 -2508 2874 -2502
rect 2868 -2514 2874 -2508
rect 2868 -2520 2874 -2514
rect 2868 -2526 2874 -2520
rect 2868 -2532 2874 -2526
rect 2868 -2538 2874 -2532
rect 2868 -2544 2874 -2538
rect 2868 -2550 2874 -2544
rect 2874 -1050 2880 -1044
rect 2874 -1056 2880 -1050
rect 2874 -1062 2880 -1056
rect 2874 -1068 2880 -1062
rect 2874 -1074 2880 -1068
rect 2874 -1080 2880 -1074
rect 2874 -1086 2880 -1080
rect 2874 -1092 2880 -1086
rect 2874 -1098 2880 -1092
rect 2874 -1104 2880 -1098
rect 2874 -1110 2880 -1104
rect 2874 -1116 2880 -1110
rect 2874 -1122 2880 -1116
rect 2874 -1128 2880 -1122
rect 2874 -1134 2880 -1128
rect 2874 -1140 2880 -1134
rect 2874 -1146 2880 -1140
rect 2874 -1152 2880 -1146
rect 2874 -1158 2880 -1152
rect 2874 -1164 2880 -1158
rect 2874 -1170 2880 -1164
rect 2874 -1176 2880 -1170
rect 2874 -1182 2880 -1176
rect 2874 -1188 2880 -1182
rect 2874 -1194 2880 -1188
rect 2874 -1200 2880 -1194
rect 2874 -1206 2880 -1200
rect 2874 -1212 2880 -1206
rect 2874 -1218 2880 -1212
rect 2874 -1224 2880 -1218
rect 2874 -1230 2880 -1224
rect 2874 -1236 2880 -1230
rect 2874 -1242 2880 -1236
rect 2874 -1248 2880 -1242
rect 2874 -1254 2880 -1248
rect 2874 -1260 2880 -1254
rect 2874 -1266 2880 -1260
rect 2874 -1272 2880 -1266
rect 2874 -1278 2880 -1272
rect 2874 -1284 2880 -1278
rect 2874 -1290 2880 -1284
rect 2874 -1296 2880 -1290
rect 2874 -1302 2880 -1296
rect 2874 -1308 2880 -1302
rect 2874 -1314 2880 -1308
rect 2874 -1320 2880 -1314
rect 2874 -1326 2880 -1320
rect 2874 -1332 2880 -1326
rect 2874 -1338 2880 -1332
rect 2874 -1344 2880 -1338
rect 2874 -1350 2880 -1344
rect 2874 -1356 2880 -1350
rect 2874 -1362 2880 -1356
rect 2874 -1368 2880 -1362
rect 2874 -1374 2880 -1368
rect 2874 -1380 2880 -1374
rect 2874 -1386 2880 -1380
rect 2874 -1392 2880 -1386
rect 2874 -1398 2880 -1392
rect 2874 -1404 2880 -1398
rect 2874 -1410 2880 -1404
rect 2874 -1416 2880 -1410
rect 2874 -1422 2880 -1416
rect 2874 -1428 2880 -1422
rect 2874 -1434 2880 -1428
rect 2874 -1440 2880 -1434
rect 2874 -1446 2880 -1440
rect 2874 -2352 2880 -2346
rect 2874 -2358 2880 -2352
rect 2874 -2364 2880 -2358
rect 2874 -2370 2880 -2364
rect 2874 -2376 2880 -2370
rect 2874 -2382 2880 -2376
rect 2874 -2388 2880 -2382
rect 2874 -2394 2880 -2388
rect 2874 -2400 2880 -2394
rect 2874 -2406 2880 -2400
rect 2874 -2412 2880 -2406
rect 2874 -2418 2880 -2412
rect 2874 -2424 2880 -2418
rect 2874 -2430 2880 -2424
rect 2874 -2436 2880 -2430
rect 2874 -2442 2880 -2436
rect 2874 -2448 2880 -2442
rect 2874 -2454 2880 -2448
rect 2874 -2460 2880 -2454
rect 2874 -2466 2880 -2460
rect 2874 -2472 2880 -2466
rect 2874 -2478 2880 -2472
rect 2874 -2484 2880 -2478
rect 2874 -2490 2880 -2484
rect 2874 -2496 2880 -2490
rect 2874 -2502 2880 -2496
rect 2874 -2508 2880 -2502
rect 2874 -2514 2880 -2508
rect 2874 -2520 2880 -2514
rect 2874 -2526 2880 -2520
rect 2874 -2532 2880 -2526
rect 2874 -2538 2880 -2532
rect 2874 -2544 2880 -2538
rect 2880 -1044 2886 -1038
rect 2880 -1050 2886 -1044
rect 2880 -1056 2886 -1050
rect 2880 -1062 2886 -1056
rect 2880 -1068 2886 -1062
rect 2880 -1074 2886 -1068
rect 2880 -1080 2886 -1074
rect 2880 -1086 2886 -1080
rect 2880 -1092 2886 -1086
rect 2880 -1098 2886 -1092
rect 2880 -1104 2886 -1098
rect 2880 -1110 2886 -1104
rect 2880 -1116 2886 -1110
rect 2880 -1122 2886 -1116
rect 2880 -1128 2886 -1122
rect 2880 -1134 2886 -1128
rect 2880 -1140 2886 -1134
rect 2880 -1146 2886 -1140
rect 2880 -1152 2886 -1146
rect 2880 -1158 2886 -1152
rect 2880 -1164 2886 -1158
rect 2880 -1170 2886 -1164
rect 2880 -1176 2886 -1170
rect 2880 -1182 2886 -1176
rect 2880 -1188 2886 -1182
rect 2880 -1194 2886 -1188
rect 2880 -1200 2886 -1194
rect 2880 -1206 2886 -1200
rect 2880 -1212 2886 -1206
rect 2880 -1218 2886 -1212
rect 2880 -1224 2886 -1218
rect 2880 -1230 2886 -1224
rect 2880 -1236 2886 -1230
rect 2880 -1242 2886 -1236
rect 2880 -1248 2886 -1242
rect 2880 -1254 2886 -1248
rect 2880 -1260 2886 -1254
rect 2880 -1266 2886 -1260
rect 2880 -1272 2886 -1266
rect 2880 -1278 2886 -1272
rect 2880 -1284 2886 -1278
rect 2880 -1290 2886 -1284
rect 2880 -1296 2886 -1290
rect 2880 -1302 2886 -1296
rect 2880 -1308 2886 -1302
rect 2880 -1314 2886 -1308
rect 2880 -1320 2886 -1314
rect 2880 -1326 2886 -1320
rect 2880 -1332 2886 -1326
rect 2880 -1338 2886 -1332
rect 2880 -1344 2886 -1338
rect 2880 -1350 2886 -1344
rect 2880 -1356 2886 -1350
rect 2880 -1362 2886 -1356
rect 2880 -1368 2886 -1362
rect 2880 -1374 2886 -1368
rect 2880 -1380 2886 -1374
rect 2880 -1386 2886 -1380
rect 2880 -1392 2886 -1386
rect 2880 -1398 2886 -1392
rect 2880 -1404 2886 -1398
rect 2880 -1410 2886 -1404
rect 2880 -1416 2886 -1410
rect 2880 -1422 2886 -1416
rect 2880 -1428 2886 -1422
rect 2880 -2352 2886 -2346
rect 2880 -2358 2886 -2352
rect 2880 -2364 2886 -2358
rect 2880 -2370 2886 -2364
rect 2880 -2376 2886 -2370
rect 2880 -2382 2886 -2376
rect 2880 -2388 2886 -2382
rect 2880 -2394 2886 -2388
rect 2880 -2400 2886 -2394
rect 2880 -2406 2886 -2400
rect 2880 -2412 2886 -2406
rect 2880 -2418 2886 -2412
rect 2880 -2424 2886 -2418
rect 2880 -2430 2886 -2424
rect 2880 -2436 2886 -2430
rect 2880 -2442 2886 -2436
rect 2880 -2448 2886 -2442
rect 2880 -2454 2886 -2448
rect 2880 -2460 2886 -2454
rect 2880 -2466 2886 -2460
rect 2880 -2472 2886 -2466
rect 2880 -2478 2886 -2472
rect 2880 -2484 2886 -2478
rect 2880 -2490 2886 -2484
rect 2880 -2496 2886 -2490
rect 2880 -2502 2886 -2496
rect 2880 -2508 2886 -2502
rect 2880 -2514 2886 -2508
rect 2880 -2520 2886 -2514
rect 2880 -2526 2886 -2520
rect 2880 -2532 2886 -2526
rect 2880 -2538 2886 -2532
rect 2886 -1038 2892 -1032
rect 2886 -1044 2892 -1038
rect 2886 -1050 2892 -1044
rect 2886 -1056 2892 -1050
rect 2886 -1062 2892 -1056
rect 2886 -1068 2892 -1062
rect 2886 -1074 2892 -1068
rect 2886 -1080 2892 -1074
rect 2886 -1086 2892 -1080
rect 2886 -1092 2892 -1086
rect 2886 -1098 2892 -1092
rect 2886 -1104 2892 -1098
rect 2886 -1110 2892 -1104
rect 2886 -1116 2892 -1110
rect 2886 -1122 2892 -1116
rect 2886 -1128 2892 -1122
rect 2886 -1134 2892 -1128
rect 2886 -1140 2892 -1134
rect 2886 -1146 2892 -1140
rect 2886 -1152 2892 -1146
rect 2886 -1158 2892 -1152
rect 2886 -1164 2892 -1158
rect 2886 -1170 2892 -1164
rect 2886 -1176 2892 -1170
rect 2886 -1182 2892 -1176
rect 2886 -1188 2892 -1182
rect 2886 -1194 2892 -1188
rect 2886 -1200 2892 -1194
rect 2886 -1206 2892 -1200
rect 2886 -1212 2892 -1206
rect 2886 -1218 2892 -1212
rect 2886 -1224 2892 -1218
rect 2886 -1230 2892 -1224
rect 2886 -1236 2892 -1230
rect 2886 -1242 2892 -1236
rect 2886 -1248 2892 -1242
rect 2886 -1254 2892 -1248
rect 2886 -1260 2892 -1254
rect 2886 -1266 2892 -1260
rect 2886 -1272 2892 -1266
rect 2886 -1278 2892 -1272
rect 2886 -1284 2892 -1278
rect 2886 -1290 2892 -1284
rect 2886 -1296 2892 -1290
rect 2886 -1302 2892 -1296
rect 2886 -1308 2892 -1302
rect 2886 -1314 2892 -1308
rect 2886 -1320 2892 -1314
rect 2886 -1326 2892 -1320
rect 2886 -1332 2892 -1326
rect 2886 -1338 2892 -1332
rect 2886 -1344 2892 -1338
rect 2886 -1350 2892 -1344
rect 2886 -1356 2892 -1350
rect 2886 -1362 2892 -1356
rect 2886 -1368 2892 -1362
rect 2886 -1374 2892 -1368
rect 2886 -1380 2892 -1374
rect 2886 -1386 2892 -1380
rect 2886 -1392 2892 -1386
rect 2886 -1398 2892 -1392
rect 2886 -1404 2892 -1398
rect 2886 -1410 2892 -1404
rect 2886 -1416 2892 -1410
rect 2886 -2352 2892 -2346
rect 2886 -2358 2892 -2352
rect 2886 -2364 2892 -2358
rect 2886 -2370 2892 -2364
rect 2886 -2376 2892 -2370
rect 2886 -2382 2892 -2376
rect 2886 -2388 2892 -2382
rect 2886 -2394 2892 -2388
rect 2886 -2400 2892 -2394
rect 2886 -2406 2892 -2400
rect 2886 -2412 2892 -2406
rect 2886 -2418 2892 -2412
rect 2886 -2424 2892 -2418
rect 2886 -2430 2892 -2424
rect 2886 -2436 2892 -2430
rect 2886 -2442 2892 -2436
rect 2886 -2448 2892 -2442
rect 2886 -2454 2892 -2448
rect 2886 -2460 2892 -2454
rect 2886 -2466 2892 -2460
rect 2886 -2472 2892 -2466
rect 2886 -2478 2892 -2472
rect 2886 -2484 2892 -2478
rect 2886 -2490 2892 -2484
rect 2886 -2496 2892 -2490
rect 2886 -2502 2892 -2496
rect 2886 -2508 2892 -2502
rect 2886 -2514 2892 -2508
rect 2886 -2520 2892 -2514
rect 2886 -2526 2892 -2520
rect 2886 -2532 2892 -2526
rect 2892 -1038 2898 -1032
rect 2892 -1044 2898 -1038
rect 2892 -1050 2898 -1044
rect 2892 -1056 2898 -1050
rect 2892 -1062 2898 -1056
rect 2892 -1068 2898 -1062
rect 2892 -1074 2898 -1068
rect 2892 -1080 2898 -1074
rect 2892 -1086 2898 -1080
rect 2892 -1092 2898 -1086
rect 2892 -1098 2898 -1092
rect 2892 -1104 2898 -1098
rect 2892 -1110 2898 -1104
rect 2892 -1116 2898 -1110
rect 2892 -1122 2898 -1116
rect 2892 -1128 2898 -1122
rect 2892 -1134 2898 -1128
rect 2892 -1140 2898 -1134
rect 2892 -1146 2898 -1140
rect 2892 -1152 2898 -1146
rect 2892 -1158 2898 -1152
rect 2892 -1164 2898 -1158
rect 2892 -1170 2898 -1164
rect 2892 -1176 2898 -1170
rect 2892 -1182 2898 -1176
rect 2892 -1188 2898 -1182
rect 2892 -1194 2898 -1188
rect 2892 -1200 2898 -1194
rect 2892 -1206 2898 -1200
rect 2892 -1212 2898 -1206
rect 2892 -1218 2898 -1212
rect 2892 -1224 2898 -1218
rect 2892 -1230 2898 -1224
rect 2892 -1236 2898 -1230
rect 2892 -1242 2898 -1236
rect 2892 -1248 2898 -1242
rect 2892 -1254 2898 -1248
rect 2892 -1260 2898 -1254
rect 2892 -1266 2898 -1260
rect 2892 -1272 2898 -1266
rect 2892 -1278 2898 -1272
rect 2892 -1284 2898 -1278
rect 2892 -1290 2898 -1284
rect 2892 -1296 2898 -1290
rect 2892 -1302 2898 -1296
rect 2892 -1308 2898 -1302
rect 2892 -1314 2898 -1308
rect 2892 -1320 2898 -1314
rect 2892 -1326 2898 -1320
rect 2892 -1332 2898 -1326
rect 2892 -1338 2898 -1332
rect 2892 -1344 2898 -1338
rect 2892 -1350 2898 -1344
rect 2892 -1356 2898 -1350
rect 2892 -1362 2898 -1356
rect 2892 -1368 2898 -1362
rect 2892 -1374 2898 -1368
rect 2892 -1380 2898 -1374
rect 2892 -1386 2898 -1380
rect 2892 -1392 2898 -1386
rect 2892 -1398 2898 -1392
rect 2892 -1404 2898 -1398
rect 2892 -2352 2898 -2346
rect 2892 -2358 2898 -2352
rect 2892 -2364 2898 -2358
rect 2892 -2370 2898 -2364
rect 2892 -2376 2898 -2370
rect 2892 -2382 2898 -2376
rect 2892 -2388 2898 -2382
rect 2892 -2394 2898 -2388
rect 2892 -2400 2898 -2394
rect 2892 -2406 2898 -2400
rect 2892 -2412 2898 -2406
rect 2892 -2418 2898 -2412
rect 2892 -2424 2898 -2418
rect 2892 -2430 2898 -2424
rect 2892 -2436 2898 -2430
rect 2892 -2442 2898 -2436
rect 2892 -2448 2898 -2442
rect 2892 -2454 2898 -2448
rect 2892 -2460 2898 -2454
rect 2892 -2466 2898 -2460
rect 2892 -2472 2898 -2466
rect 2892 -2478 2898 -2472
rect 2892 -2484 2898 -2478
rect 2892 -2490 2898 -2484
rect 2892 -2496 2898 -2490
rect 2892 -2502 2898 -2496
rect 2892 -2508 2898 -2502
rect 2892 -2514 2898 -2508
rect 2892 -2520 2898 -2514
rect 2898 -1032 2904 -1026
rect 2898 -1038 2904 -1032
rect 2898 -1044 2904 -1038
rect 2898 -1050 2904 -1044
rect 2898 -1056 2904 -1050
rect 2898 -1062 2904 -1056
rect 2898 -1068 2904 -1062
rect 2898 -1074 2904 -1068
rect 2898 -1080 2904 -1074
rect 2898 -1086 2904 -1080
rect 2898 -1092 2904 -1086
rect 2898 -1098 2904 -1092
rect 2898 -1104 2904 -1098
rect 2898 -1110 2904 -1104
rect 2898 -1116 2904 -1110
rect 2898 -1122 2904 -1116
rect 2898 -1128 2904 -1122
rect 2898 -1134 2904 -1128
rect 2898 -1140 2904 -1134
rect 2898 -1146 2904 -1140
rect 2898 -1152 2904 -1146
rect 2898 -1158 2904 -1152
rect 2898 -1164 2904 -1158
rect 2898 -1170 2904 -1164
rect 2898 -1176 2904 -1170
rect 2898 -1182 2904 -1176
rect 2898 -1188 2904 -1182
rect 2898 -1194 2904 -1188
rect 2898 -1200 2904 -1194
rect 2898 -1206 2904 -1200
rect 2898 -1212 2904 -1206
rect 2898 -1218 2904 -1212
rect 2898 -1224 2904 -1218
rect 2898 -1230 2904 -1224
rect 2898 -1236 2904 -1230
rect 2898 -1242 2904 -1236
rect 2898 -1248 2904 -1242
rect 2898 -1254 2904 -1248
rect 2898 -1260 2904 -1254
rect 2898 -1266 2904 -1260
rect 2898 -1272 2904 -1266
rect 2898 -1278 2904 -1272
rect 2898 -1284 2904 -1278
rect 2898 -1290 2904 -1284
rect 2898 -1296 2904 -1290
rect 2898 -1302 2904 -1296
rect 2898 -1308 2904 -1302
rect 2898 -1314 2904 -1308
rect 2898 -1320 2904 -1314
rect 2898 -1326 2904 -1320
rect 2898 -1332 2904 -1326
rect 2898 -1338 2904 -1332
rect 2898 -1344 2904 -1338
rect 2898 -1350 2904 -1344
rect 2898 -1356 2904 -1350
rect 2898 -1362 2904 -1356
rect 2898 -1368 2904 -1362
rect 2898 -1374 2904 -1368
rect 2898 -1380 2904 -1374
rect 2898 -2352 2904 -2346
rect 2898 -2358 2904 -2352
rect 2898 -2364 2904 -2358
rect 2898 -2370 2904 -2364
rect 2898 -2376 2904 -2370
rect 2898 -2382 2904 -2376
rect 2898 -2388 2904 -2382
rect 2898 -2394 2904 -2388
rect 2898 -2400 2904 -2394
rect 2898 -2406 2904 -2400
rect 2898 -2412 2904 -2406
rect 2898 -2418 2904 -2412
rect 2898 -2424 2904 -2418
rect 2898 -2430 2904 -2424
rect 2898 -2436 2904 -2430
rect 2898 -2442 2904 -2436
rect 2898 -2448 2904 -2442
rect 2898 -2454 2904 -2448
rect 2898 -2460 2904 -2454
rect 2898 -2466 2904 -2460
rect 2898 -2472 2904 -2466
rect 2898 -2478 2904 -2472
rect 2898 -2484 2904 -2478
rect 2898 -2490 2904 -2484
rect 2898 -2496 2904 -2490
rect 2898 -2502 2904 -2496
rect 2898 -2508 2904 -2502
rect 2898 -2514 2904 -2508
rect 2904 -1026 2910 -1020
rect 2904 -1032 2910 -1026
rect 2904 -1038 2910 -1032
rect 2904 -1044 2910 -1038
rect 2904 -1050 2910 -1044
rect 2904 -1056 2910 -1050
rect 2904 -1062 2910 -1056
rect 2904 -1068 2910 -1062
rect 2904 -1074 2910 -1068
rect 2904 -1080 2910 -1074
rect 2904 -1086 2910 -1080
rect 2904 -1092 2910 -1086
rect 2904 -1098 2910 -1092
rect 2904 -1104 2910 -1098
rect 2904 -1110 2910 -1104
rect 2904 -1116 2910 -1110
rect 2904 -1122 2910 -1116
rect 2904 -1128 2910 -1122
rect 2904 -1134 2910 -1128
rect 2904 -1140 2910 -1134
rect 2904 -1146 2910 -1140
rect 2904 -1152 2910 -1146
rect 2904 -1158 2910 -1152
rect 2904 -1164 2910 -1158
rect 2904 -1170 2910 -1164
rect 2904 -1176 2910 -1170
rect 2904 -1182 2910 -1176
rect 2904 -1188 2910 -1182
rect 2904 -1194 2910 -1188
rect 2904 -1200 2910 -1194
rect 2904 -1206 2910 -1200
rect 2904 -1212 2910 -1206
rect 2904 -1218 2910 -1212
rect 2904 -1224 2910 -1218
rect 2904 -1230 2910 -1224
rect 2904 -1236 2910 -1230
rect 2904 -1242 2910 -1236
rect 2904 -1248 2910 -1242
rect 2904 -1254 2910 -1248
rect 2904 -1260 2910 -1254
rect 2904 -1266 2910 -1260
rect 2904 -1272 2910 -1266
rect 2904 -1278 2910 -1272
rect 2904 -1284 2910 -1278
rect 2904 -1290 2910 -1284
rect 2904 -1296 2910 -1290
rect 2904 -1302 2910 -1296
rect 2904 -1308 2910 -1302
rect 2904 -1314 2910 -1308
rect 2904 -1320 2910 -1314
rect 2904 -1326 2910 -1320
rect 2904 -1332 2910 -1326
rect 2904 -1338 2910 -1332
rect 2904 -1344 2910 -1338
rect 2904 -1350 2910 -1344
rect 2904 -1356 2910 -1350
rect 2904 -2346 2910 -2340
rect 2904 -2352 2910 -2346
rect 2904 -2358 2910 -2352
rect 2904 -2364 2910 -2358
rect 2904 -2370 2910 -2364
rect 2904 -2376 2910 -2370
rect 2904 -2382 2910 -2376
rect 2904 -2388 2910 -2382
rect 2904 -2394 2910 -2388
rect 2904 -2400 2910 -2394
rect 2904 -2406 2910 -2400
rect 2904 -2412 2910 -2406
rect 2904 -2418 2910 -2412
rect 2904 -2424 2910 -2418
rect 2904 -2430 2910 -2424
rect 2904 -2436 2910 -2430
rect 2904 -2442 2910 -2436
rect 2904 -2448 2910 -2442
rect 2904 -2454 2910 -2448
rect 2904 -2460 2910 -2454
rect 2904 -2466 2910 -2460
rect 2904 -2472 2910 -2466
rect 2904 -2478 2910 -2472
rect 2904 -2484 2910 -2478
rect 2904 -2490 2910 -2484
rect 2904 -2496 2910 -2490
rect 2904 -2502 2910 -2496
rect 2904 -2508 2910 -2502
rect 2910 -1026 2916 -1020
rect 2910 -1032 2916 -1026
rect 2910 -1038 2916 -1032
rect 2910 -1044 2916 -1038
rect 2910 -1050 2916 -1044
rect 2910 -1056 2916 -1050
rect 2910 -1062 2916 -1056
rect 2910 -1068 2916 -1062
rect 2910 -1074 2916 -1068
rect 2910 -1080 2916 -1074
rect 2910 -1086 2916 -1080
rect 2910 -1092 2916 -1086
rect 2910 -1098 2916 -1092
rect 2910 -1104 2916 -1098
rect 2910 -1110 2916 -1104
rect 2910 -1116 2916 -1110
rect 2910 -1122 2916 -1116
rect 2910 -1128 2916 -1122
rect 2910 -1134 2916 -1128
rect 2910 -1140 2916 -1134
rect 2910 -1146 2916 -1140
rect 2910 -1152 2916 -1146
rect 2910 -1158 2916 -1152
rect 2910 -1164 2916 -1158
rect 2910 -1170 2916 -1164
rect 2910 -1176 2916 -1170
rect 2910 -1182 2916 -1176
rect 2910 -1188 2916 -1182
rect 2910 -1194 2916 -1188
rect 2910 -1200 2916 -1194
rect 2910 -1206 2916 -1200
rect 2910 -1212 2916 -1206
rect 2910 -1218 2916 -1212
rect 2910 -1224 2916 -1218
rect 2910 -1230 2916 -1224
rect 2910 -1236 2916 -1230
rect 2910 -1242 2916 -1236
rect 2910 -1248 2916 -1242
rect 2910 -1254 2916 -1248
rect 2910 -1260 2916 -1254
rect 2910 -1266 2916 -1260
rect 2910 -1272 2916 -1266
rect 2910 -1278 2916 -1272
rect 2910 -1284 2916 -1278
rect 2910 -1290 2916 -1284
rect 2910 -1296 2916 -1290
rect 2910 -1302 2916 -1296
rect 2910 -1308 2916 -1302
rect 2910 -1314 2916 -1308
rect 2910 -1320 2916 -1314
rect 2910 -1326 2916 -1320
rect 2910 -1332 2916 -1326
rect 2910 -2346 2916 -2340
rect 2910 -2352 2916 -2346
rect 2910 -2358 2916 -2352
rect 2910 -2364 2916 -2358
rect 2910 -2370 2916 -2364
rect 2910 -2376 2916 -2370
rect 2910 -2382 2916 -2376
rect 2910 -2388 2916 -2382
rect 2910 -2394 2916 -2388
rect 2910 -2400 2916 -2394
rect 2910 -2406 2916 -2400
rect 2910 -2412 2916 -2406
rect 2910 -2418 2916 -2412
rect 2910 -2424 2916 -2418
rect 2910 -2430 2916 -2424
rect 2910 -2436 2916 -2430
rect 2910 -2442 2916 -2436
rect 2910 -2448 2916 -2442
rect 2910 -2454 2916 -2448
rect 2910 -2460 2916 -2454
rect 2910 -2466 2916 -2460
rect 2910 -2472 2916 -2466
rect 2910 -2478 2916 -2472
rect 2910 -2484 2916 -2478
rect 2910 -2490 2916 -2484
rect 2910 -2496 2916 -2490
rect 2910 -2502 2916 -2496
rect 2916 -1020 2922 -1014
rect 2916 -1026 2922 -1020
rect 2916 -1032 2922 -1026
rect 2916 -1038 2922 -1032
rect 2916 -1044 2922 -1038
rect 2916 -1050 2922 -1044
rect 2916 -1056 2922 -1050
rect 2916 -1062 2922 -1056
rect 2916 -1068 2922 -1062
rect 2916 -1074 2922 -1068
rect 2916 -1080 2922 -1074
rect 2916 -1086 2922 -1080
rect 2916 -1092 2922 -1086
rect 2916 -1098 2922 -1092
rect 2916 -1104 2922 -1098
rect 2916 -1110 2922 -1104
rect 2916 -1116 2922 -1110
rect 2916 -1122 2922 -1116
rect 2916 -1128 2922 -1122
rect 2916 -1134 2922 -1128
rect 2916 -1140 2922 -1134
rect 2916 -1146 2922 -1140
rect 2916 -1152 2922 -1146
rect 2916 -1158 2922 -1152
rect 2916 -1164 2922 -1158
rect 2916 -1170 2922 -1164
rect 2916 -1176 2922 -1170
rect 2916 -1182 2922 -1176
rect 2916 -1188 2922 -1182
rect 2916 -1194 2922 -1188
rect 2916 -1200 2922 -1194
rect 2916 -1206 2922 -1200
rect 2916 -1212 2922 -1206
rect 2916 -1218 2922 -1212
rect 2916 -1224 2922 -1218
rect 2916 -1230 2922 -1224
rect 2916 -1236 2922 -1230
rect 2916 -1242 2922 -1236
rect 2916 -1248 2922 -1242
rect 2916 -1254 2922 -1248
rect 2916 -1260 2922 -1254
rect 2916 -1266 2922 -1260
rect 2916 -1272 2922 -1266
rect 2916 -1278 2922 -1272
rect 2916 -1284 2922 -1278
rect 2916 -1290 2922 -1284
rect 2916 -1296 2922 -1290
rect 2916 -1302 2922 -1296
rect 2916 -2346 2922 -2340
rect 2916 -2352 2922 -2346
rect 2916 -2358 2922 -2352
rect 2916 -2364 2922 -2358
rect 2916 -2370 2922 -2364
rect 2916 -2376 2922 -2370
rect 2916 -2382 2922 -2376
rect 2916 -2388 2922 -2382
rect 2916 -2394 2922 -2388
rect 2916 -2400 2922 -2394
rect 2916 -2406 2922 -2400
rect 2916 -2412 2922 -2406
rect 2916 -2418 2922 -2412
rect 2916 -2424 2922 -2418
rect 2916 -2430 2922 -2424
rect 2916 -2436 2922 -2430
rect 2916 -2442 2922 -2436
rect 2916 -2448 2922 -2442
rect 2916 -2454 2922 -2448
rect 2916 -2460 2922 -2454
rect 2916 -2466 2922 -2460
rect 2916 -2472 2922 -2466
rect 2916 -2478 2922 -2472
rect 2916 -2484 2922 -2478
rect 2916 -2490 2922 -2484
rect 2922 -1014 2928 -1008
rect 2922 -1020 2928 -1014
rect 2922 -1026 2928 -1020
rect 2922 -1032 2928 -1026
rect 2922 -1038 2928 -1032
rect 2922 -1044 2928 -1038
rect 2922 -1050 2928 -1044
rect 2922 -1056 2928 -1050
rect 2922 -1062 2928 -1056
rect 2922 -1068 2928 -1062
rect 2922 -1074 2928 -1068
rect 2922 -1080 2928 -1074
rect 2922 -1086 2928 -1080
rect 2922 -1092 2928 -1086
rect 2922 -1098 2928 -1092
rect 2922 -1104 2928 -1098
rect 2922 -1110 2928 -1104
rect 2922 -1116 2928 -1110
rect 2922 -1122 2928 -1116
rect 2922 -1128 2928 -1122
rect 2922 -1134 2928 -1128
rect 2922 -1140 2928 -1134
rect 2922 -1146 2928 -1140
rect 2922 -1152 2928 -1146
rect 2922 -1158 2928 -1152
rect 2922 -1164 2928 -1158
rect 2922 -1170 2928 -1164
rect 2922 -1176 2928 -1170
rect 2922 -1182 2928 -1176
rect 2922 -1188 2928 -1182
rect 2922 -1194 2928 -1188
rect 2922 -1200 2928 -1194
rect 2922 -1206 2928 -1200
rect 2922 -1212 2928 -1206
rect 2922 -1218 2928 -1212
rect 2922 -1224 2928 -1218
rect 2922 -1230 2928 -1224
rect 2922 -1236 2928 -1230
rect 2922 -1242 2928 -1236
rect 2922 -1248 2928 -1242
rect 2922 -1254 2928 -1248
rect 2922 -2346 2928 -2340
rect 2922 -2352 2928 -2346
rect 2922 -2358 2928 -2352
rect 2922 -2364 2928 -2358
rect 2922 -2370 2928 -2364
rect 2922 -2376 2928 -2370
rect 2922 -2382 2928 -2376
rect 2922 -2388 2928 -2382
rect 2922 -2394 2928 -2388
rect 2922 -2400 2928 -2394
rect 2922 -2406 2928 -2400
rect 2922 -2412 2928 -2406
rect 2922 -2418 2928 -2412
rect 2922 -2424 2928 -2418
rect 2922 -2430 2928 -2424
rect 2922 -2436 2928 -2430
rect 2922 -2442 2928 -2436
rect 2922 -2448 2928 -2442
rect 2922 -2454 2928 -2448
rect 2922 -2460 2928 -2454
rect 2922 -2466 2928 -2460
rect 2922 -2472 2928 -2466
rect 2922 -2478 2928 -2472
rect 2928 -2340 2934 -2334
rect 2928 -2346 2934 -2340
rect 2928 -2352 2934 -2346
rect 2928 -2358 2934 -2352
rect 2928 -2364 2934 -2358
rect 2928 -2370 2934 -2364
rect 2928 -2376 2934 -2370
rect 2928 -2382 2934 -2376
rect 2928 -2388 2934 -2382
rect 2928 -2394 2934 -2388
rect 2928 -2400 2934 -2394
rect 2928 -2406 2934 -2400
rect 2928 -2412 2934 -2406
rect 2928 -2418 2934 -2412
rect 2928 -2424 2934 -2418
rect 2928 -2430 2934 -2424
rect 2928 -2436 2934 -2430
rect 2928 -2442 2934 -2436
rect 2928 -2448 2934 -2442
rect 2928 -2454 2934 -2448
rect 2928 -2460 2934 -2454
rect 2928 -2466 2934 -2460
rect 2928 -2472 2934 -2466
rect 2934 -2340 2940 -2334
rect 2934 -2346 2940 -2340
rect 2934 -2352 2940 -2346
rect 2934 -2358 2940 -2352
rect 2934 -2364 2940 -2358
rect 2934 -2370 2940 -2364
rect 2934 -2376 2940 -2370
rect 2934 -2382 2940 -2376
rect 2934 -2388 2940 -2382
rect 2934 -2394 2940 -2388
rect 2934 -2400 2940 -2394
rect 2934 -2406 2940 -2400
rect 2934 -2412 2940 -2406
rect 2934 -2418 2940 -2412
rect 2934 -2424 2940 -2418
rect 2934 -2430 2940 -2424
rect 2934 -2436 2940 -2430
rect 2934 -2442 2940 -2436
rect 2934 -2448 2940 -2442
rect 2934 -2454 2940 -2448
rect 2934 -2460 2940 -2454
rect 2940 -2340 2946 -2334
rect 2940 -2346 2946 -2340
rect 2940 -2352 2946 -2346
rect 2940 -2358 2946 -2352
rect 2940 -2364 2946 -2358
rect 2940 -2370 2946 -2364
rect 2940 -2376 2946 -2370
rect 2940 -2382 2946 -2376
rect 2940 -2388 2946 -2382
rect 2940 -2394 2946 -2388
rect 2940 -2400 2946 -2394
rect 2940 -2406 2946 -2400
rect 2940 -2412 2946 -2406
rect 2940 -2418 2946 -2412
rect 2940 -2424 2946 -2418
rect 2940 -2430 2946 -2424
rect 2940 -2436 2946 -2430
rect 2940 -2442 2946 -2436
rect 2940 -2448 2946 -2442
rect 2946 -2340 2952 -2334
rect 2946 -2346 2952 -2340
rect 2946 -2352 2952 -2346
rect 2946 -2358 2952 -2352
rect 2946 -2364 2952 -2358
rect 2946 -2370 2952 -2364
rect 2946 -2376 2952 -2370
rect 2946 -2382 2952 -2376
rect 2946 -2388 2952 -2382
rect 2946 -2394 2952 -2388
rect 2946 -2400 2952 -2394
rect 2946 -2406 2952 -2400
rect 2946 -2412 2952 -2406
rect 2946 -2418 2952 -2412
rect 2946 -2424 2952 -2418
rect 2946 -2430 2952 -2424
rect 2946 -2436 2952 -2430
rect 2952 -2334 2958 -2328
rect 2952 -2340 2958 -2334
rect 2952 -2346 2958 -2340
rect 2952 -2352 2958 -2346
rect 2952 -2358 2958 -2352
rect 2952 -2364 2958 -2358
rect 2952 -2370 2958 -2364
rect 2952 -2376 2958 -2370
rect 2952 -2382 2958 -2376
rect 2952 -2388 2958 -2382
rect 2952 -2394 2958 -2388
rect 2952 -2400 2958 -2394
rect 2952 -2406 2958 -2400
rect 2952 -2412 2958 -2406
rect 2952 -2418 2958 -2412
rect 2952 -2424 2958 -2418
rect 2958 -2334 2964 -2328
rect 2958 -2340 2964 -2334
rect 2958 -2346 2964 -2340
rect 2958 -2352 2964 -2346
rect 2958 -2358 2964 -2352
rect 2958 -2364 2964 -2358
rect 2958 -2370 2964 -2364
rect 2958 -2376 2964 -2370
rect 2958 -2382 2964 -2376
rect 2958 -2388 2964 -2382
rect 2958 -2394 2964 -2388
rect 2958 -2400 2964 -2394
rect 2958 -2406 2964 -2400
rect 2958 -2412 2964 -2406
rect 2964 -2334 2970 -2328
rect 2964 -2340 2970 -2334
rect 2964 -2346 2970 -2340
rect 2964 -2352 2970 -2346
rect 2964 -2358 2970 -2352
rect 2964 -2364 2970 -2358
rect 2964 -2370 2970 -2364
rect 2964 -2376 2970 -2370
rect 2964 -2382 2970 -2376
rect 2964 -2388 2970 -2382
rect 2964 -2394 2970 -2388
rect 2964 -2400 2970 -2394
rect 2970 -2334 2976 -2328
rect 2970 -2340 2976 -2334
rect 2970 -2346 2976 -2340
rect 2970 -2352 2976 -2346
rect 2970 -2358 2976 -2352
rect 2970 -2364 2976 -2358
rect 2970 -2370 2976 -2364
rect 2970 -2376 2976 -2370
rect 2970 -2382 2976 -2376
rect 2970 -2388 2976 -2382
rect 2976 -2328 2982 -2322
rect 2976 -2334 2982 -2328
rect 2976 -2340 2982 -2334
rect 2976 -2346 2982 -2340
rect 2976 -2352 2982 -2346
rect 2976 -2358 2982 -2352
rect 2976 -2364 2982 -2358
rect 2976 -2370 2982 -2364
rect 2982 -2328 2988 -2322
rect 2982 -2334 2988 -2328
rect 2982 -2340 2988 -2334
rect 2982 -2346 2988 -2340
rect 2982 -2352 2988 -2346
rect 2982 -2358 2988 -2352
rect 2988 -2328 2994 -2322
rect 2988 -2334 2994 -2328
rect 2988 -2340 2994 -2334
rect 2994 -2328 3000 -2322
<< end >>
