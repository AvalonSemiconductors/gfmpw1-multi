magic
tech gf180mcuD
magscale 1 10
timestamp 1702379971
<< nwell >>
rect 1258 19168 22710 20032
rect 1258 17600 22710 18464
rect 1258 16032 22710 16896
rect 1258 14464 22710 15328
rect 1258 12896 22710 13760
rect 1258 11328 22710 12192
rect 1258 10599 13207 10624
rect 1258 9760 22710 10599
rect 1258 8217 22710 9056
rect 1258 8192 6032 8217
rect 1258 6624 22710 7488
rect 1258 5056 22710 5920
rect 1258 3488 22710 4352
<< pwell >>
rect 1258 20032 22710 20470
rect 1258 18464 22710 19168
rect 1258 16896 22710 17600
rect 1258 15328 22710 16032
rect 1258 13760 22710 14464
rect 1258 12192 22710 12896
rect 1258 10624 22710 11328
rect 1258 9056 22710 9760
rect 1258 7488 22710 8192
rect 1258 5920 22710 6624
rect 1258 4352 22710 5056
rect 1258 3050 22710 3488
<< obsm1 >>
rect 1344 3076 22784 20444
<< metal2 >>
rect 1792 23200 1904 24000
rect 4032 23200 4144 24000
rect 6272 23200 6384 24000
rect 8512 23200 8624 24000
rect 10752 23200 10864 24000
rect 12992 23200 13104 24000
rect 15232 23200 15344 24000
rect 17472 23200 17584 24000
rect 19712 23200 19824 24000
rect 21952 23200 22064 24000
<< obsm2 >>
rect 1964 23140 3972 23268
rect 4204 23140 6212 23268
rect 6444 23140 8452 23268
rect 8684 23140 10692 23268
rect 10924 23140 12932 23268
rect 13164 23140 15172 23268
rect 15404 23140 17412 23268
rect 17644 23140 19652 23268
rect 19884 23140 21892 23268
rect 22124 23140 22756 23268
rect 1820 1586 22756 23140
<< metal3 >>
rect 23200 21952 24000 22064
rect 23200 19040 24000 19152
rect 23200 16128 24000 16240
rect 23200 13216 24000 13328
rect 23200 10304 24000 10416
rect 23200 7392 24000 7504
rect 23200 4480 24000 4592
rect 23200 1568 24000 1680
<< obsm3 >>
rect 2258 21892 23140 22036
rect 2258 19212 23200 21892
rect 2258 18980 23140 19212
rect 2258 16300 23200 18980
rect 2258 16068 23140 16300
rect 2258 13388 23200 16068
rect 2258 13156 23140 13388
rect 2258 10476 23200 13156
rect 2258 10244 23140 10476
rect 2258 7564 23200 10244
rect 2258 7332 23140 7564
rect 2258 4652 23200 7332
rect 2258 4420 23140 4652
rect 2258 1740 23200 4420
rect 2258 1596 23140 1740
<< metal4 >>
rect 3844 3076 4164 20444
rect 6504 3076 6824 20444
rect 9164 3076 9484 20444
rect 11824 3076 12144 20444
rect 14484 3076 14804 20444
rect 17144 3076 17464 20444
rect 19804 3076 20124 20444
rect 22464 3076 22784 20444
<< obsm4 >>
rect 4396 11890 6444 18462
rect 6884 11890 9104 18462
rect 9544 11890 11764 18462
rect 12204 11890 14424 18462
rect 14864 11890 17084 18462
rect 17524 11890 19744 18462
rect 20184 11890 20244 18462
<< labels >>
rlabel metal3 s 23200 1568 24000 1680 6 clk
port 1 nsew signal input
rlabel metal3 s 23200 7392 24000 7504 6 io_in[0]
port 2 nsew signal input
rlabel metal3 s 23200 10304 24000 10416 6 io_in[1]
port 3 nsew signal input
rlabel metal3 s 23200 13216 24000 13328 6 io_in[2]
port 4 nsew signal input
rlabel metal3 s 23200 16128 24000 16240 6 io_in[3]
port 5 nsew signal input
rlabel metal3 s 23200 19040 24000 19152 6 io_in[4]
port 6 nsew signal input
rlabel metal3 s 23200 21952 24000 22064 6 io_oeb
port 7 nsew signal output
rlabel metal2 s 1792 23200 1904 24000 6 io_out[0]
port 8 nsew signal output
rlabel metal2 s 4032 23200 4144 24000 6 io_out[1]
port 9 nsew signal output
rlabel metal2 s 6272 23200 6384 24000 6 io_out[2]
port 10 nsew signal output
rlabel metal2 s 8512 23200 8624 24000 6 io_out[3]
port 11 nsew signal output
rlabel metal2 s 10752 23200 10864 24000 6 io_out[4]
port 12 nsew signal output
rlabel metal2 s 12992 23200 13104 24000 6 io_out[5]
port 13 nsew signal output
rlabel metal2 s 15232 23200 15344 24000 6 io_out[6]
port 14 nsew signal output
rlabel metal2 s 17472 23200 17584 24000 6 io_out[7]
port 15 nsew signal output
rlabel metal2 s 19712 23200 19824 24000 6 io_out[8]
port 16 nsew signal output
rlabel metal2 s 21952 23200 22064 24000 6 io_out[9]
port 17 nsew signal output
rlabel metal3 s 23200 4480 24000 4592 6 rst_n
port 18 nsew signal input
rlabel metal4 s 3844 3076 4164 20444 6 vdd
port 19 nsew power bidirectional
rlabel metal4 s 9164 3076 9484 20444 6 vdd
port 19 nsew power bidirectional
rlabel metal4 s 14484 3076 14804 20444 6 vdd
port 19 nsew power bidirectional
rlabel metal4 s 19804 3076 20124 20444 6 vdd
port 19 nsew power bidirectional
rlabel metal4 s 6504 3076 6824 20444 6 vss
port 20 nsew ground bidirectional
rlabel metal4 s 11824 3076 12144 20444 6 vss
port 20 nsew ground bidirectional
rlabel metal4 s 17144 3076 17464 20444 6 vss
port 20 nsew ground bidirectional
rlabel metal4 s 22464 3076 22784 20444 6 vss
port 20 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 24000 24000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 422560
string GDS_FILE /media/lucah/fbc90f8f-67e9-406d-9872-54f02ad6a2d8/gfmpw1-multi/openlane/ue1/runs/23_12_12_12_11/results/signoff/ue1.magic.gds
string GDS_START 126424
<< end >>

