VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO wrapped_tholin_riscv
  CLASS BLOCK ;
  FOREIGN wrapped_tholin_riscv ;
  ORIGIN 0.000 0.000 ;
  SIZE 1225.000 BY 1225.000 ;
  PIN custom_settings[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 91.840 4.000 92.400 ;
    END
  END custom_settings[0]
  PIN custom_settings[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 124.320 4.000 124.880 ;
    END
  END custom_settings[1]
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 156.800 4.000 157.360 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.588000 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 481.600 4.000 482.160 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.588000 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 514.080 4.000 514.640 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 546.560 4.000 547.120 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.588000 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 579.040 4.000 579.600 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.588000 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 611.520 4.000 612.080 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 644.000 4.000 644.560 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 676.480 4.000 677.040 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 708.960 4.000 709.520 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 741.440 4.000 742.000 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 773.920 4.000 774.480 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 189.280 4.000 189.840 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 806.400 4.000 806.960 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 838.880 4.000 839.440 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 871.360 4.000 871.920 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 903.840 4.000 904.400 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 936.320 4.000 936.880 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 968.800 4.000 969.360 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1001.280 4.000 1001.840 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1033.760 4.000 1034.320 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1066.240 4.000 1066.800 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1098.720 4.000 1099.280 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 221.760 4.000 222.320 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1131.200 4.000 1131.760 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1163.680 4.000 1164.240 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1196.160 4.000 1196.720 ;
    END
  END io_in[32]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.588000 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 254.240 4.000 254.800 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.588000 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 286.720 4.000 287.280 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.588000 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 319.200 4.000 319.760 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.666400 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 351.680 4.000 352.240 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.588000 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 384.160 4.000 384.720 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.588000 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 416.640 4.000 417.200 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.588000 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 449.120 4.000 449.680 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal2 ;
        RECT 20.160 1221.000 20.720 1225.000 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal2 ;
        RECT 389.760 1221.000 390.320 1225.000 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal2 ;
        RECT 426.720 1221.000 427.280 1225.000 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal2 ;
        RECT 463.680 1221.000 464.240 1225.000 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal2 ;
        RECT 500.640 1221.000 501.200 1225.000 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal2 ;
        RECT 537.600 1221.000 538.160 1225.000 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal2 ;
        RECT 574.560 1221.000 575.120 1225.000 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.440000 ;
    PORT
      LAYER Metal2 ;
        RECT 611.520 1221.000 612.080 1225.000 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.440000 ;
    PORT
      LAYER Metal2 ;
        RECT 648.480 1221.000 649.040 1225.000 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.440000 ;
    PORT
      LAYER Metal2 ;
        RECT 685.440 1221.000 686.000 1225.000 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.440000 ;
    PORT
      LAYER Metal2 ;
        RECT 722.400 1221.000 722.960 1225.000 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal2 ;
        RECT 57.120 1221.000 57.680 1225.000 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.440000 ;
    PORT
      LAYER Metal2 ;
        RECT 759.360 1221.000 759.920 1225.000 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.440000 ;
    PORT
      LAYER Metal2 ;
        RECT 796.320 1221.000 796.880 1225.000 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.440000 ;
    PORT
      LAYER Metal2 ;
        RECT 833.280 1221.000 833.840 1225.000 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.607200 ;
    PORT
      LAYER Metal2 ;
        RECT 870.240 1221.000 870.800 1225.000 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.440000 ;
    PORT
      LAYER Metal2 ;
        RECT 907.200 1221.000 907.760 1225.000 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.440000 ;
    PORT
      LAYER Metal2 ;
        RECT 944.160 1221.000 944.720 1225.000 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.607200 ;
    PORT
      LAYER Metal2 ;
        RECT 981.120 1221.000 981.680 1225.000 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal2 ;
        RECT 1018.080 1221.000 1018.640 1225.000 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal2 ;
        RECT 1055.040 1221.000 1055.600 1225.000 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal2 ;
        RECT 1092.000 1221.000 1092.560 1225.000 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal2 ;
        RECT 94.080 1221.000 94.640 1225.000 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal2 ;
        RECT 1128.960 1221.000 1129.520 1225.000 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal2 ;
        RECT 1165.920 1221.000 1166.480 1225.000 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal2 ;
        RECT 1202.880 1221.000 1203.440 1225.000 ;
    END
  END io_oeb[32]
  PIN io_oeb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal2 ;
        RECT 131.040 1221.000 131.600 1225.000 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal2 ;
        RECT 168.000 1221.000 168.560 1225.000 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal2 ;
        RECT 204.960 1221.000 205.520 1225.000 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal2 ;
        RECT 241.920 1221.000 242.480 1225.000 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal2 ;
        RECT 278.880 1221.000 279.440 1225.000 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal2 ;
        RECT 315.840 1221.000 316.400 1225.000 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal2 ;
        RECT 352.800 1221.000 353.360 1225.000 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal2 ;
        RECT 20.160 0.000 20.720 4.000 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal2 ;
        RECT 389.760 0.000 390.320 4.000 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal2 ;
        RECT 426.720 0.000 427.280 4.000 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal2 ;
        RECT 463.680 0.000 464.240 4.000 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal2 ;
        RECT 500.640 0.000 501.200 4.000 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal2 ;
        RECT 537.600 0.000 538.160 4.000 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal2 ;
        RECT 574.560 0.000 575.120 4.000 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.237600 ;
    PORT
      LAYER Metal2 ;
        RECT 611.520 0.000 612.080 4.000 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.237600 ;
    PORT
      LAYER Metal2 ;
        RECT 648.480 0.000 649.040 4.000 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal2 ;
        RECT 685.440 0.000 686.000 4.000 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal2 ;
        RECT 722.400 0.000 722.960 4.000 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal2 ;
        RECT 57.120 0.000 57.680 4.000 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.237600 ;
    PORT
      LAYER Metal2 ;
        RECT 759.360 0.000 759.920 4.000 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.237600 ;
    PORT
      LAYER Metal2 ;
        RECT 796.320 0.000 796.880 4.000 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal2 ;
        RECT 833.280 0.000 833.840 4.000 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.440000 ;
    PORT
      LAYER Metal2 ;
        RECT 870.240 0.000 870.800 4.000 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal2 ;
        RECT 907.200 0.000 907.760 4.000 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal2 ;
        RECT 944.160 0.000 944.720 4.000 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.440000 ;
    PORT
      LAYER Metal2 ;
        RECT 981.120 0.000 981.680 4.000 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal2 ;
        RECT 1018.080 0.000 1018.640 4.000 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal2 ;
        RECT 1055.040 0.000 1055.600 4.000 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal2 ;
        RECT 1092.000 0.000 1092.560 4.000 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal2 ;
        RECT 94.080 0.000 94.640 4.000 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal2 ;
        RECT 1128.960 0.000 1129.520 4.000 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal2 ;
        RECT 1165.920 0.000 1166.480 4.000 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal2 ;
        RECT 1202.880 0.000 1203.440 4.000 ;
    END
  END io_out[32]
  PIN io_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal2 ;
        RECT 131.040 0.000 131.600 4.000 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal2 ;
        RECT 168.000 0.000 168.560 4.000 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal2 ;
        RECT 204.960 0.000 205.520 4.000 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal2 ;
        RECT 241.920 0.000 242.480 4.000 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal2 ;
        RECT 278.880 0.000 279.440 4.000 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal2 ;
        RECT 315.840 0.000 316.400 4.000 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.583500 ;
    PORT
      LAYER Metal2 ;
        RECT 352.800 0.000 353.360 4.000 ;
    END
  END io_out[9]
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.999200 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 59.360 4.000 59.920 ;
    END
  END rst_n
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 22.240 15.380 23.840 1207.660 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 175.840 15.380 177.440 1207.660 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 329.440 15.380 331.040 1207.660 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 483.040 15.380 484.640 1207.660 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 636.640 15.380 638.240 1207.660 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 790.240 15.380 791.840 1207.660 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 943.840 15.380 945.440 1207.660 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1097.440 15.380 1099.040 1207.660 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 99.040 15.380 100.640 1207.660 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 252.640 15.380 254.240 1207.660 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 406.240 15.380 407.840 1207.660 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 559.840 15.380 561.440 1207.660 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 713.440 15.380 715.040 1207.660 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 867.040 15.380 868.640 1207.660 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1020.640 15.380 1022.240 1207.660 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1174.240 15.380 1175.840 1207.660 ;
    END
  END vss
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.352000 ;
    ANTENNADIFFAREA 0.438500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 26.880 4.000 27.440 ;
    END
  END wb_clk_i
  OBS
      LAYER Nwell ;
        RECT 6.290 15.250 1218.430 1207.790 ;
      LAYER Metal1 ;
        RECT 6.720 4.070 1218.000 1209.450 ;
      LAYER Metal2 ;
        RECT 5.740 1220.700 19.860 1221.000 ;
        RECT 21.020 1220.700 56.820 1221.000 ;
        RECT 57.980 1220.700 93.780 1221.000 ;
        RECT 94.940 1220.700 130.740 1221.000 ;
        RECT 131.900 1220.700 167.700 1221.000 ;
        RECT 168.860 1220.700 204.660 1221.000 ;
        RECT 205.820 1220.700 241.620 1221.000 ;
        RECT 242.780 1220.700 278.580 1221.000 ;
        RECT 279.740 1220.700 315.540 1221.000 ;
        RECT 316.700 1220.700 352.500 1221.000 ;
        RECT 353.660 1220.700 389.460 1221.000 ;
        RECT 390.620 1220.700 426.420 1221.000 ;
        RECT 427.580 1220.700 463.380 1221.000 ;
        RECT 464.540 1220.700 500.340 1221.000 ;
        RECT 501.500 1220.700 537.300 1221.000 ;
        RECT 538.460 1220.700 574.260 1221.000 ;
        RECT 575.420 1220.700 611.220 1221.000 ;
        RECT 612.380 1220.700 648.180 1221.000 ;
        RECT 649.340 1220.700 685.140 1221.000 ;
        RECT 686.300 1220.700 722.100 1221.000 ;
        RECT 723.260 1220.700 759.060 1221.000 ;
        RECT 760.220 1220.700 796.020 1221.000 ;
        RECT 797.180 1220.700 832.980 1221.000 ;
        RECT 834.140 1220.700 869.940 1221.000 ;
        RECT 871.100 1220.700 906.900 1221.000 ;
        RECT 908.060 1220.700 943.860 1221.000 ;
        RECT 945.020 1220.700 980.820 1221.000 ;
        RECT 981.980 1220.700 1017.780 1221.000 ;
        RECT 1018.940 1220.700 1054.740 1221.000 ;
        RECT 1055.900 1220.700 1091.700 1221.000 ;
        RECT 1092.860 1220.700 1128.660 1221.000 ;
        RECT 1129.820 1220.700 1165.620 1221.000 ;
        RECT 1166.780 1220.700 1202.580 1221.000 ;
        RECT 1203.740 1220.700 1217.300 1221.000 ;
        RECT 5.740 4.300 1217.300 1220.700 ;
        RECT 5.740 4.000 19.860 4.300 ;
        RECT 21.020 4.000 56.820 4.300 ;
        RECT 57.980 4.000 93.780 4.300 ;
        RECT 94.940 4.000 130.740 4.300 ;
        RECT 131.900 4.000 167.700 4.300 ;
        RECT 168.860 4.000 204.660 4.300 ;
        RECT 205.820 4.000 241.620 4.300 ;
        RECT 242.780 4.000 278.580 4.300 ;
        RECT 279.740 4.000 315.540 4.300 ;
        RECT 316.700 4.000 352.500 4.300 ;
        RECT 353.660 4.000 389.460 4.300 ;
        RECT 390.620 4.000 426.420 4.300 ;
        RECT 427.580 4.000 463.380 4.300 ;
        RECT 464.540 4.000 500.340 4.300 ;
        RECT 501.500 4.000 537.300 4.300 ;
        RECT 538.460 4.000 574.260 4.300 ;
        RECT 575.420 4.000 611.220 4.300 ;
        RECT 612.380 4.000 648.180 4.300 ;
        RECT 649.340 4.000 685.140 4.300 ;
        RECT 686.300 4.000 722.100 4.300 ;
        RECT 723.260 4.000 759.060 4.300 ;
        RECT 760.220 4.000 796.020 4.300 ;
        RECT 797.180 4.000 832.980 4.300 ;
        RECT 834.140 4.000 869.940 4.300 ;
        RECT 871.100 4.000 906.900 4.300 ;
        RECT 908.060 4.000 943.860 4.300 ;
        RECT 945.020 4.000 980.820 4.300 ;
        RECT 981.980 4.000 1017.780 4.300 ;
        RECT 1018.940 4.000 1054.740 4.300 ;
        RECT 1055.900 4.000 1091.700 4.300 ;
        RECT 1092.860 4.000 1128.660 4.300 ;
        RECT 1129.820 4.000 1165.620 4.300 ;
        RECT 1166.780 4.000 1202.580 4.300 ;
        RECT 1203.740 4.000 1217.300 4.300 ;
      LAYER Metal3 ;
        RECT 4.000 1197.020 1217.350 1210.580 ;
        RECT 4.300 1195.860 1217.350 1197.020 ;
        RECT 4.000 1164.540 1217.350 1195.860 ;
        RECT 4.300 1163.380 1217.350 1164.540 ;
        RECT 4.000 1132.060 1217.350 1163.380 ;
        RECT 4.300 1130.900 1217.350 1132.060 ;
        RECT 4.000 1099.580 1217.350 1130.900 ;
        RECT 4.300 1098.420 1217.350 1099.580 ;
        RECT 4.000 1067.100 1217.350 1098.420 ;
        RECT 4.300 1065.940 1217.350 1067.100 ;
        RECT 4.000 1034.620 1217.350 1065.940 ;
        RECT 4.300 1033.460 1217.350 1034.620 ;
        RECT 4.000 1002.140 1217.350 1033.460 ;
        RECT 4.300 1000.980 1217.350 1002.140 ;
        RECT 4.000 969.660 1217.350 1000.980 ;
        RECT 4.300 968.500 1217.350 969.660 ;
        RECT 4.000 937.180 1217.350 968.500 ;
        RECT 4.300 936.020 1217.350 937.180 ;
        RECT 4.000 904.700 1217.350 936.020 ;
        RECT 4.300 903.540 1217.350 904.700 ;
        RECT 4.000 872.220 1217.350 903.540 ;
        RECT 4.300 871.060 1217.350 872.220 ;
        RECT 4.000 839.740 1217.350 871.060 ;
        RECT 4.300 838.580 1217.350 839.740 ;
        RECT 4.000 807.260 1217.350 838.580 ;
        RECT 4.300 806.100 1217.350 807.260 ;
        RECT 4.000 774.780 1217.350 806.100 ;
        RECT 4.300 773.620 1217.350 774.780 ;
        RECT 4.000 742.300 1217.350 773.620 ;
        RECT 4.300 741.140 1217.350 742.300 ;
        RECT 4.000 709.820 1217.350 741.140 ;
        RECT 4.300 708.660 1217.350 709.820 ;
        RECT 4.000 677.340 1217.350 708.660 ;
        RECT 4.300 676.180 1217.350 677.340 ;
        RECT 4.000 644.860 1217.350 676.180 ;
        RECT 4.300 643.700 1217.350 644.860 ;
        RECT 4.000 612.380 1217.350 643.700 ;
        RECT 4.300 611.220 1217.350 612.380 ;
        RECT 4.000 579.900 1217.350 611.220 ;
        RECT 4.300 578.740 1217.350 579.900 ;
        RECT 4.000 547.420 1217.350 578.740 ;
        RECT 4.300 546.260 1217.350 547.420 ;
        RECT 4.000 514.940 1217.350 546.260 ;
        RECT 4.300 513.780 1217.350 514.940 ;
        RECT 4.000 482.460 1217.350 513.780 ;
        RECT 4.300 481.300 1217.350 482.460 ;
        RECT 4.000 449.980 1217.350 481.300 ;
        RECT 4.300 448.820 1217.350 449.980 ;
        RECT 4.000 417.500 1217.350 448.820 ;
        RECT 4.300 416.340 1217.350 417.500 ;
        RECT 4.000 385.020 1217.350 416.340 ;
        RECT 4.300 383.860 1217.350 385.020 ;
        RECT 4.000 352.540 1217.350 383.860 ;
        RECT 4.300 351.380 1217.350 352.540 ;
        RECT 4.000 320.060 1217.350 351.380 ;
        RECT 4.300 318.900 1217.350 320.060 ;
        RECT 4.000 287.580 1217.350 318.900 ;
        RECT 4.300 286.420 1217.350 287.580 ;
        RECT 4.000 255.100 1217.350 286.420 ;
        RECT 4.300 253.940 1217.350 255.100 ;
        RECT 4.000 222.620 1217.350 253.940 ;
        RECT 4.300 221.460 1217.350 222.620 ;
        RECT 4.000 190.140 1217.350 221.460 ;
        RECT 4.300 188.980 1217.350 190.140 ;
        RECT 4.000 157.660 1217.350 188.980 ;
        RECT 4.300 156.500 1217.350 157.660 ;
        RECT 4.000 125.180 1217.350 156.500 ;
        RECT 4.300 124.020 1217.350 125.180 ;
        RECT 4.000 92.700 1217.350 124.020 ;
        RECT 4.300 91.540 1217.350 92.700 ;
        RECT 4.000 60.220 1217.350 91.540 ;
        RECT 4.300 59.060 1217.350 60.220 ;
        RECT 4.000 27.740 1217.350 59.060 ;
        RECT 4.300 26.580 1217.350 27.740 ;
        RECT 4.000 6.300 1217.350 26.580 ;
      LAYER Metal4 ;
        RECT 8.540 15.080 21.940 1204.470 ;
        RECT 24.140 15.080 98.740 1204.470 ;
        RECT 100.940 15.080 175.540 1204.470 ;
        RECT 177.740 15.080 252.340 1204.470 ;
        RECT 254.540 15.080 329.140 1204.470 ;
        RECT 331.340 15.080 405.940 1204.470 ;
        RECT 408.140 15.080 482.740 1204.470 ;
        RECT 484.940 15.080 559.540 1204.470 ;
        RECT 561.740 15.080 636.340 1204.470 ;
        RECT 638.540 15.080 713.140 1204.470 ;
        RECT 715.340 15.080 789.940 1204.470 ;
        RECT 792.140 15.080 866.740 1204.470 ;
        RECT 868.940 15.080 943.540 1204.470 ;
        RECT 945.740 15.080 1020.340 1204.470 ;
        RECT 1022.540 15.080 1097.140 1204.470 ;
        RECT 1099.340 15.080 1173.940 1204.470 ;
        RECT 1176.140 15.080 1208.340 1204.470 ;
        RECT 8.540 7.370 1208.340 15.080 ;
  END
END wrapped_tholin_riscv
END LIBRARY

