VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO wrapped_tholin_riscv
  CLASS BLOCK ;
  FOREIGN wrapped_tholin_riscv ;
  ORIGIN 0.000 0.000 ;
  SIZE 1000.000 BY 1100.000 ;
  PIN custom_settings[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 82.880 4.000 83.440 ;
    END
  END custom_settings[0]
  PIN custom_settings[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 112.000 4.000 112.560 ;
    END
  END custom_settings[1]
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 141.120 4.000 141.680 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 432.320 4.000 432.880 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 461.440 4.000 462.000 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 490.560 4.000 491.120 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 519.680 4.000 520.240 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 548.800 4.000 549.360 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 577.920 4.000 578.480 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 607.040 4.000 607.600 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 636.160 4.000 636.720 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 665.280 4.000 665.840 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 694.400 4.000 694.960 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 170.240 4.000 170.800 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 723.520 4.000 724.080 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 752.640 4.000 753.200 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 781.760 4.000 782.320 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 810.880 4.000 811.440 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 840.000 4.000 840.560 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 869.120 4.000 869.680 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 898.240 4.000 898.800 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 927.360 4.000 927.920 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 956.480 4.000 957.040 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 985.600 4.000 986.160 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 199.360 4.000 199.920 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1014.720 4.000 1015.280 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1043.840 4.000 1044.400 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1072.960 4.000 1073.520 ;
    END
  END io_in[32]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 228.480 4.000 229.040 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 257.600 4.000 258.160 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 286.720 4.000 287.280 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 315.840 4.000 316.400 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 344.960 4.000 345.520 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 374.080 4.000 374.640 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 403.200 4.000 403.760 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 15.680 1096.000 16.240 1100.000 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 318.080 1096.000 318.640 1100.000 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 348.320 1096.000 348.880 1100.000 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 378.560 1096.000 379.120 1100.000 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 408.800 1096.000 409.360 1100.000 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 439.040 1096.000 439.600 1100.000 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 469.280 1096.000 469.840 1100.000 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 499.520 1096.000 500.080 1100.000 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 529.760 1096.000 530.320 1100.000 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 560.000 1096.000 560.560 1100.000 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 590.240 1096.000 590.800 1100.000 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 45.920 1096.000 46.480 1100.000 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 620.480 1096.000 621.040 1100.000 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 650.720 1096.000 651.280 1100.000 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 680.960 1096.000 681.520 1100.000 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 711.200 1096.000 711.760 1100.000 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 741.440 1096.000 742.000 1100.000 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 771.680 1096.000 772.240 1100.000 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 801.920 1096.000 802.480 1100.000 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 832.160 1096.000 832.720 1100.000 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 862.400 1096.000 862.960 1100.000 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 892.640 1096.000 893.200 1100.000 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 76.160 1096.000 76.720 1100.000 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 922.880 1096.000 923.440 1100.000 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 953.120 1096.000 953.680 1100.000 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 983.360 1096.000 983.920 1100.000 ;
    END
  END io_oeb[32]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 106.400 1096.000 106.960 1100.000 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 136.640 1096.000 137.200 1100.000 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 166.880 1096.000 167.440 1100.000 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 197.120 1096.000 197.680 1100.000 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 227.360 1096.000 227.920 1100.000 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 257.600 1096.000 258.160 1100.000 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 287.840 1096.000 288.400 1100.000 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 15.680 0.000 16.240 4.000 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 318.080 0.000 318.640 4.000 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 348.320 0.000 348.880 4.000 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 378.560 0.000 379.120 4.000 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 408.800 0.000 409.360 4.000 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 439.040 0.000 439.600 4.000 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 469.280 0.000 469.840 4.000 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 499.520 0.000 500.080 4.000 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 529.760 0.000 530.320 4.000 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 560.000 0.000 560.560 4.000 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 590.240 0.000 590.800 4.000 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 45.920 0.000 46.480 4.000 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 620.480 0.000 621.040 4.000 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal2 ;
        RECT 650.720 0.000 651.280 4.000 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 680.960 0.000 681.520 4.000 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 711.200 0.000 711.760 4.000 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 741.440 0.000 742.000 4.000 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 771.680 0.000 772.240 4.000 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 801.920 0.000 802.480 4.000 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 832.160 0.000 832.720 4.000 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 862.400 0.000 862.960 4.000 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 892.640 0.000 893.200 4.000 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 76.160 0.000 76.720 4.000 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 922.880 0.000 923.440 4.000 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 953.120 0.000 953.680 4.000 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 983.360 0.000 983.920 4.000 ;
    END
  END io_out[32]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 106.400 0.000 106.960 4.000 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 136.640 0.000 137.200 4.000 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 166.880 0.000 167.440 4.000 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 197.120 0.000 197.680 4.000 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 227.360 0.000 227.920 4.000 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 257.600 0.000 258.160 4.000 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 287.840 0.000 288.400 4.000 ;
    END
  END io_out[9]
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 53.760 4.000 54.320 ;
    END
  END rst_n
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 22.240 15.380 23.840 1082.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 175.840 15.380 177.440 1082.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 329.440 15.380 331.040 1082.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 483.040 15.380 484.640 1082.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 636.640 15.380 638.240 1082.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 790.240 15.380 791.840 1082.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 943.840 15.380 945.440 1082.220 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 99.040 15.380 100.640 1082.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 252.640 15.380 254.240 1082.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 406.240 15.380 407.840 1082.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 559.840 15.380 561.440 1082.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 713.440 15.380 715.040 1082.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 867.040 15.380 868.640 1082.220 ;
    END
  END vss
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.738000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 24.640 4.000 25.200 ;
    END
  END wb_clk_i
  OBS
      LAYER Metal1 ;
        RECT 6.720 15.380 992.880 1082.220 ;
      LAYER Metal2 ;
        RECT 0.140 1095.700 15.380 1096.000 ;
        RECT 16.540 1095.700 45.620 1096.000 ;
        RECT 46.780 1095.700 75.860 1096.000 ;
        RECT 77.020 1095.700 106.100 1096.000 ;
        RECT 107.260 1095.700 136.340 1096.000 ;
        RECT 137.500 1095.700 166.580 1096.000 ;
        RECT 167.740 1095.700 196.820 1096.000 ;
        RECT 197.980 1095.700 227.060 1096.000 ;
        RECT 228.220 1095.700 257.300 1096.000 ;
        RECT 258.460 1095.700 287.540 1096.000 ;
        RECT 288.700 1095.700 317.780 1096.000 ;
        RECT 318.940 1095.700 348.020 1096.000 ;
        RECT 349.180 1095.700 378.260 1096.000 ;
        RECT 379.420 1095.700 408.500 1096.000 ;
        RECT 409.660 1095.700 438.740 1096.000 ;
        RECT 439.900 1095.700 468.980 1096.000 ;
        RECT 470.140 1095.700 499.220 1096.000 ;
        RECT 500.380 1095.700 529.460 1096.000 ;
        RECT 530.620 1095.700 559.700 1096.000 ;
        RECT 560.860 1095.700 589.940 1096.000 ;
        RECT 591.100 1095.700 620.180 1096.000 ;
        RECT 621.340 1095.700 650.420 1096.000 ;
        RECT 651.580 1095.700 680.660 1096.000 ;
        RECT 681.820 1095.700 710.900 1096.000 ;
        RECT 712.060 1095.700 741.140 1096.000 ;
        RECT 742.300 1095.700 771.380 1096.000 ;
        RECT 772.540 1095.700 801.620 1096.000 ;
        RECT 802.780 1095.700 831.860 1096.000 ;
        RECT 833.020 1095.700 862.100 1096.000 ;
        RECT 863.260 1095.700 892.340 1096.000 ;
        RECT 893.500 1095.700 922.580 1096.000 ;
        RECT 923.740 1095.700 952.820 1096.000 ;
        RECT 953.980 1095.700 983.060 1096.000 ;
        RECT 984.220 1095.700 993.860 1096.000 ;
        RECT 0.140 4.300 993.860 1095.700 ;
        RECT 0.140 2.890 15.380 4.300 ;
        RECT 16.540 2.890 45.620 4.300 ;
        RECT 46.780 2.890 75.860 4.300 ;
        RECT 77.020 2.890 106.100 4.300 ;
        RECT 107.260 2.890 136.340 4.300 ;
        RECT 137.500 2.890 166.580 4.300 ;
        RECT 167.740 2.890 196.820 4.300 ;
        RECT 197.980 2.890 227.060 4.300 ;
        RECT 228.220 2.890 257.300 4.300 ;
        RECT 258.460 2.890 287.540 4.300 ;
        RECT 288.700 2.890 317.780 4.300 ;
        RECT 318.940 2.890 348.020 4.300 ;
        RECT 349.180 2.890 378.260 4.300 ;
        RECT 379.420 2.890 408.500 4.300 ;
        RECT 409.660 2.890 438.740 4.300 ;
        RECT 439.900 2.890 468.980 4.300 ;
        RECT 470.140 2.890 499.220 4.300 ;
        RECT 500.380 2.890 529.460 4.300 ;
        RECT 530.620 2.890 559.700 4.300 ;
        RECT 560.860 2.890 589.940 4.300 ;
        RECT 591.100 2.890 620.180 4.300 ;
        RECT 621.340 2.890 650.420 4.300 ;
        RECT 651.580 2.890 680.660 4.300 ;
        RECT 681.820 2.890 710.900 4.300 ;
        RECT 712.060 2.890 741.140 4.300 ;
        RECT 742.300 2.890 771.380 4.300 ;
        RECT 772.540 2.890 801.620 4.300 ;
        RECT 802.780 2.890 831.860 4.300 ;
        RECT 833.020 2.890 862.100 4.300 ;
        RECT 863.260 2.890 892.340 4.300 ;
        RECT 893.500 2.890 922.580 4.300 ;
        RECT 923.740 2.890 952.820 4.300 ;
        RECT 953.980 2.890 983.060 4.300 ;
        RECT 984.220 2.890 993.860 4.300 ;
      LAYER Metal3 ;
        RECT 0.090 1073.820 993.910 1085.700 ;
        RECT 4.300 1072.660 993.910 1073.820 ;
        RECT 0.090 1044.700 993.910 1072.660 ;
        RECT 4.300 1043.540 993.910 1044.700 ;
        RECT 0.090 1015.580 993.910 1043.540 ;
        RECT 4.300 1014.420 993.910 1015.580 ;
        RECT 0.090 986.460 993.910 1014.420 ;
        RECT 4.300 985.300 993.910 986.460 ;
        RECT 0.090 957.340 993.910 985.300 ;
        RECT 4.300 956.180 993.910 957.340 ;
        RECT 0.090 928.220 993.910 956.180 ;
        RECT 4.300 927.060 993.910 928.220 ;
        RECT 0.090 899.100 993.910 927.060 ;
        RECT 4.300 897.940 993.910 899.100 ;
        RECT 0.090 869.980 993.910 897.940 ;
        RECT 4.300 868.820 993.910 869.980 ;
        RECT 0.090 840.860 993.910 868.820 ;
        RECT 4.300 839.700 993.910 840.860 ;
        RECT 0.090 811.740 993.910 839.700 ;
        RECT 4.300 810.580 993.910 811.740 ;
        RECT 0.090 782.620 993.910 810.580 ;
        RECT 4.300 781.460 993.910 782.620 ;
        RECT 0.090 753.500 993.910 781.460 ;
        RECT 4.300 752.340 993.910 753.500 ;
        RECT 0.090 724.380 993.910 752.340 ;
        RECT 4.300 723.220 993.910 724.380 ;
        RECT 0.090 695.260 993.910 723.220 ;
        RECT 4.300 694.100 993.910 695.260 ;
        RECT 0.090 666.140 993.910 694.100 ;
        RECT 4.300 664.980 993.910 666.140 ;
        RECT 0.090 637.020 993.910 664.980 ;
        RECT 4.300 635.860 993.910 637.020 ;
        RECT 0.090 607.900 993.910 635.860 ;
        RECT 4.300 606.740 993.910 607.900 ;
        RECT 0.090 578.780 993.910 606.740 ;
        RECT 4.300 577.620 993.910 578.780 ;
        RECT 0.090 549.660 993.910 577.620 ;
        RECT 4.300 548.500 993.910 549.660 ;
        RECT 0.090 520.540 993.910 548.500 ;
        RECT 4.300 519.380 993.910 520.540 ;
        RECT 0.090 491.420 993.910 519.380 ;
        RECT 4.300 490.260 993.910 491.420 ;
        RECT 0.090 462.300 993.910 490.260 ;
        RECT 4.300 461.140 993.910 462.300 ;
        RECT 0.090 433.180 993.910 461.140 ;
        RECT 4.300 432.020 993.910 433.180 ;
        RECT 0.090 404.060 993.910 432.020 ;
        RECT 4.300 402.900 993.910 404.060 ;
        RECT 0.090 374.940 993.910 402.900 ;
        RECT 4.300 373.780 993.910 374.940 ;
        RECT 0.090 345.820 993.910 373.780 ;
        RECT 4.300 344.660 993.910 345.820 ;
        RECT 0.090 316.700 993.910 344.660 ;
        RECT 4.300 315.540 993.910 316.700 ;
        RECT 0.090 287.580 993.910 315.540 ;
        RECT 4.300 286.420 993.910 287.580 ;
        RECT 0.090 258.460 993.910 286.420 ;
        RECT 4.300 257.300 993.910 258.460 ;
        RECT 0.090 229.340 993.910 257.300 ;
        RECT 4.300 228.180 993.910 229.340 ;
        RECT 0.090 200.220 993.910 228.180 ;
        RECT 4.300 199.060 993.910 200.220 ;
        RECT 0.090 171.100 993.910 199.060 ;
        RECT 4.300 169.940 993.910 171.100 ;
        RECT 0.090 141.980 993.910 169.940 ;
        RECT 4.300 140.820 993.910 141.980 ;
        RECT 0.090 112.860 993.910 140.820 ;
        RECT 4.300 111.700 993.910 112.860 ;
        RECT 0.090 83.740 993.910 111.700 ;
        RECT 4.300 82.580 993.910 83.740 ;
        RECT 0.090 54.620 993.910 82.580 ;
        RECT 4.300 53.460 993.910 54.620 ;
        RECT 0.090 25.500 993.910 53.460 ;
        RECT 4.300 24.340 993.910 25.500 ;
        RECT 0.090 2.940 993.910 24.340 ;
      LAYER Metal4 ;
        RECT 11.340 1082.520 989.380 1084.630 ;
        RECT 11.340 15.080 21.940 1082.520 ;
        RECT 24.140 15.080 98.740 1082.520 ;
        RECT 100.940 15.080 175.540 1082.520 ;
        RECT 177.740 15.080 252.340 1082.520 ;
        RECT 254.540 15.080 329.140 1082.520 ;
        RECT 331.340 15.080 405.940 1082.520 ;
        RECT 408.140 15.080 482.740 1082.520 ;
        RECT 484.940 15.080 559.540 1082.520 ;
        RECT 561.740 15.080 636.340 1082.520 ;
        RECT 638.540 15.080 713.140 1082.520 ;
        RECT 715.340 15.080 789.940 1082.520 ;
        RECT 792.140 15.080 866.740 1082.520 ;
        RECT 868.940 15.080 943.540 1082.520 ;
        RECT 945.740 15.080 989.380 1082.520 ;
        RECT 11.340 2.890 989.380 15.080 ;
  END
END wrapped_tholin_riscv
END LIBRARY

