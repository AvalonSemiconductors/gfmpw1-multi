VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO wrapped_ay8913
  CLASS BLOCK ;
  FOREIGN wrapped_ay8913 ;
  ORIGIN 0.000 0.000 ;
  SIZE 240.000 BY 240.000 ;
  PIN custom_settings[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 236.000 201.600 240.000 202.160 ;
    END
  END custom_settings[0]
  PIN custom_settings[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 236.000 225.120 240.000 225.680 ;
    END
  END custom_settings[1]
  PIN io_in_1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 236.000 13.440 240.000 14.000 ;
    END
  END io_in_1[0]
  PIN io_in_1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 236.000 36.960 240.000 37.520 ;
    END
  END io_in_1[1]
  PIN io_in_1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 236.000 60.480 240.000 61.040 ;
    END
  END io_in_1[2]
  PIN io_in_1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 236.000 84.000 240.000 84.560 ;
    END
  END io_in_1[3]
  PIN io_in_1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 236.000 107.520 240.000 108.080 ;
    END
  END io_in_1[4]
  PIN io_in_1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 236.000 131.040 240.000 131.600 ;
    END
  END io_in_1[5]
  PIN io_in_1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 236.000 154.560 240.000 155.120 ;
    END
  END io_in_1[6]
  PIN io_in_1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 236.000 178.080 240.000 178.640 ;
    END
  END io_in_1[7]
  PIN io_in_2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 148.960 236.000 149.520 240.000 ;
    END
  END io_in_2[0]
  PIN io_in_2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 208.320 236.000 208.880 240.000 ;
    END
  END io_in_2[1]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 13.440 0.000 14.000 4.000 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 91.840 0.000 92.400 4.000 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 99.680 0.000 100.240 4.000 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 107.520 0.000 108.080 4.000 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 115.360 0.000 115.920 4.000 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 123.200 0.000 123.760 4.000 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 131.040 0.000 131.600 4.000 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 138.880 0.000 139.440 4.000 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 146.720 0.000 147.280 4.000 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 154.560 0.000 155.120 4.000 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 162.400 0.000 162.960 4.000 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 21.280 0.000 21.840 4.000 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 170.240 0.000 170.800 4.000 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 178.080 0.000 178.640 4.000 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 185.920 0.000 186.480 4.000 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 193.760 0.000 194.320 4.000 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 201.600 0.000 202.160 4.000 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 209.440 0.000 210.000 4.000 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 217.280 0.000 217.840 4.000 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 225.120 0.000 225.680 4.000 ;
    END
  END io_out[27]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 29.120 0.000 29.680 4.000 ;
    END
  END io_out[2]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 36.960 0.000 37.520 4.000 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 44.800 0.000 45.360 4.000 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 52.640 0.000 53.200 4.000 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 60.480 0.000 61.040 4.000 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 68.320 0.000 68.880 4.000 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 76.160 0.000 76.720 4.000 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 84.000 0.000 84.560 4.000 ;
    END
  END io_out[9]
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 89.600 236.000 90.160 240.000 ;
    END
  END rst_n
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 22.240 15.380 23.840 223.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 175.840 15.380 177.440 223.740 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 99.040 15.380 100.640 223.740 ;
    END
  END vss
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.738000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 30.240 236.000 30.800 240.000 ;
    END
  END wb_clk_i
  OBS
      LAYER Nwell ;
        RECT 6.290 221.405 233.390 223.870 ;
        RECT 6.290 221.280 128.625 221.405 ;
      LAYER Pwell ;
        RECT 6.290 217.760 233.390 221.280 ;
      LAYER Nwell ;
        RECT 6.290 217.635 33.425 217.760 ;
        RECT 6.290 213.565 233.390 217.635 ;
        RECT 6.290 213.440 82.705 213.565 ;
      LAYER Pwell ;
        RECT 6.290 209.920 233.390 213.440 ;
      LAYER Nwell ;
        RECT 6.290 209.795 33.425 209.920 ;
        RECT 6.290 205.725 233.390 209.795 ;
        RECT 6.290 205.600 54.145 205.725 ;
      LAYER Pwell ;
        RECT 6.290 202.080 233.390 205.600 ;
      LAYER Nwell ;
        RECT 6.290 201.955 34.545 202.080 ;
        RECT 6.290 197.885 233.390 201.955 ;
        RECT 6.290 197.760 12.705 197.885 ;
      LAYER Pwell ;
        RECT 6.290 194.240 233.390 197.760 ;
      LAYER Nwell ;
        RECT 6.290 194.115 30.625 194.240 ;
        RECT 6.290 190.045 233.390 194.115 ;
        RECT 6.290 189.920 106.975 190.045 ;
      LAYER Pwell ;
        RECT 6.290 186.400 233.390 189.920 ;
      LAYER Nwell ;
        RECT 6.290 186.275 17.960 186.400 ;
        RECT 6.290 182.205 233.390 186.275 ;
        RECT 6.290 182.080 37.560 182.205 ;
      LAYER Pwell ;
        RECT 6.290 178.560 233.390 182.080 ;
      LAYER Nwell ;
        RECT 6.290 178.435 12.705 178.560 ;
        RECT 6.290 174.365 233.390 178.435 ;
        RECT 6.290 174.240 42.985 174.365 ;
      LAYER Pwell ;
        RECT 6.290 170.720 233.390 174.240 ;
      LAYER Nwell ;
        RECT 6.290 170.595 116.960 170.720 ;
        RECT 6.290 166.525 233.390 170.595 ;
        RECT 6.290 166.400 12.705 166.525 ;
      LAYER Pwell ;
        RECT 6.290 162.880 233.390 166.400 ;
      LAYER Nwell ;
        RECT 6.290 162.755 68.920 162.880 ;
        RECT 6.290 158.685 233.390 162.755 ;
        RECT 6.290 158.560 12.705 158.685 ;
      LAYER Pwell ;
        RECT 6.290 155.040 233.390 158.560 ;
      LAYER Nwell ;
        RECT 6.290 154.915 61.640 155.040 ;
        RECT 6.290 150.845 233.390 154.915 ;
        RECT 6.290 150.720 17.960 150.845 ;
      LAYER Pwell ;
        RECT 6.290 147.200 233.390 150.720 ;
      LAYER Nwell ;
        RECT 6.290 147.075 22.225 147.200 ;
        RECT 6.290 143.005 233.390 147.075 ;
        RECT 6.290 142.880 17.960 143.005 ;
      LAYER Pwell ;
        RECT 6.290 139.360 233.390 142.880 ;
      LAYER Nwell ;
        RECT 6.290 139.235 73.745 139.360 ;
        RECT 6.290 135.165 233.390 139.235 ;
        RECT 6.290 135.040 12.705 135.165 ;
      LAYER Pwell ;
        RECT 6.290 131.520 233.390 135.040 ;
      LAYER Nwell ;
        RECT 6.290 131.395 32.305 131.520 ;
        RECT 6.290 127.325 233.390 131.395 ;
        RECT 6.290 127.200 17.960 127.325 ;
      LAYER Pwell ;
        RECT 6.290 123.680 233.390 127.200 ;
      LAYER Nwell ;
        RECT 6.290 123.555 59.185 123.680 ;
        RECT 6.290 119.485 233.390 123.555 ;
        RECT 6.290 119.360 52.680 119.485 ;
      LAYER Pwell ;
        RECT 6.290 115.840 233.390 119.360 ;
      LAYER Nwell ;
        RECT 6.290 115.715 12.705 115.840 ;
        RECT 6.290 111.645 233.390 115.715 ;
        RECT 6.290 111.520 43.160 111.645 ;
      LAYER Pwell ;
        RECT 6.290 108.000 233.390 111.520 ;
      LAYER Nwell ;
        RECT 6.290 107.875 12.705 108.000 ;
        RECT 6.290 103.805 233.390 107.875 ;
        RECT 6.290 103.680 33.425 103.805 ;
      LAYER Pwell ;
        RECT 6.290 100.160 233.390 103.680 ;
      LAYER Nwell ;
        RECT 6.290 100.035 106.225 100.160 ;
        RECT 6.290 95.965 233.390 100.035 ;
        RECT 6.290 95.840 12.705 95.965 ;
      LAYER Pwell ;
        RECT 6.290 92.320 233.390 95.840 ;
      LAYER Nwell ;
        RECT 6.290 92.195 12.705 92.320 ;
        RECT 6.290 88.125 233.390 92.195 ;
        RECT 6.290 88.000 54.145 88.125 ;
      LAYER Pwell ;
        RECT 6.290 84.480 233.390 88.000 ;
      LAYER Nwell ;
        RECT 6.290 84.355 12.705 84.480 ;
        RECT 6.290 80.285 233.390 84.355 ;
        RECT 6.290 80.160 123.585 80.285 ;
      LAYER Pwell ;
        RECT 6.290 76.640 233.390 80.160 ;
      LAYER Nwell ;
        RECT 6.290 76.515 12.705 76.640 ;
        RECT 6.290 72.445 233.390 76.515 ;
        RECT 6.290 72.320 39.025 72.445 ;
      LAYER Pwell ;
        RECT 6.290 68.800 233.390 72.320 ;
      LAYER Nwell ;
        RECT 6.290 68.675 12.705 68.800 ;
        RECT 6.290 64.605 233.390 68.675 ;
        RECT 6.290 64.480 85.505 64.605 ;
      LAYER Pwell ;
        RECT 6.290 60.960 233.390 64.480 ;
      LAYER Nwell ;
        RECT 6.290 60.835 12.705 60.960 ;
        RECT 6.290 56.765 233.390 60.835 ;
        RECT 6.290 56.640 39.800 56.765 ;
      LAYER Pwell ;
        RECT 6.290 53.120 233.390 56.640 ;
      LAYER Nwell ;
        RECT 6.290 52.995 14.385 53.120 ;
        RECT 6.290 48.925 233.390 52.995 ;
        RECT 6.290 48.800 12.705 48.925 ;
      LAYER Pwell ;
        RECT 6.290 45.280 233.390 48.800 ;
      LAYER Nwell ;
        RECT 6.290 45.155 91.105 45.280 ;
        RECT 6.290 41.085 233.390 45.155 ;
        RECT 6.290 40.960 32.305 41.085 ;
      LAYER Pwell ;
        RECT 6.290 37.440 233.390 40.960 ;
      LAYER Nwell ;
        RECT 6.290 37.315 17.960 37.440 ;
        RECT 6.290 33.245 233.390 37.315 ;
        RECT 6.290 33.120 44.625 33.245 ;
      LAYER Pwell ;
        RECT 6.290 29.600 233.390 33.120 ;
      LAYER Nwell ;
        RECT 6.290 29.475 12.705 29.600 ;
        RECT 6.290 25.405 233.390 29.475 ;
        RECT 6.290 25.280 54.145 25.405 ;
      LAYER Pwell ;
        RECT 6.290 21.760 233.390 25.280 ;
      LAYER Nwell ;
        RECT 6.290 21.635 30.280 21.760 ;
        RECT 6.290 17.565 233.390 21.635 ;
        RECT 6.290 17.440 52.465 17.565 ;
      LAYER Pwell ;
        RECT 6.290 15.250 233.390 17.440 ;
      LAYER Metal1 ;
        RECT 6.720 15.380 232.960 224.410 ;
      LAYER Metal2 ;
        RECT 8.540 235.700 29.940 236.000 ;
        RECT 31.100 235.700 89.300 236.000 ;
        RECT 90.460 235.700 148.660 236.000 ;
        RECT 149.820 235.700 208.020 236.000 ;
        RECT 209.180 235.700 234.500 236.000 ;
        RECT 8.540 4.300 234.500 235.700 ;
        RECT 8.540 4.000 13.140 4.300 ;
        RECT 14.300 4.000 20.980 4.300 ;
        RECT 22.140 4.000 28.820 4.300 ;
        RECT 29.980 4.000 36.660 4.300 ;
        RECT 37.820 4.000 44.500 4.300 ;
        RECT 45.660 4.000 52.340 4.300 ;
        RECT 53.500 4.000 60.180 4.300 ;
        RECT 61.340 4.000 68.020 4.300 ;
        RECT 69.180 4.000 75.860 4.300 ;
        RECT 77.020 4.000 83.700 4.300 ;
        RECT 84.860 4.000 91.540 4.300 ;
        RECT 92.700 4.000 99.380 4.300 ;
        RECT 100.540 4.000 107.220 4.300 ;
        RECT 108.380 4.000 115.060 4.300 ;
        RECT 116.220 4.000 122.900 4.300 ;
        RECT 124.060 4.000 130.740 4.300 ;
        RECT 131.900 4.000 138.580 4.300 ;
        RECT 139.740 4.000 146.420 4.300 ;
        RECT 147.580 4.000 154.260 4.300 ;
        RECT 155.420 4.000 162.100 4.300 ;
        RECT 163.260 4.000 169.940 4.300 ;
        RECT 171.100 4.000 177.780 4.300 ;
        RECT 178.940 4.000 185.620 4.300 ;
        RECT 186.780 4.000 193.460 4.300 ;
        RECT 194.620 4.000 201.300 4.300 ;
        RECT 202.460 4.000 209.140 4.300 ;
        RECT 210.300 4.000 216.980 4.300 ;
        RECT 218.140 4.000 224.820 4.300 ;
        RECT 225.980 4.000 234.500 4.300 ;
      LAYER Metal3 ;
        RECT 8.490 224.820 235.700 225.540 ;
        RECT 8.490 202.460 236.740 224.820 ;
        RECT 8.490 201.300 235.700 202.460 ;
        RECT 8.490 178.940 236.740 201.300 ;
        RECT 8.490 177.780 235.700 178.940 ;
        RECT 8.490 155.420 236.740 177.780 ;
        RECT 8.490 154.260 235.700 155.420 ;
        RECT 8.490 131.900 236.740 154.260 ;
        RECT 8.490 130.740 235.700 131.900 ;
        RECT 8.490 108.380 236.740 130.740 ;
        RECT 8.490 107.220 235.700 108.380 ;
        RECT 8.490 84.860 236.740 107.220 ;
        RECT 8.490 83.700 235.700 84.860 ;
        RECT 8.490 61.340 236.740 83.700 ;
        RECT 8.490 60.180 235.700 61.340 ;
        RECT 8.490 37.820 236.740 60.180 ;
        RECT 8.490 36.660 235.700 37.820 ;
        RECT 8.490 14.300 236.740 36.660 ;
        RECT 8.490 13.580 235.700 14.300 ;
      LAYER Metal4 ;
        RECT 42.140 18.010 98.740 221.670 ;
        RECT 100.940 18.010 175.540 221.670 ;
        RECT 177.740 18.010 229.460 221.670 ;
  END
END wrapped_ay8913
END LIBRARY

